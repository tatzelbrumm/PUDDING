* NGSPICE file created from heichips25_pudding.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for analog_wires abstract view
.subckt analog_wires Iout VcascP[1] VcascP[0] i_in i_out
.ends

* Black-box entry subcircuit for dac128module abstract view
.subckt dac128module VbiasP[1] IOUT VbiasP[0] ON[64] ONB[64] ON[65] ONB[65] ON[66]
+ ONB[66] ON[67] ONB[67] ON[68] ONB[68] ON[69] ONB[69] ON[70] ONB[70] ON[71] ONB[71]
+ ON[72] ONB[72] EN[2] ENB[2] ON[73] ONB[73] ON[74] ONB[74] ON[75] ONB[75] ON[76]
+ ONB[76] ON[77] ONB[77] ON[78] ONB[78] ON[79] ONB[79] ON[80] ONB[80] ON[81] ONB[81]
+ ON[82] ONB[82] ON[83] ONB[83] ON[84] ONB[84] ON[85] ONB[85] ON[86] ONB[86] ON[87]
+ ONB[87] ON[88] ONB[88] ON[89] ONB[89] ON[90] ONB[90] ON[91] ONB[91] ON[92] ONB[92]
+ ON[93] ONB[93] ON[94] ONB[94] ON[95] ONB[95] ON[96] ONB[96] ON[97] ONB[97] ON[98]
+ ONB[98] ON[99] ONB[99] ON[100] ONB[100] ON[101] ONB[101] ON[102] ONB[102] ON[103]
+ ONB[103] ON[104] ONB[104] ON[105] ONB[105] ON[106] ONB[106] ON[107] ONB[107] ON[108]
+ ONB[108] ON[109] ONB[109] ON[110] ONB[110] ON[111] ONB[111] ON[112] ONB[112] ON[113]
+ ONB[113] ON[114] ONB[114] ON[115] ONB[115] ON[116] ONB[116] ON[117] ONB[117] ON[118]
+ ONB[118] ON[119] ONB[119] ON[120] ONB[120] ON[121] ONB[121] ON[122] ONB[122] EN[3]
+ ENB[3] ON[123] ONB[123] ON[124] ONB[124] ON[125] ONB[125] ON[126] ONB[126] ON[127]
+ ONB[127] ON[0] ONB[0] ON[1] ONB[1] ON[2] ONB[2] ON[3] ONB[3] ON[4] ONB[4] ON[5]
+ ONB[5] ON[6] EN[0] ENB[0] ONB[6] ON[7] ONB[7] ON[8] ONB[8] ON[9] ONB[9] ON[10] ONB[10]
+ ON[11] ONB[11] ON[12] ONB[12] ON[13] ONB[13] ON[14] ONB[14] ON[15] ONB[15] ON[16]
+ ONB[16] ON[17] ONB[17] ON[18] ONB[18] ON[19] ONB[19] ON[20] ONB[20] ON[21] ONB[21]
+ ON[22] ONB[22] ON[23] ONB[23] ON[24] ONB[24] ON[25] ONB[25] ON[26] ONB[26] ON[27]
+ ONB[27] ON[28] ONB[28] ON[29] ONB[29] ON[30] ONB[30] ON[31] ONB[31] ON[33] ONB[33]
+ ON[32] ONB[32] ON[34] ONB[34] ON[35] ONB[35] ON[36] ONB[36] ON[37] ONB[37] ON[38]
+ ONB[38] ON[39] ONB[39] ON[40] ONB[40] ON[41] ONB[41] ON[42] ONB[42] ON[43] ONB[43]
+ ON[44] ONB[44] ON[45] ONB[45] ON[46] ONB[46] ON[47] ONB[47] ON[48] ONB[48] ON[49]
+ ONB[49] ON[50] ONB[50] ON[51] ONB[51] ON[52] ONB[52] ON[53] ONB[53] ON[54] ONB[54]
+ ON[55] ONB[55] ON[56] ONB[56] ON[57] ONB[57] ON[58] ONB[58] ON[59] ONB[59] ON[60]
+ ONB[60] ON[61] ONB[61] ON[62] ONB[62] ON[63] ONB[63] EN[1] ENB[1] VcascP[1] VcascP[0]
+ VSS VDD
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

.subckt heichips25_pudding VGND VPWR clk ena i_in i_out rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_233 VPWR VGND sg13g2_decap_8
X_2106_ _0743_ net104 state\[25\] VPWR VGND sg13g2_nand2_1
X_2037_ _0703_ net154 _0702_ VPWR VGND sg13g2_nand2_1
XFILLER_10_328 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_35_483 VPWR VGND sg13g2_decap_8
X_2537__318 VPWR VGND net317 sg13g2_tiehi
XFILLER_41_431 VPWR VGND sg13g2_fill_2
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_41_497 VPWR VGND sg13g2_fill_1
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_5_321 VPWR VGND sg13g2_decap_8
XFILLER_9_148 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_5_398 VPWR VGND sg13g2_decap_8
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_37_726 VPWR VGND sg13g2_fill_1
XFILLER_37_737 VPWR VGND sg13g2_fill_1
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_20_615 VPWR VGND sg13g2_fill_1
XFILLER_20_648 VPWR VGND sg13g2_fill_1
XFILLER_32_475 VPWR VGND sg13g2_decap_4
XFILLER_44_280 VPWR VGND sg13g2_decap_8
X_1606_ state\[38\] daisychain\[38\] net139 _1002_ VPWR VGND sg13g2_mux2_1
X_1399_ VPWR _0032_ state\[13\] VGND sg13g2_inv_1
X_1468_ VGND VPWR net91 daisychain\[9\] _0892_ net45 sg13g2_a21oi_1
X_1537_ _0947_ net161 _0946_ VPWR VGND sg13g2_nand2_1
Xfanout105 net106 net105 VPWR VGND sg13g2_buf_1
Xfanout116 net118 net116 VPWR VGND sg13g2_buf_1
Xfanout127 net129 net127 VPWR VGND sg13g2_buf_1
Xfanout138 net140 net138 VPWR VGND sg13g2_buf_1
Xfanout149 net152 net149 VPWR VGND sg13g2_buf_1
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_10_125 VPWR VGND sg13g2_decap_8
XFILLER_11_604 VPWR VGND sg13g2_decap_8
XFILLER_11_615 VPWR VGND sg13g2_fill_2
XFILLER_23_475 VPWR VGND sg13g2_decap_8
XFILLER_23_486 VPWR VGND sg13g2_decap_8
XFILLER_2_357 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_fill_2
X_2504__328 VPWR VGND net327 sg13g2_tiehi
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_19_715 VPWR VGND sg13g2_decap_8
XFILLER_19_726 VPWR VGND sg13g2_fill_2
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_46_523 VPWR VGND sg13g2_fill_1
XFILLER_14_486 VPWR VGND sg13g2_fill_2
XFILLER_33_228 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
X_2440_ net326 VGND VPWR _0256_ state\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_5_195 VPWR VGND sg13g2_decap_8
X_1322_ VPWR _0117_ state\[90\] VGND sg13g2_inv_1
X_2371_ net208 VGND VPWR _0187_ daisychain\[59\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_33_773 VPWR VGND sg13g2_fill_1
XFILLER_0_806 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_4
XFILLER_23_53 VPWR VGND sg13g2_decap_8
X_2467__220 VPWR VGND net219 sg13g2_tiehi
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_3_666 VPWR VGND sg13g2_fill_2
X_2521__450 VPWR VGND net449 sg13g2_tiehi
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_589 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
X_2370__211 VPWR VGND net210 sg13g2_tiehi
XFILLER_14_294 VPWR VGND sg13g2_decap_8
XFILLER_15_740 VPWR VGND sg13g2_fill_2
XFILLER_30_710 VPWR VGND sg13g2_fill_1
XFILLER_30_743 VPWR VGND sg13g2_fill_1
XFILLER_30_776 VPWR VGND sg13g2_fill_2
XFILLER_9_99 VPWR VGND sg13g2_decap_8
X_2446__304 VPWR VGND net303 sg13g2_tiehi
X_1940_ VGND VPWR _0623_ _0624_ _0232_ _0625_ sg13g2_a21oi_1
X_1871_ state\[91\] daisychain\[91\] net148 _0570_ VPWR VGND sg13g2_mux2_1
X_2423_ net360 VGND VPWR _0239_ daisychain\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1305_ VPWR _0008_ state\[107\] VGND sg13g2_inv_1
X_2354_ net242 VGND VPWR _0170_ daisychain\[42\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2285_ VGND VPWR _0663_ _0832_ _0370_ net69 sg13g2_a21oi_1
XFILLER_25_504 VPWR VGND sg13g2_decap_8
XFILLER_37_364 VPWR VGND sg13g2_decap_8
X_2533__354 VPWR VGND net353 sg13g2_tiehi
XFILLER_33_592 VPWR VGND sg13g2_decap_8
X_2347__257 VPWR VGND net256 sg13g2_tiehi
XFILLER_0_636 VPWR VGND sg13g2_fill_2
XFILLER_18_42 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_11_264 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_8
XFILLER_7_235 VPWR VGND sg13g2_decap_8
X_2070_ _0725_ net92 state\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_19_397 VPWR VGND sg13g2_decap_8
XFILLER_22_507 VPWR VGND sg13g2_decap_8
XFILLER_34_301 VPWR VGND sg13g2_decap_8
XFILLER_34_356 VPWR VGND sg13g2_decap_4
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_47_673 VPWR VGND sg13g2_decap_8
XFILLER_30_584 VPWR VGND sg13g2_fill_2
X_1923_ VGND VPWR net112 daisychain\[100\] _0612_ net54 sg13g2_a21oi_1
X_1854_ net187 VPWR _0557_ VGND daisychain\[87\] net32 sg13g2_o21ai_1
X_1785_ VGND VPWR _0499_ _0500_ _0201_ _0501_ sg13g2_a21oi_1
X_2406_ net394 VGND VPWR _0222_ daisychain\[94\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_25_312 VPWR VGND sg13g2_fill_1
XFILLER_37_161 VPWR VGND sg13g2_decap_8
XFILLER_38_640 VPWR VGND sg13g2_decap_8
X_2337_ net276 VGND VPWR _0153_ daisychain\[25\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2268_ _0824_ net108 state\[106\] VPWR VGND sg13g2_nand2_1
X_2199_ VGND VPWR _0491_ _0789_ _0327_ net86 sg13g2_a21oi_1
XFILLER_25_367 VPWR VGND sg13g2_decap_4
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_4_227 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_29_52 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_17_813 VPWR VGND sg13g2_decap_8
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_decap_4
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_12_551 VPWR VGND sg13g2_decap_4
XFILLER_12_562 VPWR VGND sg13g2_fill_1
XFILLER_31_359 VPWR VGND sg13g2_fill_1
XFILLER_4_750 VPWR VGND sg13g2_decap_8
XFILLER_6_89 VPWR VGND sg13g2_decap_8
X_1570_ VGND VPWR _0971_ _0972_ _0158_ _0973_ sg13g2_a21oi_1
XFILLER_19_183 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_2122_ _0751_ net106 state\[33\] VPWR VGND sg13g2_nand2_1
X_2053_ VGND VPWR net90 daisychain\[126\] _0716_ net48 sg13g2_a21oi_1
XFILLER_22_304 VPWR VGND sg13g2_decap_8
XFILLER_34_175 VPWR VGND sg13g2_decap_8
XFILLER_35_665 VPWR VGND sg13g2_fill_2
X_1906_ state\[98\] daisychain\[98\] net143 _0598_ VPWR VGND sg13g2_mux2_1
X_1837_ _0543_ net172 _0542_ VPWR VGND sg13g2_nand2_1
X_1768_ VGND VPWR net128 daisychain\[69\] _0488_ net64 sg13g2_a21oi_1
X_2498__352 VPWR VGND net351 sg13g2_tiehi
X_1699_ net192 VPWR _0433_ VGND daisychain\[56\] net37 sg13g2_o21ai_1
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_13_337 VPWR VGND sg13g2_fill_2
XFILLER_15_65 VPWR VGND sg13g2_decap_8
XFILLER_31_53 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_41_657 VPWR VGND sg13g2_fill_1
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_49_702 VPWR VGND sg13g2_fill_2
X_2477__436 VPWR VGND net435 sg13g2_tiehi
XFILLER_16_142 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_fill_2
XFILLER_31_123 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_8
XFILLER_40_690 VPWR VGND sg13g2_fill_2
XFILLER_8_396 VPWR VGND sg13g2_decap_8
X_1622_ _1015_ net168 _1014_ VPWR VGND sg13g2_nand2_1
XFILLER_39_212 VPWR VGND sg13g2_decap_8
X_1484_ net179 VPWR _0905_ VGND daisychain\[13\] net23 sg13g2_o21ai_1
X_1553_ VGND VPWR net100 daisychain\[26\] _0960_ net49 sg13g2_a21oi_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
XFILLER_35_462 VPWR VGND sg13g2_fill_1
XFILLER_39_289 VPWR VGND sg13g2_decap_8
X_2105_ VGND VPWR _0947_ _0742_ _0280_ net72 sg13g2_a21oi_1
X_2036_ state\[124\] daisychain\[124\] net136 _0702_ VPWR VGND sg13g2_mux2_1
XFILLER_10_307 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_7_8 VPWR VGND sg13g2_fill_1
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_14_657 VPWR VGND sg13g2_decap_8
XFILLER_14_668 VPWR VGND sg13g2_fill_1
XFILLER_26_451 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_5_300 VPWR VGND sg13g2_decap_8
XFILLER_9_127 VPWR VGND sg13g2_decap_8
XFILLER_5_377 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_49_587 VPWR VGND sg13g2_fill_2
XFILLER_20_627 VPWR VGND sg13g2_fill_1
XFILLER_32_498 VPWR VGND sg13g2_fill_2
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_1536_ state\[24\] daisychain\[24\] net139 _0946_ VPWR VGND sg13g2_mux2_1
X_1605_ VGND VPWR _0999_ _1000_ _0165_ _1001_ sg13g2_a21oi_1
X_1398_ VPWR _0033_ state\[14\] VGND sg13g2_inv_1
X_1467_ _0891_ net155 _0890_ VPWR VGND sg13g2_nand2_1
X_2536__330 VPWR VGND net329 sg13g2_tiehi
Xfanout106 net132 net106 VPWR VGND sg13g2_buf_1
Xfanout117 net118 net117 VPWR VGND sg13g2_buf_1
Xfanout128 net129 net128 VPWR VGND sg13g2_buf_1
Xfanout139 net140 net139 VPWR VGND sg13g2_buf_1
XFILLER_27_259 VPWR VGND sg13g2_decap_4
XFILLER_43_708 VPWR VGND sg13g2_fill_2
X_2019_ net199 VPWR _0689_ VGND daisychain\[120\] net26 sg13g2_o21ai_1
XFILLER_10_104 VPWR VGND sg13g2_decap_8
XFILLER_12_99 VPWR VGND sg13g2_decap_8
XFILLER_2_336 VPWR VGND sg13g2_decap_8
XFILLER_33_207 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_46_568 VPWR VGND sg13g2_decap_8
X_2357__237 VPWR VGND net236 sg13g2_tiehi
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_5_174 VPWR VGND sg13g2_decap_8
XFILLER_6_653 VPWR VGND sg13g2_decap_4
XFILLER_49_340 VPWR VGND sg13g2_decap_8
X_1321_ VPWR _0118_ state\[91\] VGND sg13g2_inv_1
X_2559__374 VPWR VGND net373 sg13g2_tiehi
X_2370_ net210 VGND VPWR _0186_ daisychain\[58\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_17_281 VPWR VGND sg13g2_fill_2
XFILLER_18_782 VPWR VGND sg13g2_decap_8
XFILLER_18_793 VPWR VGND sg13g2_fill_1
XFILLER_33_752 VPWR VGND sg13g2_fill_2
XFILLER_37_579 VPWR VGND sg13g2_decap_8
XFILLER_20_468 VPWR VGND sg13g2_decap_8
XFILLER_20_479 VPWR VGND sg13g2_decap_8
XFILLER_32_284 VPWR VGND sg13g2_decap_8
X_1519_ net182 VPWR _0933_ VGND daisychain\[20\] net27 sg13g2_o21ai_1
X_2499_ net347 VGND VPWR _0315_ state\[59\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_16_708 VPWR VGND sg13g2_decap_8
XFILLER_28_524 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_7_417 VPWR VGND sg13g2_decap_8
XFILLER_7_428 VPWR VGND sg13g2_fill_1
XFILLER_19_513 VPWR VGND sg13g2_fill_1
XFILLER_2_133 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_557 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_14_273 VPWR VGND sg13g2_decap_8
XFILLER_30_755 VPWR VGND sg13g2_fill_2
XFILLER_42_571 VPWR VGND sg13g2_fill_2
XFILLER_9_78 VPWR VGND sg13g2_decap_8
X_1870_ VGND VPWR _0567_ _0568_ _0218_ _0569_ sg13g2_a21oi_1
X_2422_ net362 VGND VPWR _0238_ daisychain\[110\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2353_ net244 VGND VPWR _0169_ daisychain\[41\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
X_1304_ VPWR _0009_ state\[108\] VGND sg13g2_inv_1
X_2284_ _0832_ net95 state\[114\] VPWR VGND sg13g2_nand2_1
XFILLER_37_398 VPWR VGND sg13g2_decap_8
XFILLER_20_243 VPWR VGND sg13g2_decap_8
XFILLER_20_287 VPWR VGND sg13g2_fill_1
XFILLER_4_409 VPWR VGND sg13g2_decap_8
X_1999_ net180 VPWR _0673_ VGND daisychain\[116\] net24 sg13g2_o21ai_1
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_11_243 VPWR VGND sg13g2_decap_8
XFILLER_12_733 VPWR VGND sg13g2_fill_2
XFILLER_12_744 VPWR VGND sg13g2_fill_2
XFILLER_12_766 VPWR VGND sg13g2_fill_1
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_7_214 VPWR VGND sg13g2_decap_8
XFILLER_3_420 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_47_641 VPWR VGND sg13g2_decap_4
XFILLER_15_582 VPWR VGND sg13g2_decap_8
X_2491__380 VPWR VGND net379 sg13g2_tiehi
X_1922_ _0611_ net165 _0610_ VPWR VGND sg13g2_nand2_1
XFILLER_30_563 VPWR VGND sg13g2_fill_1
X_1853_ VGND VPWR net111 daisychain\[86\] _0556_ net54 sg13g2_a21oi_1
X_1784_ net195 VPWR _0501_ VGND daisychain\[73\] net40 sg13g2_o21ai_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_2405_ net396 VGND VPWR _0221_ daisychain\[93\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2336_ net278 VGND VPWR _0152_ daisychain\[24\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_29_129 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
X_2267_ VGND VPWR _0627_ _0823_ _0361_ net75 sg13g2_a21oi_1
X_2198_ _0789_ net129 state\[71\] VPWR VGND sg13g2_nand2_1
XFILLER_4_206 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_29_31 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_44_633 VPWR VGND sg13g2_fill_1
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_39_405 VPWR VGND sg13g2_fill_1
XFILLER_39_416 VPWR VGND sg13g2_fill_1
XFILLER_3_294 VPWR VGND sg13g2_decap_8
XFILLER_6_68 VPWR VGND sg13g2_decap_8
X_2558__406 VPWR VGND net405 sg13g2_tiehi
XFILLER_19_162 VPWR VGND sg13g2_decap_8
XFILLER_35_611 VPWR VGND sg13g2_fill_1
XFILLER_35_644 VPWR VGND sg13g2_decap_8
XFILLER_39_427 VPWR VGND sg13g2_fill_1
X_2121_ VGND VPWR _0979_ _0750_ _0288_ net73 sg13g2_a21oi_1
X_2052_ _0715_ net154 _0714_ VPWR VGND sg13g2_nand2_1
XFILLER_34_154 VPWR VGND sg13g2_decap_8
X_1905_ VGND VPWR _0595_ _0596_ _0225_ _0597_ sg13g2_a21oi_1
X_1836_ state\[84\] daisychain\[84\] net148 _0542_ VPWR VGND sg13g2_mux2_1
X_1767_ _0487_ net175 _0486_ VPWR VGND sg13g2_nand2_1
X_1698_ VGND VPWR net119 daisychain\[55\] _0432_ net59 sg13g2_a21oi_1
X_2319_ net312 VGND VPWR _0135_ daisychain\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_33 VPWR VGND sg13g2_decap_8
XFILLER_25_187 VPWR VGND sg13g2_decap_8
XFILLER_38_482 VPWR VGND sg13g2_decap_8
XFILLER_38_493 VPWR VGND sg13g2_fill_1
X_2316__319 VPWR VGND net318 sg13g2_tiehi
XFILLER_21_382 VPWR VGND sg13g2_fill_1
XFILLER_31_32 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_9_309 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_5_559 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_16_121 VPWR VGND sg13g2_decap_8
XFILLER_29_493 VPWR VGND sg13g2_decap_8
XFILLER_36_419 VPWR VGND sg13g2_fill_2
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_49_736 VPWR VGND sg13g2_decap_8
XFILLER_12_360 VPWR VGND sg13g2_decap_8
XFILLER_16_198 VPWR VGND sg13g2_decap_8
XFILLER_31_102 VPWR VGND sg13g2_decap_8
XFILLER_31_179 VPWR VGND sg13g2_decap_8
XFILLER_32_658 VPWR VGND sg13g2_fill_1
X_2484__408 VPWR VGND net407 sg13g2_tiehi
X_2367__217 VPWR VGND net216 sg13g2_tiehi
XFILLER_8_375 VPWR VGND sg13g2_decap_8
X_1552_ _0959_ net160 _0958_ VPWR VGND sg13g2_nand2_1
X_1621_ state\[41\] daisychain\[41\] net144 _1014_ VPWR VGND sg13g2_mux2_1
XFILLER_39_268 VPWR VGND sg13g2_decap_8
X_1483_ VGND VPWR net93 daisychain\[12\] _0904_ net45 sg13g2_a21oi_1
X_2104_ _0742_ net104 state\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_22_102 VPWR VGND sg13g2_decap_8
X_2035_ VGND VPWR _0699_ _0700_ _0251_ _0701_ sg13g2_a21oi_1
XFILLER_22_179 VPWR VGND sg13g2_decap_8
X_1819_ net194 VPWR _0529_ VGND daisychain\[80\] net39 sg13g2_o21ai_1
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_26_76 VPWR VGND sg13g2_decap_8
XFILLER_41_444 VPWR VGND sg13g2_decap_4
XFILLER_41_466 VPWR VGND sg13g2_decap_8
XFILLER_41_488 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_9_106 VPWR VGND sg13g2_decap_8
XFILLER_5_356 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_12_190 VPWR VGND sg13g2_decap_8
XFILLER_13_680 VPWR VGND sg13g2_decap_8
XFILLER_20_639 VPWR VGND sg13g2_fill_1
XFILLER_8_172 VPWR VGND sg13g2_decap_8
X_1535_ VGND VPWR _0943_ _0944_ _0151_ _0945_ sg13g2_a21oi_1
Xfanout107 net109 net107 VPWR VGND sg13g2_buf_1
Xfanout118 net132 net118 VPWR VGND sg13g2_buf_1
Xfanout129 net131 net129 VPWR VGND sg13g2_buf_1
X_1604_ net183 VPWR _1001_ VGND daisychain\[37\] net28 sg13g2_o21ai_1
XFILLER_27_238 VPWR VGND sg13g2_decap_8
X_1397_ VPWR _0034_ state\[15\] VGND sg13g2_inv_1
X_1466_ state\[10\] daisychain\[10\] net133 _0890_ VPWR VGND sg13g2_mux2_1
X_2018_ VGND VPWR net97 daisychain\[119\] _0688_ net47 sg13g2_a21oi_1
XFILLER_12_34 VPWR VGND sg13g2_decap_4
XFILLER_12_78 VPWR VGND sg13g2_decap_8
XFILLER_2_315 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_19_739 VPWR VGND sg13g2_decap_8
XFILLER_26_260 VPWR VGND sg13g2_fill_2
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_14_466 VPWR VGND sg13g2_fill_1
XFILLER_14_499 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_6_621 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_153 VPWR VGND sg13g2_decap_8
X_1320_ VPWR _0119_ state\[92\] VGND sg13g2_inv_1
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_17_260 VPWR VGND sg13g2_decap_8
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_33_764 VPWR VGND sg13g2_decap_8
XFILLER_37_569 VPWR VGND sg13g2_fill_2
X_1449_ net182 VPWR _0877_ VGND daisychain\[6\] net27 sg13g2_o21ai_1
X_1518_ VGND VPWR net99 daisychain\[19\] _0932_ net49 sg13g2_a21oi_1
X_2567_ net453 VGND VPWR _0383_ state\[127\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2498_ net351 VGND VPWR _0314_ state\[58\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_15_219 VPWR VGND sg13g2_decap_8
XFILLER_43_517 VPWR VGND sg13g2_fill_1
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_14_252 VPWR VGND sg13g2_decap_8
XFILLER_15_742 VPWR VGND sg13g2_fill_1
XFILLER_15_775 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_30_789 VPWR VGND sg13g2_decap_4
XFILLER_2_690 VPWR VGND sg13g2_decap_8
X_1303_ VPWR _0010_ state\[109\] VGND sg13g2_inv_1
X_2421_ net364 VGND VPWR _0237_ daisychain\[109\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2352_ net246 VGND VPWR _0168_ daisychain\[40\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2283_ VGND VPWR _0659_ _0831_ _0369_ net69 sg13g2_a21oi_1
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_38_812 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_20_222 VPWR VGND sg13g2_decap_8
XFILLER_33_561 VPWR VGND sg13g2_fill_2
X_1998_ VGND VPWR net94 daisychain\[115\] _0672_ net46 sg13g2_a21oi_1
XFILLER_0_616 VPWR VGND sg13g2_fill_1
XFILLER_0_638 VPWR VGND sg13g2_fill_1
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_fill_1
XFILLER_16_539 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_28_366 VPWR VGND sg13g2_decap_4
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_11_222 VPWR VGND sg13g2_decap_8
XFILLER_11_299 VPWR VGND sg13g2_decap_8
XFILLER_12_778 VPWR VGND sg13g2_fill_2
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_19_300 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_decap_8
X_2376__455 VPWR VGND net454 sg13g2_tiehi
XFILLER_46_196 VPWR VGND sg13g2_decap_8
X_1921_ state\[101\] daisychain\[101\] net142 _0610_ VPWR VGND sg13g2_mux2_1
X_1852_ _0555_ net165 _0554_ VPWR VGND sg13g2_nand2_1
XFILLER_30_597 VPWR VGND sg13g2_fill_1
XFILLER_6_281 VPWR VGND sg13g2_decap_8
XFILLER_7_771 VPWR VGND sg13g2_decap_8
X_1783_ VGND VPWR net127 daisychain\[72\] _0500_ net63 sg13g2_a21oi_1
XFILLER_29_108 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_2500__344 VPWR VGND net343 sg13g2_tiehi
X_2404_ net398 VGND VPWR _0220_ daisychain\[92\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2335_ net280 VGND VPWR _0151_ daisychain\[23\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2266_ _0823_ net107 state\[105\] VPWR VGND sg13g2_nand2_1
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_38_653 VPWR VGND sg13g2_decap_8
XFILLER_41_807 VPWR VGND sg13g2_decap_8
X_2197_ VGND VPWR _0487_ _0788_ _0326_ net86 sg13g2_a21oi_1
XFILLER_5_708 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_20_89 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_29_87 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_16_369 VPWR VGND sg13g2_fill_1
XFILLER_24_391 VPWR VGND sg13g2_decap_4
XFILLER_32_818 VPWR VGND sg13g2_decap_4
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_44_645 VPWR VGND sg13g2_fill_2
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_6_47 VPWR VGND sg13g2_fill_2
XFILLER_3_273 VPWR VGND sg13g2_decap_8
XFILLER_4_796 VPWR VGND sg13g2_fill_2
X_2120_ _0750_ net106 state\[32\] VPWR VGND sg13g2_nand2_1
XFILLER_19_141 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
X_2051_ state\[127\] daisychain\[127\] net136 _0714_ VPWR VGND sg13g2_mux2_1
X_1904_ net187 VPWR _0597_ VGND daisychain\[97\] net32 sg13g2_o21ai_1
X_1835_ VGND VPWR _0539_ _0540_ _0211_ _0541_ sg13g2_a21oi_1
X_1766_ state\[70\] daisychain\[70\] net151 _0486_ VPWR VGND sg13g2_mux2_1
X_1697_ _0431_ net170 _0430_ VPWR VGND sg13g2_nand2_1
X_2318_ net314 VGND VPWR _0134_ daisychain\[6\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2249_ VGND VPWR _0591_ _0814_ _0352_ net77 sg13g2_a21oi_1
XFILLER_25_111 VPWR VGND sg13g2_fill_1
XFILLER_25_166 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_41_637 VPWR VGND sg13g2_decap_8
XFILLER_41_648 VPWR VGND sg13g2_fill_2
XFILLER_31_11 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_decap_8
X_2507__306 VPWR VGND net305 sg13g2_tiehi
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_49_759 VPWR VGND sg13g2_fill_2
Xoutput9 net9 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_out[4] VPWR VGND sg13g2_buf_1
X_2442__320 VPWR VGND net319 sg13g2_tiehi
XFILLER_16_100 VPWR VGND sg13g2_decap_8
XFILLER_29_472 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_16_177 VPWR VGND sg13g2_decap_8
XFILLER_31_158 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
X_1482_ _0903_ net155 _0902_ VPWR VGND sg13g2_nand2_1
X_1551_ state\[27\] daisychain\[27\] net138 _0958_ VPWR VGND sg13g2_mux2_1
X_1620_ VGND VPWR _1011_ _1012_ _0168_ _1013_ sg13g2_a21oi_1
XFILLER_27_409 VPWR VGND sg13g2_fill_1
XFILLER_39_247 VPWR VGND sg13g2_decap_8
X_2103_ VGND VPWR _0943_ _0741_ _0279_ net72 sg13g2_a21oi_1
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_35_453 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
X_2034_ net178 VPWR _0701_ VGND daisychain\[123\] net26 sg13g2_o21ai_1
XFILLER_31_681 VPWR VGND sg13g2_decap_8
X_1818_ VGND VPWR net126 daisychain\[79\] _0528_ net62 sg13g2_a21oi_1
X_1749_ net195 VPWR _0473_ VGND daisychain\[66\] net40 sg13g2_o21ai_1
XFILLER_14_604 VPWR VGND sg13g2_fill_1
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_55 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_46_718 VPWR VGND sg13g2_fill_2
XFILLER_46_729 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_26_475 VPWR VGND sg13g2_decap_8
XFILLER_26_486 VPWR VGND sg13g2_fill_2
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_41_401 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_5_335 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_20_607 VPWR VGND sg13g2_fill_1
XFILLER_32_401 VPWR VGND sg13g2_decap_4
XFILLER_32_434 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_fill_1
XFILLER_8_151 VPWR VGND sg13g2_decap_8
X_1465_ VGND VPWR _0887_ _0888_ _0137_ _0889_ sg13g2_a21oi_1
X_1534_ net183 VPWR _0945_ VGND daisychain\[23\] net28 sg13g2_o21ai_1
Xfanout108 net109 net108 VPWR VGND sg13g2_buf_1
Xfanout119 net122 net119 VPWR VGND sg13g2_buf_1
X_1603_ VGND VPWR net105 daisychain\[36\] _1000_ net57 sg13g2_a21oi_1
XFILLER_27_217 VPWR VGND sg13g2_decap_8
XFILLER_36_751 VPWR VGND sg13g2_decap_4
X_1396_ VPWR _0035_ state\[16\] VGND sg13g2_inv_1
X_2017_ _0687_ net158 _0686_ VPWR VGND sg13g2_nand2_1
XFILLER_10_139 VPWR VGND sg13g2_decap_8
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_46_515 VPWR VGND sg13g2_fill_2
XFILLER_18_228 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_10_684 VPWR VGND sg13g2_fill_2
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_5_132 VPWR VGND sg13g2_decap_8
XFILLER_6_699 VPWR VGND sg13g2_decap_8
XFILLER_24_209 VPWR VGND sg13g2_decap_8
XFILLER_37_537 VPWR VGND sg13g2_decap_4
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_33_754 VPWR VGND sg13g2_fill_1
X_2386__435 VPWR VGND net434 sg13g2_tiehi
XFILLER_4_80 VPWR VGND sg13g2_decap_8
X_1448_ VGND VPWR net101 daisychain\[5\] _0876_ net49 sg13g2_a21oi_1
X_1517_ _0931_ net159 _0930_ VPWR VGND sg13g2_nand2_1
X_2566_ net389 VGND VPWR _0382_ state\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2497_ net355 VGND VPWR _0313_ state\[57\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1379_ VPWR _0054_ state\[33\] VGND sg13g2_inv_1
X_2473__452 VPWR VGND net451 sg13g2_tiehi
XFILLER_11_426 VPWR VGND sg13g2_decap_8
XFILLER_23_242 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_14_231 VPWR VGND sg13g2_decap_8
XFILLER_15_754 VPWR VGND sg13g2_decap_8
XFILLER_15_787 VPWR VGND sg13g2_decap_8
XFILLER_30_702 VPWR VGND sg13g2_fill_1
XFILLER_30_735 VPWR VGND sg13g2_fill_1
XFILLER_34_529 VPWR VGND sg13g2_fill_2
XFILLER_42_573 VPWR VGND sg13g2_fill_1
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_30_768 VPWR VGND sg13g2_fill_1
XFILLER_6_485 VPWR VGND sg13g2_fill_2
Xfanout90 net98 net90 VPWR VGND sg13g2_buf_1
X_2420_ net366 VGND VPWR _0236_ daisychain\[108\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_1302_ VPWR _0012_ state\[110\] VGND sg13g2_inv_1
X_2351_ net248 VGND VPWR _0167_ daisychain\[39\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2282_ _0831_ net107 state\[113\] VPWR VGND sg13g2_nand2_1
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_25_518 VPWR VGND sg13g2_decap_8
XFILLER_25_529 VPWR VGND sg13g2_fill_2
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_20_201 VPWR VGND sg13g2_decap_8
X_1997_ _0671_ net157 _0670_ VPWR VGND sg13g2_nand2_1
X_2549_ net381 VGND VPWR _0365_ state\[109\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_28_301 VPWR VGND sg13g2_fill_2
XFILLER_11_201 VPWR VGND sg13g2_decap_8
XFILLER_12_735 VPWR VGND sg13g2_fill_1
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_11_278 VPWR VGND sg13g2_decap_8
XFILLER_12_757 VPWR VGND sg13g2_decap_8
XFILLER_7_249 VPWR VGND sg13g2_decap_8
XFILLER_3_455 VPWR VGND sg13g2_decap_8
XFILLER_34_315 VPWR VGND sg13g2_decap_8
XFILLER_34_348 VPWR VGND sg13g2_fill_2
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_47_654 VPWR VGND sg13g2_decap_4
XFILLER_15_551 VPWR VGND sg13g2_fill_2
XFILLER_30_543 VPWR VGND sg13g2_fill_1
XFILLER_30_554 VPWR VGND sg13g2_fill_2
XFILLER_42_392 VPWR VGND sg13g2_decap_8
X_1920_ VGND VPWR _0607_ _0608_ _0228_ _0609_ sg13g2_a21oi_1
X_1851_ state\[87\] daisychain\[87\] net142 _0554_ VPWR VGND sg13g2_mux2_1
XFILLER_6_260 VPWR VGND sg13g2_decap_8
X_2403_ net400 VGND VPWR _0219_ daisychain\[91\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1782_ _0499_ net174 _0498_ VPWR VGND sg13g2_nand2_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_38_621 VPWR VGND sg13g2_fill_1
X_2334_ net282 VGND VPWR _0150_ daisychain\[22\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2265_ VGND VPWR _0623_ _0822_ _0360_ net75 sg13g2_a21oi_1
X_2196_ _0788_ net129 state\[70\] VPWR VGND sg13g2_nand2_1
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_21_510 VPWR VGND sg13g2_decap_8
XFILLER_25_326 VPWR VGND sg13g2_decap_4
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_38_687 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_20_68 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_29_66 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_44_624 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv1 VPWR digitalen.g\[2\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_12_510 VPWR VGND sg13g2_fill_2
XFILLER_12_576 VPWR VGND sg13g2_decap_8
XFILLER_12_587 VPWR VGND sg13g2_fill_2
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_44_668 VPWR VGND sg13g2_fill_1
XFILLER_45_98 VPWR VGND sg13g2_decap_8
X_2412__383 VPWR VGND net382 sg13g2_tiehi
XFILLER_3_252 VPWR VGND sg13g2_decap_8
XFILLER_4_731 VPWR VGND sg13g2_decap_8
XFILLER_4_764 VPWR VGND sg13g2_fill_2
XFILLER_4_786 VPWR VGND sg13g2_decap_4
XFILLER_8_547 VPWR VGND sg13g2_decap_8
XFILLER_10_90 VPWR VGND sg13g2_decap_8
XFILLER_19_120 VPWR VGND sg13g2_decap_8
X_2050_ VGND VPWR _0711_ _0712_ _0254_ _0713_ sg13g2_a21oi_1
XFILLER_19_197 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_34_189 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_15_392 VPWR VGND sg13g2_decap_4
X_1903_ VGND VPWR net112 daisychain\[96\] _0596_ net55 sg13g2_a21oi_1
X_1834_ net194 VPWR _0541_ VGND daisychain\[83\] net39 sg13g2_o21ai_1
X_1765_ VGND VPWR _0483_ _0484_ _0197_ _0485_ sg13g2_a21oi_1
X_1696_ state\[56\] daisychain\[56\] net146 _0430_ VPWR VGND sg13g2_mux2_1
X_2317_ net316 VGND VPWR _0133_ daisychain\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2248_ _0814_ net111 state\[96\] VPWR VGND sg13g2_nand2_1
X_2179_ VGND VPWR _0451_ _0779_ _0317_ net82 sg13g2_a21oi_1
XFILLER_14_808 VPWR VGND sg13g2_decap_8
XFILLER_15_13 VPWR VGND sg13g2_fill_2
XFILLER_15_79 VPWR VGND sg13g2_decap_8
XFILLER_25_145 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_31_67 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_16_156 VPWR VGND sg13g2_decap_8
XFILLER_44_476 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_31_137 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
X_2525__418 VPWR VGND net417 sg13g2_tiehi
X_1481_ state\[13\] daisychain\[13\] net134 _0902_ VPWR VGND sg13g2_mux2_1
X_1550_ VGND VPWR _0955_ _0956_ _0154_ _0957_ sg13g2_a21oi_1
XFILLER_39_226 VPWR VGND sg13g2_decap_8
X_2102_ _0741_ net105 state\[23\] VPWR VGND sg13g2_nand2_1
X_2033_ VGND VPWR net89 daisychain\[122\] _0700_ net48 sg13g2_a21oi_1
XFILLER_22_137 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_8
X_2315__321 VPWR VGND net320 sg13g2_tiehi
X_1817_ _0527_ net173 _0526_ VPWR VGND sg13g2_nand2_1
X_1748_ VGND VPWR net130 daisychain\[65\] _0472_ net64 sg13g2_a21oi_1
X_2396__415 VPWR VGND net414 sg13g2_tiehi
X_1679_ net192 VPWR _0417_ VGND daisychain\[52\] net37 sg13g2_o21ai_1
XFILLER_14_627 VPWR VGND sg13g2_decap_4
XFILLER_26_432 VPWR VGND sg13g2_fill_2
XFILLER_26_443 VPWR VGND sg13g2_decap_4
XFILLER_26_465 VPWR VGND sg13g2_decap_4
XFILLER_26_498 VPWR VGND sg13g2_fill_1
XFILLER_10_822 VPWR VGND sg13g2_fill_1
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_21_192 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_3_38 VPWR VGND sg13g2_decap_8
XFILLER_5_314 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_17_454 VPWR VGND sg13g2_fill_1
XFILLER_17_487 VPWR VGND sg13g2_decap_4
XFILLER_20_619 VPWR VGND sg13g2_fill_1
XFILLER_32_424 VPWR VGND sg13g2_fill_2
XFILLER_32_446 VPWR VGND sg13g2_decap_8
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_45_763 VPWR VGND sg13g2_decap_4
XFILLER_40_490 VPWR VGND sg13g2_fill_2
XFILLER_8_130 VPWR VGND sg13g2_decap_8
X_1602_ _0999_ net161 _0998_ VPWR VGND sg13g2_nand2_1
X_1395_ VPWR _0036_ state\[17\] VGND sg13g2_inv_1
X_1464_ net179 VPWR _0889_ VGND daisychain\[9\] net23 sg13g2_o21ai_1
X_1533_ VGND VPWR net104 daisychain\[22\] _0944_ net51 sg13g2_a21oi_1
Xfanout109 net114 net109 VPWR VGND sg13g2_buf_1
XFILLER_35_273 VPWR VGND sg13g2_decap_8
X_2016_ state\[120\] daisychain\[120\] net136 _0686_ VPWR VGND sg13g2_mux2_1
XFILLER_10_118 VPWR VGND sg13g2_decap_8
XFILLER_23_468 VPWR VGND sg13g2_decap_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_19_708 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_5_111 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_5_188 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_9_461 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_1516_ state\[20\] daisychain\[20\] net137 _0930_ VPWR VGND sg13g2_mux2_1
X_2565_ net261 VGND VPWR _0381_ state\[125\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2503__332 VPWR VGND net331 sg13g2_tiehi
XFILLER_28_505 VPWR VGND sg13g2_decap_4
X_1378_ VPWR _0055_ state\[34\] VGND sg13g2_inv_1
X_1447_ _0875_ net159 _0874_ VPWR VGND sg13g2_nand2_1
X_2496_ net359 VGND VPWR _0312_ state\[56\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_11_405 VPWR VGND sg13g2_decap_8
XFILLER_23_221 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
X_2480__424 VPWR VGND net423 sg13g2_tiehi
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_3_604 VPWR VGND sg13g2_decap_8
XFILLER_3_637 VPWR VGND sg13g2_decap_4
XFILLER_48_21 VPWR VGND sg13g2_decap_8
X_2508__298 VPWR VGND net297 sg13g2_tiehi
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_14_210 VPWR VGND sg13g2_decap_8
XFILLER_14_287 VPWR VGND sg13g2_decap_8
XFILLER_15_733 VPWR VGND sg13g2_decap_8
XFILLER_30_747 VPWR VGND sg13g2_fill_1
Xfanout91 net93 net91 VPWR VGND sg13g2_buf_1
Xfanout80 net87 net80 VPWR VGND sg13g2_buf_1
XFILLER_10_471 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_49_151 VPWR VGND sg13g2_decap_8
X_1301_ VPWR _0013_ state\[111\] VGND sg13g2_inv_1
Xclkbuf_leaf_1_clk clknet_2_1__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_2422__363 VPWR VGND net362 sg13g2_tiehi
X_2350_ net250 VGND VPWR _0166_ daisychain\[38\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2281_ VGND VPWR _0655_ _0830_ _0368_ net75 sg13g2_a21oi_1
XFILLER_18_571 VPWR VGND sg13g2_decap_8
XFILLER_33_530 VPWR VGND sg13g2_fill_1
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_20_257 VPWR VGND sg13g2_decap_4
XFILLER_33_585 VPWR VGND sg13g2_decap_8
X_1996_ state\[116\] daisychain\[116\] net135 _0670_ VPWR VGND sg13g2_mux2_1
XFILLER_0_607 VPWR VGND sg13g2_decap_4
XFILLER_0_629 VPWR VGND sg13g2_decap_8
X_2548_ net397 VGND VPWR _0364_ state\[108\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_18_13 VPWR VGND sg13g2_fill_1
XFILLER_44_817 VPWR VGND sg13g2_decap_4
X_2479_ net427 VGND VPWR _0295_ state\[39\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_11_257 VPWR VGND sg13g2_decap_8
XFILLER_24_530 VPWR VGND sg13g2_fill_1
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_7_228 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_2_3__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_19_313 VPWR VGND sg13g2_fill_1
XFILLER_47_600 VPWR VGND sg13g2_decap_4
XFILLER_15_530 VPWR VGND sg13g2_fill_2
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_47_633 VPWR VGND sg13g2_fill_2
XFILLER_15_574 VPWR VGND sg13g2_decap_4
XFILLER_15_596 VPWR VGND sg13g2_decap_4
XFILLER_30_511 VPWR VGND sg13g2_fill_1
XFILLER_42_371 VPWR VGND sg13g2_decap_8
X_2567__454 VPWR VGND net453 sg13g2_tiehi
X_1850_ VGND VPWR _0551_ _0552_ _0214_ _0553_ sg13g2_a21oi_1
X_1781_ state\[73\] daisychain\[73\] net150 _0498_ VPWR VGND sg13g2_mux2_1
X_2402_ net402 VGND VPWR _0218_ daisychain\[90\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2333_ net284 VGND VPWR _0149_ daisychain\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_38_611 VPWR VGND sg13g2_decap_4
X_2264_ _0822_ net108 state\[104\] VPWR VGND sg13g2_nand2_1
X_2195_ VGND VPWR _0483_ _0787_ _0325_ net86 sg13g2_a21oi_1
XFILLER_33_382 VPWR VGND sg13g2_fill_2
XFILLER_40_308 VPWR VGND sg13g2_decap_8
X_2325__301 VPWR VGND net300 sg13g2_tiehi
X_1979_ net186 VPWR _0657_ VGND daisychain\[112\] net31 sg13g2_o21ai_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_45 VPWR VGND sg13g2_decap_8
XFILLER_28_165 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_44_647 VPWR VGND sg13g2_fill_1
XFILLER_45_77 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv2 VPWR digitalen.g\[2\].u.OUTP digitalen.g\[2\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_3_231 VPWR VGND sg13g2_decap_8
XFILLER_4_743 VPWR VGND sg13g2_decap_8
XFILLER_6_49 VPWR VGND sg13g2_fill_1
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_176 VPWR VGND sg13g2_decap_8
XFILLER_30_330 VPWR VGND sg13g2_fill_2
XFILLER_34_168 VPWR VGND sg13g2_decap_8
XFILLER_35_658 VPWR VGND sg13g2_decap_8
X_1902_ _0595_ net166 _0594_ VPWR VGND sg13g2_nand2_1
X_1833_ VGND VPWR net125 daisychain\[82\] _0540_ net61 sg13g2_a21oi_1
X_1764_ net196 VPWR _0485_ VGND daisychain\[69\] net41 sg13g2_o21ai_1
X_2316_ net318 VGND VPWR _0132_ daisychain\[4\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1695_ VGND VPWR _0427_ _0428_ _0183_ _0429_ sg13g2_a21oi_1
X_2247_ VGND VPWR _0587_ _0813_ _0351_ net77 sg13g2_a21oi_1
X_2178_ _0779_ net123 state\[61\] VPWR VGND sg13g2_nand2_1
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_58 VPWR VGND sg13g2_decap_8
XFILLER_21_330 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_31_46 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_12_330 VPWR VGND sg13g2_decap_8
XFILLER_16_135 VPWR VGND sg13g2_decap_8
XFILLER_31_116 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_8_389 VPWR VGND sg13g2_decap_8
XFILLER_39_205 VPWR VGND sg13g2_decap_8
XFILLER_4_584 VPWR VGND sg13g2_decap_8
X_1480_ VGND VPWR _0899_ _0900_ _0140_ _0901_ sg13g2_a21oi_1
XFILLER_48_750 VPWR VGND sg13g2_fill_1
X_2101_ VGND VPWR _0939_ _0740_ _0278_ net72 sg13g2_a21oi_1
X_2032_ _0699_ net154 _0698_ VPWR VGND sg13g2_nand2_1
XFILLER_16_680 VPWR VGND sg13g2_fill_1
XFILLER_16_691 VPWR VGND sg13g2_fill_2
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_30_193 VPWR VGND sg13g2_decap_8
X_2541__254 VPWR VGND net253 sg13g2_tiehi
X_1816_ state\[80\] daisychain\[80\] net148 _0526_ VPWR VGND sg13g2_mux2_1
X_1747_ _0471_ net174 _0470_ VPWR VGND sg13g2_nand2_1
X_1678_ VGND VPWR net120 daisychain\[51\] _0416_ net59 sg13g2_a21oi_1
X_2476__440 VPWR VGND net439 sg13g2_tiehi
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_fill_1
XFILLER_21_171 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_fill_1
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_13_661 VPWR VGND sg13g2_fill_1
XFILLER_13_694 VPWR VGND sg13g2_decap_8
XFILLER_44_252 VPWR VGND sg13g2_decap_8
XFILLER_9_632 VPWR VGND sg13g2_decap_8
XFILLER_9_643 VPWR VGND sg13g2_fill_1
XFILLER_8_186 VPWR VGND sg13g2_decap_8
X_1532_ _0943_ net161 _0942_ VPWR VGND sg13g2_nand2_1
X_1601_ state\[37\] daisychain\[37\] net139 _0998_ VPWR VGND sg13g2_mux2_1
XFILLER_4_381 VPWR VGND sg13g2_decap_8
X_1394_ VPWR _0037_ state\[18\] VGND sg13g2_inv_1
X_1463_ VGND VPWR net92 daisychain\[8\] _0888_ net45 sg13g2_a21oi_1
XFILLER_23_425 VPWR VGND sg13g2_fill_1
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_36_731 VPWR VGND sg13g2_decap_4
X_2432__343 VPWR VGND net342 sg13g2_tiehi
X_2015_ VGND VPWR _0683_ _0684_ _0247_ _0685_ sg13g2_a21oi_1
XFILLER_23_458 VPWR VGND sg13g2_decap_8
XFILLER_2_329 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_42_778 VPWR VGND sg13g2_fill_2
X_2333__285 VPWR VGND net284 sg13g2_tiehi
XFILLER_10_675 VPWR VGND sg13g2_fill_1
XFILLER_10_686 VPWR VGND sg13g2_fill_1
XFILLER_5_167 VPWR VGND sg13g2_decap_8
XFILLER_6_646 VPWR VGND sg13g2_decap_8
XFILLER_6_657 VPWR VGND sg13g2_fill_1
X_2409__389 VPWR VGND net388 sg13g2_tiehi
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_17_274 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_745 VPWR VGND sg13g2_decap_8
XFILLER_32_277 VPWR VGND sg13g2_decap_8
XFILLER_33_789 VPWR VGND sg13g2_decap_4
X_1515_ VGND VPWR _0927_ _0928_ _0147_ _0929_ sg13g2_a21oi_1
X_2564_ net357 VGND VPWR _0380_ state\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2495_ net363 VGND VPWR _0311_ state\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_28_517 VPWR VGND sg13g2_decap_8
X_1377_ VPWR _0056_ state\[35\] VGND sg13g2_inv_1
X_1446_ state\[6\] daisychain\[6\] net138 _0874_ VPWR VGND sg13g2_mux2_1
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_14_266 VPWR VGND sg13g2_decap_8
Xfanout92 net93 net92 VPWR VGND sg13g2_buf_1
Xfanout81 net82 net81 VPWR VGND sg13g2_buf_1
Xfanout70 net88 net70 VPWR VGND sg13g2_buf_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_6_421 VPWR VGND sg13g2_decap_8
XFILLER_6_465 VPWR VGND sg13g2_decap_4
XFILLER_6_498 VPWR VGND sg13g2_fill_2
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
X_1300_ VPWR _0014_ state\[112\] VGND sg13g2_inv_1
X_2280_ _0830_ net107 state\[112\] VPWR VGND sg13g2_nand2_1
XFILLER_20_236 VPWR VGND sg13g2_decap_8
XFILLER_9_281 VPWR VGND sg13g2_decap_8
X_1995_ VGND VPWR _0667_ _0668_ _0243_ _0669_ sg13g2_a21oi_1
X_1429_ net180 VPWR _0861_ VGND daisychain\[2\] net24 sg13g2_o21ai_1
X_2547_ net413 VGND VPWR _0363_ state\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2478_ net431 VGND VPWR _0294_ state\[38\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_16_509 VPWR VGND sg13g2_fill_2
XFILLER_11_236 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_decap_8
XFILLER_7_207 VPWR VGND sg13g2_decap_8
Xclkload1 clkload1/Y clknet_leaf_10_clk VPWR VGND sg13g2_inv_2
XFILLER_20_781 VPWR VGND sg13g2_fill_1
XFILLER_3_413 VPWR VGND sg13g2_decap_8
XFILLER_19_325 VPWR VGND sg13g2_fill_2
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_24_90 VPWR VGND sg13g2_decap_4
XFILLER_30_567 VPWR VGND sg13g2_fill_1
XFILLER_30_589 VPWR VGND sg13g2_fill_1
XFILLER_7_741 VPWR VGND sg13g2_fill_1
XFILLER_7_785 VPWR VGND sg13g2_fill_2
X_1780_ VGND VPWR _0495_ _0496_ _0200_ _0497_ sg13g2_a21oi_1
XFILLER_6_295 VPWR VGND sg13g2_decap_8
X_2401_ net404 VGND VPWR _0217_ daisychain\[89\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2332_ net286 VGND VPWR _0148_ daisychain\[20\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_37_133 VPWR VGND sg13g2_decap_8
X_2263_ VGND VPWR _0619_ _0821_ _0359_ net75 sg13g2_a21oi_1
X_2194_ _0787_ net129 state\[69\] VPWR VGND sg13g2_nand2_1
XFILLER_20_15 VPWR VGND sg13g2_fill_2
X_1978_ VGND VPWR net96 daisychain\[111\] _0656_ net47 sg13g2_a21oi_1
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_24 VPWR VGND sg13g2_decap_8
XFILLER_12_501 VPWR VGND sg13g2_fill_1
XFILLER_16_328 VPWR VGND sg13g2_decap_4
XFILLER_24_372 VPWR VGND sg13g2_decap_4
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_8_538 VPWR VGND sg13g2_decap_4
XFILLER_3_210 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_8
XFILLER_19_155 VPWR VGND sg13g2_decap_8
XFILLER_35_604 VPWR VGND sg13g2_fill_2
XFILLER_35_637 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_34_147 VPWR VGND sg13g2_decap_8
X_1901_ state\[97\] daisychain\[97\] net143 _0594_ VPWR VGND sg13g2_mux2_1
X_1832_ _0539_ net172 _0538_ VPWR VGND sg13g2_nand2_1
X_1763_ VGND VPWR net128 daisychain\[68\] _0484_ net64 sg13g2_a21oi_1
X_1694_ net192 VPWR _0429_ VGND daisychain\[55\] net37 sg13g2_o21ai_1
X_2315_ net320 VGND VPWR _0131_ daisychain\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2246_ _0813_ net111 state\[95\] VPWR VGND sg13g2_nand2_1
XFILLER_15_15 VPWR VGND sg13g2_fill_1
XFILLER_15_26 VPWR VGND sg13g2_decap_8
XFILLER_38_475 VPWR VGND sg13g2_decap_8
X_2177_ VGND VPWR _0447_ _0778_ _0316_ net82 sg13g2_a21oi_1
XFILLER_31_25 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_1_758 VPWR VGND sg13g2_fill_2
Xoutput14 net14 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_16_114 VPWR VGND sg13g2_decap_8
XFILLER_29_486 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_12_353 VPWR VGND sg13g2_decap_8
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_21_80 VPWR VGND sg13g2_decap_8
XFILLER_8_368 VPWR VGND sg13g2_decap_8
X_2343__265 VPWR VGND net264 sg13g2_tiehi
X_2100_ _0740_ net104 state\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_47_294 VPWR VGND sg13g2_decap_8
X_2419__369 VPWR VGND net368 sg13g2_tiehi
X_2031_ state\[123\] daisychain\[123\] net136 _0698_ VPWR VGND sg13g2_mux2_1
XFILLER_15_191 VPWR VGND sg13g2_decap_8
XFILLER_30_172 VPWR VGND sg13g2_decap_8
XFILLER_31_695 VPWR VGND sg13g2_decap_8
X_1815_ VGND VPWR _0523_ _0524_ _0207_ _0525_ sg13g2_a21oi_1
XFILLER_7_93 VPWR VGND sg13g2_fill_2
X_1746_ state\[66\] daisychain\[66\] net150 _0470_ VPWR VGND sg13g2_mux2_1
X_1677_ _0415_ net170 _0414_ VPWR VGND sg13g2_nand2_1
XFILLER_39_751 VPWR VGND sg13g2_decap_8
XFILLER_39_773 VPWR VGND sg13g2_fill_1
XFILLER_39_784 VPWR VGND sg13g2_fill_2
X_2229_ VGND VPWR _0551_ _0804_ _0342_ net84 sg13g2_a21oi_1
XFILLER_10_802 VPWR VGND sg13g2_fill_2
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_26_434 VPWR VGND sg13g2_fill_1
XFILLER_26_69 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_41_415 VPWR VGND sg13g2_decap_4
XFILLER_41_437 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_fill_2
XFILLER_41_459 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_21_150 VPWR VGND sg13g2_decap_8
XFILLER_5_349 VPWR VGND sg13g2_decap_8
X_2483__412 VPWR VGND net411 sg13g2_tiehi
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_12_183 VPWR VGND sg13g2_decap_8
XFILLER_13_673 VPWR VGND sg13g2_decap_8
XFILLER_40_492 VPWR VGND sg13g2_fill_1
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
X_1462_ _0887_ net155 _0886_ VPWR VGND sg13g2_nand2_1
X_1531_ state\[23\] daisychain\[23\] net139 _0942_ VPWR VGND sg13g2_mux2_1
X_2529__386 VPWR VGND net385 sg13g2_tiehi
X_1600_ VGND VPWR _0995_ _0996_ _0164_ _0997_ sg13g2_a21oi_1
XFILLER_36_710 VPWR VGND sg13g2_fill_2
XFILLER_48_581 VPWR VGND sg13g2_fill_1
X_1393_ VPWR _0038_ state\[19\] VGND sg13g2_inv_1
XFILLER_35_231 VPWR VGND sg13g2_decap_8
XFILLER_36_787 VPWR VGND sg13g2_decap_4
X_2014_ net180 VPWR _0685_ VGND daisychain\[119\] net24 sg13g2_o21ai_1
XFILLER_12_38 VPWR VGND sg13g2_fill_2
X_2847_ daisychain\[127\] net22 VPWR VGND sg13g2_buf_1
XFILLER_2_308 VPWR VGND sg13g2_decap_8
X_1729_ net193 VPWR _0457_ VGND daisychain\[62\] net38 sg13g2_o21ai_1
XFILLER_26_253 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_10_698 VPWR VGND sg13g2_decap_8
XFILLER_5_146 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_17_253 VPWR VGND sg13g2_decap_8
XFILLER_18_754 VPWR VGND sg13g2_fill_1
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_fill_1
XFILLER_33_779 VPWR VGND sg13g2_decap_4
XFILLER_45_595 VPWR VGND sg13g2_decap_8
XFILLER_9_463 VPWR VGND sg13g2_fill_1
X_2312__326 VPWR VGND net325 sg13g2_tiehi
XFILLER_4_94 VPWR VGND sg13g2_decap_8
X_1445_ VGND VPWR _0871_ _0872_ _0133_ _0873_ sg13g2_a21oi_1
X_1514_ net182 VPWR _0929_ VGND daisychain\[19\] net27 sg13g2_o21ai_1
X_2563_ net421 VGND VPWR _0379_ state\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2494_ net367 VGND VPWR _0310_ state\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_551 VPWR VGND sg13g2_decap_4
X_1376_ VPWR _0057_ state\[36\] VGND sg13g2_inv_1
XFILLER_23_256 VPWR VGND sg13g2_decap_8
XFILLER_32_790 VPWR VGND sg13g2_fill_1
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_14_245 VPWR VGND sg13g2_decap_8
XFILLER_15_768 VPWR VGND sg13g2_decap_8
XFILLER_42_532 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_30_727 VPWR VGND sg13g2_fill_1
XFILLER_6_400 VPWR VGND sg13g2_decap_8
Xfanout93 net98 net93 VPWR VGND sg13g2_buf_1
Xfanout82 net87 net82 VPWR VGND sg13g2_buf_1
Xfanout71 net74 net71 VPWR VGND sg13g2_buf_1
Xfanout60 net65 net60 VPWR VGND sg13g2_buf_1
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_38_805 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_20_215 VPWR VGND sg13g2_decap_8
XFILLER_33_554 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
X_1994_ net180 VPWR _0669_ VGND daisychain\[115\] net24 sg13g2_o21ai_1
XFILLER_9_260 VPWR VGND sg13g2_decap_8
X_1428_ VGND VPWR net94 daisychain\[1\] _0860_ net46 sg13g2_a21oi_1
X_2546_ net429 VGND VPWR _0362_ state\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2477_ net435 VGND VPWR _0293_ state\[37\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2401__405 VPWR VGND net404 sg13g2_tiehi
XFILLER_24_510 VPWR VGND sg13g2_fill_2
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
X_1359_ VPWR _0076_ state\[53\] VGND sg13g2_inv_1
XFILLER_11_215 VPWR VGND sg13g2_decap_8
XFILLER_20_760 VPWR VGND sg13g2_fill_1
XFILLER_20_793 VPWR VGND sg13g2_fill_1
Xclkload2 VPWR clkload2/Y clknet_leaf_14_clk VGND sg13g2_inv_1
XFILLER_35_819 VPWR VGND sg13g2_decap_4
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_47_635 VPWR VGND sg13g2_fill_1
XFILLER_15_510 VPWR VGND sg13g2_decap_8
XFILLER_34_329 VPWR VGND sg13g2_decap_4
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_6_274 VPWR VGND sg13g2_decap_8
XFILLER_7_764 VPWR VGND sg13g2_decap_8
X_2400_ net406 VGND VPWR _0216_ daisychain\[88\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2331_ net288 VGND VPWR _0147_ daisychain\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2262_ _0821_ net110 state\[103\] VPWR VGND sg13g2_nand2_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
X_2353__245 VPWR VGND net244 sg13g2_tiehi
X_2193_ VGND VPWR _0479_ _0786_ _0324_ net85 sg13g2_a21oi_1
XFILLER_21_524 VPWR VGND sg13g2_decap_8
XFILLER_33_384 VPWR VGND sg13g2_fill_1
X_2429__349 VPWR VGND net348 sg13g2_tiehi
X_1977_ _0655_ net164 _0654_ VPWR VGND sg13g2_nand2_1
XFILLER_0_406 VPWR VGND sg13g2_decap_8
X_2529_ net385 VGND VPWR _0345_ state\[89\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_24_340 VPWR VGND sg13g2_fill_1
XFILLER_40_822 VPWR VGND sg13g2_fill_1
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_44_638 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_3_266 VPWR VGND sg13g2_decap_8
XFILLER_19_134 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_30_332 VPWR VGND sg13g2_fill_1
XFILLER_31_800 VPWR VGND sg13g2_decap_8
XFILLER_43_671 VPWR VGND sg13g2_decap_8
X_1900_ VGND VPWR _0591_ _0592_ _0224_ _0593_ sg13g2_a21oi_1
X_1831_ state\[83\] daisychain\[83\] net148 _0538_ VPWR VGND sg13g2_mux2_1
XFILLER_7_594 VPWR VGND sg13g2_decap_8
X_1762_ _0483_ net175 _0482_ VPWR VGND sg13g2_nand2_1
X_1693_ VGND VPWR net119 daisychain\[54\] _0428_ net59 sg13g2_a21oi_1
XFILLER_38_432 VPWR VGND sg13g2_decap_8
XFILLER_38_443 VPWR VGND sg13g2_fill_1
XFILLER_38_465 VPWR VGND sg13g2_decap_4
X_2314_ net322 VGND VPWR _0130_ daisychain\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2245_ VGND VPWR _0583_ _0812_ _0350_ net77 sg13g2_a21oi_1
X_2176_ _0778_ net122 state\[60\] VPWR VGND sg13g2_nand2_1
XFILLER_25_159 VPWR VGND sg13g2_decap_8
X_2511__274 VPWR VGND net273 sg13g2_tiehi
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_29_465 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_13_822 VPWR VGND sg13g2_fill_1
XFILLER_24_181 VPWR VGND sg13g2_decap_8
XFILLER_40_652 VPWR VGND sg13g2_decap_8
XFILLER_8_347 VPWR VGND sg13g2_decap_8
XFILLER_48_741 VPWR VGND sg13g2_decap_8
X_2030_ VGND VPWR _0695_ _0696_ _0250_ _0697_ sg13g2_a21oi_1
XFILLER_15_170 VPWR VGND sg13g2_decap_8
XFILLER_35_446 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_30_151 VPWR VGND sg13g2_decap_8
XFILLER_31_663 VPWR VGND sg13g2_fill_1
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_7_72 VPWR VGND sg13g2_decap_8
X_1814_ net196 VPWR _0525_ VGND daisychain\[79\] net41 sg13g2_o21ai_1
X_1745_ VGND VPWR _0467_ _0468_ _0193_ _0469_ sg13g2_a21oi_1
X_1676_ state\[52\] daisychain\[52\] net146 _0414_ VPWR VGND sg13g2_mux2_1
XFILLER_38_273 VPWR VGND sg13g2_decap_8
X_2228_ _0804_ net124 state\[86\] VPWR VGND sg13g2_nand2_1
X_2159_ VGND VPWR _0411_ _0769_ _0307_ net81 sg13g2_a21oi_1
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_5_328 VPWR VGND sg13g2_decap_8
XFILLER_1_512 VPWR VGND sg13g2_fill_1
XFILLER_29_262 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_12_162 VPWR VGND sg13g2_decap_8
XFILLER_25_490 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
X_1392_ VPWR _0040_ state\[20\] VGND sg13g2_inv_1
X_1461_ state\[9\] daisychain\[9\] net134 _0886_ VPWR VGND sg13g2_mux2_1
X_1530_ VGND VPWR _0939_ _0940_ _0150_ _0941_ sg13g2_a21oi_1
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_36_744 VPWR VGND sg13g2_decap_8
X_2013_ VGND VPWR net97 daisychain\[118\] _0684_ net47 sg13g2_a21oi_1
XFILLER_35_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_2_0__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_12_17 VPWR VGND sg13g2_fill_2
X_2846_ daisychain\[126\] net21 VPWR VGND sg13g2_buf_1
X_1728_ VGND VPWR net123 daisychain\[61\] _0456_ net60 sg13g2_a21oi_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
X_1659_ net191 VPWR _0401_ VGND daisychain\[48\] net36 sg13g2_o21ai_1
XFILLER_26_232 VPWR VGND sg13g2_decap_8
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_42_736 VPWR VGND sg13g2_fill_1
XFILLER_10_611 VPWR VGND sg13g2_fill_2
XFILLER_10_644 VPWR VGND sg13g2_decap_4
XFILLER_10_655 VPWR VGND sg13g2_fill_2
XFILLER_22_493 VPWR VGND sg13g2_decap_8
XFILLER_2_810 VPWR VGND sg13g2_decap_8
XFILLER_2_821 VPWR VGND sg13g2_fill_2
XFILLER_5_125 VPWR VGND sg13g2_decap_8
XFILLER_18_744 VPWR VGND sg13g2_fill_1
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_17_232 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
X_2562_ net229 VGND VPWR _0378_ state\[122\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_4_40 VPWR VGND sg13g2_fill_1
XFILLER_4_73 VPWR VGND sg13g2_decap_8
XFILLER_5_692 VPWR VGND sg13g2_decap_8
X_1375_ VPWR _0058_ state\[37\] VGND sg13g2_inv_1
X_1444_ net182 VPWR _0873_ VGND daisychain\[5\] net27 sg13g2_o21ai_1
X_1513_ VGND VPWR net99 daisychain\[18\] _0928_ net49 sg13g2_a21oi_1
Xclkbuf_leaf_4_clk clknet_2_3__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_2493_ net371 VGND VPWR _0309_ state\[53\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_23_235 VPWR VGND sg13g2_decap_8
X_2408__391 VPWR VGND net390 sg13g2_tiehi
X_2363__225 VPWR VGND net224 sg13g2_tiehi
XFILLER_48_35 VPWR VGND sg13g2_decap_8
X_2439__329 VPWR VGND net328 sg13g2_tiehi
XFILLER_14_224 VPWR VGND sg13g2_decap_8
XFILLER_15_747 VPWR VGND sg13g2_decap_8
XFILLER_27_530 VPWR VGND sg13g2_fill_1
XFILLER_30_706 VPWR VGND sg13g2_fill_1
XFILLER_30_739 VPWR VGND sg13g2_fill_1
XFILLER_42_511 VPWR VGND sg13g2_fill_2
XFILLER_9_18 VPWR VGND sg13g2_fill_2
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_22_290 VPWR VGND sg13g2_decap_8
Xfanout94 net96 net94 VPWR VGND sg13g2_buf_1
Xfanout83 net87 net83 VPWR VGND sg13g2_buf_1
Xfanout72 net74 net72 VPWR VGND sg13g2_buf_1
Xfanout61 net62 net61 VPWR VGND sg13g2_buf_1
Xfanout50 net52 net50 VPWR VGND sg13g2_buf_1
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
XFILLER_33_599 VPWR VGND sg13g2_fill_1
X_1993_ VGND VPWR net95 daisychain\[114\] _0668_ net46 sg13g2_a21oi_1
X_2545_ net445 VGND VPWR _0361_ state\[105\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1358_ VPWR _0077_ state\[54\] VGND sg13g2_inv_1
X_1427_ _0859_ net155 _0858_ VPWR VGND sg13g2_nand2_1
X_2476_ net439 VGND VPWR _0292_ state\[36\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_36_393 VPWR VGND sg13g2_decap_4
XFILLER_43_308 VPWR VGND sg13g2_decap_8
X_1289_ VPWR _0026_ state\[123\] VGND sg13g2_inv_1
X_2514__250 VPWR VGND net249 sg13g2_tiehi
Xclkload3 clknet_leaf_15_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_3_448 VPWR VGND sg13g2_decap_8
XFILLER_19_327 VPWR VGND sg13g2_fill_1
XFILLER_34_308 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_fill_1
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_10_293 VPWR VGND sg13g2_decap_8
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_6_253 VPWR VGND sg13g2_decap_8
XFILLER_7_787 VPWR VGND sg13g2_fill_1
XFILLER_7_798 VPWR VGND sg13g2_fill_2
XFILLER_2_492 VPWR VGND sg13g2_decap_4
XFILLER_38_647 VPWR VGND sg13g2_fill_2
X_2330_ net290 VGND VPWR _0146_ daisychain\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2261_ VGND VPWR _0615_ _0820_ _0358_ net77 sg13g2_a21oi_1
X_2192_ _0786_ net128 state\[68\] VPWR VGND sg13g2_nand2_1
XFILLER_18_393 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_21_503 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_46_680 VPWR VGND sg13g2_decap_8
XFILLER_46_691 VPWR VGND sg13g2_fill_1
X_1976_ state\[112\] daisychain\[112\] net141 _0654_ VPWR VGND sg13g2_mux2_1
X_2528_ net393 VGND VPWR _0344_ state\[88\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_29_59 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_44_617 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
X_2459_ net251 VGND VPWR _0275_ state\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2486__400 VPWR VGND net399 sg13g2_tiehi
XFILLER_3_245 VPWR VGND sg13g2_decap_8
XFILLER_4_757 VPWR VGND sg13g2_decap_8
XFILLER_10_83 VPWR VGND sg13g2_decap_8
XFILLER_19_113 VPWR VGND sg13g2_decap_8
XFILLER_4_779 VPWR VGND sg13g2_decap_8
XFILLER_15_341 VPWR VGND sg13g2_fill_1
XFILLER_19_92 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_fill_1
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_fill_2
XFILLER_30_311 VPWR VGND sg13g2_fill_1
XFILLER_30_344 VPWR VGND sg13g2_fill_2
XFILLER_30_388 VPWR VGND sg13g2_decap_4
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
X_1830_ VGND VPWR _0535_ _0536_ _0210_ _0537_ sg13g2_a21oi_1
X_1761_ state\[69\] daisychain\[69\] net151 _0482_ VPWR VGND sg13g2_mux2_1
X_2313_ net324 VGND VPWR _0129_ daisychain\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1692_ _0427_ net170 _0426_ VPWR VGND sg13g2_nand2_1
X_2244_ _0812_ net113 state\[94\] VPWR VGND sg13g2_nand2_1
X_2175_ VGND VPWR _0443_ _0777_ _0315_ net82 sg13g2_a21oi_1
XFILLER_19_691 VPWR VGND sg13g2_decap_4
XFILLER_21_344 VPWR VGND sg13g2_fill_2
XFILLER_33_193 VPWR VGND sg13g2_decap_8
XFILLER_34_672 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
X_1959_ net186 VPWR _0641_ VGND daisychain\[108\] net31 sg13g2_o21ai_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_16_149 VPWR VGND sg13g2_decap_8
XFILLER_44_469 VPWR VGND sg13g2_decap_8
XFILLER_24_160 VPWR VGND sg13g2_decap_8
XFILLER_40_664 VPWR VGND sg13g2_decap_4
XFILLER_40_686 VPWR VGND sg13g2_decap_4
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_4_521 VPWR VGND sg13g2_fill_1
XFILLER_39_219 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
XFILLER_31_642 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_7_40 VPWR VGND sg13g2_decap_4
XFILLER_7_95 VPWR VGND sg13g2_fill_1
X_1813_ VGND VPWR net130 daisychain\[78\] _0524_ net64 sg13g2_a21oi_1
X_1744_ net196 VPWR _0469_ VGND daisychain\[65\] net41 sg13g2_o21ai_1
X_2322__307 VPWR VGND net306 sg13g2_tiehi
X_1675_ VGND VPWR _0411_ _0412_ _0179_ _0413_ sg13g2_a21oi_1
XFILLER_26_458 VPWR VGND sg13g2_decap_8
XFILLER_26_469 VPWR VGND sg13g2_fill_2
XFILLER_38_252 VPWR VGND sg13g2_decap_8
X_2227_ VGND VPWR _0547_ _0803_ _0341_ net84 sg13g2_a21oi_1
X_2158_ _0769_ net120 state\[51\] VPWR VGND sg13g2_nand2_1
X_2089_ VGND VPWR _0915_ _0734_ _0272_ net67 sg13g2_a21oi_1
XFILLER_10_815 VPWR VGND sg13g2_decap_8
XFILLER_21_185 VPWR VGND sg13g2_decap_8
XFILLER_5_307 VPWR VGND sg13g2_decap_8
XFILLER_29_241 VPWR VGND sg13g2_decap_8
X_2373__205 VPWR VGND net204 sg13g2_tiehi
XFILLER_16_93 VPWR VGND sg13g2_decap_8
XFILLER_17_447 VPWR VGND sg13g2_decap_8
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_45_767 VPWR VGND sg13g2_fill_1
X_2418__371 VPWR VGND net370 sg13g2_tiehi
XFILLER_12_141 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_4_395 VPWR VGND sg13g2_decap_8
X_1391_ VPWR _0041_ state\[21\] VGND sg13g2_inv_1
X_1460_ VGND VPWR _0883_ _0884_ _0136_ _0885_ sg13g2_a21oi_1
XFILLER_36_712 VPWR VGND sg13g2_fill_1
X_2012_ _0683_ net157 _0682_ VPWR VGND sg13g2_nand2_1
XFILLER_16_480 VPWR VGND sg13g2_fill_2
XFILLER_35_266 VPWR VGND sg13g2_decap_8
X_2845_ daisychain\[125\] net20 VPWR VGND sg13g2_buf_1
XFILLER_8_690 VPWR VGND sg13g2_decap_8
X_1727_ _0455_ net171 _0454_ VPWR VGND sg13g2_nand2_1
X_1658_ VGND VPWR net117 daisychain\[47\] _0400_ net58 sg13g2_a21oi_1
X_1589_ net183 VPWR _0989_ VGND daisychain\[34\] net28 sg13g2_o21ai_1
XFILLER_26_211 VPWR VGND sg13g2_decap_8
XFILLER_26_299 VPWR VGND sg13g2_decap_4
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_22_472 VPWR VGND sg13g2_decap_8
XFILLER_5_104 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_17_211 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_18_789 VPWR VGND sg13g2_decap_4
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_9_454 VPWR VGND sg13g2_decap_8
X_1512_ _0927_ net159 _0926_ VPWR VGND sg13g2_nand2_1
X_2561_ net293 VGND VPWR _0377_ state\[121\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2492_ net375 VGND VPWR _0308_ state\[52\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_4_192 VPWR VGND sg13g2_decap_8
X_1374_ VPWR _0059_ state\[38\] VGND sg13g2_inv_1
X_1443_ VGND VPWR net101 daisychain\[4\] _0872_ net53 sg13g2_a21oi_1
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_36_520 VPWR VGND sg13g2_fill_1
XFILLER_36_575 VPWR VGND sg13g2_fill_2
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_31_291 VPWR VGND sg13g2_fill_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_39_380 VPWR VGND sg13g2_decap_8
X_2554__278 VPWR VGND net277 sg13g2_tiehi
XFILLER_14_203 VPWR VGND sg13g2_decap_8
XFILLER_15_726 VPWR VGND sg13g2_decap_8
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_1
Xfanout62 net65 net62 VPWR VGND sg13g2_buf_1
Xfanout51 net52 net51 VPWR VGND sg13g2_buf_1
Xfanout40 net41 net40 VPWR VGND sg13g2_buf_1
XFILLER_10_464 VPWR VGND sg13g2_decap_8
XFILLER_6_435 VPWR VGND sg13g2_decap_8
Xfanout95 net96 net95 VPWR VGND sg13g2_buf_1
Xfanout84 net87 net84 VPWR VGND sg13g2_buf_1
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_2_630 VPWR VGND sg13g2_decap_8
XFILLER_2_663 VPWR VGND sg13g2_decap_4
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_13_291 VPWR VGND sg13g2_decap_8
XFILLER_33_578 VPWR VGND sg13g2_decap_8
XFILLER_9_295 VPWR VGND sg13g2_decap_8
Xclkload10 VPWR clkload10/Y clknet_leaf_11_clk VGND sg13g2_inv_1
X_1992_ _0667_ net157 _0666_ VPWR VGND sg13g2_nand2_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2544_ net205 VGND VPWR _0360_ state\[104\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2475_ net443 VGND VPWR _0291_ state\[35\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1288_ VPWR _0027_ state\[124\] VGND sg13g2_inv_1
X_1357_ VPWR _0078_ state\[55\] VGND sg13g2_inv_1
X_1426_ state\[2\] daisychain\[2\] net133 _0858_ VPWR VGND sg13g2_mux2_1
XFILLER_24_512 VPWR VGND sg13g2_fill_1
XFILLER_24_523 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_20_740 VPWR VGND sg13g2_fill_1
XFILLER_20_773 VPWR VGND sg13g2_fill_1
XFILLER_3_427 VPWR VGND sg13g2_decap_8
Xclkload4 VPWR clkload4/Y clknet_leaf_16_clk VGND sg13g2_inv_1
XFILLER_47_604 VPWR VGND sg13g2_fill_1
XFILLER_46_147 VPWR VGND sg13g2_decap_8
X_2532__362 VPWR VGND net361 sg13g2_tiehi
XFILLER_11_740 VPWR VGND sg13g2_fill_1
XFILLER_15_567 VPWR VGND sg13g2_decap_8
XFILLER_15_589 VPWR VGND sg13g2_decap_8
XFILLER_30_559 VPWR VGND sg13g2_fill_1
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_10_272 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_6_232 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
XFILLER_38_604 VPWR VGND sg13g2_decap_8
XFILLER_38_615 VPWR VGND sg13g2_fill_1
XFILLER_38_626 VPWR VGND sg13g2_fill_1
X_2260_ _0820_ net110 state\[102\] VPWR VGND sg13g2_nand2_1
X_2191_ VGND VPWR _0475_ _0785_ _0323_ net85 sg13g2_a21oi_1
XFILLER_33_375 VPWR VGND sg13g2_decap_8
X_1975_ VGND VPWR _0651_ _0652_ _0239_ _0653_ sg13g2_a21oi_1
XFILLER_29_38 VPWR VGND sg13g2_decap_8
X_1409_ VPWR _0061_ state\[3\] VGND sg13g2_inv_1
X_2527_ net401 VGND VPWR _0343_ state\[87\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2458_ net255 VGND VPWR _0274_ state\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_28_158 VPWR VGND sg13g2_decap_8
XFILLER_37_692 VPWR VGND sg13g2_decap_8
X_2389_ net428 VGND VPWR _0205_ daisychain\[77\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_20_570 VPWR VGND sg13g2_decap_8
XFILLER_24_331 VPWR VGND sg13g2_decap_8
XFILLER_10_62 VPWR VGND sg13g2_decap_8
XFILLER_3_224 VPWR VGND sg13g2_decap_8
X_2382__443 VPWR VGND net442 sg13g2_tiehi
XFILLER_19_71 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_15_353 VPWR VGND sg13g2_decap_8
XFILLER_16_821 VPWR VGND sg13g2_fill_2
XFILLER_19_169 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_43_662 VPWR VGND sg13g2_decap_4
XFILLER_7_585 VPWR VGND sg13g2_decap_4
X_2428__351 VPWR VGND net350 sg13g2_tiehi
X_1760_ VGND VPWR _0479_ _0480_ _0196_ _0481_ sg13g2_a21oi_1
X_1691_ state\[55\] daisychain\[55\] net146 _0426_ VPWR VGND sg13g2_mux2_1
X_2312_ net325 VGND VPWR _0128_ daisychain\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_25_117 VPWR VGND sg13g2_fill_1
XFILLER_38_423 VPWR VGND sg13g2_fill_1
XFILLER_38_489 VPWR VGND sg13g2_decap_4
X_2243_ VGND VPWR _0579_ _0811_ _0349_ net77 sg13g2_a21oi_1
X_2174_ _0777_ net122 state\[59\] VPWR VGND sg13g2_nand2_1
XFILLER_33_172 VPWR VGND sg13g2_decap_8
XFILLER_31_39 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[2] VPWR VGND sg13g2_buf_1
X_2329__293 VPWR VGND net292 sg13g2_tiehi
X_1958_ VGND VPWR net108 daisychain\[107\] _0640_ net53 sg13g2_a21oi_1
X_1889_ net187 VPWR _0585_ VGND daisychain\[94\] net32 sg13g2_o21ai_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_434 VPWR VGND sg13g2_decap_4
XFILLER_16_128 VPWR VGND sg13g2_decap_8
XFILLER_31_109 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_12_323 VPWR VGND sg13g2_decap_8
XFILLER_12_367 VPWR VGND sg13g2_fill_1
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_0_750 VPWR VGND sg13g2_decap_8
XFILLER_21_94 VPWR VGND sg13g2_decap_8
XFILLER_4_577 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_16_673 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_30_186 VPWR VGND sg13g2_decap_8
XFILLER_7_382 VPWR VGND sg13g2_decap_8
X_1812_ _0523_ net175 _0522_ VPWR VGND sg13g2_nand2_1
X_1743_ VGND VPWR net130 daisychain\[64\] _0468_ net64 sg13g2_a21oi_1
X_1674_ net192 VPWR _0413_ VGND daisychain\[51\] net37 sg13g2_o21ai_1
X_2226_ _0803_ net125 state\[85\] VPWR VGND sg13g2_nand2_1
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_38_231 VPWR VGND sg13g2_decap_8
X_2157_ VGND VPWR _0407_ _0768_ _0306_ net81 sg13g2_a21oi_1
X_2088_ _0734_ net99 state\[16\] VPWR VGND sg13g2_nand2_1
XFILLER_21_164 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_29_220 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_12_120 VPWR VGND sg13g2_decap_8
XFILLER_16_72 VPWR VGND sg13g2_decap_8
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_12_197 VPWR VGND sg13g2_decap_8
XFILLER_13_687 VPWR VGND sg13g2_fill_2
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_5_820 VPWR VGND sg13g2_fill_2
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
X_1390_ VPWR _0042_ state\[22\] VGND sg13g2_inv_1
XFILLER_35_245 VPWR VGND sg13g2_decap_8
X_2011_ state\[119\] daisychain\[119\] net153 _0682_ VPWR VGND sg13g2_mux2_1
XFILLER_12_19 VPWR VGND sg13g2_fill_1
X_2844_ daisychain\[124\] net19 VPWR VGND sg13g2_buf_1
X_1726_ state\[62\] daisychain\[62\] net147 _0454_ VPWR VGND sg13g2_mux2_1
X_1657_ _0399_ net169 _0398_ VPWR VGND sg13g2_nand2_1
X_1588_ VGND VPWR net105 daisychain\[33\] _0988_ net51 sg13g2_a21oi_1
XFILLER_37_49 VPWR VGND sg13g2_decap_8
X_2209_ VGND VPWR _0511_ _0794_ _0332_ net85 sg13g2_a21oi_1
XFILLER_22_451 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_42_716 VPWR VGND sg13g2_fill_2
XFILLER_6_628 VPWR VGND sg13g2_decap_4
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_17_267 VPWR VGND sg13g2_decap_8
XFILLER_45_587 VPWR VGND sg13g2_fill_2
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_9_400 VPWR VGND sg13g2_decap_8
XFILLER_9_411 VPWR VGND sg13g2_fill_1
XFILLER_4_171 VPWR VGND sg13g2_decap_8
XFILLER_5_661 VPWR VGND sg13g2_fill_2
X_1442_ _0871_ net159 _0870_ VPWR VGND sg13g2_nand2_1
X_1511_ state\[19\] daisychain\[19\] net137 _0926_ VPWR VGND sg13g2_mux2_1
X_2560_ net341 VGND VPWR _0376_ state\[120\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2491_ net379 VGND VPWR _0307_ state\[51\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1373_ VPWR _0060_ state\[39\] VGND sg13g2_inv_1
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_36_532 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_31_270 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
X_1709_ net192 VPWR _0441_ VGND daisychain\[58\] net37 sg13g2_o21ai_1
XFILLER_42_513 VPWR VGND sg13g2_fill_1
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_14_259 VPWR VGND sg13g2_decap_8
Xfanout30 net44 net30 VPWR VGND sg13g2_buf_1
Xfanout96 net97 net96 VPWR VGND sg13g2_buf_1
Xfanout85 net86 net85 VPWR VGND sg13g2_buf_1
Xfanout74 net88 net74 VPWR VGND sg13g2_buf_1
Xfanout63 net64 net63 VPWR VGND sg13g2_buf_1
Xfanout52 net66 net52 VPWR VGND sg13g2_buf_1
Xfanout41 net42 net41 VPWR VGND sg13g2_buf_1
X_2450__288 VPWR VGND net287 sg13g2_tiehi
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_6_414 VPWR VGND sg13g2_decap_8
XFILLER_6_447 VPWR VGND sg13g2_decap_4
XFILLER_6_469 VPWR VGND sg13g2_fill_1
XFILLER_18_510 VPWR VGND sg13g2_fill_1
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_fill_2
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_38_819 VPWR VGND sg13g2_decap_4
XFILLER_49_123 VPWR VGND sg13g2_decap_8
X_2392__423 VPWR VGND net422 sg13g2_tiehi
XFILLER_13_270 VPWR VGND sg13g2_decap_8
XFILLER_20_229 VPWR VGND sg13g2_decap_8
XFILLER_41_590 VPWR VGND sg13g2_decap_4
XFILLER_9_274 VPWR VGND sg13g2_decap_8
Xclkload11 VPWR clkload11/Y clknet_leaf_13_clk VGND sg13g2_inv_1
X_1991_ state\[115\] daisychain\[115\] net135 _0666_ VPWR VGND sg13g2_mux2_1
X_1425_ VGND VPWR _0855_ _0856_ _0129_ _0857_ sg13g2_a21oi_1
X_2543_ net221 VGND VPWR _0359_ state\[103\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2474_ net447 VGND VPWR _0290_ state\[34\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1287_ VPWR _0028_ state\[125\] VGND sg13g2_inv_1
X_1356_ VPWR _0079_ state\[56\] VGND sg13g2_inv_1
X_2438__331 VPWR VGND net330 sg13g2_tiehi
XFILLER_11_229 VPWR VGND sg13g2_decap_8
XFILLER_20_752 VPWR VGND sg13g2_fill_1
XFILLER_34_28 VPWR VGND sg13g2_decap_8
Xclkload5 clkload5/Y clknet_leaf_0_clk VPWR VGND sg13g2_inv_8
XFILLER_20_785 VPWR VGND sg13g2_fill_1
XFILLER_3_406 VPWR VGND sg13g2_decap_8
XFILLER_19_307 VPWR VGND sg13g2_fill_1
XFILLER_19_318 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_15_524 VPWR VGND sg13g2_fill_1
XFILLER_27_362 VPWR VGND sg13g2_decap_8
XFILLER_27_373 VPWR VGND sg13g2_fill_2
XFILLER_27_395 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_43_822 VPWR VGND sg13g2_fill_1
XFILLER_46_126 VPWR VGND sg13g2_decap_8
X_2339__273 VPWR VGND net272 sg13g2_tiehi
XFILLER_10_251 VPWR VGND sg13g2_decap_8
XFILLER_24_83 VPWR VGND sg13g2_decap_8
XFILLER_24_94 VPWR VGND sg13g2_fill_1
XFILLER_6_211 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_6_288 VPWR VGND sg13g2_decap_8
XFILLER_7_778 VPWR VGND sg13g2_decap_8
XFILLER_18_351 VPWR VGND sg13g2_decap_4
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
X_2190_ _0785_ net128 state\[67\] VPWR VGND sg13g2_nand2_1
X_1974_ net189 VPWR _0653_ VGND daisychain\[111\] net34 sg13g2_o21ai_1
XFILLER_29_17 VPWR VGND sg13g2_decap_8
X_1408_ VPWR _0072_ state\[4\] VGND sg13g2_inv_1
X_2526_ net409 VGND VPWR _0342_ state\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2457_ net259 VGND VPWR _0273_ state\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2388_ net430 VGND VPWR _0204_ daisychain\[76\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
X_1339_ VPWR _0098_ state\[73\] VGND sg13g2_inv_1
XFILLER_24_365 VPWR VGND sg13g2_decap_8
XFILLER_24_376 VPWR VGND sg13g2_fill_1
XFILLER_10_41 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
XFILLER_19_148 VPWR VGND sg13g2_decap_8
XFILLER_19_50 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_30_302 VPWR VGND sg13g2_decap_8
XFILLER_30_346 VPWR VGND sg13g2_fill_1
XFILLER_31_814 VPWR VGND sg13g2_decap_4
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_43_685 VPWR VGND sg13g2_fill_1
XFILLER_30_379 VPWR VGND sg13g2_decap_4
X_1690_ VGND VPWR _0423_ _0424_ _0182_ _0425_ sg13g2_a21oi_1
XFILLER_2_280 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
X_2311_ VGND VPWR _0715_ _0845_ _0383_ net70 sg13g2_a21oi_1
X_2242_ _0811_ net110 state\[93\] VPWR VGND sg13g2_nand2_1
XFILLER_46_490 VPWR VGND sg13g2_decap_8
X_2173_ VGND VPWR _0439_ _0776_ _0314_ net82 sg13g2_a21oi_1
XFILLER_21_302 VPWR VGND sg13g2_decap_4
XFILLER_31_18 VPWR VGND sg13g2_decap_8
XFILLER_33_151 VPWR VGND sg13g2_decap_8
X_1957_ _0639_ net164 _0638_ VPWR VGND sg13g2_nand2_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[3] VPWR VGND sg13g2_buf_1
X_2509_ net289 VGND VPWR _0325_ state\[69\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1888_ VGND VPWR net110 daisychain\[93\] _0584_ net55 sg13g2_a21oi_1
XFILLER_29_479 VPWR VGND sg13g2_decap_8
XFILLER_12_302 VPWR VGND sg13g2_decap_8
XFILLER_16_107 VPWR VGND sg13g2_decap_8
XFILLER_24_195 VPWR VGND sg13g2_decap_8
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_21_73 VPWR VGND sg13g2_decap_8
XFILLER_4_512 VPWR VGND sg13g2_decap_8
XFILLER_16_652 VPWR VGND sg13g2_decap_8
XFILLER_35_416 VPWR VGND sg13g2_fill_1
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_15_184 VPWR VGND sg13g2_decap_8
XFILLER_30_165 VPWR VGND sg13g2_decap_8
XFILLER_31_688 VPWR VGND sg13g2_decap_8
X_1811_ state\[79\] daisychain\[79\] net151 _0522_ VPWR VGND sg13g2_mux2_1
XFILLER_7_361 VPWR VGND sg13g2_decap_8
XFILLER_7_86 VPWR VGND sg13g2_decap_8
X_1742_ _0467_ net175 _0466_ VPWR VGND sg13g2_nand2_1
X_1673_ VGND VPWR net119 daisychain\[50\] _0412_ net59 sg13g2_a21oi_1
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_39_744 VPWR VGND sg13g2_decap_8
X_2225_ VGND VPWR _0543_ _0802_ _0340_ net83 sg13g2_a21oi_1
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_38_287 VPWR VGND sg13g2_decap_8
XFILLER_41_408 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_2_1__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_2156_ _0768_ net120 state\[50\] VPWR VGND sg13g2_nand2_1
X_2087_ VGND VPWR _0911_ _0733_ _0271_ net68 sg13g2_a21oi_1
XFILLER_21_143 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_fill_2
XFILLER_1_537 VPWR VGND sg13g2_fill_2
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_12_176 VPWR VGND sg13g2_decap_8
XFILLER_13_666 VPWR VGND sg13g2_decap_8
XFILLER_16_51 VPWR VGND sg13g2_decap_8
XFILLER_4_353 VPWR VGND sg13g2_decap_8
XFILLER_8_158 VPWR VGND sg13g2_decap_8
X_2540__270 VPWR VGND net269 sg13g2_tiehi
X_2010_ VGND VPWR _0679_ _0680_ _0246_ _0681_ sg13g2_a21oi_1
XFILLER_16_482 VPWR VGND sg13g2_fill_1
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_31_430 VPWR VGND sg13g2_decap_8
XFILLER_31_496 VPWR VGND sg13g2_fill_1
X_2843_ daisychain\[123\] net18 VPWR VGND sg13g2_buf_1
X_1725_ VGND VPWR _0451_ _0452_ _0189_ _0453_ sg13g2_a21oi_1
Xclkbuf_leaf_7_clk clknet_2_3__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_1656_ state\[48\] daisychain\[48\] net145 _0398_ VPWR VGND sg13g2_mux2_1
X_1587_ _0987_ net161 _0986_ VPWR VGND sg13g2_nand2_1
XFILLER_26_246 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_39_530 VPWR VGND sg13g2_fill_2
X_2208_ _0794_ net127 state\[76\] VPWR VGND sg13g2_nand2_1
X_2139_ VGND VPWR _1015_ _0759_ _0297_ net79 sg13g2_a21oi_1
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_fill_1
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
X_2379__449 VPWR VGND net448 sg13g2_tiehi
XFILLER_17_246 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_fill_1
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_13_485 VPWR VGND sg13g2_decap_4
XFILLER_32_249 VPWR VGND sg13g2_decap_8
X_2349__253 VPWR VGND net252 sg13g2_tiehi
XFILLER_4_150 VPWR VGND sg13g2_decap_8
X_1441_ state\[5\] daisychain\[5\] net137 _0870_ VPWR VGND sg13g2_mux2_1
X_1510_ VGND VPWR _0923_ _0924_ _0146_ _0925_ sg13g2_a21oi_1
X_2490_ net383 VGND VPWR _0306_ state\[50\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_4_87 VPWR VGND sg13g2_decap_8
X_1372_ VPWR _0062_ state\[40\] VGND sg13g2_inv_1
XFILLER_23_249 VPWR VGND sg13g2_decap_8
XFILLER_36_577 VPWR VGND sg13g2_fill_1
X_1708_ VGND VPWR net121 daisychain\[57\] _0440_ net59 sg13g2_a21oi_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_1639_ net190 VPWR _0385_ VGND daisychain\[44\] net35 sg13g2_o21ai_1
XFILLER_14_238 VPWR VGND sg13g2_decap_8
XFILLER_42_525 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_13_41 VPWR VGND sg13g2_fill_1
XFILLER_13_74 VPWR VGND sg13g2_decap_8
Xfanout31 net34 net31 VPWR VGND sg13g2_buf_1
Xfanout97 net98 net97 VPWR VGND sg13g2_buf_1
Xfanout86 net87 net86 VPWR VGND sg13g2_buf_1
Xfanout75 net78 net75 VPWR VGND sg13g2_buf_1
Xfanout64 net65 net64 VPWR VGND sg13g2_buf_1
Xfanout53 net56 net53 VPWR VGND sg13g2_buf_1
Xfanout42 net43 net42 VPWR VGND sg13g2_buf_1
XFILLER_2_643 VPWR VGND sg13g2_fill_1
XFILLER_18_500 VPWR VGND sg13g2_fill_2
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_46_820 VPWR VGND sg13g2_fill_2
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_fill_2
XFILLER_20_208 VPWR VGND sg13g2_decap_8
XFILLER_45_385 VPWR VGND sg13g2_decap_8
X_1990_ VGND VPWR _0663_ _0664_ _0242_ _0665_ sg13g2_a21oi_1
XFILLER_9_253 VPWR VGND sg13g2_decap_8
X_2542_ net237 VGND VPWR _0358_ state\[102\] clknet_leaf_9_clk sg13g2_dfrbpq_1
Xclkload12 clkload12/Y clknet_leaf_4_clk VPWR VGND sg13g2_inv_2
X_1355_ VPWR _0080_ state\[57\] VGND sg13g2_inv_1
X_1424_ net180 VPWR _0857_ VGND daisychain\[1\] net24 sg13g2_o21ai_1
X_2473_ net451 VGND VPWR _0289_ state\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_24_503 VPWR VGND sg13g2_decap_8
XFILLER_36_385 VPWR VGND sg13g2_decap_4
X_1286_ VPWR _0029_ state\[126\] VGND sg13g2_inv_1
XFILLER_11_208 VPWR VGND sg13g2_decap_8
XFILLER_20_731 VPWR VGND sg13g2_fill_1
XFILLER_20_764 VPWR VGND sg13g2_fill_2
Xclkload6 VPWR clkload6/Y clknet_leaf_2_clk VGND sg13g2_inv_1
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_43_801 VPWR VGND sg13g2_fill_2
XFILLER_10_230 VPWR VGND sg13g2_decap_8
XFILLER_24_62 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_4
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_6_267 VPWR VGND sg13g2_decap_8
XFILLER_7_746 VPWR VGND sg13g2_fill_2
XFILLER_7_757 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_2_462 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_fill_1
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_21_517 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_decap_8
X_1973_ VGND VPWR net96 daisychain\[110\] _0652_ net56 sg13g2_a21oi_1
X_2525_ net417 VGND VPWR _0341_ state\[85\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_116 VPWR VGND sg13g2_decap_8
X_1338_ VPWR _0099_ state\[74\] VGND sg13g2_inv_1
X_1407_ VPWR _0083_ state\[5\] VGND sg13g2_inv_1
X_2456_ net263 VGND VPWR _0272_ state\[16\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2405__397 VPWR VGND net396 sg13g2_tiehi
X_2387_ net432 VGND VPWR _0203_ daisychain\[75\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_12_506 VPWR VGND sg13g2_decap_4
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_40_815 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_10_97 VPWR VGND sg13g2_decap_8
XFILLER_3_259 VPWR VGND sg13g2_decap_8
XFILLER_4_738 VPWR VGND sg13g2_fill_1
XFILLER_15_311 VPWR VGND sg13g2_fill_1
XFILLER_19_127 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_38_414 VPWR VGND sg13g2_fill_1
X_2310_ _0845_ state\[127\] net90 VPWR VGND sg13g2_nand2_1
X_2241_ VGND VPWR _0575_ _0810_ _0348_ net83 sg13g2_a21oi_1
X_2172_ _0776_ net121 state\[58\] VPWR VGND sg13g2_nand2_1
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_19_661 VPWR VGND sg13g2_decap_8
XFILLER_19_672 VPWR VGND sg13g2_fill_1
XFILLER_33_130 VPWR VGND sg13g2_decap_8
XFILLER_34_686 VPWR VGND sg13g2_decap_8
XFILLER_38_469 VPWR VGND sg13g2_fill_1
XFILLER_34_697 VPWR VGND sg13g2_decap_4
X_1956_ state\[108\] daisychain\[108\] net143 _0638_ VPWR VGND sg13g2_mux2_1
X_1887_ _0583_ net165 _0582_ VPWR VGND sg13g2_nand2_1
Xoutput19 net19 uo_out[4] VPWR VGND sg13g2_buf_1
X_2508_ net297 VGND VPWR _0324_ state\[68\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_44_406 VPWR VGND sg13g2_decap_8
X_2439_ net328 VGND VPWR _0255_ daisychain\[127\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_13_815 VPWR VGND sg13g2_decap_8
XFILLER_24_174 VPWR VGND sg13g2_decap_8
XFILLER_37_480 VPWR VGND sg13g2_fill_1
XFILLER_21_52 VPWR VGND sg13g2_decap_8
XFILLER_0_785 VPWR VGND sg13g2_decap_8
XFILLER_48_734 VPWR VGND sg13g2_decap_8
XFILLER_16_642 VPWR VGND sg13g2_fill_1
XFILLER_35_439 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_fill_1
XFILLER_15_163 VPWR VGND sg13g2_decap_8
XFILLER_30_144 VPWR VGND sg13g2_decap_8
XFILLER_31_656 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_7_340 VPWR VGND sg13g2_decap_8
X_2389__429 VPWR VGND net428 sg13g2_tiehi
X_1810_ VGND VPWR _0519_ _0520_ _0206_ _0521_ sg13g2_a21oi_1
X_1741_ state\[65\] daisychain\[65\] net151 _0466_ VPWR VGND sg13g2_mux2_1
X_2506__314 VPWR VGND net313 sg13g2_tiehi
X_1672_ _0411_ net170 _0410_ VPWR VGND sg13g2_nand2_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_39_712 VPWR VGND sg13g2_decap_4
X_2552__334 VPWR VGND net333 sg13g2_tiehi
X_2359__233 VPWR VGND net232 sg13g2_tiehi
X_2224_ _0802_ net125 state\[84\] VPWR VGND sg13g2_nand2_1
X_2155_ VGND VPWR _0403_ _0767_ _0305_ net80 sg13g2_a21oi_1
XFILLER_21_122 VPWR VGND sg13g2_decap_8
XFILLER_34_483 VPWR VGND sg13g2_fill_2
X_2086_ _0733_ net92 state\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_21_199 VPWR VGND sg13g2_decap_8
X_1939_ net186 VPWR _0625_ VGND daisychain\[104\] net31 sg13g2_o21ai_1
XFILLER_29_255 VPWR VGND sg13g2_fill_2
XFILLER_44_203 VPWR VGND sg13g2_decap_8
X_2518__218 VPWR VGND net217 sg13g2_tiehi
X_2453__276 VPWR VGND net275 sg13g2_tiehi
XFILLER_12_155 VPWR VGND sg13g2_decap_8
XFILLER_25_483 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_5_822 VPWR VGND sg13g2_fill_1
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_fill_1
XFILLER_43_280 VPWR VGND sg13g2_decap_8
XFILLER_8_660 VPWR VGND sg13g2_decap_8
X_2547__414 VPWR VGND net413 sg13g2_tiehi
X_2842_ daisychain\[122\] net17 VPWR VGND sg13g2_buf_1
X_1724_ net193 VPWR _0453_ VGND daisychain\[61\] net38 sg13g2_o21ai_1
X_1655_ VGND VPWR _0395_ _0396_ _0175_ _0397_ sg13g2_a21oi_1
X_1586_ state\[34\] daisychain\[34\] net139 _0986_ VPWR VGND sg13g2_mux2_1
XFILLER_26_225 VPWR VGND sg13g2_decap_8
XFILLER_42_718 VPWR VGND sg13g2_fill_1
XFILLER_42_729 VPWR VGND sg13g2_decap_8
X_2207_ VGND VPWR _0507_ _0793_ _0331_ net85 sg13g2_a21oi_1
X_2138_ _0759_ net116 state\[41\] VPWR VGND sg13g2_nand2_1
X_2069_ VGND VPWR _0875_ _0724_ _0262_ net71 sg13g2_a21oi_1
XFILLER_10_604 VPWR VGND sg13g2_fill_2
XFILLER_10_648 VPWR VGND sg13g2_fill_2
XFILLER_22_486 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_5_118 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_17_225 VPWR VGND sg13g2_decap_8
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_45_534 VPWR VGND sg13g2_decap_8
XFILLER_45_589 VPWR VGND sg13g2_fill_1
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_5_641 VPWR VGND sg13g2_fill_2
XFILLER_5_674 VPWR VGND sg13g2_fill_2
X_1371_ VPWR _0063_ state\[41\] VGND sg13g2_inv_1
X_1440_ VGND VPWR _0867_ _0868_ _0132_ _0869_ sg13g2_a21oi_1
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_23_228 VPWR VGND sg13g2_decap_8
X_1707_ _0439_ net171 _0438_ VPWR VGND sg13g2_nand2_1
X_1638_ VGND VPWR net116 daisychain\[43\] _0384_ net58 sg13g2_a21oi_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_1569_ net185 VPWR _0973_ VGND daisychain\[30\] net30 sg13g2_o21ai_1
XFILLER_14_217 VPWR VGND sg13g2_decap_8
XFILLER_39_394 VPWR VGND sg13g2_decap_8
X_2415__377 VPWR VGND net376 sg13g2_tiehi
XFILLER_10_478 VPWR VGND sg13g2_fill_1
XFILLER_13_53 VPWR VGND sg13g2_decap_8
Xfanout32 net33 net32 VPWR VGND sg13g2_buf_1
Xfanout98 _0846_ net98 VPWR VGND sg13g2_buf_1
Xfanout87 net88 net87 VPWR VGND sg13g2_buf_1
Xfanout76 net78 net76 VPWR VGND sg13g2_buf_1
Xfanout65 net66 net65 VPWR VGND sg13g2_buf_1
Xfanout54 net55 net54 VPWR VGND sg13g2_buf_1
Xfanout43 net44 net43 VPWR VGND sg13g2_buf_1
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_2_611 VPWR VGND sg13g2_fill_2
XFILLER_2_699 VPWR VGND sg13g2_fill_1
XFILLER_18_578 VPWR VGND sg13g2_decap_4
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_33_548 VPWR VGND sg13g2_fill_2
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_9_232 VPWR VGND sg13g2_decap_8
X_2541_ net253 VGND VPWR _0357_ state\[101\] clknet_leaf_4_clk sg13g2_dfrbpq_1
Xclkload13 VPWR clkload13/Y clknet_leaf_7_clk VGND sg13g2_inv_1
X_2472_ net VGND VPWR _0288_ state\[32\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1285_ VPWR _0846_ net154 VGND sg13g2_inv_1
X_1354_ VPWR _0081_ state\[58\] VGND sg13g2_inv_1
X_1423_ VGND VPWR net97 daisychain\[0\] _0856_ net47 sg13g2_a21oi_1
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_36_397 VPWR VGND sg13g2_fill_2
XFILLER_20_710 VPWR VGND sg13g2_fill_2
Xclkload7 VPWR clkload7/Y clknet_leaf_17_clk VGND sg13g2_inv_1
XFILLER_39_191 VPWR VGND sg13g2_decap_8
XFILLER_24_41 VPWR VGND sg13g2_decap_8
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_10_286 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_6_246 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
XFILLER_2_485 VPWR VGND sg13g2_decap_8
XFILLER_2_496 VPWR VGND sg13g2_fill_2
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_19_810 VPWR VGND sg13g2_fill_1
XFILLER_19_821 VPWR VGND sg13g2_fill_2
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_33_312 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_46_673 VPWR VGND sg13g2_decap_8
X_2318__315 VPWR VGND net314 sg13g2_tiehi
X_1972_ _0651_ net167 _0650_ VPWR VGND sg13g2_nand2_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2524_ net425 VGND VPWR _0340_ state\[84\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2455_ net267 VGND VPWR _0271_ state\[15\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2399__409 VPWR VGND net408 sg13g2_tiehi
X_1337_ VPWR _0100_ state\[75\] VGND sg13g2_inv_1
X_1406_ VPWR _0094_ state\[6\] VGND sg13g2_inv_1
X_2386_ net434 VGND VPWR _0202_ daisychain\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_161 VPWR VGND sg13g2_decap_8
X_2369__213 VPWR VGND net212 sg13g2_tiehi
XFILLER_10_10 VPWR VGND sg13g2_fill_1
XFILLER_10_21 VPWR VGND sg13g2_fill_2
XFILLER_20_584 VPWR VGND sg13g2_decap_4
X_2449__292 VPWR VGND net291 sg13g2_tiehi
XFILLER_10_76 VPWR VGND sg13g2_decap_8
XFILLER_3_238 VPWR VGND sg13g2_decap_8
XFILLER_19_106 VPWR VGND sg13g2_decap_8
XFILLER_19_85 VPWR VGND sg13g2_decap_8
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_43_643 VPWR VGND sg13g2_decap_4
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_30_337 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_3_761 VPWR VGND sg13g2_fill_2
XFILLER_38_448 VPWR VGND sg13g2_decap_8
X_2240_ _0810_ net126 state\[92\] VPWR VGND sg13g2_nand2_1
X_2171_ VGND VPWR _0435_ _0775_ _0313_ net81 sg13g2_a21oi_1
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_19_684 VPWR VGND sg13g2_decap_8
XFILLER_21_337 VPWR VGND sg13g2_decap_8
XFILLER_33_186 VPWR VGND sg13g2_decap_8
X_1955_ VGND VPWR _0635_ _0636_ _0235_ _0637_ sg13g2_a21oi_1
X_1886_ state\[94\] daisychain\[94\] net142 _0582_ VPWR VGND sg13g2_mux2_1
X_2557__438 VPWR VGND net437 sg13g2_tiehi
X_2507_ net305 VGND VPWR _0323_ state\[67\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2438_ net330 VGND VPWR _0254_ daisychain\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_37_492 VPWR VGND sg13g2_decap_8
X_2369_ net212 VGND VPWR _0185_ daisychain\[57\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_12_337 VPWR VGND sg13g2_decap_8
XFILLER_24_153 VPWR VGND sg13g2_decap_8
XFILLER_40_668 VPWR VGND sg13g2_fill_2
XFILLER_40_679 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_20_392 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_15_142 VPWR VGND sg13g2_decap_8
XFILLER_31_602 VPWR VGND sg13g2_decap_8
XFILLER_35_429 VPWR VGND sg13g2_fill_2
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_30_123 VPWR VGND sg13g2_decap_8
XFILLER_7_33 VPWR VGND sg13g2_decap_8
XFILLER_7_44 VPWR VGND sg13g2_fill_1
X_1740_ VGND VPWR _0463_ _0464_ _0192_ _0465_ sg13g2_a21oi_1
X_1671_ state\[51\] daisychain\[51\] net146 _0410_ VPWR VGND sg13g2_mux2_1
XFILLER_7_396 VPWR VGND sg13g2_decap_8
XFILLER_38_245 VPWR VGND sg13g2_decap_8
X_2223_ VGND VPWR _0539_ _0801_ _0339_ net83 sg13g2_a21oi_1
X_2154_ _0767_ net118 state\[49\] VPWR VGND sg13g2_nand2_1
X_2085_ VGND VPWR _0907_ _0732_ _0270_ net67 sg13g2_a21oi_1
XFILLER_10_808 VPWR VGND sg13g2_decap_8
XFILLER_21_101 VPWR VGND sg13g2_decap_8
XFILLER_21_178 VPWR VGND sg13g2_decap_8
XFILLER_1_506 VPWR VGND sg13g2_fill_1
X_2524__426 VPWR VGND net425 sg13g2_tiehi
X_1938_ VGND VPWR net107 daisychain\[103\] _0624_ net53 sg13g2_a21oi_1
X_1869_ net197 VPWR _0569_ VGND daisychain\[90\] net42 sg13g2_o21ai_1
XFILLER_29_234 VPWR VGND sg13g2_decap_8
XFILLER_16_86 VPWR VGND sg13g2_decap_8
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_12_134 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_9_639 VPWR VGND sg13g2_decap_4
XFILLER_4_311 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_decap_8
X_2460__248 VPWR VGND net247 sg13g2_tiehi
X_2425__357 VPWR VGND net356 sg13g2_tiehi
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_16_462 VPWR VGND sg13g2_fill_2
XFILLER_16_473 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
X_2841_ daisychain\[121\] net16 VPWR VGND sg13g2_buf_1
XFILLER_7_193 VPWR VGND sg13g2_decap_8
XFILLER_8_672 VPWR VGND sg13g2_decap_4
XFILLER_8_683 VPWR VGND sg13g2_decap_8
X_1723_ VGND VPWR net121 daisychain\[60\] _0452_ net60 sg13g2_a21oi_1
X_1654_ net191 VPWR _0397_ VGND daisychain\[47\] net36 sg13g2_o21ai_1
X_2326__299 VPWR VGND net298 sg13g2_tiehi
X_2206_ _0793_ net127 state\[75\] VPWR VGND sg13g2_nand2_1
X_1585_ VGND VPWR _0983_ _0984_ _0161_ _0985_ sg13g2_a21oi_1
XFILLER_26_204 VPWR VGND sg13g2_decap_8
X_2137_ VGND VPWR _1011_ _0758_ _0296_ net79 sg13g2_a21oi_1
X_2068_ _0724_ net101 state\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_22_465 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_17_204 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_13_443 VPWR VGND sg13g2_fill_1
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_41_763 VPWR VGND sg13g2_fill_2
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_9_447 VPWR VGND sg13g2_decap_8
XFILLER_4_185 VPWR VGND sg13g2_decap_8
XFILLER_4_23 VPWR VGND sg13g2_fill_2
X_1370_ VPWR _0064_ state\[42\] VGND sg13g2_inv_1
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_36_546 VPWR VGND sg13g2_fill_1
XFILLER_31_284 VPWR VGND sg13g2_decap_8
XFILLER_8_480 VPWR VGND sg13g2_fill_2
X_1706_ state\[58\] daisychain\[58\] net147 _0438_ VPWR VGND sg13g2_mux2_1
X_1637_ _1027_ net168 _1026_ VPWR VGND sg13g2_nand2_1
XFILLER_39_373 VPWR VGND sg13g2_decap_8
X_1499_ net181 VPWR _0917_ VGND daisychain\[16\] net25 sg13g2_o21ai_1
X_2378__451 VPWR VGND net450 sg13g2_tiehi
X_1568_ VGND VPWR net102 daisychain\[29\] _0972_ net50 sg13g2_a21oi_1
Xfanout33 net34 net33 VPWR VGND sg13g2_buf_1
Xfanout55 net56 net55 VPWR VGND sg13g2_buf_1
Xfanout44 _0851_ net44 VPWR VGND sg13g2_buf_1
XFILLER_10_435 VPWR VGND sg13g2_fill_2
XFILLER_10_457 VPWR VGND sg13g2_decap_8
XFILLER_6_428 VPWR VGND sg13g2_decap_8
Xfanout99 net103 net99 VPWR VGND sg13g2_buf_1
Xfanout88 _0847_ net88 VPWR VGND sg13g2_buf_1
Xfanout77 net78 net77 VPWR VGND sg13g2_buf_1
Xfanout66 _0850_ net66 VPWR VGND sg13g2_buf_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_623 VPWR VGND sg13g2_decap_8
XFILLER_2_656 VPWR VGND sg13g2_decap_8
XFILLER_2_667 VPWR VGND sg13g2_fill_2
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_18_502 VPWR VGND sg13g2_fill_1
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_fill_1
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_9_211 VPWR VGND sg13g2_decap_8
XFILLER_5_483 VPWR VGND sg13g2_decap_8
XFILLER_9_288 VPWR VGND sg13g2_decap_8
X_1422_ _0855_ net155 _0854_ VPWR VGND sg13g2_nand2_1
X_2540_ net269 VGND VPWR _0356_ state\[100\] clknet_leaf_4_clk sg13g2_dfrbpq_1
Xclkload14 VPWR clkload14/Y clknet_leaf_8_clk VGND sg13g2_inv_1
X_2471_ net203 VGND VPWR _0287_ state\[31\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1284_ VPWR _0030_ state\[127\] VGND sg13g2_inv_1
X_1353_ VPWR _0082_ state\[59\] VGND sg13g2_inv_1
XFILLER_24_516 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_20_744 VPWR VGND sg13g2_fill_1
XFILLER_20_777 VPWR VGND sg13g2_fill_1
Xclkload8 clkload8/Y clknet_leaf_18_clk VPWR VGND sg13g2_inv_8
XFILLER_27_343 VPWR VGND sg13g2_fill_2
XFILLER_39_170 VPWR VGND sg13g2_decap_8
XFILLER_43_803 VPWR VGND sg13g2_fill_1
XFILLER_11_711 VPWR VGND sg13g2_fill_1
XFILLER_24_20 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_10_265 VPWR VGND sg13g2_decap_8
XFILLER_2_420 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_fill_1
XFILLER_6_225 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_18_343 VPWR VGND sg13g2_fill_2
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_14_571 VPWR VGND sg13g2_fill_1
X_1971_ state\[111\] daisychain\[111\] net135 _0650_ VPWR VGND sg13g2_mux2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_1405_ VPWR _0105_ state\[7\] VGND sg13g2_inv_1
X_2523_ net433 VGND VPWR _0339_ state\[83\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2454_ net271 VGND VPWR _0270_ state\[14\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2385_ net436 VGND VPWR _0201_ daisychain\[73\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_37_685 VPWR VGND sg13g2_fill_2
X_1336_ VPWR _0101_ state\[76\] VGND sg13g2_inv_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
XFILLER_20_541 VPWR VGND sg13g2_fill_2
XFILLER_10_55 VPWR VGND sg13g2_decap_8
XFILLER_20_563 VPWR VGND sg13g2_decap_8
XFILLER_20_596 VPWR VGND sg13g2_fill_2
XFILLER_3_217 VPWR VGND sg13g2_decap_8
X_2527__402 VPWR VGND net401 sg13g2_tiehi
XFILLER_19_64 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_15_346 VPWR VGND sg13g2_decap_8
XFILLER_16_814 VPWR VGND sg13g2_decap_8
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_43_666 VPWR VGND sg13g2_fill_1
X_2456__264 VPWR VGND net263 sg13g2_tiehi
XFILLER_7_578 VPWR VGND sg13g2_decap_8
XFILLER_7_589 VPWR VGND sg13g2_fill_1
XFILLER_18_151 VPWR VGND sg13g2_decap_8
XFILLER_2_294 VPWR VGND sg13g2_decap_8
X_2435__337 VPWR VGND net336 sg13g2_tiehi
X_2170_ _0775_ net121 state\[57\] VPWR VGND sg13g2_nand2_1
XFILLER_33_165 VPWR VGND sg13g2_decap_8
XFILLER_34_666 VPWR VGND sg13g2_fill_1
X_1954_ net186 VPWR _0637_ VGND daisychain\[107\] net31 sg13g2_o21ai_1
X_1885_ VGND VPWR _0579_ _0580_ _0221_ _0581_ sg13g2_a21oi_1
X_2506_ net313 VGND VPWR _0322_ state\[66\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2437_ net332 VGND VPWR _0253_ daisychain\[125\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2368_ net214 VGND VPWR _0184_ daisychain\[56\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_24_132 VPWR VGND sg13g2_decap_8
XFILLER_40_603 VPWR VGND sg13g2_fill_1
X_1319_ VPWR _0120_ state\[93\] VGND sg13g2_inv_1
X_2336__279 VPWR VGND net278 sg13g2_tiehi
X_2299_ VGND VPWR _0691_ _0839_ _0377_ net70 sg13g2_a21oi_1
XFILLER_12_316 VPWR VGND sg13g2_decap_8
XFILLER_20_360 VPWR VGND sg13g2_decap_8
XFILLER_40_614 VPWR VGND sg13g2_fill_1
XFILLER_21_87 VPWR VGND sg13g2_decap_8
XFILLER_4_526 VPWR VGND sg13g2_fill_2
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_15_121 VPWR VGND sg13g2_decap_8
XFILLER_15_198 VPWR VGND sg13g2_decap_8
XFILLER_16_622 VPWR VGND sg13g2_decap_4
XFILLER_16_633 VPWR VGND sg13g2_decap_4
XFILLER_16_666 VPWR VGND sg13g2_decap_8
XFILLER_30_102 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_30_179 VPWR VGND sg13g2_decap_8
XFILLER_7_375 VPWR VGND sg13g2_decap_8
X_1670_ VGND VPWR _0407_ _0408_ _0178_ _0409_ sg13g2_a21oi_1
XFILLER_30_4 VPWR VGND sg13g2_decap_4
X_2222_ _0801_ net125 state\[83\] VPWR VGND sg13g2_nand2_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
XFILLER_38_224 VPWR VGND sg13g2_decap_8
XFILLER_39_758 VPWR VGND sg13g2_decap_8
XFILLER_39_769 VPWR VGND sg13g2_decap_4
X_2153_ VGND VPWR _0399_ _0766_ _0304_ net80 sg13g2_a21oi_1
X_2084_ _0732_ net92 state\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_21_157 VPWR VGND sg13g2_decap_8
XFILLER_34_496 VPWR VGND sg13g2_decap_8
X_1937_ _0623_ net164 _0622_ VPWR VGND sg13g2_nand2_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
X_1868_ VGND VPWR net124 daisychain\[89\] _0568_ net61 sg13g2_a21oi_1
X_1799_ net195 VPWR _0513_ VGND daisychain\[76\] net40 sg13g2_o21ai_1
XFILLER_29_213 VPWR VGND sg13g2_decap_8
XFILLER_29_257 VPWR VGND sg13g2_fill_1
XFILLER_12_113 VPWR VGND sg13g2_decap_8
XFILLER_16_65 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_5_813 VPWR VGND sg13g2_decap_8
X_2388__431 VPWR VGND net430 sg13g2_tiehi
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
X_2840_ daisychain\[120\] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_172 VPWR VGND sg13g2_decap_8
X_1722_ _0451_ net171 _0450_ VPWR VGND sg13g2_nand2_1
X_1653_ VGND VPWR net117 daisychain\[46\] _0396_ net58 sg13g2_a21oi_1
X_1584_ net184 VPWR _0985_ VGND daisychain\[33\] net29 sg13g2_o21ai_1
XFILLER_39_577 VPWR VGND sg13g2_fill_1
X_2205_ VGND VPWR _0503_ _0792_ _0330_ net83 sg13g2_a21oi_1
XFILLER_22_444 VPWR VGND sg13g2_decap_8
XFILLER_35_761 VPWR VGND sg13g2_fill_1
X_2136_ _0758_ net115 state\[40\] VPWR VGND sg13g2_nand2_1
X_2067_ VGND VPWR _0871_ _0723_ _0261_ net71 sg13g2_a21oi_1
XFILLER_10_606 VPWR VGND sg13g2_fill_1
X_2487__396 VPWR VGND net395 sg13g2_tiehi
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_45_525 VPWR VGND sg13g2_decap_4
XFILLER_13_411 VPWR VGND sg13g2_decap_4
XFILLER_25_271 VPWR VGND sg13g2_fill_1
XFILLER_25_293 VPWR VGND sg13g2_decap_4
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_41_731 VPWR VGND sg13g2_decap_8
XFILLER_41_742 VPWR VGND sg13g2_fill_1
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_4_13 VPWR VGND sg13g2_decap_4
XFILLER_4_164 VPWR VGND sg13g2_decap_8
XFILLER_5_610 VPWR VGND sg13g2_decap_8
XFILLER_5_621 VPWR VGND sg13g2_fill_2
XFILLER_5_643 VPWR VGND sg13g2_fill_1
XFILLER_5_676 VPWR VGND sg13g2_fill_1
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_16_282 VPWR VGND sg13g2_fill_2
XFILLER_32_720 VPWR VGND sg13g2_fill_1
XFILLER_36_525 VPWR VGND sg13g2_fill_2
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_31_263 VPWR VGND sg13g2_decap_8
X_1705_ VGND VPWR _0435_ _0436_ _0185_ _0437_ sg13g2_a21oi_1
X_1636_ state\[44\] daisychain\[44\] net144 _1026_ VPWR VGND sg13g2_mux2_1
X_1567_ _0971_ net162 _0970_ VPWR VGND sg13g2_nand2_1
XFILLER_39_352 VPWR VGND sg13g2_decap_8
X_1498_ VGND VPWR net93 daisychain\[15\] _0916_ net66 sg13g2_a21oi_1
X_2119_ VGND VPWR _0975_ _0749_ _0287_ net73 sg13g2_a21oi_1
XFILLER_22_263 VPWR VGND sg13g2_decap_4
XFILLER_35_591 VPWR VGND sg13g2_fill_2
Xfanout23 net25 net23 VPWR VGND sg13g2_buf_1
Xfanout34 net44 net34 VPWR VGND sg13g2_buf_1
Xfanout89 net90 net89 VPWR VGND sg13g2_buf_1
Xfanout78 net88 net78 VPWR VGND sg13g2_buf_1
Xfanout67 net68 net67 VPWR VGND sg13g2_buf_1
Xfanout56 net66 net56 VPWR VGND sg13g2_buf_1
Xfanout45 net66 net45 VPWR VGND sg13g2_buf_1
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_fill_1
XFILLER_6_407 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_fill_2
XFILLER_33_528 VPWR VGND sg13g2_fill_2
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_41_550 VPWR VGND sg13g2_decap_8
XFILLER_41_583 VPWR VGND sg13g2_decap_8
XFILLER_9_267 VPWR VGND sg13g2_decap_8
XFILLER_5_440 VPWR VGND sg13g2_decap_8
X_1421_ state\[1\] daisychain\[1\] net133 _0854_ VPWR VGND sg13g2_mux2_1
X_2470_ net207 VGND VPWR _0286_ state\[30\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
X_1352_ VPWR _0084_ state\[60\] VGND sg13g2_inv_1
XFILLER_20_723 VPWR VGND sg13g2_fill_1
XFILLER_20_756 VPWR VGND sg13g2_fill_1
XFILLER_20_789 VPWR VGND sg13g2_decap_4
Xclkload9 clknet_leaf_9_clk clkload9/Y VPWR VGND sg13g2_inv_4
X_1619_ net190 VPWR _1013_ VGND daisychain\[40\] net35 sg13g2_o21ai_1
XFILLER_15_517 VPWR VGND sg13g2_decap_8
XFILLER_27_355 VPWR VGND sg13g2_decap_8
XFILLER_27_388 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_43_815 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_10_244 VPWR VGND sg13g2_decap_8
XFILLER_11_701 VPWR VGND sg13g2_fill_1
XFILLER_24_76 VPWR VGND sg13g2_decap_8
XFILLER_30_509 VPWR VGND sg13g2_fill_2
XFILLER_6_204 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
X_2346__259 VPWR VGND net258 sg13g2_tiehi
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_18_355 VPWR VGND sg13g2_fill_1
XFILLER_45_196 VPWR VGND sg13g2_decap_8
X_1970_ VGND VPWR _0647_ _0648_ _0238_ _0649_ sg13g2_a21oi_1
XFILLER_6_782 VPWR VGND sg13g2_decap_4
X_2522_ net441 VGND VPWR _0338_ state\[82\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1335_ VPWR _0102_ state\[77\] VGND sg13g2_inv_1
X_1404_ VPWR _0116_ state\[8\] VGND sg13g2_inv_1
X_2453_ net275 VGND VPWR _0269_ state\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2384_ net438 VGND VPWR _0200_ daisychain\[72\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_24_303 VPWR VGND sg13g2_fill_1
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_37_664 VPWR VGND sg13g2_decap_4
XFILLER_49_480 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
XFILLER_24_358 VPWR VGND sg13g2_decap_8
XFILLER_10_23 VPWR VGND sg13g2_fill_1
XFILLER_10_34 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_15_303 VPWR VGND sg13g2_fill_2
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_31_807 VPWR VGND sg13g2_decap_8
XFILLER_31_818 VPWR VGND sg13g2_fill_2
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_43_678 VPWR VGND sg13g2_decap_8
X_2463__236 VPWR VGND net235 sg13g2_tiehi
XFILLER_2_273 VPWR VGND sg13g2_decap_8
XFILLER_3_763 VPWR VGND sg13g2_fill_1
X_2398__411 VPWR VGND net410 sg13g2_tiehi
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_38_439 VPWR VGND sg13g2_decap_4
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_21_306 VPWR VGND sg13g2_fill_1
XFILLER_33_144 VPWR VGND sg13g2_decap_8
X_1953_ VGND VPWR net107 daisychain\[106\] _0636_ net53 sg13g2_a21oi_1
X_1884_ net188 VPWR _0581_ VGND daisychain\[93\] net33 sg13g2_o21ai_1
X_2505_ net321 VGND VPWR _0321_ state\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1318_ VPWR _0121_ state\[94\] VGND sg13g2_inv_1
X_2436_ net334 VGND VPWR _0252_ daisychain\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2367_ net216 VGND VPWR _0183_ daisychain\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2298_ _0839_ net89 state\[121\] VPWR VGND sg13g2_nand2_1
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_33 VPWR VGND sg13g2_decap_4
XFILLER_24_188 VPWR VGND sg13g2_decap_8
XFILLER_4_505 VPWR VGND sg13g2_decap_8
XFILLER_21_66 VPWR VGND sg13g2_decap_8
XFILLER_15_100 VPWR VGND sg13g2_decap_8
XFILLER_28_483 VPWR VGND sg13g2_fill_1
XFILLER_28_494 VPWR VGND sg13g2_fill_2
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_48_748 VPWR VGND sg13g2_fill_2
XFILLER_15_177 VPWR VGND sg13g2_decap_8
XFILLER_30_158 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_8_811 VPWR VGND sg13g2_decap_8
XFILLER_8_822 VPWR VGND sg13g2_fill_1
XFILLER_7_13 VPWR VGND sg13g2_fill_2
XFILLER_7_354 VPWR VGND sg13g2_decap_8
XFILLER_7_79 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_39_737 VPWR VGND sg13g2_fill_2
X_2221_ VGND VPWR _0535_ _0800_ _0338_ net83 sg13g2_a21oi_1
X_2152_ _0766_ net118 state\[48\] VPWR VGND sg13g2_nand2_1
XFILLER_46_280 VPWR VGND sg13g2_decap_8
X_2083_ VGND VPWR _0903_ _0731_ _0269_ net67 sg13g2_a21oi_1
XFILLER_21_136 VPWR VGND sg13g2_decap_8
XFILLER_30_681 VPWR VGND sg13g2_fill_1
X_2563__422 VPWR VGND net421 sg13g2_tiehi
X_1936_ state\[104\] daisychain\[104\] net141 _0622_ VPWR VGND sg13g2_mux2_1
X_1867_ _0567_ net172 _0566_ VPWR VGND sg13g2_nand2_1
X_1798_ VGND VPWR net127 daisychain\[75\] _0512_ net63 sg13g2_a21oi_1
XFILLER_17_409 VPWR VGND sg13g2_fill_2
XFILLER_29_269 VPWR VGND sg13g2_fill_1
XFILLER_44_217 VPWR VGND sg13g2_decap_8
X_2419_ net368 VGND VPWR _0235_ daisychain\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_12_169 VPWR VGND sg13g2_decap_8
XFILLER_13_604 VPWR VGND sg13g2_fill_2
XFILLER_13_648 VPWR VGND sg13g2_fill_1
XFILLER_25_497 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_fill_2
XFILLER_40_445 VPWR VGND sg13g2_fill_2
XFILLER_40_478 VPWR VGND sg13g2_fill_1
XFILLER_20_180 VPWR VGND sg13g2_decap_8
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_fill_1
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_11_180 VPWR VGND sg13g2_decap_8
XFILLER_31_423 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
X_1721_ state\[61\] daisychain\[61\] net147 _0450_ VPWR VGND sg13g2_mux2_1
XFILLER_7_151 VPWR VGND sg13g2_decap_8
X_1652_ _0395_ net169 _0394_ VPWR VGND sg13g2_nand2_1
X_1583_ VGND VPWR net106 daisychain\[32\] _0984_ net52 sg13g2_a21oi_1
XFILLER_39_501 VPWR VGND sg13g2_fill_2
X_2204_ _0792_ net125 state\[74\] VPWR VGND sg13g2_nand2_1
X_2135_ VGND VPWR _1007_ _0757_ _0295_ net79 sg13g2_a21oi_1
XFILLER_19_291 VPWR VGND sg13g2_decap_4
XFILLER_22_434 VPWR VGND sg13g2_fill_2
XFILLER_26_239 VPWR VGND sg13g2_decap_8
XFILLER_34_294 VPWR VGND sg13g2_decap_8
X_2066_ _0723_ net101 state\[5\] VPWR VGND sg13g2_nand2_1
X_2528__394 VPWR VGND net393 sg13g2_tiehi
X_1919_ net187 VPWR _0609_ VGND daisychain\[100\] net32 sg13g2_o21ai_1
XFILLER_2_817 VPWR VGND sg13g2_decap_4
XFILLER_17_239 VPWR VGND sg13g2_decap_8
XFILLER_25_250 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
X_2494__368 VPWR VGND net367 sg13g2_tiehi
XFILLER_13_489 VPWR VGND sg13g2_fill_1
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_41_765 VPWR VGND sg13g2_fill_1
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_4_143 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_fill_1
XFILLER_5_699 VPWR VGND sg13g2_decap_4
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
X_2356__239 VPWR VGND net238 sg13g2_tiehi
XFILLER_16_261 VPWR VGND sg13g2_decap_8
XFILLER_17_740 VPWR VGND sg13g2_decap_8
XFILLER_17_762 VPWR VGND sg13g2_decap_4
XFILLER_31_242 VPWR VGND sg13g2_decap_8
X_1704_ net192 VPWR _0437_ VGND daisychain\[57\] net37 sg13g2_o21ai_1
X_1497_ _0915_ net159 _0914_ VPWR VGND sg13g2_nand2_1
X_1635_ VGND VPWR _1023_ _1024_ _0171_ _1025_ sg13g2_a21oi_1
X_1566_ state\[30\] daisychain\[30\] net138 _0970_ VPWR VGND sg13g2_mux2_1
XFILLER_39_331 VPWR VGND sg13g2_decap_8
XFILLER_42_518 VPWR VGND sg13g2_decap_8
X_2118_ _0749_ net106 state\[31\] VPWR VGND sg13g2_nand2_1
X_2049_ net178 VPWR _0713_ VGND daisychain\[126\] net26 sg13g2_o21ai_1
XFILLER_10_437 VPWR VGND sg13g2_fill_1
XFILLER_22_242 VPWR VGND sg13g2_decap_8
XFILLER_22_297 VPWR VGND sg13g2_decap_8
Xfanout24 net25 net24 VPWR VGND sg13g2_buf_1
Xfanout79 net87 net79 VPWR VGND sg13g2_buf_1
Xfanout68 net69 net68 VPWR VGND sg13g2_buf_1
Xfanout57 net58 net57 VPWR VGND sg13g2_buf_1
Xfanout46 net47 net46 VPWR VGND sg13g2_buf_1
Xfanout35 net43 net35 VPWR VGND sg13g2_buf_1
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_46_813 VPWR VGND sg13g2_decap_8
X_2459__252 VPWR VGND net251 sg13g2_tiehi
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_fill_1
XFILLER_33_507 VPWR VGND sg13g2_fill_1
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_9_246 VPWR VGND sg13g2_decap_8
X_1351_ VPWR _0085_ state\[61\] VGND sg13g2_inv_1
X_1420_ VGND VPWR _0849_ _0852_ _0128_ _0853_ sg13g2_a21oi_1
Xdigitalen.g\[1\].u.inv1 VPWR digitalen.g\[1\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_49_695 VPWR VGND sg13g2_decap_8
XFILLER_17_581 VPWR VGND sg13g2_decap_8
XFILLER_20_702 VPWR VGND sg13g2_fill_1
XFILLER_20_735 VPWR VGND sg13g2_fill_2
XFILLER_9_780 VPWR VGND sg13g2_fill_1
X_1618_ VGND VPWR net115 daisychain\[39\] _1012_ net57 sg13g2_a21oi_1
XFILLER_5_90 VPWR VGND sg13g2_decap_8
X_1549_ net182 VPWR _0957_ VGND daisychain\[26\] net27 sg13g2_o21ai_1
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_10_223 VPWR VGND sg13g2_decap_8
XFILLER_24_55 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_2_455 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_18_345 VPWR VGND sg13g2_fill_1
XFILLER_46_643 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_33_326 VPWR VGND sg13g2_fill_2
XFILLER_41_392 VPWR VGND sg13g2_decap_4
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_46_687 VPWR VGND sg13g2_decap_4
X_2521_ net449 VGND VPWR _0337_ state\[81\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2544__206 VPWR VGND net205 sg13g2_tiehi
XFILLER_28_109 VPWR VGND sg13g2_decap_8
XFILLER_5_293 VPWR VGND sg13g2_decap_8
X_1334_ VPWR _0103_ state\[78\] VGND sg13g2_inv_1
X_1403_ VPWR _0127_ state\[9\] VGND sg13g2_inv_1
X_2452_ net279 VGND VPWR _0268_ state\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2383_ net440 VGND VPWR _0199_ daisychain\[71\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_37_687 VPWR VGND sg13g2_fill_1
XFILLER_40_808 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_19_33 VPWR VGND sg13g2_fill_2
XFILLER_19_44 VPWR VGND sg13g2_fill_2
XFILLER_19_99 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_11_554 VPWR VGND sg13g2_decap_4
XFILLER_2_252 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_19_621 VPWR VGND sg13g2_decap_8
XFILLER_19_632 VPWR VGND sg13g2_fill_1
XFILLER_19_654 VPWR VGND sg13g2_decap_8
XFILLER_33_123 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
X_2470__208 VPWR VGND net207 sg13g2_tiehi
XFILLER_14_392 VPWR VGND sg13g2_fill_2
XFILLER_34_679 VPWR VGND sg13g2_decap_8
X_1952_ _0635_ net164 _0634_ VPWR VGND sg13g2_nand2_1
X_1883_ VGND VPWR net110 daisychain\[92\] _0580_ net55 sg13g2_a21oi_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_2504_ net327 VGND VPWR _0320_ state\[64\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2435_ net336 VGND VPWR _0251_ daisychain\[123\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
X_1317_ VPWR _0122_ state\[95\] VGND sg13g2_inv_1
X_2366_ net218 VGND VPWR _0182_ daisychain\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2297_ VGND VPWR _0687_ _0838_ _0376_ net70 sg13g2_a21oi_1
XFILLER_13_808 VPWR VGND sg13g2_decap_8
XFILLER_24_167 VPWR VGND sg13g2_decap_8
XFILLER_21_45 VPWR VGND sg13g2_decap_8
XFILLER_4_528 VPWR VGND sg13g2_fill_1
XFILLER_4_539 VPWR VGND sg13g2_fill_2
XFILLER_0_767 VPWR VGND sg13g2_fill_1
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_11_362 VPWR VGND sg13g2_decap_8
XFILLER_11_384 VPWR VGND sg13g2_decap_8
XFILLER_15_156 VPWR VGND sg13g2_decap_8
XFILLER_30_137 VPWR VGND sg13g2_decap_8
XFILLER_31_649 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_7_333 VPWR VGND sg13g2_decap_8
X_2510__282 VPWR VGND net281 sg13g2_tiehi
XFILLER_3_550 VPWR VGND sg13g2_fill_1
XFILLER_38_259 VPWR VGND sg13g2_decap_8
XFILLER_39_705 VPWR VGND sg13g2_decap_8
X_2220_ _0800_ net125 state\[82\] VPWR VGND sg13g2_nand2_1
X_2151_ VGND VPWR _0395_ _0765_ _0303_ net80 sg13g2_a21oi_1
X_2082_ _0731_ net91 state\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_21_115 VPWR VGND sg13g2_decap_8
X_2335__281 VPWR VGND net280 sg13g2_tiehi
XFILLER_30_660 VPWR VGND sg13g2_fill_1
XFILLER_30_693 VPWR VGND sg13g2_fill_1
X_2366__219 VPWR VGND net218 sg13g2_tiehi
X_1935_ VGND VPWR _0619_ _0620_ _0231_ _0621_ sg13g2_a21oi_1
X_1866_ state\[90\] daisychain\[90\] net149 _0566_ VPWR VGND sg13g2_mux2_1
X_1797_ _0511_ net174 _0510_ VPWR VGND sg13g2_nand2_1
X_2418_ net370 VGND VPWR _0234_ daisychain\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_16_34 VPWR VGND sg13g2_fill_2
XFILLER_29_248 VPWR VGND sg13g2_decap_8
XFILLER_38_771 VPWR VGND sg13g2_decap_8
X_2349_ net252 VGND VPWR _0165_ daisychain\[37\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_12_148 VPWR VGND sg13g2_decap_8
XFILLER_25_476 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_decap_8
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_16_421 VPWR VGND sg13g2_fill_1
XFILLER_31_402 VPWR VGND sg13g2_fill_1
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_44_785 VPWR VGND sg13g2_fill_1
XFILLER_7_130 VPWR VGND sg13g2_decap_8
XFILLER_8_642 VPWR VGND sg13g2_fill_2
XFILLER_8_653 VPWR VGND sg13g2_decap_8
X_1720_ VGND VPWR _0447_ _0448_ _0188_ _0449_ sg13g2_a21oi_1
X_1651_ state\[47\] daisychain\[47\] net145 _0394_ VPWR VGND sg13g2_mux2_1
X_1582_ _0983_ net162 _0982_ VPWR VGND sg13g2_nand2_1
XFILLER_26_218 VPWR VGND sg13g2_decap_8
XFILLER_35_741 VPWR VGND sg13g2_fill_2
X_2203_ VGND VPWR _0499_ _0791_ _0329_ net85 sg13g2_a21oi_1
X_2134_ _0757_ net115 state\[39\] VPWR VGND sg13g2_nand2_1
X_2065_ VGND VPWR _0867_ _0722_ _0260_ net75 sg13g2_a21oi_1
XFILLER_22_479 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
X_2452__280 VPWR VGND net279 sg13g2_tiehi
X_1918_ VGND VPWR net109 daisychain\[99\] _0608_ net54 sg13g2_a21oi_1
X_1849_ net197 VPWR _0553_ VGND daisychain\[86\] net42 sg13g2_o21ai_1
XFILLER_17_218 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_9_439 VPWR VGND sg13g2_decap_4
XFILLER_4_122 VPWR VGND sg13g2_decap_8
XFILLER_4_199 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_decap_8
XFILLER_5_667 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_36_516 VPWR VGND sg13g2_decap_4
XFILLER_36_527 VPWR VGND sg13g2_fill_1
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_16_240 VPWR VGND sg13g2_decap_8
XFILLER_31_221 VPWR VGND sg13g2_decap_8
XFILLER_32_777 VPWR VGND sg13g2_fill_1
XFILLER_32_788 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_1703_ VGND VPWR net121 daisychain\[56\] _0436_ net59 sg13g2_a21oi_1
X_1634_ net190 VPWR _1025_ VGND daisychain\[43\] net35 sg13g2_o21ai_1
XFILLER_39_310 VPWR VGND sg13g2_decap_8
X_1496_ state\[16\] daisychain\[16\] net137 _0914_ VPWR VGND sg13g2_mux2_1
X_1565_ VGND VPWR _0967_ _0968_ _0157_ _0969_ sg13g2_a21oi_1
XFILLER_35_582 VPWR VGND sg13g2_fill_1
XFILLER_39_387 VPWR VGND sg13g2_decap_8
X_2117_ VGND VPWR _0971_ _0748_ _0286_ net74 sg13g2_a21oi_1
X_2048_ VGND VPWR net90 daisychain\[125\] _0712_ net48 sg13g2_a21oi_1
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_22_221 VPWR VGND sg13g2_decap_8
Xfanout25 net44 net25 VPWR VGND sg13g2_buf_1
Xfanout69 net88 net69 VPWR VGND sg13g2_buf_1
Xfanout58 net65 net58 VPWR VGND sg13g2_buf_1
Xfanout47 net48 net47 VPWR VGND sg13g2_buf_1
Xfanout36 net43 net36 VPWR VGND sg13g2_buf_1
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_2_604 VPWR VGND sg13g2_decap_8
XFILLER_2_637 VPWR VGND sg13g2_fill_1
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_46_803 VPWR VGND sg13g2_fill_2
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_9_225 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[1\].u.inv2 VPWR digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN VGND
+ sg13g2_inv_1
X_2466__224 VPWR VGND net223 sg13g2_tiehi
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_49_652 VPWR VGND sg13g2_decap_8
X_1350_ VPWR _0086_ state\[62\] VGND sg13g2_inv_1
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_49_663 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_0_clk clknet_2_1__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_20_769 VPWR VGND sg13g2_fill_1
X_2445__308 VPWR VGND net307 sg13g2_tiehi
XFILLER_8_291 VPWR VGND sg13g2_decap_8
X_1617_ _1011_ net168 _1010_ VPWR VGND sg13g2_nand2_1
XFILLER_39_184 VPWR VGND sg13g2_decap_8
X_1479_ net179 VPWR _0901_ VGND daisychain\[12\] net23 sg13g2_o21ai_1
X_1548_ VGND VPWR net99 daisychain\[25\] _0956_ net49 sg13g2_a21oi_1
XFILLER_23_530 VPWR VGND sg13g2_fill_1
XFILLER_24_34 VPWR VGND sg13g2_decap_8
XFILLER_27_379 VPWR VGND sg13g2_fill_1
XFILLER_10_202 VPWR VGND sg13g2_decap_8
XFILLER_10_279 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_6_239 VPWR VGND sg13g2_decap_8
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_2_478 VPWR VGND sg13g2_fill_2
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_18_302 VPWR VGND sg13g2_decap_4
XFILLER_19_803 VPWR VGND sg13g2_decap_8
XFILLER_19_814 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_46_600 VPWR VGND sg13g2_decap_8
XFILLER_46_655 VPWR VGND sg13g2_fill_2
XFILLER_46_666 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_decap_8
XFILLER_5_272 VPWR VGND sg13g2_decap_8
XFILLER_6_740 VPWR VGND sg13g2_fill_1
X_1402_ VPWR _0011_ state\[10\] VGND sg13g2_inv_1
X_2520_ net201 VGND VPWR _0336_ state\[80\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2548__398 VPWR VGND net397 sg13g2_tiehi
X_2451_ net283 VGND VPWR _0267_ state\[11\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1333_ VPWR _0104_ state\[79\] VGND sg13g2_inv_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_2382_ net442 VGND VPWR _0198_ daisychain\[70\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_24_338 VPWR VGND sg13g2_fill_2
XFILLER_32_360 VPWR VGND sg13g2_fill_1
XFILLER_36_154 VPWR VGND sg13g2_decap_8
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_20_577 VPWR VGND sg13g2_decap_8
XFILLER_20_588 VPWR VGND sg13g2_fill_2
XFILLER_10_69 VPWR VGND sg13g2_decap_8
X_2345__261 VPWR VGND net260 sg13g2_tiehi
XFILLER_15_305 VPWR VGND sg13g2_fill_1
XFILLER_19_78 VPWR VGND sg13g2_decap_8
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_43_636 VPWR VGND sg13g2_decap_8
XFILLER_43_647 VPWR VGND sg13g2_fill_1
XFILLER_2_231 VPWR VGND sg13g2_decap_8
XFILLER_3_721 VPWR VGND sg13g2_decap_8
XFILLER_18_8 VPWR VGND sg13g2_fill_1
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_19_677 VPWR VGND sg13g2_decap_8
XFILLER_33_102 VPWR VGND sg13g2_decap_8
XFILLER_33_179 VPWR VGND sg13g2_decap_8
XFILLER_34_625 VPWR VGND sg13g2_fill_2
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_14_371 VPWR VGND sg13g2_decap_8
X_1951_ state\[107\] daisychain\[107\] net141 _0634_ VPWR VGND sg13g2_mux2_1
X_1882_ _0579_ net165 _0578_ VPWR VGND sg13g2_nand2_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_6_581 VPWR VGND sg13g2_decap_4
X_2503_ net331 VGND VPWR _0319_ state\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2434_ net338 VGND VPWR _0250_ daisychain\[122\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2365_ net220 VGND VPWR _0181_ daisychain\[53\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XFILLER_37_485 VPWR VGND sg13g2_decap_8
X_1316_ VPWR _0123_ state\[96\] VGND sg13g2_inv_1
X_2296_ _0838_ net98 state\[120\] VPWR VGND sg13g2_nand2_1
XFILLER_24_113 VPWR VGND sg13g2_fill_1
XFILLER_24_146 VPWR VGND sg13g2_decap_8
XFILLER_33_680 VPWR VGND sg13g2_fill_2
XFILLER_20_374 VPWR VGND sg13g2_fill_2
X_2497__356 VPWR VGND net355 sg13g2_tiehi
XFILLER_15_135 VPWR VGND sg13g2_decap_8
XFILLER_16_647 VPWR VGND sg13g2_fill_1
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_11_341 VPWR VGND sg13g2_decap_8
XFILLER_30_116 VPWR VGND sg13g2_decap_8
XFILLER_7_15 VPWR VGND sg13g2_fill_1
XFILLER_7_26 VPWR VGND sg13g2_decap_8
XFILLER_7_312 VPWR VGND sg13g2_decap_8
XFILLER_3_562 VPWR VGND sg13g2_fill_2
XFILLER_7_389 VPWR VGND sg13g2_decap_8
XFILLER_19_452 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
XFILLER_39_739 VPWR VGND sg13g2_fill_1
XFILLER_47_772 VPWR VGND sg13g2_fill_2
X_2150_ _0765_ net117 state\[47\] VPWR VGND sg13g2_nand2_1
X_2081_ VGND VPWR _0899_ _0730_ _0268_ net68 sg13g2_a21oi_1
X_1934_ net188 VPWR _0621_ VGND daisychain\[103\] net33 sg13g2_o21ai_1
XFILLER_30_672 VPWR VGND sg13g2_fill_1
X_1865_ VGND VPWR _0563_ _0564_ _0217_ _0565_ sg13g2_a21oi_1
X_1796_ state\[76\] daisychain\[76\] net150 _0510_ VPWR VGND sg13g2_mux2_1
XFILLER_29_227 VPWR VGND sg13g2_decap_8
X_2417_ net372 VGND VPWR _0233_ daisychain\[105\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2348_ net254 VGND VPWR _0164_ daisychain\[36\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_13_606 VPWR VGND sg13g2_fill_1
XFILLER_38_750 VPWR VGND sg13g2_decap_8
XFILLER_38_794 VPWR VGND sg13g2_fill_2
X_2279_ VGND VPWR _0651_ _0829_ _0367_ net76 sg13g2_a21oi_1
XFILLER_12_127 VPWR VGND sg13g2_decap_8
XFILLER_16_79 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_4_304 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_44_731 VPWR VGND sg13g2_fill_2
X_2551__350 VPWR VGND net349 sg13g2_tiehi
XFILLER_7_186 VPWR VGND sg13g2_decap_8
XFILLER_8_621 VPWR VGND sg13g2_decap_8
XFILLER_8_632 VPWR VGND sg13g2_fill_1
XFILLER_8_676 VPWR VGND sg13g2_fill_2
X_1650_ VGND VPWR _0391_ _0392_ _0174_ _0393_ sg13g2_a21oi_1
X_1581_ state\[33\] daisychain\[33\] net140 _0982_ VPWR VGND sg13g2_mux2_1
XFILLER_3_392 VPWR VGND sg13g2_decap_8
X_2202_ _0791_ net129 state\[73\] VPWR VGND sg13g2_nand2_1
XFILLER_34_252 VPWR VGND sg13g2_decap_8
X_2133_ VGND VPWR _1003_ _0756_ _0294_ net72 sg13g2_a21oi_1
X_2064_ _0722_ net107 state\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_22_458 VPWR VGND sg13g2_decap_8
X_1917_ _0607_ net166 _0606_ VPWR VGND sg13g2_nand2_1
XFILLER_1_329 VPWR VGND sg13g2_decap_8
X_1848_ VGND VPWR net124 daisychain\[85\] _0552_ net61 sg13g2_a21oi_1
X_1779_ net195 VPWR _0497_ VGND daisychain\[72\] net40 sg13g2_o21ai_1
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_41_701 VPWR VGND sg13g2_decap_8
XFILLER_41_756 VPWR VGND sg13g2_decap_8
XFILLER_9_407 VPWR VGND sg13g2_decap_4
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_4_101 VPWR VGND sg13g2_decap_8
XFILLER_5_657 VPWR VGND sg13g2_decap_4
X_2546__430 VPWR VGND net429 sg13g2_tiehi
XFILLER_4_178 VPWR VGND sg13g2_decap_8
X_2403__401 VPWR VGND net400 sg13g2_tiehi
XFILLER_36_539 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_31_200 VPWR VGND sg13g2_decap_8
XFILLER_31_277 VPWR VGND sg13g2_decap_8
XFILLER_44_561 VPWR VGND sg13g2_fill_1
XFILLER_8_473 VPWR VGND sg13g2_decap_8
X_1702_ _0435_ net170 _0434_ VPWR VGND sg13g2_nand2_1
X_1633_ VGND VPWR net116 daisychain\[42\] _1024_ net57 sg13g2_a21oi_1
X_1564_ net185 VPWR _0969_ VGND daisychain\[29\] net30 sg13g2_o21ai_1
XFILLER_39_366 VPWR VGND sg13g2_decap_8
X_1495_ VGND VPWR _0911_ _0912_ _0143_ _0913_ sg13g2_a21oi_1
XFILLER_22_200 VPWR VGND sg13g2_decap_8
XFILLER_27_528 VPWR VGND sg13g2_fill_2
XFILLER_35_561 VPWR VGND sg13g2_decap_8
XFILLER_35_572 VPWR VGND sg13g2_fill_1
Xfanout26 net44 net26 VPWR VGND sg13g2_buf_1
Xfanout37 net38 net37 VPWR VGND sg13g2_buf_1
X_2116_ _0748_ net102 state\[30\] VPWR VGND sg13g2_nand2_1
X_2047_ _0711_ net154 _0710_ VPWR VGND sg13g2_nand2_1
XFILLER_10_428 VPWR VGND sg13g2_decap_8
Xfanout59 net60 net59 VPWR VGND sg13g2_buf_1
Xfanout48 net66 net48 VPWR VGND sg13g2_buf_1
X_2385__437 VPWR VGND net436 sg13g2_tiehi
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_2_649 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
X_2355__241 VPWR VGND net240 sg13g2_tiehi
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_14_734 VPWR VGND sg13g2_decap_4
XFILLER_9_204 VPWR VGND sg13g2_decap_8
XFILLER_17_561 VPWR VGND sg13g2_decap_8
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_20_715 VPWR VGND sg13g2_fill_1
XFILLER_20_748 VPWR VGND sg13g2_fill_1
XFILLER_32_564 VPWR VGND sg13g2_fill_2
XFILLER_8_270 VPWR VGND sg13g2_decap_8
X_1547_ _0955_ net159 _0954_ VPWR VGND sg13g2_nand2_1
X_1616_ state\[40\] daisychain\[40\] net144 _1010_ VPWR VGND sg13g2_mux2_1
XFILLER_27_325 VPWR VGND sg13g2_decap_4
XFILLER_27_369 VPWR VGND sg13g2_decap_4
XFILLER_39_163 VPWR VGND sg13g2_decap_8
X_1478_ VGND VPWR net93 daisychain\[11\] _0900_ net45 sg13g2_a21oi_1
XFILLER_24_13 VPWR VGND sg13g2_decap_8
XFILLER_10_258 VPWR VGND sg13g2_decap_8
XFILLER_2_413 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_6_218 VPWR VGND sg13g2_decap_8
XFILLER_7_719 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_33_328 VPWR VGND sg13g2_fill_1
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_10_770 VPWR VGND sg13g2_decap_8
XFILLER_14_564 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_5_251 VPWR VGND sg13g2_decap_8
X_1401_ VPWR _0022_ state\[11\] VGND sg13g2_inv_1
X_2450_ net287 VGND VPWR _0266_ state\[10\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2381_ net444 VGND VPWR _0197_ daisychain\[69\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_49_494 VPWR VGND sg13g2_decap_8
X_1332_ VPWR _0106_ state\[80\] VGND sg13g2_inv_1
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_20_501 VPWR VGND sg13g2_decap_4
XFILLER_32_372 VPWR VGND sg13g2_fill_2
XFILLER_37_678 VPWR VGND sg13g2_decap_8
X_2531__370 VPWR VGND net369 sg13g2_tiehi
X_2490__384 VPWR VGND net383 sg13g2_tiehi
XFILLER_20_556 VPWR VGND sg13g2_decap_8
XFILLER_32_394 VPWR VGND sg13g2_decap_8
XFILLER_10_48 VPWR VGND sg13g2_decap_8
XFILLER_19_35 VPWR VGND sg13g2_fill_1
XFILLER_15_339 VPWR VGND sg13g2_fill_2
XFILLER_16_807 VPWR VGND sg13g2_decap_8
XFILLER_19_57 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_30_309 VPWR VGND sg13g2_fill_2
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_7_516 VPWR VGND sg13g2_decap_8
XFILLER_2_210 VPWR VGND sg13g2_decap_8
XFILLER_3_700 VPWR VGND sg13g2_decap_4
XFILLER_2_287 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_30_810 VPWR VGND sg13g2_fill_1
XFILLER_30_821 VPWR VGND sg13g2_fill_2
XFILLER_33_158 VPWR VGND sg13g2_decap_8
XFILLER_34_659 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
X_1950_ VGND VPWR _0631_ _0632_ _0234_ _0633_ sg13g2_a21oi_1
X_2502_ net335 VGND VPWR _0318_ state\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2411__385 VPWR VGND net384 sg13g2_tiehi
X_1881_ state\[93\] daisychain\[93\] net142 _0578_ VPWR VGND sg13g2_mux2_1
X_1315_ VPWR _0124_ state\[97\] VGND sg13g2_inv_1
X_2433_ net340 VGND VPWR _0249_ daisychain\[121\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2364_ net222 VGND VPWR _0180_ daisychain\[52\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_24_125 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
X_2295_ VGND VPWR _0683_ _0837_ _0375_ net69 sg13g2_a21oi_1
XFILLER_12_309 VPWR VGND sg13g2_decap_8
XFILLER_20_386 VPWR VGND sg13g2_fill_2
XFILLER_4_519 VPWR VGND sg13g2_fill_2
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_15_114 VPWR VGND sg13g2_decap_8
XFILLER_16_626 VPWR VGND sg13g2_fill_2
XFILLER_16_637 VPWR VGND sg13g2_fill_1
XFILLER_16_659 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_11_320 VPWR VGND sg13g2_decap_8
XFILLER_7_368 VPWR VGND sg13g2_decap_8
XFILLER_30_8 VPWR VGND sg13g2_fill_2
XFILLER_3_541 VPWR VGND sg13g2_decap_8
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
X_2080_ _0730_ net91 state\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_30_651 VPWR VGND sg13g2_fill_2
XFILLER_34_489 VPWR VGND sg13g2_decap_8
X_1933_ VGND VPWR net107 daisychain\[102\] _0620_ net55 sg13g2_a21oi_1
X_1864_ net197 VPWR _0565_ VGND daisychain\[89\] net42 sg13g2_o21ai_1
X_1795_ VGND VPWR _0507_ _0508_ _0203_ _0509_ sg13g2_a21oi_1
XFILLER_29_206 VPWR VGND sg13g2_decap_8
X_2416_ net374 VGND VPWR _0232_ daisychain\[104\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2347_ net256 VGND VPWR _0163_ daisychain\[35\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2278_ _0829_ net114 state\[111\] VPWR VGND sg13g2_nand2_1
XFILLER_12_106 VPWR VGND sg13g2_decap_8
XFILLER_16_36 VPWR VGND sg13g2_fill_1
XFILLER_16_58 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
X_2314__323 VPWR VGND net322 sg13g2_tiehi
XFILLER_20_194 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_5_806 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_16_412 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
X_2395__417 VPWR VGND net416 sg13g2_tiehi
XFILLER_16_456 VPWR VGND sg13g2_fill_1
XFILLER_28_294 VPWR VGND sg13g2_fill_2
XFILLER_43_231 VPWR VGND sg13g2_decap_8
X_2469__212 VPWR VGND net211 sg13g2_tiehi
XFILLER_11_194 VPWR VGND sg13g2_decap_8
XFILLER_7_165 VPWR VGND sg13g2_decap_8
X_2365__221 VPWR VGND net220 sg13g2_tiehi
X_1580_ VGND VPWR _0979_ _0980_ _0160_ _0981_ sg13g2_a21oi_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_3_371 VPWR VGND sg13g2_decap_8
X_2201_ VGND VPWR _0495_ _0790_ _0328_ net85 sg13g2_a21oi_1
X_2132_ _0756_ net105 state\[38\] VPWR VGND sg13g2_nand2_1
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_35_754 VPWR VGND sg13g2_decap_8
XFILLER_47_570 VPWR VGND sg13g2_decap_4
X_2063_ VGND VPWR _0863_ _0721_ _0259_ net67 sg13g2_a21oi_1
XFILLER_8_81 VPWR VGND sg13g2_decap_8
X_1916_ state\[100\] daisychain\[100\] net143 _0606_ VPWR VGND sg13g2_mux2_1
X_1847_ _0551_ net172 _0550_ VPWR VGND sg13g2_nand2_1
XFILLER_1_308 VPWR VGND sg13g2_decap_8
X_1778_ VGND VPWR net127 daisychain\[71\] _0496_ net63 sg13g2_a21oi_1
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_13_404 VPWR VGND sg13g2_decap_8
XFILLER_13_415 VPWR VGND sg13g2_fill_1
XFILLER_25_264 VPWR VGND sg13g2_decap_8
XFILLER_25_286 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_4_157 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_4_17 VPWR VGND sg13g2_fill_1
XFILLER_16_275 VPWR VGND sg13g2_decap_8
XFILLER_36_507 VPWR VGND sg13g2_decap_4
XFILLER_44_573 VPWR VGND sg13g2_decap_4
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_31_256 VPWR VGND sg13g2_decap_8
XFILLER_8_430 VPWR VGND sg13g2_fill_2
X_1701_ state\[57\] daisychain\[57\] net146 _0434_ VPWR VGND sg13g2_mux2_1
X_1494_ net181 VPWR _0913_ VGND daisychain\[15\] net25 sg13g2_o21ai_1
X_1632_ _1023_ net168 _1022_ VPWR VGND sg13g2_nand2_1
X_1563_ VGND VPWR net101 daisychain\[28\] _0968_ net50 sg13g2_a21oi_1
XFILLER_39_345 VPWR VGND sg13g2_decap_8
X_2115_ VGND VPWR _0967_ _0747_ _0285_ net74 sg13g2_a21oi_1
XFILLER_22_256 VPWR VGND sg13g2_decap_8
XFILLER_22_267 VPWR VGND sg13g2_fill_2
Xfanout27 net30 net27 VPWR VGND sg13g2_buf_1
Xfanout49 net52 net49 VPWR VGND sg13g2_buf_1
Xfanout38 net43 net38 VPWR VGND sg13g2_buf_1
X_2046_ state\[126\] daisychain\[126\] net136 _0710_ VPWR VGND sg13g2_mux2_1
XFILLER_13_37 VPWR VGND sg13g2_decap_4
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_5_433 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_1_694 VPWR VGND sg13g2_fill_1
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_17_595 VPWR VGND sg13g2_fill_2
XFILLER_44_392 VPWR VGND sg13g2_decap_8
XFILLER_20_727 VPWR VGND sg13g2_fill_1
X_1477_ _0899_ net155 _0898_ VPWR VGND sg13g2_nand2_1
X_1546_ state\[26\] daisychain\[26\] net137 _0954_ VPWR VGND sg13g2_mux2_1
X_2421__365 VPWR VGND net364 sg13g2_tiehi
X_1615_ VGND VPWR _1007_ _1008_ _0167_ _1009_ sg13g2_a21oi_1
XFILLER_39_142 VPWR VGND sg13g2_decap_8
XFILLER_43_808 VPWR VGND sg13g2_decap_8
XFILLER_10_237 VPWR VGND sg13g2_decap_8
XFILLER_24_69 VPWR VGND sg13g2_decap_8
XFILLER_35_381 VPWR VGND sg13g2_fill_2
XFILLER_42_329 VPWR VGND sg13g2_decap_8
X_2029_ net178 VPWR _0697_ VGND daisychain\[122\] net26 sg13g2_o21ai_1
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_2_469 VPWR VGND sg13g2_decap_4
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_14_521 VPWR VGND sg13g2_decap_4
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_14_91 VPWR VGND sg13g2_decap_8
XFILLER_5_230 VPWR VGND sg13g2_decap_8
XFILLER_6_720 VPWR VGND sg13g2_decap_4
X_1331_ VPWR _0107_ state\[81\] VGND sg13g2_inv_1
X_1400_ VPWR _0031_ state\[12\] VGND sg13g2_inv_1
Xwires dac/IOUT dac/VcascP[1] dac/VcascP[0] i_in i_out analog_wires
X_2479__428 VPWR VGND net427 sg13g2_tiehi
X_2380_ net446 VGND VPWR _0196_ daisychain\[68\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_37_657 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_32_351 VPWR VGND sg13g2_decap_4
XFILLER_36_189 VPWR VGND sg13g2_decap_8
X_1529_ net183 VPWR _0941_ VGND daisychain\[22\] net28 sg13g2_o21ai_1
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_11_524 VPWR VGND sg13g2_fill_1
XFILLER_2_266 VPWR VGND sg13g2_decap_8
X_2324__303 VPWR VGND net302 sg13g2_tiehi
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_19_668 VPWR VGND sg13g2_decap_4
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_33_137 VPWR VGND sg13g2_decap_8
XFILLER_34_627 VPWR VGND sg13g2_fill_1
X_1880_ VGND VPWR _0575_ _0576_ _0220_ _0577_ sg13g2_a21oi_1
XFILLER_10_590 VPWR VGND sg13g2_decap_8
X_2501_ net339 VGND VPWR _0317_ state\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1314_ VPWR _0125_ state\[98\] VGND sg13g2_inv_1
X_2432_ net342 VGND VPWR _0248_ daisychain\[120\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2375__201 VPWR VGND net200 sg13g2_tiehi
X_2363_ net224 VGND VPWR _0179_ daisychain\[51\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2294_ _0837_ net97 state\[119\] VPWR VGND sg13g2_nand2_1
XFILLER_37_432 VPWR VGND sg13g2_decap_8
XFILLER_37_476 VPWR VGND sg13g2_decap_4
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_20_376 VPWR VGND sg13g2_fill_1
XFILLER_33_682 VPWR VGND sg13g2_fill_1
XFILLER_21_59 VPWR VGND sg13g2_decap_8
X_2462__240 VPWR VGND net239 sg13g2_tiehi
XFILLER_28_454 VPWR VGND sg13g2_fill_2
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_11_376 VPWR VGND sg13g2_fill_2
XFILLER_3_520 VPWR VGND sg13g2_decap_8
XFILLER_7_347 VPWR VGND sg13g2_decap_8
XFILLER_3_564 VPWR VGND sg13g2_fill_1
XFILLER_3_597 VPWR VGND sg13g2_decap_8
X_2441__324 VPWR VGND net323 sg13g2_tiehi
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_47_774 VPWR VGND sg13g2_fill_1
XFILLER_47_785 VPWR VGND sg13g2_fill_1
XFILLER_21_129 VPWR VGND sg13g2_decap_8
XFILLER_30_685 VPWR VGND sg13g2_fill_1
X_1932_ _0619_ net165 _0618_ VPWR VGND sg13g2_nand2_1
X_1863_ VGND VPWR net111 daisychain\[88\] _0564_ net61 sg13g2_a21oi_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_2415_ net376 VGND VPWR _0231_ daisychain\[103\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1794_ net195 VPWR _0509_ VGND daisychain\[75\] net40 sg13g2_o21ai_1
X_2346_ net258 VGND VPWR _0162_ daisychain\[34\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2277_ VGND VPWR _0647_ _0828_ _0366_ net76 sg13g2_a21oi_1
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_20_173 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_28_251 VPWR VGND sg13g2_fill_1
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_44_733 VPWR VGND sg13g2_fill_1
XFILLER_11_173 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_3_350 VPWR VGND sg13g2_decap_8
XFILLER_7_144 VPWR VGND sg13g2_decap_8
X_2200_ _0790_ net129 state\[72\] VPWR VGND sg13g2_nand2_1
X_2131_ VGND VPWR _0999_ _0755_ _0293_ net72 sg13g2_a21oi_1
X_2062_ _0721_ net92 state\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_2_0__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_1915_ VGND VPWR _0603_ _0604_ _0227_ _0605_ sg13g2_a21oi_1
X_1846_ state\[86\] daisychain\[86\] net149 _0550_ VPWR VGND sg13g2_mux2_1
X_1777_ _0495_ net174 _0494_ VPWR VGND sg13g2_nand2_1
XFILLER_27_14 VPWR VGND sg13g2_decap_8
X_2329_ net292 VGND VPWR _0145_ daisychain\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_21_482 VPWR VGND sg13g2_decap_8
XFILLER_25_243 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
X_2431__345 VPWR VGND net344 sg13g2_tiehi
XFILLER_4_136 VPWR VGND sg13g2_decap_8
XFILLER_5_604 VPWR VGND sg13g2_fill_1
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_16_254 VPWR VGND sg13g2_decap_8
XFILLER_17_733 VPWR VGND sg13g2_decap_8
XFILLER_17_755 VPWR VGND sg13g2_decap_8
XFILLER_17_766 VPWR VGND sg13g2_fill_1
XFILLER_31_235 VPWR VGND sg13g2_decap_8
X_2332__287 VPWR VGND net286 sg13g2_tiehi
X_1700_ VGND VPWR _0431_ _0432_ _0184_ _0433_ sg13g2_a21oi_1
X_1631_ state\[43\] daisychain\[43\] net144 _1022_ VPWR VGND sg13g2_mux2_1
XFILLER_4_692 VPWR VGND sg13g2_decap_8
X_1493_ VGND VPWR net92 daisychain\[14\] _0912_ net45 sg13g2_a21oi_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_1562_ _0967_ net160 _0966_ VPWR VGND sg13g2_nand2_1
XFILLER_39_324 VPWR VGND sg13g2_decap_8
X_2493__372 VPWR VGND net371 sg13g2_tiehi
X_2114_ _0747_ net102 state\[29\] VPWR VGND sg13g2_nand2_1
X_2045_ VGND VPWR _0707_ _0708_ _0253_ _0709_ sg13g2_a21oi_1
XFILLER_22_235 VPWR VGND sg13g2_decap_8
Xfanout28 net29 net28 VPWR VGND sg13g2_buf_1
Xfanout39 net42 net39 VPWR VGND sg13g2_buf_1
X_1829_ net194 VPWR _0537_ VGND daisychain\[82\] net39 sg13g2_o21ai_1
XFILLER_18_508 VPWR VGND sg13g2_fill_2
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_5_412 VPWR VGND sg13g2_decap_8
XFILLER_9_239 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_49_622 VPWR VGND sg13g2_decap_8
XFILLER_17_574 VPWR VGND sg13g2_decap_8
XFILLER_20_706 VPWR VGND sg13g2_fill_1
XFILLER_32_500 VPWR VGND sg13g2_fill_1
XFILLER_44_371 VPWR VGND sg13g2_decap_8
X_1614_ net190 VPWR _1009_ VGND daisychain\[39\] net35 sg13g2_o21ai_1
XFILLER_39_121 VPWR VGND sg13g2_decap_8
XFILLER_5_50 VPWR VGND sg13g2_fill_1
XFILLER_5_83 VPWR VGND sg13g2_decap_8
X_1476_ state\[12\] daisychain\[12\] net133 _0898_ VPWR VGND sg13g2_mux2_1
X_1545_ VGND VPWR _0951_ _0952_ _0153_ _0953_ sg13g2_a21oi_1
XFILLER_23_500 VPWR VGND sg13g2_fill_2
XFILLER_27_349 VPWR VGND sg13g2_fill_2
XFILLER_39_198 VPWR VGND sg13g2_decap_8
XFILLER_42_308 VPWR VGND sg13g2_decap_8
X_2028_ VGND VPWR net89 daisychain\[121\] _0696_ net48 sg13g2_a21oi_1
XFILLER_10_216 VPWR VGND sg13g2_decap_8
XFILLER_24_48 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_2_448 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_33_319 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_14_70 VPWR VGND sg13g2_decap_8
XFILLER_41_396 VPWR VGND sg13g2_fill_1
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_5_286 VPWR VGND sg13g2_decap_8
X_1330_ VPWR _0108_ state\[82\] VGND sg13g2_inv_1
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_32_374 VPWR VGND sg13g2_fill_1
XFILLER_9_570 VPWR VGND sg13g2_decap_8
X_1459_ net179 VPWR _0885_ VGND daisychain\[8\] net23 sg13g2_o21ai_1
X_1528_ VGND VPWR net104 daisychain\[21\] _0940_ net51 sg13g2_a21oi_1
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_11_547 VPWR VGND sg13g2_decap_8
XFILLER_3_713 VPWR VGND sg13g2_fill_2
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_decap_8
XFILLER_19_603 VPWR VGND sg13g2_fill_2
XFILLER_19_614 VPWR VGND sg13g2_decap_8
XFILLER_33_116 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_14_385 VPWR VGND sg13g2_decap_8
XFILLER_26_190 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
X_2500_ net343 VGND VPWR _0316_ state\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2431_ net344 VGND VPWR _0247_ daisychain\[119\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_1313_ VPWR _0126_ state\[99\] VGND sg13g2_inv_1
X_2362_ net226 VGND VPWR _0178_ daisychain\[50\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2293_ VGND VPWR _0679_ _0836_ _0374_ net69 sg13g2_a21oi_1
XFILLER_17_190 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_decap_4
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_0_716 VPWR VGND sg13g2_fill_2
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_11_355 VPWR VGND sg13g2_decap_8
XFILLER_15_149 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_31_609 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_decap_8
XFILLER_7_326 VPWR VGND sg13g2_decap_8
XFILLER_21_108 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_14_182 VPWR VGND sg13g2_decap_8
XFILLER_30_664 VPWR VGND sg13g2_fill_1
XFILLER_30_697 VPWR VGND sg13g2_fill_2
X_1931_ state\[103\] daisychain\[103\] net141 _0618_ VPWR VGND sg13g2_mux2_1
X_1862_ _0563_ net172 _0562_ VPWR VGND sg13g2_nand2_1
X_1793_ VGND VPWR net129 daisychain\[74\] _0508_ net63 sg13g2_a21oi_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
X_2414_ net378 VGND VPWR _0230_ daisychain\[102\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2342__267 VPWR VGND net266 sg13g2_tiehi
XFILLER_37_252 VPWR VGND sg13g2_decap_8
XFILLER_38_764 VPWR VGND sg13g2_decap_8
X_2345_ net260 VGND VPWR _0161_ daisychain\[33\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2276_ _0828_ net114 state\[110\] VPWR VGND sg13g2_nand2_1
XFILLER_25_469 VPWR VGND sg13g2_decap_8
XFILLER_20_152 VPWR VGND sg13g2_decap_8
XFILLER_4_318 VPWR VGND sg13g2_decap_8
X_2505__322 VPWR VGND net321 sg13g2_tiehi
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_44_701 VPWR VGND sg13g2_decap_8
XFILLER_44_778 VPWR VGND sg13g2_decap_8
XFILLER_11_152 VPWR VGND sg13g2_decap_8
XFILLER_12_631 VPWR VGND sg13g2_decap_8
XFILLER_7_123 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_35_701 VPWR VGND sg13g2_decap_8
X_2517__226 VPWR VGND net225 sg13g2_tiehi
X_2130_ _0755_ net105 state\[37\] VPWR VGND sg13g2_nand2_1
X_2061_ VGND VPWR _0859_ _0720_ _0258_ net67 sg13g2_a21oi_1
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_35_789 VPWR VGND sg13g2_decap_8
XFILLER_47_594 VPWR VGND sg13g2_fill_1
X_1914_ net187 VPWR _0605_ VGND daisychain\[99\] net32 sg13g2_o21ai_1
XFILLER_7_690 VPWR VGND sg13g2_fill_2
X_1845_ VGND VPWR _0547_ _0548_ _0213_ _0549_ sg13g2_a21oi_1
X_1776_ state\[72\] daisychain\[72\] net150 _0494_ VPWR VGND sg13g2_mux2_1
X_2328_ net294 VGND VPWR _0144_ daisychain\[16\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_25_222 VPWR VGND sg13g2_decap_8
XFILLER_38_561 VPWR VGND sg13g2_fill_2
XFILLER_38_583 VPWR VGND sg13g2_fill_1
XFILLER_41_715 VPWR VGND sg13g2_fill_2
XFILLER_43_14 VPWR VGND sg13g2_decap_8
X_2259_ VGND VPWR _0611_ _0819_ _0357_ net77 sg13g2_a21oi_1
XFILLER_21_461 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_1_822 VPWR VGND sg13g2_fill_1
XFILLER_4_115 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_16_233 VPWR VGND sg13g2_decap_8
XFILLER_17_92 VPWR VGND sg13g2_decap_8
XFILLER_31_214 VPWR VGND sg13g2_decap_8
XFILLER_32_748 VPWR VGND sg13g2_fill_2
XFILLER_44_542 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_8_432 VPWR VGND sg13g2_fill_1
X_1630_ VGND VPWR _1019_ _1020_ _0170_ _1021_ sg13g2_a21oi_1
XFILLER_39_303 VPWR VGND sg13g2_decap_8
X_1492_ _0911_ net156 _0910_ VPWR VGND sg13g2_nand2_1
X_1561_ state\[29\] daisychain\[29\] net138 _0966_ VPWR VGND sg13g2_mux2_1
X_2113_ VGND VPWR _0963_ _0746_ _0284_ net74 sg13g2_a21oi_1
X_2044_ net178 VPWR _0709_ VGND daisychain\[125\] net26 sg13g2_o21ai_1
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_35_597 VPWR VGND sg13g2_decap_8
Xfanout29 net30 net29 VPWR VGND sg13g2_buf_1
X_2502__336 VPWR VGND net335 sg13g2_tiehi
X_1828_ VGND VPWR net125 daisychain\[81\] _0536_ net61 sg13g2_a21oi_1
X_1759_ net195 VPWR _0481_ VGND daisychain\[68\] net40 sg13g2_o21ai_1
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_41_578 VPWR VGND sg13g2_fill_1
XFILLER_9_218 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_29_380 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_32_589 VPWR VGND sg13g2_fill_1
XFILLER_5_62 VPWR VGND sg13g2_decap_8
XFILLER_8_284 VPWR VGND sg13g2_decap_8
X_1544_ net183 VPWR _0953_ VGND daisychain\[25\] net28 sg13g2_o21ai_1
X_1613_ VGND VPWR net115 daisychain\[38\] _1008_ net57 sg13g2_a21oi_1
XFILLER_27_306 VPWR VGND sg13g2_fill_2
XFILLER_39_100 VPWR VGND sg13g2_decap_8
XFILLER_39_177 VPWR VGND sg13g2_decap_8
X_1475_ VGND VPWR _0895_ _0896_ _0139_ _0897_ sg13g2_a21oi_1
XFILLER_23_512 VPWR VGND sg13g2_decap_8
XFILLER_24_27 VPWR VGND sg13g2_decap_8
XFILLER_27_339 VPWR VGND sg13g2_decap_4
XFILLER_35_350 VPWR VGND sg13g2_decap_8
XFILLER_35_383 VPWR VGND sg13g2_fill_1
X_2027_ _0695_ net154 _0694_ VPWR VGND sg13g2_nand2_1
XFILLER_11_729 VPWR VGND sg13g2_fill_1
XFILLER_2_427 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
X_2400__407 VPWR VGND net406 sg13g2_tiehi
XFILLER_18_306 VPWR VGND sg13g2_fill_2
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_30_81 VPWR VGND sg13g2_decap_8
XFILLER_5_265 VPWR VGND sg13g2_decap_8
XFILLER_6_733 VPWR VGND sg13g2_decap_8
X_2444__312 VPWR VGND net311 sg13g2_tiehi
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_32_386 VPWR VGND sg13g2_decap_4
XFILLER_9_560 VPWR VGND sg13g2_decap_4
X_1527_ _0939_ net161 _0938_ VPWR VGND sg13g2_nand2_1
XFILLER_27_147 VPWR VGND sg13g2_decap_8
X_1389_ VPWR _0043_ state\[23\] VGND sg13g2_inv_1
X_1458_ VGND VPWR net92 daisychain\[7\] _0884_ net45 sg13g2_a21oi_1
XFILLER_23_342 VPWR VGND sg13g2_fill_2
X_2352__247 VPWR VGND net246 sg13g2_tiehi
X_2543__222 VPWR VGND net221 sg13g2_tiehi
XFILLER_2_224 VPWR VGND sg13g2_decap_8
XFILLER_18_158 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_574 VPWR VGND sg13g2_decap_8
X_2430_ net346 VGND VPWR _0246_ daisychain\[118\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2361_ net228 VGND VPWR _0177_ daisychain\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_1312_ VPWR _0001_ state\[100\] VGND sg13g2_inv_1
X_2292_ _0836_ net94 state\[118\] VPWR VGND sg13g2_nand2_1
XFILLER_24_139 VPWR VGND sg13g2_decap_8
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_33_640 VPWR VGND sg13g2_fill_2
XFILLER_20_367 VPWR VGND sg13g2_decap_8
X_2538__302 VPWR VGND net301 sg13g2_tiehi
X_2559_ net373 VGND VPWR _0375_ state\[119\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_15_128 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_11_334 VPWR VGND sg13g2_decap_8
XFILLER_11_378 VPWR VGND sg13g2_fill_1
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_30_109 VPWR VGND sg13g2_decap_8
XFILLER_7_305 VPWR VGND sg13g2_decap_8
XFILLER_11_61 VPWR VGND sg13g2_decap_8
XFILLER_3_500 VPWR VGND sg13g2_decap_8
XFILLER_3_533 VPWR VGND sg13g2_decap_4
XFILLER_3_555 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_14_161 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_decap_8
X_1930_ VGND VPWR _0615_ _0616_ _0230_ _0617_ sg13g2_a21oi_1
XFILLER_30_643 VPWR VGND sg13g2_fill_1
XFILLER_30_676 VPWR VGND sg13g2_fill_2
X_1861_ state\[89\] daisychain\[89\] net149 _0562_ VPWR VGND sg13g2_mux2_1
X_1792_ _0507_ net174 _0506_ VPWR VGND sg13g2_nand2_1
XFILLER_6_393 VPWR VGND sg13g2_decap_8
X_2496__360 VPWR VGND net359 sg13g2_tiehi
X_2413_ net380 VGND VPWR _0229_ daisychain\[101\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2344_ net262 VGND VPWR _0160_ daisychain\[32\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_37_231 VPWR VGND sg13g2_decap_8
X_2275_ VGND VPWR _0643_ _0827_ _0365_ net76 sg13g2_a21oi_1
XFILLER_20_131 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
X_2475__444 VPWR VGND net443 sg13g2_tiehi
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_44_724 VPWR VGND sg13g2_decap_8
XFILLER_11_131 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_4_820 VPWR VGND sg13g2_fill_2
XFILLER_7_179 VPWR VGND sg13g2_decap_8
XFILLER_3_385 VPWR VGND sg13g2_decap_8
X_2523__434 VPWR VGND net433 sg13g2_tiehi
XFILLER_19_253 VPWR VGND sg13g2_decap_8
XFILLER_47_540 VPWR VGND sg13g2_decap_8
X_2060_ _0720_ net91 state\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_30_473 VPWR VGND sg13g2_fill_1
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_8_40 VPWR VGND sg13g2_fill_2
X_1913_ VGND VPWR net109 daisychain\[98\] _0604_ net54 sg13g2_a21oi_1
XFILLER_6_190 VPWR VGND sg13g2_decap_8
XFILLER_7_680 VPWR VGND sg13g2_decap_4
XFILLER_8_95 VPWR VGND sg13g2_decap_8
X_1844_ net194 VPWR _0549_ VGND daisychain\[85\] net39 sg13g2_o21ai_1
X_1775_ VGND VPWR _0491_ _0492_ _0199_ _0493_ sg13g2_a21oi_1
X_2327_ net296 VGND VPWR _0143_ daisychain\[15\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2258_ _0819_ net110 state\[101\] VPWR VGND sg13g2_nand2_1
XFILLER_25_201 VPWR VGND sg13g2_decap_8
XFILLER_27_49 VPWR VGND sg13g2_decap_8
XFILLER_38_573 VPWR VGND sg13g2_fill_1
XFILLER_38_595 VPWR VGND sg13g2_decap_4
XFILLER_41_738 VPWR VGND sg13g2_decap_4
X_2535__338 VPWR VGND net337 sg13g2_tiehi
X_2189_ VGND VPWR _0471_ _0784_ _0322_ net85 sg13g2_a21oi_1
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_5_617 VPWR VGND sg13g2_decap_4
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_16_212 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_17_71 VPWR VGND sg13g2_decap_8
XFILLER_33_81 VPWR VGND sg13g2_decap_8
X_1560_ VGND VPWR _0963_ _0964_ _0156_ _0965_ sg13g2_a21oi_1
XFILLER_39_359 VPWR VGND sg13g2_decap_8
XFILLER_3_182 VPWR VGND sg13g2_decap_8
X_1491_ state\[15\] daisychain\[15\] net134 _0910_ VPWR VGND sg13g2_mux2_1
X_2112_ _0746_ net101 state\[28\] VPWR VGND sg13g2_nand2_1
XFILLER_35_521 VPWR VGND sg13g2_fill_1
XFILLER_35_554 VPWR VGND sg13g2_decap_8
XFILLER_35_587 VPWR VGND sg13g2_decap_4
XFILLER_47_392 VPWR VGND sg13g2_decap_8
X_2043_ VGND VPWR net89 daisychain\[124\] _0708_ net48 sg13g2_a21oi_1
XFILLER_16_790 VPWR VGND sg13g2_decap_4
XFILLER_30_270 VPWR VGND sg13g2_decap_8
X_1827_ _0535_ net172 _0534_ VPWR VGND sg13g2_nand2_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
X_1758_ VGND VPWR net128 daisychain\[67\] _0480_ net63 sg13g2_a21oi_1
X_1689_ net192 VPWR _0425_ VGND daisychain\[54\] net37 sg13g2_o21ai_1
XFILLER_26_510 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_14_705 VPWR VGND sg13g2_decap_4
XFILLER_14_727 VPWR VGND sg13g2_decap_8
XFILLER_41_557 VPWR VGND sg13g2_fill_2
XFILLER_5_447 VPWR VGND sg13g2_fill_1
X_2362__227 VPWR VGND net226 sg13g2_tiehi
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
X_2407__393 VPWR VGND net392 sg13g2_tiehi
XFILLER_17_554 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_12_281 VPWR VGND sg13g2_decap_8
XFILLER_20_719 VPWR VGND sg13g2_fill_1
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
XFILLER_9_731 VPWR VGND sg13g2_decap_8
XFILLER_9_742 VPWR VGND sg13g2_fill_1
X_1474_ net179 VPWR _0897_ VGND daisychain\[11\] net23 sg13g2_o21ai_1
X_1543_ VGND VPWR net104 daisychain\[24\] _0952_ net51 sg13g2_a21oi_1
X_1612_ _1007_ net168 _1006_ VPWR VGND sg13g2_nand2_1
XFILLER_27_318 VPWR VGND sg13g2_decap_8
XFILLER_39_156 VPWR VGND sg13g2_decap_8
X_2026_ state\[122\] daisychain\[122\] net136 _0694_ VPWR VGND sg13g2_mux2_1
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_2_406 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_26_373 VPWR VGND sg13g2_decap_4
XFILLER_45_126 VPWR VGND sg13g2_decap_8
X_2472__200 VPWR VGND net sg13g2_tiehi
XFILLER_10_763 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_10_796 VPWR VGND sg13g2_fill_1
XFILLER_30_60 VPWR VGND sg13g2_decap_8
XFILLER_5_244 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_37_627 VPWR VGND sg13g2_fill_2
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_20_505 VPWR VGND sg13g2_fill_1
XFILLER_32_365 VPWR VGND sg13g2_decap_8
XFILLER_33_811 VPWR VGND sg13g2_decap_8
XFILLER_33_822 VPWR VGND sg13g2_fill_1
X_1457_ _0883_ net155 _0882_ VPWR VGND sg13g2_nand2_1
X_1526_ state\[22\] daisychain\[22\] net139 _0938_ VPWR VGND sg13g2_mux2_1
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
X_1388_ VPWR _0044_ state\[24\] VGND sg13g2_inv_1
XFILLER_23_310 VPWR VGND sg13g2_fill_1
XFILLER_7_509 VPWR VGND sg13g2_decap_8
X_2009_ net181 VPWR _0681_ VGND daisychain\[118\] net25 sg13g2_o21ai_1
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_3_715 VPWR VGND sg13g2_fill_1
XFILLER_19_605 VPWR VGND sg13g2_fill_1
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_30_803 VPWR VGND sg13g2_fill_1
XFILLER_30_814 VPWR VGND sg13g2_fill_1
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_542 VPWR VGND sg13g2_decap_8
X_2526__410 VPWR VGND net409 sg13g2_tiehi
X_1311_ VPWR _0002_ state\[101\] VGND sg13g2_inv_1
X_2360_ net230 VGND VPWR _0176_ daisychain\[48\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2291_ VGND VPWR _0675_ _0835_ _0373_ net69 sg13g2_a21oi_1
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_20 VPWR VGND sg13g2_decap_4
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_20_324 VPWR VGND sg13g2_decap_4
XFILLER_24_118 VPWR VGND sg13g2_decap_8
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_0_718 VPWR VGND sg13g2_fill_1
XFILLER_28_402 VPWR VGND sg13g2_fill_2
X_1509_ net182 VPWR _0925_ VGND daisychain\[18\] net27 sg13g2_o21ai_1
X_2558_ net405 VGND VPWR _0374_ state\[118\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2489_ net387 VGND VPWR _0305_ state\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_15_107 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_11_313 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_8_818 VPWR VGND sg13g2_decap_4
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_14_140 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
X_1860_ VGND VPWR _0559_ _0560_ _0216_ _0561_ sg13g2_a21oi_1
XFILLER_6_372 VPWR VGND sg13g2_decap_8
X_1791_ state\[75\] daisychain\[75\] net150 _0506_ VPWR VGND sg13g2_mux2_1
X_2412_ net382 VGND VPWR _0228_ daisychain\[100\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2343_ net264 VGND VPWR _0159_ daisychain\[31\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2274_ _0827_ net109 state\[109\] VPWR VGND sg13g2_nand2_1
XFILLER_37_210 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_38_733 VPWR VGND sg13g2_fill_1
XFILLER_38_788 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_17_clk clknet_2_1__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_20_110 VPWR VGND sg13g2_decap_8
XFILLER_20_187 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
X_1989_ net180 VPWR _0665_ VGND daisychain\[114\] net24 sg13g2_o21ai_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
X_2321__309 VPWR VGND net308 sg13g2_tiehi
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_11_110 VPWR VGND sg13g2_decap_8
XFILLER_12_622 VPWR VGND sg13g2_decap_4
XFILLER_16_449 VPWR VGND sg13g2_decap_8
XFILLER_24_482 VPWR VGND sg13g2_decap_8
XFILLER_31_408 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_11_187 VPWR VGND sg13g2_decap_8
XFILLER_7_158 VPWR VGND sg13g2_decap_8
XFILLER_8_648 VPWR VGND sg13g2_fill_1
X_2482__416 VPWR VGND net415 sg13g2_tiehi
XFILLER_3_364 VPWR VGND sg13g2_decap_8
XFILLER_19_232 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_35_736 VPWR VGND sg13g2_fill_1
XFILLER_35_747 VPWR VGND sg13g2_decap_8
XFILLER_47_563 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
X_2417__373 VPWR VGND net372 sg13g2_tiehi
X_2372__207 VPWR VGND net206 sg13g2_tiehi
XFILLER_8_74 VPWR VGND sg13g2_decap_8
X_1912_ _0603_ net166 _0602_ VPWR VGND sg13g2_nand2_1
X_1843_ VGND VPWR net124 daisychain\[84\] _0548_ net62 sg13g2_a21oi_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_6_clk clknet_2_3__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_1774_ net196 VPWR _0493_ VGND daisychain\[71\] net41 sg13g2_o21ai_1
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_38_563 VPWR VGND sg13g2_fill_1
X_2326_ net298 VGND VPWR _0142_ daisychain\[14\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2257_ VGND VPWR _0607_ _0818_ _0356_ net78 sg13g2_a21oi_1
XFILLER_25_257 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
X_2188_ _0784_ net128 state\[66\] VPWR VGND sg13g2_nand2_1
XFILLER_21_496 VPWR VGND sg13g2_decap_8
X_2509__290 VPWR VGND net289 sg13g2_tiehi
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_17_747 VPWR VGND sg13g2_decap_4
XFILLER_29_530 VPWR VGND sg13g2_fill_1
XFILLER_44_566 VPWR VGND sg13g2_decap_8
XFILLER_12_496 VPWR VGND sg13g2_fill_1
XFILLER_16_268 VPWR VGND sg13g2_decap_8
XFILLER_31_249 VPWR VGND sg13g2_decap_8
XFILLER_33_60 VPWR VGND sg13g2_decap_8
X_2447__300 VPWR VGND net299 sg13g2_tiehi
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_1490_ VGND VPWR _0907_ _0908_ _0142_ _0909_ sg13g2_a21oi_1
XFILLER_39_338 VPWR VGND sg13g2_decap_8
X_2111_ VGND VPWR _0959_ _0745_ _0283_ net71 sg13g2_a21oi_1
X_2042_ _0707_ net154 _0706_ VPWR VGND sg13g2_nand2_1
XFILLER_22_249 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_31_783 VPWR VGND sg13g2_decap_4
X_1826_ state\[82\] daisychain\[82\] net148 _0534_ VPWR VGND sg13g2_mux2_1
X_1757_ _0479_ net174 _0478_ VPWR VGND sg13g2_nand2_1
X_1688_ VGND VPWR net119 daisychain\[53\] _0424_ net59 sg13g2_a21oi_1
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
X_2309_ VGND VPWR _0711_ _0844_ _0382_ net70 sg13g2_a21oi_1
XFILLER_13_249 VPWR VGND sg13g2_decap_8
XFILLER_21_293 VPWR VGND sg13g2_decap_4
XFILLER_5_426 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_49_636 VPWR VGND sg13g2_decap_8
XFILLER_17_588 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_12_260 VPWR VGND sg13g2_decap_8
XFILLER_13_794 VPWR VGND sg13g2_fill_2
XFILLER_40_591 VPWR VGND sg13g2_decap_8
XFILLER_8_242 VPWR VGND sg13g2_decap_8
X_1611_ state\[39\] daisychain\[39\] net144 _1006_ VPWR VGND sg13g2_mux2_1
XFILLER_5_20 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_fill_2
XFILLER_5_97 VPWR VGND sg13g2_decap_8
X_1473_ VGND VPWR net93 daisychain\[10\] _0896_ net45 sg13g2_a21oi_1
X_1542_ _0951_ net161 _0950_ VPWR VGND sg13g2_nand2_1
XFILLER_27_308 VPWR VGND sg13g2_fill_1
XFILLER_39_135 VPWR VGND sg13g2_decap_8
X_2025_ VGND VPWR _0691_ _0692_ _0249_ _0693_ sg13g2_a21oi_1
XFILLER_35_374 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
X_1809_ net196 VPWR _0521_ VGND daisychain\[78\] net41 sg13g2_o21ai_1
XFILLER_14_514 VPWR VGND sg13g2_decap_8
XFILLER_14_525 VPWR VGND sg13g2_fill_2
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_10_742 VPWR VGND sg13g2_decap_8
XFILLER_14_84 VPWR VGND sg13g2_decap_8
XFILLER_6_713 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_5_223 VPWR VGND sg13g2_decap_8
X_2520__202 VPWR VGND net201 sg13g2_tiehi
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_32_311 VPWR VGND sg13g2_fill_1
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_45_661 VPWR VGND sg13g2_fill_2
X_1387_ VPWR _0045_ state\[25\] VGND sg13g2_inv_1
X_1456_ state\[8\] daisychain\[8\] net134 _0882_ VPWR VGND sg13g2_mux2_1
X_1525_ VGND VPWR _0935_ _0936_ _0149_ _0937_ sg13g2_a21oi_1
XFILLER_27_105 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
X_2008_ VGND VPWR net94 daisychain\[117\] _0680_ net46 sg13g2_a21oi_1
XFILLER_2_259 VPWR VGND sg13g2_decap_8
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_19_628 VPWR VGND sg13g2_decap_4
X_2478__432 VPWR VGND net431 sg13g2_tiehi
XFILLER_14_322 VPWR VGND sg13g2_fill_1
XFILLER_14_355 VPWR VGND sg13g2_fill_2
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_10_583 VPWR VGND sg13g2_fill_2
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
X_1310_ VPWR _0003_ state\[102\] VGND sg13g2_inv_1
Xheichips25_pudding VPWR VGND uio_oe[0] sg13g2_tiehi
X_2381__445 VPWR VGND net444 sg13g2_tiehi
X_2290_ _0835_ net94 state\[117\] VPWR VGND sg13g2_nand2_1
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_32_130 VPWR VGND sg13g2_decap_8
XFILLER_33_642 VPWR VGND sg13g2_fill_1
X_2557_ net437 VGND VPWR _0373_ state\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2427__353 VPWR VGND net352 sg13g2_tiehi
XFILLER_46_49 VPWR VGND sg13g2_decap_8
X_1439_ net186 VPWR _0869_ VGND daisychain\[4\] net31 sg13g2_o21ai_1
X_1508_ VGND VPWR net99 daisychain\[17\] _0924_ net49 sg13g2_a21oi_1
X_2488_ net391 VGND VPWR _0304_ state\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_11_369 VPWR VGND sg13g2_decap_8
XFILLER_11_96 VPWR VGND sg13g2_decap_8
XFILLER_3_513 VPWR VGND sg13g2_decap_8
X_2328__295 VPWR VGND net294 sg13g2_tiehi
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_14_196 VPWR VGND sg13g2_decap_8
XFILLER_15_642 VPWR VGND sg13g2_fill_1
XFILLER_15_697 VPWR VGND sg13g2_fill_2
XFILLER_30_601 VPWR VGND sg13g2_fill_1
XFILLER_30_656 VPWR VGND sg13g2_fill_1
XFILLER_30_689 VPWR VGND sg13g2_fill_1
X_1790_ VGND VPWR _0503_ _0504_ _0202_ _0505_ sg13g2_a21oi_1
XFILLER_6_351 VPWR VGND sg13g2_decap_8
X_2411_ net384 VGND VPWR _0227_ daisychain\[99\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_38_701 VPWR VGND sg13g2_fill_2
XFILLER_38_712 VPWR VGND sg13g2_fill_2
X_2342_ net266 VGND VPWR _0158_ daisychain\[30\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2273_ VGND VPWR _0639_ _0826_ _0364_ net75 sg13g2_a21oi_1
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_38_778 VPWR VGND sg13g2_fill_1
XFILLER_20_166 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
X_1988_ VGND VPWR net95 daisychain\[113\] _0664_ net46 sg13g2_a21oi_1
XFILLER_28_200 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_decap_4
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_24_461 VPWR VGND sg13g2_decap_8
XFILLER_8_605 VPWR VGND sg13g2_fill_2
XFILLER_11_166 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_343 VPWR VGND sg13g2_decap_8
XFILLER_4_822 VPWR VGND sg13g2_fill_1
XFILLER_7_137 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_19_211 VPWR VGND sg13g2_decap_8
Xfanout190 net198 net190 VPWR VGND sg13g2_buf_1
XFILLER_34_203 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_30_420 VPWR VGND sg13g2_fill_1
XFILLER_42_280 VPWR VGND sg13g2_decap_8
XFILLER_8_42 VPWR VGND sg13g2_fill_1
XFILLER_8_53 VPWR VGND sg13g2_decap_8
X_1911_ state\[99\] daisychain\[99\] net141 _0602_ VPWR VGND sg13g2_mux2_1
X_1842_ _0547_ net173 _0546_ VPWR VGND sg13g2_nand2_1
X_1773_ VGND VPWR net128 daisychain\[70\] _0492_ net64 sg13g2_a21oi_1
X_2325_ net300 VGND VPWR _0141_ daisychain\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2256_ _0818_ net112 state\[100\] VPWR VGND sg13g2_nand2_1
X_2187_ VGND VPWR _0467_ _0783_ _0321_ net86 sg13g2_a21oi_1
XFILLER_25_236 VPWR VGND sg13g2_decap_8
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_21_475 VPWR VGND sg13g2_decap_8
XFILLER_4_129 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_16_247 VPWR VGND sg13g2_decap_8
XFILLER_17_726 VPWR VGND sg13g2_decap_8
XFILLER_32_718 VPWR VGND sg13g2_fill_2
XFILLER_31_228 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_fill_1
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_4_685 VPWR VGND sg13g2_decap_8
XFILLER_39_317 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
X_2110_ _0745_ net102 state\[27\] VPWR VGND sg13g2_nand2_1
X_2041_ state\[125\] daisychain\[125\] net136 _0706_ VPWR VGND sg13g2_mux2_1
XFILLER_22_228 VPWR VGND sg13g2_decap_8
XFILLER_31_751 VPWR VGND sg13g2_decap_4
XFILLER_31_762 VPWR VGND sg13g2_fill_2
XFILLER_35_578 VPWR VGND sg13g2_decap_4
X_1825_ VGND VPWR _0531_ _0532_ _0209_ _0533_ sg13g2_a21oi_1
X_1756_ state\[68\] daisychain\[68\] net151 _0478_ VPWR VGND sg13g2_mux2_1
XFILLER_38_28 VPWR VGND sg13g2_decap_4
X_2308_ _0844_ net90 state\[126\] VPWR VGND sg13g2_nand2_1
X_1687_ _0423_ net170 _0422_ VPWR VGND sg13g2_nand2_1
XFILLER_38_350 VPWR VGND sg13g2_decap_8
X_2239_ VGND VPWR _0571_ _0809_ _0347_ net83 sg13g2_a21oi_1
XFILLER_13_228 VPWR VGND sg13g2_decap_8
XFILLER_5_405 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_49_659 VPWR VGND sg13g2_decap_4
XFILLER_13_751 VPWR VGND sg13g2_decap_8
XFILLER_29_394 VPWR VGND sg13g2_decap_4
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
XFILLER_8_298 VPWR VGND sg13g2_decap_8
X_1610_ VGND VPWR _1003_ _1004_ _0166_ _1005_ sg13g2_a21oi_1
XFILLER_39_114 VPWR VGND sg13g2_decap_8
XFILLER_4_471 VPWR VGND sg13g2_fill_1
XFILLER_4_482 VPWR VGND sg13g2_decap_4
XFILLER_5_76 VPWR VGND sg13g2_decap_8
X_1472_ _0895_ net156 _0894_ VPWR VGND sg13g2_nand2_1
X_1541_ state\[25\] daisychain\[25\] net137 _0950_ VPWR VGND sg13g2_mux2_1
XFILLER_35_364 VPWR VGND sg13g2_decap_4
X_2391__425 VPWR VGND net424 sg13g2_tiehi
X_2024_ net178 VPWR _0693_ VGND daisychain\[121\] net26 sg13g2_o21ai_1
XFILLER_10_209 VPWR VGND sg13g2_decap_8
XFILLER_23_526 VPWR VGND sg13g2_decap_4
X_1808_ VGND VPWR net127 daisychain\[77\] _0520_ net63 sg13g2_a21oi_1
X_1739_ net196 VPWR _0465_ VGND daisychain\[64\] net41 sg13g2_o21ai_1
XFILLER_46_607 VPWR VGND sg13g2_decap_4
X_2437__333 VPWR VGND net332 sg13g2_tiehi
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_decap_4
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_5_202 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_30_95 VPWR VGND sg13g2_decap_8
XFILLER_5_279 VPWR VGND sg13g2_decap_8
XFILLER_17_320 VPWR VGND sg13g2_fill_1
XFILLER_17_342 VPWR VGND sg13g2_fill_1
XFILLER_18_821 VPWR VGND sg13g2_fill_2
XFILLER_37_629 VPWR VGND sg13g2_fill_1
XFILLER_39_93 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
X_2338__275 VPWR VGND net274 sg13g2_tiehi
XFILLER_44_161 VPWR VGND sg13g2_decap_8
X_1524_ net183 VPWR _0937_ VGND daisychain\[21\] net28 sg13g2_o21ai_1
XFILLER_4_290 VPWR VGND sg13g2_decap_8
X_1386_ VPWR _0046_ state\[26\] VGND sg13g2_inv_1
X_1455_ VGND VPWR _0879_ _0880_ _0135_ _0881_ sg13g2_a21oi_1
XFILLER_35_161 VPWR VGND sg13g2_decap_8
X_2007_ _0679_ net157 _0678_ VPWR VGND sg13g2_nand2_1
XFILLER_11_529 VPWR VGND sg13g2_decap_8
XFILLER_2_238 VPWR VGND sg13g2_decap_8
XFILLER_3_728 VPWR VGND sg13g2_fill_2
XFILLER_33_109 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_14_301 VPWR VGND sg13g2_decap_8
XFILLER_14_378 VPWR VGND sg13g2_decap_8
XFILLER_25_73 VPWR VGND sg13g2_decap_4
XFILLER_26_183 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
X_2485__404 VPWR VGND net403 sg13g2_tiehi
XFILLER_6_511 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_17_183 VPWR VGND sg13g2_decap_8
XFILLER_18_695 VPWR VGND sg13g2_fill_2
XFILLER_24_109 VPWR VGND sg13g2_decap_4
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_9_393 VPWR VGND sg13g2_decap_8
X_1507_ _0923_ net159 _0922_ VPWR VGND sg13g2_nand2_1
X_2556_ net213 VGND VPWR _0372_ state\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2487_ net395 VGND VPWR _0303_ state\[47\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_404 VPWR VGND sg13g2_fill_1
XFILLER_46_28 VPWR VGND sg13g2_decap_8
X_1369_ VPWR _0065_ state\[43\] VGND sg13g2_inv_1
X_1438_ VGND VPWR net94 daisychain\[3\] _0868_ net46 sg13g2_a21oi_1
XFILLER_11_348 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_11_75 VPWR VGND sg13g2_decap_8
XFILLER_7_319 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_fill_1
Xdac dac/VbiasP[1] dac/IOUT dac/VbiasP[0] state\[64\] _0088_ state\[65\] _0089_ state\[66\]
+ _0090_ state\[67\] _0091_ state\[68\] _0092_ state\[69\] _0093_ state\[70\] _0095_
+ state\[71\] _0096_ state\[72\] _0097_ digitalen.g\[2\].u.OUTP digitalen.g\[2\].u.OUTN
+ state\[73\] _0098_ state\[74\] _0099_ state\[75\] _0100_ state\[76\] _0101_ state\[77\]
+ _0102_ state\[78\] _0103_ state\[79\] _0104_ state\[80\] _0106_ state\[81\] _0107_
+ state\[82\] _0108_ state\[83\] _0109_ state\[84\] _0110_ state\[85\] _0111_ state\[86\]
+ _0112_ state\[87\] _0113_ state\[88\] _0114_ state\[89\] _0115_ state\[90\] _0117_
+ state\[91\] _0118_ state\[92\] _0119_ state\[93\] _0120_ state\[94\] _0121_ state\[95\]
+ _0122_ state\[96\] _0123_ state\[97\] _0124_ state\[98\] _0125_ state\[99\] _0126_
+ state\[100\] _0001_ state\[101\] _0002_ state\[102\] _0003_ state\[103\] _0004_
+ state\[104\] _0005_ state\[105\] _0006_ state\[106\] _0007_ state\[107\] _0008_
+ state\[108\] _0009_ state\[109\] _0010_ state\[110\] _0012_ state\[111\] _0013_
+ state\[112\] _0014_ state\[113\] _0015_ state\[114\] _0016_ state\[115\] _0017_
+ state\[116\] _0018_ state\[117\] _0019_ state\[118\] _0020_ state\[119\] _0021_
+ state\[120\] _0023_ state\[121\] _0024_ state\[122\] _0025_ digitalen.g\[3\].u.OUTP
+ digitalen.g\[3\].u.OUTN state\[123\] _0026_ state\[124\] _0027_ state\[125\] _0028_
+ state\[126\] _0029_ state\[127\] _0030_ state\[0\] _0000_ state\[1\] _0039_ state\[2\]
+ _0050_ state\[3\] _0061_ state\[4\] _0072_ state\[5\] _0083_ state\[6\] digitalen.g\[0\].u.OUTP
+ digitalen.g\[0\].u.OUTN _0094_ state\[7\] _0105_ state\[8\] _0116_ state\[9\] _0127_
+ state\[10\] _0011_ state\[11\] _0022_ state\[12\] _0031_ state\[13\] _0032_ state\[14\]
+ _0033_ state\[15\] _0034_ state\[16\] _0035_ state\[17\] _0036_ state\[18\] _0037_
+ state\[19\] _0038_ state\[20\] _0040_ state\[21\] _0041_ state\[22\] _0042_ state\[23\]
+ _0043_ state\[24\] _0044_ state\[25\] _0045_ state\[26\] _0046_ state\[27\] _0047_
+ state\[28\] _0048_ state\[29\] _0049_ state\[30\] _0051_ state\[31\] _0052_ state\[33\]
+ _0054_ state\[32\] _0053_ state\[34\] _0055_ state\[35\] _0056_ state\[36\] _0057_
+ state\[37\] _0058_ state\[38\] _0059_ state\[39\] _0060_ state\[40\] _0062_ state\[41\]
+ _0063_ state\[42\] _0064_ state\[43\] _0065_ state\[44\] _0066_ state\[45\] _0067_
+ state\[46\] _0068_ state\[47\] _0069_ state\[48\] _0070_ state\[49\] _0071_ state\[50\]
+ _0073_ state\[51\] _0074_ state\[52\] _0075_ state\[53\] _0076_ state\[54\] _0077_
+ state\[55\] _0078_ state\[56\] _0079_ state\[57\] _0080_ state\[58\] _0081_ state\[59\]
+ _0082_ state\[60\] _0084_ state\[61\] _0085_ state\[62\] _0086_ state\[63\] _0087_
+ digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN dac/VcascP[1] dac/VcascP[0] VGND
+ VPWR dac128module
XFILLER_19_415 VPWR VGND sg13g2_fill_1
XFILLER_19_459 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_10_370 VPWR VGND sg13g2_decap_8
XFILLER_14_175 VPWR VGND sg13g2_decap_8
XFILLER_30_635 VPWR VGND sg13g2_fill_1
XFILLER_30_668 VPWR VGND sg13g2_fill_1
XFILLER_42_462 VPWR VGND sg13g2_decap_8
XFILLER_6_330 VPWR VGND sg13g2_decap_8
X_2410_ net386 VGND VPWR _0226_ daisychain\[98\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2341_ net268 VGND VPWR _0157_ daisychain\[29\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_37_245 VPWR VGND sg13g2_decap_8
XFILLER_38_757 VPWR VGND sg13g2_fill_2
X_2272_ _0826_ net109 state\[108\] VPWR VGND sg13g2_nand2_1
XFILLER_20_145 VPWR VGND sg13g2_decap_8
XFILLER_9_190 VPWR VGND sg13g2_decap_8
X_1987_ _0663_ net157 _0662_ VPWR VGND sg13g2_nand2_1
XFILLER_0_539 VPWR VGND sg13g2_decap_8
X_2539_ net285 VGND VPWR _0355_ state\[99\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_11_145 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_decap_8
XFILLER_8_628 VPWR VGND sg13g2_decap_4
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_3_322 VPWR VGND sg13g2_decap_8
XFILLER_3_399 VPWR VGND sg13g2_decap_8
XFILLER_47_554 VPWR VGND sg13g2_decap_4
Xfanout180 net181 net180 VPWR VGND sg13g2_buf_1
Xfanout191 net198 net191 VPWR VGND sg13g2_buf_1
XFILLER_15_462 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_43_782 VPWR VGND sg13g2_decap_4
X_1910_ VGND VPWR _0599_ _0600_ _0226_ _0601_ sg13g2_a21oi_1
X_1841_ state\[85\] daisychain\[85\] net149 _0546_ VPWR VGND sg13g2_mux2_1
X_1772_ _0491_ net175 _0490_ VPWR VGND sg13g2_nand2_1
X_2324_ net302 VGND VPWR _0140_ daisychain\[12\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2320__311 VPWR VGND net310 sg13g2_tiehi
XFILLER_25_215 VPWR VGND sg13g2_decap_8
XFILLER_38_521 VPWR VGND sg13g2_fill_1
XFILLER_38_554 VPWR VGND sg13g2_decap_8
X_2255_ VGND VPWR _0603_ _0817_ _0355_ net76 sg13g2_a21oi_1
X_2186_ _0783_ net130 state\[65\] VPWR VGND sg13g2_nand2_1
XFILLER_21_410 VPWR VGND sg13g2_fill_2
XFILLER_21_454 VPWR VGND sg13g2_decap_8
XFILLER_33_270 VPWR VGND sg13g2_decap_8
XFILLER_34_771 VPWR VGND sg13g2_fill_2
XFILLER_41_708 VPWR VGND sg13g2_decap_8
XFILLER_4_108 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_16_226 VPWR VGND sg13g2_decap_8
XFILLER_17_85 VPWR VGND sg13g2_decap_8
XFILLER_31_207 VPWR VGND sg13g2_decap_8
XFILLER_44_535 VPWR VGND sg13g2_decap_8
XFILLER_12_443 VPWR VGND sg13g2_decap_8
XFILLER_12_454 VPWR VGND sg13g2_decap_4
XFILLER_33_95 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_8_447 VPWR VGND sg13g2_decap_8
XFILLER_3_196 VPWR VGND sg13g2_decap_8
X_2040_ VGND VPWR _0703_ _0704_ _0252_ _0705_ sg13g2_a21oi_1
XFILLER_16_771 VPWR VGND sg13g2_fill_2
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_31_730 VPWR VGND sg13g2_decap_8
XFILLER_35_568 VPWR VGND sg13g2_decap_4
XFILLER_30_295 VPWR VGND sg13g2_decap_8
X_2348__255 VPWR VGND net254 sg13g2_tiehi
X_1824_ net194 VPWR _0533_ VGND daisychain\[81\] net39 sg13g2_o21ai_1
X_1755_ VGND VPWR _0475_ _0476_ _0195_ _0477_ sg13g2_a21oi_1
X_1686_ state\[54\] daisychain\[54\] net146 _0422_ VPWR VGND sg13g2_mux2_1
X_2307_ VGND VPWR _0707_ _0843_ _0381_ net70 sg13g2_a21oi_1
X_2238_ _0809_ net126 state\[91\] VPWR VGND sg13g2_nand2_1
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_26_524 VPWR VGND sg13g2_decap_8
X_2169_ VGND VPWR _0431_ _0774_ _0312_ net81 sg13g2_a21oi_1
XFILLER_21_262 VPWR VGND sg13g2_decap_4
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_656 VPWR VGND sg13g2_fill_2
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_29_362 VPWR VGND sg13g2_decap_4
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_17_568 VPWR VGND sg13g2_fill_2
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_12_295 VPWR VGND sg13g2_decap_8
XFILLER_5_55 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
XFILLER_9_778 VPWR VGND sg13g2_fill_2
X_1540_ VGND VPWR _0947_ _0948_ _0152_ _0949_ sg13g2_a21oi_1
X_1471_ state\[11\] daisychain\[11\] net133 _0894_ VPWR VGND sg13g2_mux2_1
X_2501__340 VPWR VGND net339 sg13g2_tiehi
XFILLER_23_505 VPWR VGND sg13g2_decap_8
XFILLER_35_343 VPWR VGND sg13g2_decap_8
X_2023_ VGND VPWR net89 daisychain\[120\] _0692_ net48 sg13g2_a21oi_1
XFILLER_31_593 VPWR VGND sg13g2_decap_4
X_1807_ _0519_ net175 _0518_ VPWR VGND sg13g2_nand2_1
XFILLER_49_39 VPWR VGND sg13g2_decap_8
X_1738_ VGND VPWR net130 daisychain\[63\] _0464_ net64 sg13g2_a21oi_1
X_1669_ net190 VPWR _0409_ VGND daisychain\[50\] net35 sg13g2_o21ai_1
XFILLER_26_332 VPWR VGND sg13g2_decap_8
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_10_777 VPWR VGND sg13g2_decap_8
XFILLER_30_74 VPWR VGND sg13g2_decap_8
XFILLER_5_258 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_39_72 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_17_332 VPWR VGND sg13g2_decap_4
XFILLER_17_387 VPWR VGND sg13g2_fill_2
XFILLER_29_192 VPWR VGND sg13g2_decap_8
XFILLER_32_302 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_45_663 VPWR VGND sg13g2_fill_1
XFILLER_32_379 VPWR VGND sg13g2_decap_8
XFILLER_9_553 VPWR VGND sg13g2_decap_8
XFILLER_9_564 VPWR VGND sg13g2_fill_2
X_1454_ net179 VPWR _0881_ VGND daisychain\[7\] net23 sg13g2_o21ai_1
X_1523_ VGND VPWR net99 daisychain\[20\] _0936_ net49 sg13g2_a21oi_1
XFILLER_48_490 VPWR VGND sg13g2_decap_8
X_1385_ VPWR _0047_ state\[27\] VGND sg13g2_inv_1
XFILLER_35_140 VPWR VGND sg13g2_decap_8
X_2006_ state\[118\] daisychain\[118\] net153 _0678_ VPWR VGND sg13g2_mux2_1
X_2839_ state\[127\] net14 VPWR VGND sg13g2_buf_1
XFILLER_2_217 VPWR VGND sg13g2_decap_8
XFILLER_4_8 VPWR VGND sg13g2_fill_1
X_2404__399 VPWR VGND net398 sg13g2_tiehi
XFILLER_26_162 VPWR VGND sg13g2_decap_8
XFILLER_42_611 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_14_335 VPWR VGND sg13g2_fill_2
XFILLER_25_52 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_6_556 VPWR VGND sg13g2_fill_1
XFILLER_6_567 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_37_405 VPWR VGND sg13g2_decap_4
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_17_162 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_9_372 VPWR VGND sg13g2_decap_8
X_1437_ _0867_ net164 _0866_ VPWR VGND sg13g2_nand2_1
X_1506_ state\[18\] daisychain\[18\] net137 _0922_ VPWR VGND sg13g2_mux2_1
X_2555_ net245 VGND VPWR _0371_ state\[115\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2486_ net399 VGND VPWR _0302_ state\[46\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_416 VPWR VGND sg13g2_fill_1
XFILLER_36_460 VPWR VGND sg13g2_fill_1
X_1299_ VPWR _0015_ state\[113\] VGND sg13g2_inv_1
X_1368_ VPWR _0066_ state\[44\] VGND sg13g2_inv_1
XFILLER_11_327 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_11_54 VPWR VGND sg13g2_decap_8
XFILLER_3_548 VPWR VGND sg13g2_fill_2
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_47_725 VPWR VGND sg13g2_fill_1
XFILLER_14_154 VPWR VGND sg13g2_decap_8
XFILLER_15_600 VPWR VGND sg13g2_fill_1
XFILLER_27_493 VPWR VGND sg13g2_fill_2
XFILLER_30_614 VPWR VGND sg13g2_fill_1
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_42_441 VPWR VGND sg13g2_decap_8
XFILLER_30_647 VPWR VGND sg13g2_fill_1
XFILLER_2_570 VPWR VGND sg13g2_decap_4
XFILLER_6_386 VPWR VGND sg13g2_decap_8
X_2340_ net270 VGND VPWR _0156_ daisychain\[28\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2271_ VGND VPWR _0635_ _0825_ _0363_ net75 sg13g2_a21oi_1
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
XFILLER_38_703 VPWR VGND sg13g2_fill_1
XFILLER_20_124 VPWR VGND sg13g2_decap_8
X_1986_ state\[114\] daisychain\[114\] net135 _0662_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
X_2538_ net301 VGND VPWR _0354_ state\[98\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2469_ net211 VGND VPWR _0285_ state\[29\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2358__235 VPWR VGND net234 sg13g2_tiehi
XFILLER_16_419 VPWR VGND sg13g2_fill_2
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_44_739 VPWR VGND sg13g2_decap_8
XFILLER_11_124 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_24_496 VPWR VGND sg13g2_decap_8
XFILLER_4_802 VPWR VGND sg13g2_fill_2
XFILLER_3_301 VPWR VGND sg13g2_decap_8
XFILLER_3_378 VPWR VGND sg13g2_decap_8
XFILLER_4_813 VPWR VGND sg13g2_decap_8
XFILLER_19_246 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_47_533 VPWR VGND sg13g2_decap_8
X_2556__214 VPWR VGND net213 sg13g2_tiehi
Xfanout170 net171 net170 VPWR VGND sg13g2_buf_1
Xfanout181 net199 net181 VPWR VGND sg13g2_buf_1
Xfanout192 net193 net192 VPWR VGND sg13g2_buf_1
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_43_761 VPWR VGND sg13g2_decap_8
XFILLER_8_33 VPWR VGND sg13g2_decap_8
X_1840_ VGND VPWR _0543_ _0544_ _0212_ _0545_ sg13g2_a21oi_1
XFILLER_6_183 VPWR VGND sg13g2_decap_8
XFILLER_7_673 VPWR VGND sg13g2_fill_2
XFILLER_7_684 VPWR VGND sg13g2_fill_2
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_1771_ state\[71\] daisychain\[71\] net150 _0490_ VPWR VGND sg13g2_mux2_1
X_2323_ net304 VGND VPWR _0139_ daisychain\[11\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2254_ _0817_ net112 state\[99\] VPWR VGND sg13g2_nand2_1
XFILLER_19_0 VPWR VGND sg13g2_fill_2
XFILLER_38_588 VPWR VGND sg13g2_decap_8
XFILLER_38_599 VPWR VGND sg13g2_fill_1
X_2185_ VGND VPWR _0463_ _0782_ _0320_ net86 sg13g2_a21oi_1
XFILLER_21_444 VPWR VGND sg13g2_fill_2
X_1969_ net189 VPWR _0649_ VGND daisychain\[110\] net34 sg13g2_o21ai_1
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_16_205 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_12_400 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_decap_8
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_15_282 VPWR VGND sg13g2_decap_8
XFILLER_16_783 VPWR VGND sg13g2_decap_8
XFILLER_30_263 VPWR VGND sg13g2_decap_8
XFILLER_43_591 VPWR VGND sg13g2_decap_4
X_1823_ VGND VPWR net126 daisychain\[80\] _0532_ net62 sg13g2_a21oi_1
XFILLER_7_481 VPWR VGND sg13g2_fill_1
X_1754_ net195 VPWR _0477_ VGND daisychain\[67\] net40 sg13g2_o21ai_1
X_1685_ VGND VPWR _0419_ _0420_ _0181_ _0421_ sg13g2_a21oi_1
XFILLER_26_503 VPWR VGND sg13g2_fill_2
X_2539__286 VPWR VGND net285 sg13g2_tiehi
X_2306_ _0843_ net90 state\[125\] VPWR VGND sg13g2_nand2_1
X_2237_ VGND VPWR _0567_ _0808_ _0346_ net84 sg13g2_a21oi_1
XFILLER_14_709 VPWR VGND sg13g2_fill_2
Xheichips25_pudding_460 VPWR VGND uio_oe[5] sg13g2_tiehi
X_2168_ _0774_ net121 state\[56\] VPWR VGND sg13g2_nand2_1
X_2099_ VGND VPWR _0935_ _0739_ _0277_ net72 sg13g2_a21oi_1
XFILLER_21_241 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_49_606 VPWR VGND sg13g2_decap_4
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_17_525 VPWR VGND sg13g2_fill_2
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_29_341 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_12_274 VPWR VGND sg13g2_decap_8
XFILLER_13_775 VPWR VGND sg13g2_decap_4
XFILLER_40_572 VPWR VGND sg13g2_fill_1
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
X_2414__379 VPWR VGND net378 sg13g2_tiehi
XFILLER_4_451 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_8
X_1470_ VGND VPWR _0891_ _0892_ _0138_ _0893_ sg13g2_a21oi_1
XFILLER_0_690 VPWR VGND sg13g2_fill_1
XFILLER_39_149 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
X_2022_ _0691_ net154 _0690_ VPWR VGND sg13g2_nand2_1
X_1806_ state\[78\] daisychain\[78\] net151 _0518_ VPWR VGND sg13g2_mux2_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
X_1737_ _0463_ net175 _0462_ VPWR VGND sg13g2_nand2_1
X_1668_ VGND VPWR net117 daisychain\[49\] _0408_ net58 sg13g2_a21oi_1
X_1599_ net190 VPWR _0997_ VGND daisychain\[36\] net35 sg13g2_o21ai_1
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_14_506 VPWR VGND sg13g2_decap_4
XFILLER_26_377 VPWR VGND sg13g2_fill_1
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_10_756 VPWR VGND sg13g2_decap_8
XFILLER_10_789 VPWR VGND sg13g2_decap_8
XFILLER_14_98 VPWR VGND sg13g2_decap_8
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_5_237 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_51 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_29_171 VPWR VGND sg13g2_decap_8
XFILLER_33_804 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
XFILLER_45_620 VPWR VGND sg13g2_decap_8
XFILLER_13_594 VPWR VGND sg13g2_decap_4
XFILLER_5_760 VPWR VGND sg13g2_decap_8
X_1453_ VGND VPWR net101 daisychain\[6\] _0880_ net50 sg13g2_a21oi_1
X_1522_ _0935_ net161 _0934_ VPWR VGND sg13g2_nand2_1
XFILLER_27_119 VPWR VGND sg13g2_decap_8
XFILLER_36_642 VPWR VGND sg13g2_decap_8
X_1384_ VPWR _0048_ state\[28\] VGND sg13g2_inv_1
X_2317__317 VPWR VGND net316 sg13g2_tiehi
X_2005_ VGND VPWR _0675_ _0676_ _0245_ _0677_ sg13g2_a21oi_1
XFILLER_35_196 VPWR VGND sg13g2_decap_8
X_2838_ state\[126\] net13 VPWR VGND sg13g2_buf_1
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_26_141 VPWR VGND sg13g2_decap_8
XFILLER_42_601 VPWR VGND sg13g2_fill_1
XFILLER_10_520 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
X_2368__215 VPWR VGND net214 sg13g2_tiehi
XFILLER_10_597 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_2_13 VPWR VGND sg13g2_decap_8
XFILLER_2_24 VPWR VGND sg13g2_fill_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_17_141 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_fill_1
XFILLER_20_328 VPWR VGND sg13g2_fill_2
XFILLER_20_339 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_decap_4
XFILLER_9_351 VPWR VGND sg13g2_decap_8
X_2554_ net277 VGND VPWR _0370_ state\[114\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1367_ VPWR _0067_ state\[45\] VGND sg13g2_inv_1
X_1436_ state\[4\] daisychain\[4\] net141 _0866_ VPWR VGND sg13g2_mux2_1
X_1505_ VGND VPWR _0919_ _0920_ _0145_ _0921_ sg13g2_a21oi_1
X_2485_ net403 VGND VPWR _0301_ state\[45\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1298_ VPWR _0016_ state\[114\] VGND sg13g2_inv_1
XFILLER_11_306 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_3_527 VPWR VGND sg13g2_fill_1
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_14_133 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_42_420 VPWR VGND sg13g2_decap_8
XFILLER_6_365 VPWR VGND sg13g2_decap_8
XFILLER_7_800 VPWR VGND sg13g2_fill_1
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_2270_ _0825_ net108 state\[107\] VPWR VGND sg13g2_nand2_1
XFILLER_18_450 VPWR VGND sg13g2_decap_8
XFILLER_18_483 VPWR VGND sg13g2_decap_4
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_38_759 VPWR VGND sg13g2_fill_1
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_46_781 VPWR VGND sg13g2_fill_1
XFILLER_46_792 VPWR VGND sg13g2_fill_2
XFILLER_20_103 VPWR VGND sg13g2_decap_8
XFILLER_33_431 VPWR VGND sg13g2_decap_8
X_1985_ VGND VPWR _0659_ _0660_ _0241_ _0661_ sg13g2_a21oi_1
X_2537_ net317 VGND VPWR _0353_ state\[97\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_214 VPWR VGND sg13g2_decap_8
X_1419_ net180 VPWR _0853_ VGND daisychain\[0\] net24 sg13g2_o21ai_1
X_2468_ net215 VGND VPWR _0284_ state\[28\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2399_ net408 VGND VPWR _0215_ daisychain\[87\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_11_103 VPWR VGND sg13g2_decap_8
XFILLER_12_626 VPWR VGND sg13g2_fill_1
XFILLER_24_475 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_37_781 VPWR VGND sg13g2_fill_2
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_20_681 VPWR VGND sg13g2_fill_1
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_3_357 VPWR VGND sg13g2_decap_8
XFILLER_19_225 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
Xfanout160 net163 net160 VPWR VGND sg13g2_buf_1
Xfanout171 net176 net171 VPWR VGND sg13g2_buf_1
Xfanout182 net185 net182 VPWR VGND sg13g2_buf_1
Xfanout193 net198 net193 VPWR VGND sg13g2_buf_1
XFILLER_30_478 VPWR VGND sg13g2_decap_4
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
X_1770_ VGND VPWR _0487_ _0488_ _0198_ _0489_ sg13g2_a21oi_1
XFILLER_6_162 VPWR VGND sg13g2_decap_8
X_2424__359 VPWR VGND net358 sg13g2_tiehi
X_2322_ net306 VGND VPWR _0138_ daisychain\[10\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2253_ VGND VPWR _0599_ _0816_ _0354_ net78 sg13g2_a21oi_1
X_2184_ _0782_ net130 state\[64\] VPWR VGND sg13g2_nand2_1
XFILLER_19_792 VPWR VGND sg13g2_decap_8
XFILLER_21_412 VPWR VGND sg13g2_fill_1
XFILLER_34_773 VPWR VGND sg13g2_fill_1
XFILLER_34_784 VPWR VGND sg13g2_fill_2
Xdigitalen.g\[0\].u.inv1 VPWR digitalen.g\[0\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_21_489 VPWR VGND sg13g2_decap_8
X_2481__420 VPWR VGND net419 sg13g2_tiehi
X_1968_ VGND VPWR net109 daisychain\[109\] _0648_ net56 sg13g2_a21oi_1
X_1899_ net188 VPWR _0593_ VGND daisychain\[96\] net33 sg13g2_o21ai_1
XFILLER_29_523 VPWR VGND sg13g2_decap_8
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_44_559 VPWR VGND sg13g2_fill_2
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_4_611 VPWR VGND sg13g2_fill_2
X_2562__230 VPWR VGND net229 sg13g2_tiehi
XFILLER_12_8 VPWR VGND sg13g2_fill_1
XFILLER_15_261 VPWR VGND sg13g2_decap_8
XFILLER_16_773 VPWR VGND sg13g2_fill_1
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_30_242 VPWR VGND sg13g2_decap_8
XFILLER_31_776 VPWR VGND sg13g2_decap_8
X_1822_ _0531_ net173 _0530_ VPWR VGND sg13g2_nand2_1
X_1753_ VGND VPWR net128 daisychain\[66\] _0476_ net63 sg13g2_a21oi_1
X_1684_ net192 VPWR _0421_ VGND daisychain\[53\] net37 sg13g2_o21ai_1
XFILLER_38_364 VPWR VGND sg13g2_decap_8
X_2305_ VGND VPWR _0703_ _0842_ _0380_ net70 sg13g2_a21oi_1
X_2236_ _0808_ net124 state\[90\] VPWR VGND sg13g2_nand2_1
X_2167_ VGND VPWR _0427_ _0773_ _0311_ net81 sg13g2_a21oi_1
XFILLER_21_220 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_461 VPWR VGND uio_oe[6] sg13g2_tiehi
X_2098_ _0739_ net104 state\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_21_297 VPWR VGND sg13g2_fill_1
XFILLER_5_419 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_29_320 VPWR VGND sg13g2_decap_8
XFILLER_49_629 VPWR VGND sg13g2_decap_8
XFILLER_13_710 VPWR VGND sg13g2_fill_2
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_29_331 VPWR VGND sg13g2_fill_1
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
X_2377__453 VPWR VGND net452 sg13g2_tiehi
XFILLER_12_253 VPWR VGND sg13g2_decap_8
XFILLER_13_765 VPWR VGND sg13g2_decap_4
XFILLER_40_584 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
X_2564__358 VPWR VGND net357 sg13g2_tiehi
XFILLER_4_430 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_36_802 VPWR VGND sg13g2_decap_8
XFILLER_39_128 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_48_695 VPWR VGND sg13g2_decap_8
X_2021_ state\[121\] daisychain\[121\] net136 _0690_ VPWR VGND sg13g2_mux2_1
XFILLER_16_592 VPWR VGND sg13g2_decap_4
X_1805_ VGND VPWR _0515_ _0516_ _0205_ _0517_ sg13g2_a21oi_1
X_1736_ state\[64\] daisychain\[64\] net151 _0462_ VPWR VGND sg13g2_mux2_1
X_1667_ _0407_ net170 _0406_ VPWR VGND sg13g2_nand2_1
X_1598_ VGND VPWR net115 daisychain\[35\] _0996_ net57 sg13g2_a21oi_1
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
X_2219_ VGND VPWR _0531_ _0799_ _0337_ net83 sg13g2_a21oi_1
XFILLER_14_22 VPWR VGND sg13g2_fill_2
XFILLER_14_77 VPWR VGND sg13g2_decap_8
XFILLER_6_706 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_5_216 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_29_150 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_fill_2
XFILLER_9_577 VPWR VGND sg13g2_fill_2
X_1383_ VPWR _0049_ state\[29\] VGND sg13g2_inv_1
X_1452_ _0879_ net160 _0878_ VPWR VGND sg13g2_nand2_1
X_1521_ state\[21\] daisychain\[21\] net139 _0934_ VPWR VGND sg13g2_mux2_1
XFILLER_36_676 VPWR VGND sg13g2_fill_2
X_2004_ net181 VPWR _0677_ VGND daisychain\[117\] net25 sg13g2_o21ai_1
XFILLER_35_175 VPWR VGND sg13g2_decap_8
X_2837_ state\[125\] net12 VPWR VGND sg13g2_buf_1
X_1719_ net193 VPWR _0449_ VGND daisychain\[60\] net38 sg13g2_o21ai_1
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_14_315 VPWR VGND sg13g2_fill_2
XFILLER_14_337 VPWR VGND sg13g2_fill_1
XFILLER_14_348 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_26_197 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_10_565 VPWR VGND sg13g2_fill_1
XFILLER_10_576 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_6_525 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_17_120 VPWR VGND sg13g2_decap_8
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_17_197 VPWR VGND sg13g2_decap_8
XFILLER_32_123 VPWR VGND sg13g2_decap_8
XFILLER_9_330 VPWR VGND sg13g2_decap_8
X_1504_ net182 VPWR _0921_ VGND daisychain\[17\] net27 sg13g2_o21ai_1
X_2553_ net309 VGND VPWR _0369_ state\[113\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1366_ VPWR _0068_ state\[46\] VGND sg13g2_inv_1
X_1435_ VGND VPWR _0863_ _0864_ _0131_ _0865_ sg13g2_a21oi_1
X_2484_ net407 VGND VPWR _0300_ state\[44\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_23_123 VPWR VGND sg13g2_decap_8
X_1297_ VPWR _0017_ state\[115\] VGND sg13g2_inv_1
X_2434__339 VPWR VGND net338 sg13g2_tiehi
XFILLER_11_45 VPWR VGND sg13g2_decap_4
XFILLER_11_89 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_14_112 VPWR VGND sg13g2_decap_8
XFILLER_14_189 VPWR VGND sg13g2_decap_8
XFILLER_15_635 VPWR VGND sg13g2_fill_2
XFILLER_27_495 VPWR VGND sg13g2_fill_1
XFILLER_30_605 VPWR VGND sg13g2_fill_1
XFILLER_42_476 VPWR VGND sg13g2_fill_2
XFILLER_10_384 VPWR VGND sg13g2_fill_2
XFILLER_6_344 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_14_690 VPWR VGND sg13g2_fill_1
XFILLER_20_159 VPWR VGND sg13g2_decap_8
XFILLER_33_465 VPWR VGND sg13g2_decap_4
X_1984_ net186 VPWR _0661_ VGND daisychain\[113\] net31 sg13g2_o21ai_1
X_2536_ net329 VGND VPWR _0352_ state\[96\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2467_ net219 VGND VPWR _0283_ state\[27\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_44_708 VPWR VGND sg13g2_decap_8
XFILLER_44_719 VPWR VGND sg13g2_fill_1
X_1349_ VPWR _0087_ state\[63\] VGND sg13g2_inv_1
X_1418_ VGND VPWR net97 net2 _0852_ net47 sg13g2_a21oi_1
X_2398_ net410 VGND VPWR _0214_ daisychain\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_24_454 VPWR VGND sg13g2_decap_8
XFILLER_37_793 VPWR VGND sg13g2_fill_2
XFILLER_11_159 VPWR VGND sg13g2_decap_8
XFILLER_20_660 VPWR VGND sg13g2_fill_1
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_3_336 VPWR VGND sg13g2_decap_8
XFILLER_4_804 VPWR VGND sg13g2_fill_1
XFILLER_19_204 VPWR VGND sg13g2_decap_8
Xfanout150 net151 net150 VPWR VGND sg13g2_buf_1
Xfanout161 net163 net161 VPWR VGND sg13g2_buf_1
Xfanout172 net173 net172 VPWR VGND sg13g2_buf_1
Xfanout183 net184 net183 VPWR VGND sg13g2_buf_1
XFILLER_27_292 VPWR VGND sg13g2_decap_8
XFILLER_35_708 VPWR VGND sg13g2_fill_1
XFILLER_47_63 VPWR VGND sg13g2_decap_8
Xfanout194 net197 net194 VPWR VGND sg13g2_buf_1
XFILLER_11_671 VPWR VGND sg13g2_decap_8
XFILLER_11_682 VPWR VGND sg13g2_fill_2
XFILLER_15_476 VPWR VGND sg13g2_fill_2
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_fill_1
X_2387__433 VPWR VGND net432 sg13g2_tiehi
XFILLER_10_181 VPWR VGND sg13g2_decap_8
XFILLER_6_141 VPWR VGND sg13g2_decap_8
X_2321_ net308 VGND VPWR _0137_ daisychain\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2252_ _0816_ net112 state\[98\] VPWR VGND sg13g2_nand2_1
X_2183_ VGND VPWR _0459_ _0781_ _0319_ net82 sg13g2_a21oi_1
XFILLER_19_771 VPWR VGND sg13g2_decap_8
XFILLER_25_229 VPWR VGND sg13g2_decap_8
XFILLER_33_284 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[0\].u.inv2 VPWR digitalen.g\[0\].u.OUTP digitalen.g\[0\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_21_468 VPWR VGND sg13g2_decap_8
X_1967_ _0647_ net167 _0646_ VPWR VGND sg13g2_nand2_1
X_1898_ VGND VPWR net111 daisychain\[95\] _0592_ net54 sg13g2_a21oi_1
X_2519_ net209 VGND VPWR _0335_ state\[79\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_17_719 VPWR VGND sg13g2_decap_8
XFILLER_17_99 VPWR VGND sg13g2_decap_8
XFILLER_44_505 VPWR VGND sg13g2_fill_2
XFILLER_24_251 VPWR VGND sg13g2_decap_8
XFILLER_33_32 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_fill_1
XFILLER_15_240 VPWR VGND sg13g2_decap_8
XFILLER_30_221 VPWR VGND sg13g2_decap_8
XFILLER_31_744 VPWR VGND sg13g2_decap_8
XFILLER_31_755 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_10_clk clknet_2_0__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_1821_ state\[81\] daisychain\[81\] net148 _0530_ VPWR VGND sg13g2_mux2_1
X_1752_ _0475_ net174 _0474_ VPWR VGND sg13g2_nand2_1
X_1683_ VGND VPWR net119 daisychain\[52\] _0420_ net59 sg13g2_a21oi_1
X_2304_ _0842_ net90 state\[124\] VPWR VGND sg13g2_nand2_1
XFILLER_26_505 VPWR VGND sg13g2_fill_1
XFILLER_38_343 VPWR VGND sg13g2_decap_8
X_2235_ VGND VPWR _0563_ _0807_ _0345_ net84 sg13g2_a21oi_1
X_2166_ _0773_ net119 state\[55\] VPWR VGND sg13g2_nand2_1
X_2097_ VGND VPWR _0931_ _0738_ _0276_ net71 sg13g2_a21oi_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_462 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_310 VPWR VGND sg13g2_fill_1
XFILLER_13_744 VPWR VGND sg13g2_decap_8
XFILLER_17_527 VPWR VGND sg13g2_fill_1
XFILLER_29_387 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_12_232 VPWR VGND sg13g2_decap_8
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_39_107 VPWR VGND sg13g2_decap_8
XFILLER_5_69 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
X_2020_ VGND VPWR _0687_ _0688_ _0248_ _0689_ sg13g2_a21oi_1
XFILLER_23_519 VPWR VGND sg13g2_decap_8
XFILLER_31_552 VPWR VGND sg13g2_decap_8
XFILLER_35_357 VPWR VGND sg13g2_decap_8
XFILLER_35_368 VPWR VGND sg13g2_fill_2
XFILLER_7_291 VPWR VGND sg13g2_decap_8
X_1804_ net195 VPWR _0517_ VGND daisychain\[77\] net40 sg13g2_o21ai_1
X_1735_ VGND VPWR _0459_ _0460_ _0191_ _0461_ sg13g2_a21oi_1
X_1666_ state\[50\] daisychain\[50\] net146 _0406_ VPWR VGND sg13g2_mux2_1
X_1597_ _0995_ net168 _0994_ VPWR VGND sg13g2_nand2_1
XFILLER_38_140 VPWR VGND sg13g2_decap_8
X_2513__258 VPWR VGND net257 sg13g2_tiehi
X_2218_ _0799_ net126 state\[81\] VPWR VGND sg13g2_nand2_1
X_2149_ VGND VPWR _0391_ _0764_ _0302_ net73 sg13g2_a21oi_1
XFILLER_10_736 VPWR VGND sg13g2_fill_1
XFILLER_22_530 VPWR VGND sg13g2_fill_1
X_2413__381 VPWR VGND net380 sg13g2_tiehi
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_30_88 VPWR VGND sg13g2_decap_8
XFILLER_39_86 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_44_154 VPWR VGND sg13g2_decap_8
X_1520_ VGND VPWR _0931_ _0932_ _0148_ _0933_ sg13g2_a21oi_1
XFILLER_4_283 VPWR VGND sg13g2_decap_8
X_1382_ VPWR _0051_ state\[30\] VGND sg13g2_inv_1
X_1451_ state\[7\] daisychain\[7\] net133 _0878_ VPWR VGND sg13g2_mux2_1
XFILLER_35_154 VPWR VGND sg13g2_decap_8
X_2003_ VGND VPWR net94 daisychain\[116\] _0676_ net46 sg13g2_a21oi_1
X_2836_ state\[124\] net11 VPWR VGND sg13g2_buf_1
X_1718_ VGND VPWR net121 daisychain\[59\] _0448_ net60 sg13g2_a21oi_1
X_1649_ net191 VPWR _0393_ VGND daisychain\[46\] net36 sg13g2_o21ai_1
XFILLER_10_511 VPWR VGND sg13g2_fill_1
XFILLER_22_371 VPWR VGND sg13g2_decap_4
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_25_66 VPWR VGND sg13g2_decap_8
XFILLER_25_77 VPWR VGND sg13g2_fill_2
XFILLER_26_176 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_6_504 VPWR VGND sg13g2_decap_8
X_2448__296 VPWR VGND net295 sg13g2_tiehi
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_17_176 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_13_371 VPWR VGND sg13g2_fill_2
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_9_386 VPWR VGND sg13g2_decap_8
XFILLER_5_581 VPWR VGND sg13g2_fill_2
X_1503_ VGND VPWR net99 daisychain\[16\] _0920_ net49 sg13g2_a21oi_1
X_2552_ net333 VGND VPWR _0368_ state\[112\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2483_ net411 VGND VPWR _0299_ state\[43\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1296_ VPWR _0018_ state\[116\] VGND sg13g2_inv_1
X_1365_ VPWR _0069_ state\[47\] VGND sg13g2_inv_1
X_1434_ net180 VPWR _0865_ VGND daisychain\[3\] net24 sg13g2_o21ai_1
X_2397__413 VPWR VGND net412 sg13g2_tiehi
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_3_507 VPWR VGND sg13g2_fill_2
XFILLER_11_68 VPWR VGND sg13g2_decap_8
XFILLER_19_408 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_fill_2
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_11_820 VPWR VGND sg13g2_fill_2
XFILLER_14_168 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_fill_1
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_42_455 VPWR VGND sg13g2_decap_8
XFILLER_10_363 VPWR VGND sg13g2_decap_8
XFILLER_6_323 VPWR VGND sg13g2_decap_8
X_2565__262 VPWR VGND net261 sg13g2_tiehi
XFILLER_2_584 VPWR VGND sg13g2_fill_1
XFILLER_37_238 VPWR VGND sg13g2_decap_8
XFILLER_18_430 VPWR VGND sg13g2_decap_8
XFILLER_46_772 VPWR VGND sg13g2_fill_1
XFILLER_14_680 VPWR VGND sg13g2_decap_4
XFILLER_20_138 VPWR VGND sg13g2_decap_8
XFILLER_9_183 VPWR VGND sg13g2_decap_8
X_1983_ VGND VPWR net95 daisychain\[112\] _0660_ net53 sg13g2_a21oi_1
X_1417_ VGND VPWR _0851_ net3 net158 sg13g2_or2_1
X_2535_ net337 VGND VPWR _0351_ state\[95\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2466_ net223 VGND VPWR _0282_ state\[26\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_28_249 VPWR VGND sg13g2_fill_2
XFILLER_3_91 VPWR VGND sg13g2_decap_8
X_1348_ VPWR _0088_ state\[64\] VGND sg13g2_inv_1
X_2397_ net412 VGND VPWR _0213_ daisychain\[85\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_11_138 VPWR VGND sg13g2_decap_8
XFILLER_7_109 VPWR VGND sg13g2_decap_8
XFILLER_20_694 VPWR VGND sg13g2_fill_1
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_3_315 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_4
XFILLER_47_547 VPWR VGND sg13g2_decap_8
Xfanout140 net153 net140 VPWR VGND sg13g2_buf_1
Xfanout151 net152 net151 VPWR VGND sg13g2_buf_1
Xfanout162 net163 net162 VPWR VGND sg13g2_buf_1
Xfanout173 net176 net173 VPWR VGND sg13g2_buf_1
Xfanout184 net185 net184 VPWR VGND sg13g2_buf_1
Xfanout195 net196 net195 VPWR VGND sg13g2_buf_1
XFILLER_15_455 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_43_742 VPWR VGND sg13g2_fill_1
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_47_558 VPWR VGND sg13g2_fill_1
XFILLER_10_160 VPWR VGND sg13g2_decap_8
XFILLER_6_120 VPWR VGND sg13g2_decap_8
XFILLER_8_47 VPWR VGND sg13g2_fill_2
XFILLER_2_392 VPWR VGND sg13g2_decap_8
XFILLER_6_197 VPWR VGND sg13g2_decap_8
X_2320_ net310 VGND VPWR _0136_ daisychain\[8\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2251_ VGND VPWR _0595_ _0815_ _0353_ net78 sg13g2_a21oi_1
XFILLER_25_208 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ _0781_ net123 state\[63\] VPWR VGND sg13g2_nand2_1
XFILLER_21_436 VPWR VGND sg13g2_fill_2
XFILLER_33_263 VPWR VGND sg13g2_decap_8
XFILLER_34_764 VPWR VGND sg13g2_fill_2
X_1966_ state\[110\] daisychain\[110\] net143 _0646_ VPWR VGND sg13g2_mux2_1
X_1897_ _0591_ net165 _0590_ VPWR VGND sg13g2_nand2_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_2518_ net217 VGND VPWR _0334_ state\[78\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2449_ net291 VGND VPWR _0265_ state\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_16_219 VPWR VGND sg13g2_decap_8
XFILLER_17_78 VPWR VGND sg13g2_decap_8
XFILLER_24_230 VPWR VGND sg13g2_decap_8
X_2516__234 VPWR VGND net233 sg13g2_tiehi
XFILLER_12_436 VPWR VGND sg13g2_decap_8
XFILLER_12_458 VPWR VGND sg13g2_fill_2
XFILLER_24_296 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_decap_8
XFILLER_40_734 VPWR VGND sg13g2_fill_1
XFILLER_40_789 VPWR VGND sg13g2_decap_8
X_2566__390 VPWR VGND net389 sg13g2_tiehi
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_fill_1
X_2423__361 VPWR VGND net360 sg13g2_tiehi
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_15_296 VPWR VGND sg13g2_decap_8
XFILLER_16_753 VPWR VGND sg13g2_decap_4
XFILLER_16_764 VPWR VGND sg13g2_decap_8
XFILLER_30_200 VPWR VGND sg13g2_decap_8
XFILLER_43_583 VPWR VGND sg13g2_fill_2
XFILLER_47_399 VPWR VGND sg13g2_decap_8
X_1820_ VGND VPWR _0527_ _0528_ _0208_ _0529_ sg13g2_a21oi_1
XFILLER_30_277 VPWR VGND sg13g2_fill_2
X_1751_ state\[67\] daisychain\[67\] net150 _0474_ VPWR VGND sg13g2_mux2_1
X_1682_ _0419_ net170 _0418_ VPWR VGND sg13g2_nand2_1
XFILLER_38_322 VPWR VGND sg13g2_decap_8
X_2303_ VGND VPWR _0699_ _0841_ _0379_ net70 sg13g2_a21oi_1
X_2234_ _0807_ net124 state\[89\] VPWR VGND sg13g2_nand2_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_4
XFILLER_26_517 VPWR VGND sg13g2_decap_8
X_2165_ VGND VPWR _0423_ _0772_ _0310_ net81 sg13g2_a21oi_1
X_2096_ _0738_ net100 state\[20\] VPWR VGND sg13g2_nand2_1
XFILLER_21_255 VPWR VGND sg13g2_decap_8
X_1949_ net186 VPWR _0633_ VGND daisychain\[106\] net31 sg13g2_o21ai_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_29_355 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_12_211 VPWR VGND sg13g2_decap_8
XFILLER_13_701 VPWR VGND sg13g2_fill_1
XFILLER_13_712 VPWR VGND sg13g2_fill_1
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_9_716 VPWR VGND sg13g2_fill_1
XFILLER_12_288 VPWR VGND sg13g2_decap_8
XFILLER_9_738 VPWR VGND sg13g2_decap_4
XFILLER_5_48 VPWR VGND sg13g2_fill_2
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
X_1803_ VGND VPWR net127 daisychain\[76\] _0516_ net63 sg13g2_a21oi_1
XFILLER_7_270 VPWR VGND sg13g2_decap_8
X_1734_ net193 VPWR _0461_ VGND daisychain\[63\] net38 sg13g2_o21ai_1
X_1665_ VGND VPWR _0403_ _0404_ _0177_ _0405_ sg13g2_a21oi_1
X_1596_ state\[36\] daisychain\[36\] net144 _0994_ VPWR VGND sg13g2_mux2_1
XFILLER_26_303 VPWR VGND sg13g2_fill_2
XFILLER_39_675 VPWR VGND sg13g2_fill_2
X_2217_ VGND VPWR _0527_ _0798_ _0336_ net83 sg13g2_a21oi_1
XFILLER_14_24 VPWR VGND sg13g2_fill_1
XFILLER_14_35 VPWR VGND sg13g2_fill_2
XFILLER_38_196 VPWR VGND sg13g2_decap_8
X_2148_ _0764_ net117 state\[46\] VPWR VGND sg13g2_nand2_1
X_2079_ VGND VPWR _0895_ _0729_ _0267_ net68 sg13g2_a21oi_1
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_30_67 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_39_32 VPWR VGND sg13g2_fill_1
XFILLER_39_65 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_17_325 VPWR VGND sg13g2_decap_8
XFILLER_17_336 VPWR VGND sg13g2_fill_2
XFILLER_29_185 VPWR VGND sg13g2_decap_8
XFILLER_33_818 VPWR VGND sg13g2_decap_4
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_9_546 VPWR VGND sg13g2_decap_8
XFILLER_4_262 VPWR VGND sg13g2_decap_8
X_1450_ VGND VPWR _0875_ _0876_ _0134_ _0877_ sg13g2_a21oi_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
X_1381_ VPWR _0052_ state\[31\] VGND sg13g2_inv_1
XFILLER_16_380 VPWR VGND sg13g2_fill_1
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_36_678 VPWR VGND sg13g2_fill_1
XFILLER_48_483 VPWR VGND sg13g2_decap_8
X_2002_ _0675_ net157 _0674_ VPWR VGND sg13g2_nand2_1
X_2835_ state\[123\] net10 VPWR VGND sg13g2_buf_1
X_1717_ _0447_ net171 _0446_ VPWR VGND sg13g2_nand2_1
X_1648_ VGND VPWR net117 daisychain\[45\] _0392_ net58 sg13g2_a21oi_1
X_1579_ net184 VPWR _0981_ VGND daisychain\[32\] net29 sg13g2_o21ai_1
XFILLER_26_111 VPWR VGND sg13g2_decap_8
XFILLER_26_122 VPWR VGND sg13g2_fill_1
XFILLER_26_155 VPWR VGND sg13g2_decap_8
XFILLER_14_328 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_6_549 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_17_155 VPWR VGND sg13g2_decap_8
XFILLER_18_667 VPWR VGND sg13g2_fill_1
XFILLER_45_420 VPWR VGND sg13g2_decap_8
X_2455__268 VPWR VGND net267 sg13g2_tiehi
XFILLER_32_158 VPWR VGND sg13g2_decap_8
XFILLER_9_365 VPWR VGND sg13g2_decap_8
X_1433_ VGND VPWR net94 daisychain\[2\] _0864_ net46 sg13g2_a21oi_1
X_1502_ _0919_ net159 _0918_ VPWR VGND sg13g2_nand2_1
X_2551_ net349 VGND VPWR _0367_ state\[111\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2482_ net415 VGND VPWR _0298_ state\[42\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_28_409 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
X_1295_ VPWR _0019_ state\[117\] VGND sg13g2_inv_1
X_1364_ VPWR _0070_ state\[48\] VGND sg13g2_inv_1
XFILLER_23_158 VPWR VGND sg13g2_decap_8
X_2519__210 VPWR VGND net209 sg13g2_tiehi
XFILLER_15_637 VPWR VGND sg13g2_fill_1
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_42_434 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_10_342 VPWR VGND sg13g2_decap_8
XFILLER_10_386 VPWR VGND sg13g2_fill_1
XFILLER_14_147 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_fill_1
XFILLER_42_478 VPWR VGND sg13g2_fill_1
XFILLER_6_302 VPWR VGND sg13g2_decap_8
XFILLER_2_574 VPWR VGND sg13g2_fill_1
XFILLER_6_379 VPWR VGND sg13g2_decap_8
XFILLER_18_420 VPWR VGND sg13g2_fill_2
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_20_117 VPWR VGND sg13g2_decap_8
XFILLER_33_445 VPWR VGND sg13g2_decap_4
XFILLER_45_294 VPWR VGND sg13g2_decap_8
X_2433__341 VPWR VGND net340 sg13g2_tiehi
X_1982_ _0659_ net164 _0658_ VPWR VGND sg13g2_nand2_1
XFILLER_9_162 VPWR VGND sg13g2_decap_8
X_2534_ net345 VGND VPWR _0350_ state\[94\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_1347_ VPWR _0089_ state\[65\] VGND sg13g2_inv_1
X_1416_ net158 net3 _0850_ VPWR VGND sg13g2_nor2_1
X_2465_ net227 VGND VPWR _0281_ state\[25\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2396_ net414 VGND VPWR _0212_ daisychain\[84\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_37_795 VPWR VGND sg13g2_fill_1
XFILLER_11_117 VPWR VGND sg13g2_decap_8
XFILLER_20_673 VPWR VGND sg13g2_fill_1
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_24_489 VPWR VGND sg13g2_decap_8
X_2334__283 VPWR VGND net282 sg13g2_tiehi
XFILLER_19_239 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
Xfanout130 net131 net130 VPWR VGND sg13g2_buf_1
Xfanout141 net143 net141 VPWR VGND sg13g2_buf_1
Xfanout152 net153 net152 VPWR VGND sg13g2_buf_1
Xfanout163 net177 net163 VPWR VGND sg13g2_buf_1
Xfanout174 net175 net174 VPWR VGND sg13g2_buf_1
Xfanout185 net199 net185 VPWR VGND sg13g2_buf_1
Xfanout196 net197 net196 VPWR VGND sg13g2_buf_1
XFILLER_15_478 VPWR VGND sg13g2_fill_1
XFILLER_27_283 VPWR VGND sg13g2_fill_1
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_43_754 VPWR VGND sg13g2_decap_8
XFILLER_30_448 VPWR VGND sg13g2_fill_2
XFILLER_6_176 VPWR VGND sg13g2_decap_8
XFILLER_7_666 VPWR VGND sg13g2_decap_8
XFILLER_2_371 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
X_2250_ _0815_ net112 state\[97\] VPWR VGND sg13g2_nand2_1
X_2181_ VGND VPWR _0455_ _0780_ _0318_ net82 sg13g2_a21oi_1
XFILLER_21_426 VPWR VGND sg13g2_fill_2
XFILLER_33_242 VPWR VGND sg13g2_decap_8
X_1965_ VGND VPWR _0643_ _0644_ _0237_ _0645_ sg13g2_a21oi_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_2517_ net225 VGND VPWR _0333_ state\[77\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2522__442 VPWR VGND net441 sg13g2_tiehi
X_1896_ state\[96\] daisychain\[96\] net142 _0590_ VPWR VGND sg13g2_mux2_1
X_2448_ net295 VGND VPWR _0264_ state\[8\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2379_ net448 VGND VPWR _0195_ daisychain\[67\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_0_820 VPWR VGND sg13g2_fill_2
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
X_2534__346 VPWR VGND net345 sg13g2_tiehi
XFILLER_15_275 VPWR VGND sg13g2_decap_8
XFILLER_30_256 VPWR VGND sg13g2_decap_8
XFILLER_31_702 VPWR VGND sg13g2_decap_8
X_1750_ VGND VPWR _0471_ _0472_ _0194_ _0473_ sg13g2_a21oi_1
XFILLER_11_492 VPWR VGND sg13g2_decap_4
XFILLER_7_474 VPWR VGND sg13g2_decap_8
X_1681_ state\[53\] daisychain\[53\] net146 _0418_ VPWR VGND sg13g2_mux2_1
XFILLER_38_301 VPWR VGND sg13g2_decap_8
X_2302_ _0841_ net89 state\[123\] VPWR VGND sg13g2_nand2_1
X_2233_ VGND VPWR _0559_ _0806_ _0344_ net77 sg13g2_a21oi_1
X_2164_ _0772_ net119 state\[54\] VPWR VGND sg13g2_nand2_1
XFILLER_19_570 VPWR VGND sg13g2_decap_8
XFILLER_34_540 VPWR VGND sg13g2_decap_4
XFILLER_34_584 VPWR VGND sg13g2_decap_4
XFILLER_38_378 VPWR VGND sg13g2_decap_4
X_2095_ VGND VPWR _0927_ _0737_ _0275_ net71 sg13g2_a21oi_1
XFILLER_21_234 VPWR VGND sg13g2_decap_8
X_1948_ VGND VPWR net107 daisychain\[105\] _0632_ net53 sg13g2_a21oi_1
X_1879_ net188 VPWR _0577_ VGND daisychain\[92\] net33 sg13g2_o21ai_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_17_518 VPWR VGND sg13g2_fill_2
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_12_267 VPWR VGND sg13g2_decap_8
XFILLER_13_779 VPWR VGND sg13g2_fill_1
XFILLER_40_510 VPWR VGND sg13g2_fill_2
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_40_598 VPWR VGND sg13g2_fill_1
XFILLER_4_444 VPWR VGND sg13g2_decap_8
XFILLER_5_27 VPWR VGND sg13g2_decap_8
XFILLER_5_38 VPWR VGND sg13g2_decap_4
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_10_8 VPWR VGND sg13g2_fill_2
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_36_816 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_8_750 VPWR VGND sg13g2_fill_2
X_1802_ _0515_ net174 _0514_ VPWR VGND sg13g2_nand2_1
X_1733_ VGND VPWR net123 daisychain\[62\] _0460_ net60 sg13g2_a21oi_1
X_1664_ net191 VPWR _0405_ VGND daisychain\[49\] net36 sg13g2_o21ai_1
X_1595_ VGND VPWR _0991_ _0992_ _0163_ _0993_ sg13g2_a21oi_1
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_39_621 VPWR VGND sg13g2_fill_1
XFILLER_39_632 VPWR VGND sg13g2_decap_8
X_2216_ _0798_ net126 state\[80\] VPWR VGND sg13g2_nand2_1
X_2147_ VGND VPWR _0387_ _0763_ _0301_ net80 sg13g2_a21oi_1
XFILLER_22_521 VPWR VGND sg13g2_decap_8
XFILLER_34_392 VPWR VGND sg13g2_decap_8
XFILLER_41_329 VPWR VGND sg13g2_decap_8
X_2078_ _0729_ net93 state\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_10_749 VPWR VGND sg13g2_decap_8
XFILLER_30_46 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_44 VPWR VGND sg13g2_decap_8
XFILLER_29_164 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_45_602 VPWR VGND sg13g2_decap_8
XFILLER_13_532 VPWR VGND sg13g2_decap_8
XFILLER_13_587 VPWR VGND sg13g2_decap_8
XFILLER_13_598 VPWR VGND sg13g2_fill_2
XFILLER_4_241 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_fill_2
X_1380_ VPWR _0053_ state\[32\] VGND sg13g2_inv_1
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
X_2001_ state\[117\] daisychain\[117\] net135 _0674_ VPWR VGND sg13g2_mux2_1
XFILLER_35_189 VPWR VGND sg13g2_decap_8
X_2834_ state\[122\] net9 VPWR VGND sg13g2_buf_1
X_1716_ state\[60\] daisychain\[60\] net147 _0446_ VPWR VGND sg13g2_mux2_1
X_1647_ _0391_ net169 _0390_ VPWR VGND sg13g2_nand2_1
X_1578_ VGND VPWR net106 daisychain\[31\] _0980_ net52 sg13g2_a21oi_1
XFILLER_26_134 VPWR VGND sg13g2_decap_8
XFILLER_22_351 VPWR VGND sg13g2_fill_2
XFILLER_22_384 VPWR VGND sg13g2_fill_2
XFILLER_22_395 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_fill_2
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
X_2344__263 VPWR VGND net262 sg13g2_tiehi
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_17_134 VPWR VGND sg13g2_decap_8
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_fill_2
XFILLER_41_671 VPWR VGND sg13g2_decap_8
XFILLER_9_344 VPWR VGND sg13g2_decap_8
X_2550_ net365 VGND VPWR _0366_ state\[110\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_49_4 VPWR VGND sg13g2_decap_8
XFILLER_5_583 VPWR VGND sg13g2_fill_1
X_1363_ VPWR _0071_ state\[49\] VGND sg13g2_inv_1
X_1432_ _0863_ net155 _0862_ VPWR VGND sg13g2_nand2_1
X_1501_ state\[17\] daisychain\[17\] net137 _0918_ VPWR VGND sg13g2_mux2_1
X_2481_ net419 VGND VPWR _0297_ state\[41\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_421 VPWR VGND sg13g2_fill_1
X_1294_ VPWR _0020_ state\[118\] VGND sg13g2_inv_1
XFILLER_17_690 VPWR VGND sg13g2_fill_1
XFILLER_20_800 VPWR VGND sg13g2_fill_1
XFILLER_20_811 VPWR VGND sg13g2_fill_1
XFILLER_23_137 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[3\].u.inv1 VPWR digitalen.g\[3\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_11_37 VPWR VGND sg13g2_fill_2
X_2560__342 VPWR VGND net341 sg13g2_tiehi
XFILLER_14_126 VPWR VGND sg13g2_decap_8
XFILLER_27_421 VPWR VGND sg13g2_fill_2
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_10_321 VPWR VGND sg13g2_decap_8
XFILLER_11_822 VPWR VGND sg13g2_fill_1
XFILLER_6_358 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_fill_2
XFILLER_18_410 VPWR VGND sg13g2_fill_2
XFILLER_18_443 VPWR VGND sg13g2_decap_8
XFILLER_38_708 VPWR VGND sg13g2_decap_4
XFILLER_46_752 VPWR VGND sg13g2_fill_2
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_9_141 VPWR VGND sg13g2_decap_8
X_1981_ state\[113\] daisychain\[113\] net135 _0658_ VPWR VGND sg13g2_mux2_1
XFILLER_5_391 VPWR VGND sg13g2_decap_8
X_2533_ net353 VGND VPWR _0349_ state\[93\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_28_207 VPWR VGND sg13g2_decap_8
X_1346_ VPWR _0090_ state\[66\] VGND sg13g2_inv_1
X_1415_ _0849_ net156 _0848_ VPWR VGND sg13g2_nand2_1
X_2464_ net231 VGND VPWR _0280_ state\[24\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2395_ net416 VGND VPWR _0211_ daisychain\[83\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_24_468 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_20_652 VPWR VGND sg13g2_fill_1
XFILLER_20_685 VPWR VGND sg13g2_fill_1
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xfanout120 net122 net120 VPWR VGND sg13g2_buf_1
Xfanout131 net132 net131 VPWR VGND sg13g2_buf_1
XFILLER_15_402 VPWR VGND sg13g2_fill_2
XFILLER_19_218 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
Xfanout142 net143 net142 VPWR VGND sg13g2_buf_1
Xfanout153 net5 net153 VPWR VGND sg13g2_buf_1
Xfanout164 net167 net164 VPWR VGND sg13g2_buf_1
Xfanout175 net176 net175 VPWR VGND sg13g2_buf_1
Xfanout186 net189 net186 VPWR VGND sg13g2_buf_1
Xfanout197 net198 net197 VPWR VGND sg13g2_buf_1
XFILLER_27_273 VPWR VGND sg13g2_fill_1
XFILLER_30_416 VPWR VGND sg13g2_decap_4
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_10_195 VPWR VGND sg13g2_decap_8
XFILLER_6_155 VPWR VGND sg13g2_decap_8
XFILLER_7_601 VPWR VGND sg13g2_decap_4
XFILLER_2_350 VPWR VGND sg13g2_decap_8
X_2180_ _0780_ net123 state\[62\] VPWR VGND sg13g2_nand2_1
XFILLER_18_295 VPWR VGND sg13g2_decap_8
XFILLER_19_785 VPWR VGND sg13g2_decap_8
XFILLER_33_221 VPWR VGND sg13g2_decap_8
XFILLER_34_766 VPWR VGND sg13g2_fill_1
XFILLER_46_582 VPWR VGND sg13g2_fill_2
XFILLER_46_593 VPWR VGND sg13g2_decap_8
XFILLER_21_438 VPWR VGND sg13g2_fill_1
XFILLER_33_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_1964_ net189 VPWR _0645_ VGND daisychain\[109\] net34 sg13g2_o21ai_1
X_1895_ VGND VPWR _0587_ _0588_ _0223_ _0589_ sg13g2_a21oi_1
X_2516_ net233 VGND VPWR _0332_ state\[76\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2447_ net299 VGND VPWR _0263_ state\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1329_ VPWR _0109_ state\[83\] VGND sg13g2_inv_1
X_2378_ net450 VGND VPWR _0194_ daisychain\[66\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_24_265 VPWR VGND sg13g2_decap_4
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_37_593 VPWR VGND sg13g2_fill_2
XFILLER_20_493 VPWR VGND sg13g2_decap_4
XFILLER_4_604 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_16_722 VPWR VGND sg13g2_decap_4
XFILLER_35_519 VPWR VGND sg13g2_fill_2
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_15_254 VPWR VGND sg13g2_decap_8
XFILLER_30_235 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_fill_2
XFILLER_31_725 VPWR VGND sg13g2_fill_1
XFILLER_31_769 VPWR VGND sg13g2_decap_8
XFILLER_43_585 VPWR VGND sg13g2_fill_1
X_2402__403 VPWR VGND net402 sg13g2_tiehi
X_2301_ VGND VPWR _0695_ _0840_ _0378_ net70 sg13g2_a21oi_1
X_1680_ VGND VPWR _0415_ _0416_ _0180_ _0417_ sg13g2_a21oi_1
XFILLER_31_4 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2232_ _0806_ net113 state\[88\] VPWR VGND sg13g2_nand2_1
X_2163_ VGND VPWR _0419_ _0771_ _0309_ net81 sg13g2_a21oi_1
XFILLER_21_213 VPWR VGND sg13g2_decap_8
X_2094_ _0737_ net100 state\[19\] VPWR VGND sg13g2_nand2_1
XFILLER_9_92 VPWR VGND sg13g2_decap_8
X_1947_ _0631_ net164 _0630_ VPWR VGND sg13g2_nand2_1
X_1878_ VGND VPWR net110 daisychain\[91\] _0576_ net62 sg13g2_a21oi_1
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_12_246 VPWR VGND sg13g2_decap_8
XFILLER_13_758 VPWR VGND sg13g2_decap_8
XFILLER_13_769 VPWR VGND sg13g2_fill_2
XFILLER_40_577 VPWR VGND sg13g2_decap_8
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_8
XFILLER_4_467 VPWR VGND sg13g2_decap_4
X_2384__439 VPWR VGND net438 sg13g2_tiehi
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_48_666 VPWR VGND sg13g2_fill_2
X_2458__256 VPWR VGND net255 sg13g2_tiehi
XFILLER_16_596 VPWR VGND sg13g2_fill_1
XFILLER_43_371 VPWR VGND sg13g2_decap_8
X_2354__243 VPWR VGND net242 sg13g2_tiehi
XFILLER_12_780 VPWR VGND sg13g2_fill_1
XFILLER_12_791 VPWR VGND sg13g2_decap_4
X_1801_ state\[77\] daisychain\[77\] net150 _0514_ VPWR VGND sg13g2_mux2_1
X_1732_ _0459_ net171 _0458_ VPWR VGND sg13g2_nand2_1
X_1663_ VGND VPWR net117 daisychain\[48\] _0404_ net58 sg13g2_a21oi_1
X_1594_ net183 VPWR _0993_ VGND daisychain\[35\] net28 sg13g2_o21ai_1
XFILLER_19_390 VPWR VGND sg13g2_decap_8
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_39_677 VPWR VGND sg13g2_fill_1
X_2215_ VGND VPWR _0523_ _0797_ _0335_ net86 sg13g2_a21oi_1
X_2146_ _0763_ net117 state\[45\] VPWR VGND sg13g2_nand2_1
X_2077_ VGND VPWR _0891_ _0728_ _0266_ net68 sg13g2_a21oi_1
XFILLER_14_15 VPWR VGND sg13g2_fill_2
XFILLER_14_37 VPWR VGND sg13g2_fill_1
XFILLER_22_500 VPWR VGND sg13g2_decap_8
XFILLER_34_360 VPWR VGND sg13g2_fill_1
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_30_25 VPWR VGND sg13g2_decap_8
XFILLER_5_209 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_29_143 VPWR VGND sg13g2_decap_8
XFILLER_25_360 VPWR VGND sg13g2_decap_8
XFILLER_25_393 VPWR VGND sg13g2_decap_4
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_4_220 VPWR VGND sg13g2_decap_8
XFILLER_4_297 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
X_2000_ VGND VPWR _0671_ _0672_ _0244_ _0673_ sg13g2_a21oi_1
XFILLER_16_360 VPWR VGND sg13g2_decap_4
XFILLER_23_308 VPWR VGND sg13g2_fill_2
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_44_680 VPWR VGND sg13g2_decap_8
XFILLER_44_691 VPWR VGND sg13g2_fill_1
X_2833_ state\[121\] net8 VPWR VGND sg13g2_buf_1
XFILLER_6_82 VPWR VGND sg13g2_decap_8
X_1715_ VGND VPWR _0443_ _0444_ _0187_ _0445_ sg13g2_a21oi_1
X_1646_ state\[46\] daisychain\[46\] net140 _0390_ VPWR VGND sg13g2_mux2_1
X_1577_ _0979_ net162 _0978_ VPWR VGND sg13g2_nand2_1
XFILLER_14_308 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
X_2129_ VGND VPWR _0995_ _0754_ _0292_ net79 sg13g2_a21oi_1
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_6_518 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_fill_1
XFILLER_17_113 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_32_116 VPWR VGND sg13g2_decap_8
XFILLER_9_323 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
X_1500_ VGND VPWR _0915_ _0916_ _0144_ _0917_ sg13g2_a21oi_1
X_2480_ net423 VGND VPWR _0296_ state\[40\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_49_750 VPWR VGND sg13g2_decap_4
XFILLER_49_761 VPWR VGND sg13g2_fill_1
X_1293_ VPWR _0021_ state\[119\] VGND sg13g2_inv_1
X_1362_ VPWR _0073_ state\[50\] VGND sg13g2_inv_1
X_1431_ state\[3\] daisychain\[3\] net133 _0862_ VPWR VGND sg13g2_mux2_1
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_36_466 VPWR VGND sg13g2_fill_1
XFILLER_31_193 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[3\].u.inv2 VPWR digitalen.g\[3\].u.OUTP digitalen.g\[3\].u.OUTN VGND
+ sg13g2_inv_1
X_2410__387 VPWR VGND net386 sg13g2_tiehi
XFILLER_11_49 VPWR VGND sg13g2_fill_1
X_1629_ net190 VPWR _1021_ VGND daisychain\[42\] net35 sg13g2_o21ai_1
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_39_282 VPWR VGND sg13g2_decap_8
XFILLER_10_300 VPWR VGND sg13g2_decap_8
XFILLER_14_105 VPWR VGND sg13g2_decap_8
XFILLER_15_628 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_fill_2
XFILLER_42_469 VPWR VGND sg13g2_decap_8
X_2489__388 VPWR VGND net387 sg13g2_tiehi
XFILLER_10_377 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_337 VPWR VGND sg13g2_decap_8
XFILLER_7_816 VPWR VGND sg13g2_decap_8
XFILLER_18_400 VPWR VGND sg13g2_fill_1
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_14_650 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_fill_2
XFILLER_41_480 VPWR VGND sg13g2_decap_4
XFILLER_9_120 VPWR VGND sg13g2_decap_8
X_1980_ VGND VPWR _0655_ _0656_ _0240_ _0657_ sg13g2_a21oi_1
XFILLER_5_370 VPWR VGND sg13g2_decap_8
XFILLER_9_197 VPWR VGND sg13g2_decap_8
X_2532_ net361 VGND VPWR _0348_ state\[92\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2463_ net235 VGND VPWR _0279_ state\[23\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1345_ VPWR _0091_ state\[67\] VGND sg13g2_inv_1
X_1414_ state\[0\] daisychain\[0\] net133 _0848_ VPWR VGND sg13g2_mux2_1
X_2394_ net418 VGND VPWR _0210_ daisychain\[82\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_24_447 VPWR VGND sg13g2_decap_8
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_20_631 VPWR VGND sg13g2_fill_1
XFILLER_20_664 VPWR VGND sg13g2_fill_1
XFILLER_32_491 VPWR VGND sg13g2_decap_8
XFILLER_3_329 VPWR VGND sg13g2_decap_8
Xfanout110 net113 net110 VPWR VGND sg13g2_buf_1
Xfanout121 net122 net121 VPWR VGND sg13g2_buf_1
Xfanout132 _0846_ net132 VPWR VGND sg13g2_buf_1
Xfanout143 net153 net143 VPWR VGND sg13g2_buf_1
Xfanout154 net158 net154 VPWR VGND sg13g2_buf_1
Xfanout165 net167 net165 VPWR VGND sg13g2_buf_1
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_27_263 VPWR VGND sg13g2_fill_2
XFILLER_47_56 VPWR VGND sg13g2_decap_8
Xfanout176 net177 net176 VPWR VGND sg13g2_buf_1
Xfanout187 net188 net187 VPWR VGND sg13g2_buf_1
Xfanout198 net199 net198 VPWR VGND sg13g2_buf_1
XFILLER_11_664 VPWR VGND sg13g2_decap_8
XFILLER_15_469 VPWR VGND sg13g2_decap_8
XFILLER_42_266 VPWR VGND sg13g2_decap_8
X_2313__325 VPWR VGND net324 sg13g2_tiehi
XFILLER_10_174 VPWR VGND sg13g2_decap_8
XFILLER_12_92 VPWR VGND sg13g2_decap_8
XFILLER_6_134 VPWR VGND sg13g2_decap_8
X_2394__419 VPWR VGND net418 sg13g2_tiehi
XFILLER_18_263 VPWR VGND sg13g2_decap_4
XFILLER_18_285 VPWR VGND sg13g2_fill_1
XFILLER_19_753 VPWR VGND sg13g2_decap_8
XFILLER_19_764 VPWR VGND sg13g2_decap_8
XFILLER_33_200 VPWR VGND sg13g2_decap_8
XFILLER_33_277 VPWR VGND sg13g2_decap_8
XFILLER_34_701 VPWR VGND sg13g2_fill_2
XFILLER_46_561 VPWR VGND sg13g2_decap_8
X_2364__223 VPWR VGND net222 sg13g2_tiehi
X_1963_ VGND VPWR net109 daisychain\[108\] _0644_ net53 sg13g2_a21oi_1
X_1894_ net187 VPWR _0589_ VGND daisychain\[95\] net32 sg13g2_o21ai_1
X_2515_ net241 VGND VPWR _0331_ state\[75\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2446_ net303 VGND VPWR _0262_ state\[6\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1328_ VPWR _0110_ state\[84\] VGND sg13g2_inv_1
X_2377_ net452 VGND VPWR _0193_ daisychain\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_24_244 VPWR VGND sg13g2_decap_8
XFILLER_33_25 VPWR VGND sg13g2_decap_8
X_2451__284 VPWR VGND net283 sg13g2_tiehi
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_0_822 VPWR VGND sg13g2_fill_1
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_15_233 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_fill_2
XFILLER_11_472 VPWR VGND sg13g2_decap_4
XFILLER_30_214 VPWR VGND sg13g2_decap_8
XFILLER_31_737 VPWR VGND sg13g2_decap_8
XFILLER_7_410 VPWR VGND sg13g2_decap_8
X_2300_ _0840_ net89 state\[122\] VPWR VGND sg13g2_nand2_1
X_2231_ VGND VPWR _0555_ _0805_ _0343_ net77 sg13g2_a21oi_1
XFILLER_24_4 VPWR VGND sg13g2_decap_4
XFILLER_38_336 VPWR VGND sg13g2_decap_8
X_2162_ _0771_ net119 state\[53\] VPWR VGND sg13g2_nand2_1
X_2093_ VGND VPWR _0923_ _0736_ _0274_ net71 sg13g2_a21oi_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_fill_1
XFILLER_9_71 VPWR VGND sg13g2_decap_8
XFILLER_30_781 VPWR VGND sg13g2_fill_1
X_1946_ state\[106\] daisychain\[106\] net141 _0630_ VPWR VGND sg13g2_mux2_1
X_1877_ _0575_ net173 _0574_ VPWR VGND sg13g2_nand2_1
XFILLER_28_25 VPWR VGND sg13g2_decap_8
X_2429_ net348 VGND VPWR _0245_ daisychain\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_37_391 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_12_225 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_16_553 VPWR VGND sg13g2_fill_2
XFILLER_31_545 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
X_1800_ VGND VPWR _0511_ _0512_ _0204_ _0513_ sg13g2_a21oi_1
XFILLER_7_284 VPWR VGND sg13g2_decap_8
XFILLER_8_763 VPWR VGND sg13g2_fill_2
X_2465__228 VPWR VGND net227 sg13g2_tiehi
X_1731_ state\[63\] daisychain\[63\] net147 _0458_ VPWR VGND sg13g2_mux2_1
X_1662_ _0403_ net169 _0402_ VPWR VGND sg13g2_nand2_1
X_2214_ _0797_ net130 state\[79\] VPWR VGND sg13g2_nand2_1
X_1593_ VGND VPWR net105 daisychain\[34\] _0992_ net51 sg13g2_a21oi_1
XFILLER_26_339 VPWR VGND sg13g2_decap_8
XFILLER_34_350 VPWR VGND sg13g2_fill_1
XFILLER_38_133 VPWR VGND sg13g2_decap_8
X_2145_ VGND VPWR _1027_ _0762_ _0300_ net79 sg13g2_a21oi_1
X_2076_ _0728_ net91 state\[10\] VPWR VGND sg13g2_nand2_1
X_1929_ net188 VPWR _0617_ VGND daisychain\[102\] net33 sg13g2_o21ai_1
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_29_122 VPWR VGND sg13g2_decap_8
XFILLER_39_79 VPWR VGND sg13g2_decap_8
X_2420__367 VPWR VGND net366 sg13g2_tiehi
XFILLER_29_199 VPWR VGND sg13g2_decap_8
XFILLER_32_309 VPWR VGND sg13g2_fill_2
XFILLER_41_821 VPWR VGND sg13g2_fill_2
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_755 VPWR VGND sg13g2_fill_1
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_4_276 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
X_2832_ state\[120\] net7 VPWR VGND sg13g2_buf_1
XFILLER_6_61 VPWR VGND sg13g2_decap_8
X_1714_ net193 VPWR _0445_ VGND daisychain\[59\] net38 sg13g2_o21ai_1
X_1645_ VGND VPWR _0387_ _0388_ _0173_ _0389_ sg13g2_a21oi_1
X_1576_ state\[32\] daisychain\[32\] net140 _0978_ VPWR VGND sg13g2_mux2_1
XFILLER_25_48 VPWR VGND sg13g2_fill_1
XFILLER_25_59 VPWR VGND sg13g2_decap_8
XFILLER_26_169 VPWR VGND sg13g2_decap_8
XFILLER_42_618 VPWR VGND sg13g2_decap_8
X_2128_ _0754_ net115 state\[36\] VPWR VGND sg13g2_nand2_1
X_2059_ VGND VPWR _0855_ _0719_ _0257_ net68 sg13g2_a21oi_1
XFILLER_22_353 VPWR VGND sg13g2_fill_1
XFILLER_22_364 VPWR VGND sg13g2_decap_8
XFILLER_22_386 VPWR VGND sg13g2_fill_1
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_17_169 VPWR VGND sg13g2_decap_8
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_25_180 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_302 VPWR VGND sg13g2_decap_8
XFILLER_5_574 VPWR VGND sg13g2_decap_8
XFILLER_9_379 VPWR VGND sg13g2_decap_8
X_1430_ VGND VPWR _0859_ _0860_ _0130_ _0861_ sg13g2_a21oi_1
X_2323__305 VPWR VGND net304 sg13g2_tiehi
XFILLER_49_773 VPWR VGND sg13g2_decap_4
X_1292_ VPWR _0023_ state\[120\] VGND sg13g2_inv_1
X_1361_ VPWR _0074_ state\[51\] VGND sg13g2_inv_1
XFILLER_16_191 VPWR VGND sg13g2_decap_8
XFILLER_36_456 VPWR VGND sg13g2_decap_4
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_fill_1
XFILLER_31_172 VPWR VGND sg13g2_decap_8
X_1559_ net185 VPWR _0965_ VGND daisychain\[28\] net30 sg13g2_o21ai_1
X_1628_ VGND VPWR net116 daisychain\[41\] _1020_ net57 sg13g2_a21oi_1
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_39_261 VPWR VGND sg13g2_decap_8
X_2374__203 VPWR VGND net202 sg13g2_tiehi
XFILLER_11_813 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_42_448 VPWR VGND sg13g2_decap_8
XFILLER_10_356 VPWR VGND sg13g2_decap_8
XFILLER_6_316 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_46_765 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_decap_8
XFILLER_14_673 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_fill_1
XFILLER_9_176 VPWR VGND sg13g2_decap_8
X_1413_ VPWR _0847_ net178 VGND sg13g2_inv_1
X_2531_ net369 VGND VPWR _0347_ state\[91\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2462_ net239 VGND VPWR _0278_ state\[22\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2393_ net420 VGND VPWR _0209_ daisychain\[81\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_36_231 VPWR VGND sg13g2_decap_8
XFILLER_37_765 VPWR VGND sg13g2_decap_4
XFILLER_3_84 VPWR VGND sg13g2_decap_8
X_1344_ VPWR _0092_ state\[68\] VGND sg13g2_inv_1
XFILLER_20_643 VPWR VGND sg13g2_fill_2
XFILLER_20_698 VPWR VGND sg13g2_fill_1
XFILLER_3_308 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
Xfanout100 net103 net100 VPWR VGND sg13g2_buf_1
Xfanout111 net112 net111 VPWR VGND sg13g2_buf_1
Xfanout122 net123 net122 VPWR VGND sg13g2_buf_1
Xfanout133 net135 net133 VPWR VGND sg13g2_buf_1
Xfanout144 net152 net144 VPWR VGND sg13g2_buf_1
Xfanout155 net156 net155 VPWR VGND sg13g2_buf_1
Xfanout166 net167 net166 VPWR VGND sg13g2_buf_1
Xfanout177 net4 net177 VPWR VGND sg13g2_buf_1
Xfanout188 net189 net188 VPWR VGND sg13g2_buf_1
Xfanout199 net1 net199 VPWR VGND sg13g2_buf_1
XFILLER_15_415 VPWR VGND sg13g2_fill_1
XFILLER_27_231 VPWR VGND sg13g2_decap_8
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_43_768 VPWR VGND sg13g2_decap_8
XFILLER_10_153 VPWR VGND sg13g2_decap_8
XFILLER_11_621 VPWR VGND sg13g2_fill_1
XFILLER_11_654 VPWR VGND sg13g2_fill_1
XFILLER_30_407 VPWR VGND sg13g2_fill_1
XFILLER_6_113 VPWR VGND sg13g2_decap_8
XFILLER_12_71 VPWR VGND sg13g2_decap_8
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_19_732 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_decap_8
XFILLER_46_551 VPWR VGND sg13g2_fill_2
XFILLER_14_492 VPWR VGND sg13g2_decap_8
XFILLER_33_256 VPWR VGND sg13g2_decap_8
X_1962_ _0643_ net167 _0642_ VPWR VGND sg13g2_nand2_1
X_1893_ VGND VPWR net111 daisychain\[94\] _0588_ net54 sg13g2_a21oi_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2514_ net249 VGND VPWR _0330_ state\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2445_ net307 VGND VPWR _0261_ state\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2376_ net454 VGND VPWR _0192_ daisychain\[64\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_24_223 VPWR VGND sg13g2_decap_8
X_1327_ VPWR _0111_ state\[85\] VGND sg13g2_inv_1
XFILLER_12_407 VPWR VGND sg13g2_fill_2
XFILLER_12_429 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_15_212 VPWR VGND sg13g2_decap_8
XFILLER_15_289 VPWR VGND sg13g2_decap_8
XFILLER_16_702 VPWR VGND sg13g2_fill_2
XFILLER_16_746 VPWR VGND sg13g2_decap_8
XFILLER_16_757 VPWR VGND sg13g2_fill_2
XFILLER_43_565 VPWR VGND sg13g2_fill_2
XFILLER_43_576 VPWR VGND sg13g2_decap_8
X_2430__347 VPWR VGND net346 sg13g2_tiehi
XFILLER_11_440 VPWR VGND sg13g2_decap_4
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_decap_8
X_2230_ _0805_ net111 state\[87\] VPWR VGND sg13g2_nand2_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_fill_2
XFILLER_19_584 VPWR VGND sg13g2_fill_2
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
X_2161_ VGND VPWR _0415_ _0770_ _0308_ net81 sg13g2_a21oi_1
X_2092_ _0736_ net100 state\[18\] VPWR VGND sg13g2_nand2_1
XFILLER_21_248 VPWR VGND sg13g2_decap_8
XFILLER_30_760 VPWR VGND sg13g2_fill_1
XFILLER_30_793 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_456 VPWR VGND uio_oe[1] sg13g2_tiehi
X_2331__289 VPWR VGND net288 sg13g2_tiehi
X_1945_ VGND VPWR _0627_ _0628_ _0233_ _0629_ sg13g2_a21oi_1
X_1876_ state\[92\] daisychain\[92\] net148 _0574_ VPWR VGND sg13g2_mux2_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_348 VPWR VGND sg13g2_decap_8
X_2428_ net350 VGND VPWR _0244_ daisychain\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2359_ net232 VGND VPWR _0175_ daisychain\[47\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_12_204 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_9_709 VPWR VGND sg13g2_fill_2
XFILLER_40_568 VPWR VGND sg13g2_decap_4
XFILLER_4_458 VPWR VGND sg13g2_decap_4
XFILLER_0_686 VPWR VGND sg13g2_decap_4
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_12_771 VPWR VGND sg13g2_decap_8
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_11_292 VPWR VGND sg13g2_decap_8
XFILLER_7_263 VPWR VGND sg13g2_decap_8
X_1730_ VGND VPWR _0455_ _0456_ _0190_ _0457_ sg13g2_a21oi_1
X_1661_ state\[49\] daisychain\[49\] net145 _0402_ VPWR VGND sg13g2_mux2_1
X_1592_ _0991_ net168 _0990_ VPWR VGND sg13g2_nand2_1
XFILLER_38_112 VPWR VGND sg13g2_decap_8
X_2213_ VGND VPWR _0519_ _0796_ _0334_ net86 sg13g2_a21oi_1
X_2144_ _0762_ net116 state\[44\] VPWR VGND sg13g2_nand2_1
XFILLER_38_189 VPWR VGND sg13g2_decap_8
X_2075_ VGND VPWR _0887_ _0727_ _0265_ net67 sg13g2_a21oi_1
X_2383__441 VPWR VGND net440 sg13g2_tiehi
X_1928_ VGND VPWR net110 daisychain\[101\] _0616_ net55 sg13g2_a21oi_1
X_1859_ net187 VPWR _0561_ VGND daisychain\[88\] net32 sg13g2_o21ai_1
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_29_101 VPWR VGND sg13g2_decap_8
XFILLER_29_178 VPWR VGND sg13g2_decap_8
XFILLER_39_58 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_45_627 VPWR VGND sg13g2_fill_2
XFILLER_13_568 VPWR VGND sg13g2_fill_1
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_9_539 VPWR VGND sg13g2_decap_8
XFILLER_4_255 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_fill_2
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_20_82 VPWR VGND sg13g2_decap_8
XFILLER_29_80 VPWR VGND sg13g2_decap_8
XFILLER_32_822 VPWR VGND sg13g2_fill_1
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_36_605 VPWR VGND sg13g2_fill_2
XFILLER_48_476 VPWR VGND sg13g2_decap_8
X_1713_ VGND VPWR net121 daisychain\[58\] _0444_ net60 sg13g2_a21oi_1
X_1644_ net191 VPWR _0389_ VGND daisychain\[45\] net36 sg13g2_o21ai_1
X_1575_ VGND VPWR _0975_ _0976_ _0159_ _0977_ sg13g2_a21oi_1
XFILLER_26_104 VPWR VGND sg13g2_decap_8
X_2127_ VGND VPWR _0991_ _0753_ _0291_ net79 sg13g2_a21oi_1
XFILLER_26_148 VPWR VGND sg13g2_decap_8
X_2058_ _0719_ net91 state\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_10_527 VPWR VGND sg13g2_fill_2
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_2_726 VPWR VGND sg13g2_decap_4
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_14_822 VPWR VGND sg13g2_fill_1
XFILLER_17_148 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_15_93 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_41_685 VPWR VGND sg13g2_fill_2
XFILLER_9_358 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_decap_8
X_1360_ VPWR _0075_ state\[52\] VGND sg13g2_inv_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_36_413 VPWR VGND sg13g2_fill_2
XFILLER_48_273 VPWR VGND sg13g2_decap_8
X_1291_ VPWR _0024_ state\[121\] VGND sg13g2_inv_1
XFILLER_16_170 VPWR VGND sg13g2_decap_8
XFILLER_31_151 VPWR VGND sg13g2_decap_8
XFILLER_44_490 VPWR VGND sg13g2_decap_4
XFILLER_32_696 VPWR VGND sg13g2_decap_8
X_1489_ net179 VPWR _0909_ VGND daisychain\[14\] net23 sg13g2_o21ai_1
X_1558_ VGND VPWR net101 daisychain\[27\] _0964_ net50 sg13g2_a21oi_1
X_1627_ _1019_ net168 _1018_ VPWR VGND sg13g2_nand2_1
XFILLER_27_402 VPWR VGND sg13g2_decap_8
XFILLER_39_240 VPWR VGND sg13g2_decap_8
XFILLER_42_427 VPWR VGND sg13g2_decap_8
X_2454__272 VPWR VGND net271 sg13g2_tiehi
XFILLER_10_335 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_35_490 VPWR VGND sg13g2_fill_2
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_18_457 VPWR VGND sg13g2_fill_2
XFILLER_33_438 VPWR VGND sg13g2_decap_8
XFILLER_33_449 VPWR VGND sg13g2_fill_2
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_4
XFILLER_42_91 VPWR VGND sg13g2_decap_8
XFILLER_9_155 VPWR VGND sg13g2_decap_8
X_2530_ net377 VGND VPWR _0346_ state\[90\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_3_63 VPWR VGND sg13g2_decap_8
X_1343_ VPWR _0093_ state\[69\] VGND sg13g2_inv_1
X_1412_ VPWR _0000_ state\[0\] VGND sg13g2_inv_1
X_2461_ net243 VGND VPWR _0277_ state\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2440__327 VPWR VGND net326 sg13g2_tiehi
X_2392_ net422 VGND VPWR _0208_ daisychain\[80\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_20_611 VPWR VGND sg13g2_fill_1
XFILLER_22_39 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_2_0__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_20_677 VPWR VGND sg13g2_fill_1
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
Xfanout101 net103 net101 VPWR VGND sg13g2_buf_1
Xfanout112 net113 net112 VPWR VGND sg13g2_buf_1
Xfanout123 net132 net123 VPWR VGND sg13g2_buf_1
Xfanout134 net135 net134 VPWR VGND sg13g2_buf_1
Xfanout145 net152 net145 VPWR VGND sg13g2_buf_1
Xfanout156 net157 net156 VPWR VGND sg13g2_buf_1
Xfanout167 net177 net167 VPWR VGND sg13g2_buf_1
Xfanout178 net199 net178 VPWR VGND sg13g2_buf_1
Xfanout189 net199 net189 VPWR VGND sg13g2_buf_1
X_2341__269 VPWR VGND net268 sg13g2_tiehi
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_43_747 VPWR VGND sg13g2_fill_2
XFILLER_10_132 VPWR VGND sg13g2_decap_8
XFILLER_11_611 VPWR VGND sg13g2_decap_4
XFILLER_11_688 VPWR VGND sg13g2_fill_1
XFILLER_11_699 VPWR VGND sg13g2_fill_2
XFILLER_23_482 VPWR VGND sg13g2_fill_1
XFILLER_23_493 VPWR VGND sg13g2_decap_8
XFILLER_2_364 VPWR VGND sg13g2_decap_8
XFILLER_6_169 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_19_722 VPWR VGND sg13g2_decap_4
XFILLER_34_725 VPWR VGND sg13g2_fill_2
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_33_235 VPWR VGND sg13g2_decap_8
XFILLER_42_780 VPWR VGND sg13g2_fill_1
X_2550__366 VPWR VGND net365 sg13g2_tiehi
X_2468__216 VPWR VGND net215 sg13g2_tiehi
X_1961_ state\[109\] daisychain\[109\] net143 _0642_ VPWR VGND sg13g2_mux2_1
X_1892_ _0587_ net165 _0586_ VPWR VGND sg13g2_nand2_1
X_2513_ net257 VGND VPWR _0329_ state\[73\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_1326_ VPWR _0112_ state\[86\] VGND sg13g2_inv_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2444_ net311 VGND VPWR _0260_ state\[4\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2375_ net200 VGND VPWR _0191_ daisychain\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_12_419 VPWR VGND sg13g2_fill_2
XFILLER_24_202 VPWR VGND sg13g2_decap_8
XFILLER_37_530 VPWR VGND sg13g2_fill_2
XFILLER_37_541 VPWR VGND sg13g2_fill_1
XFILLER_0_813 VPWR VGND sg13g2_decap_8
X_2393__421 VPWR VGND net420 sg13g2_tiehi
XFILLER_15_268 VPWR VGND sg13g2_decap_8
XFILLER_30_249 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_7_456 VPWR VGND sg13g2_fill_2
XFILLER_7_467 VPWR VGND sg13g2_decap_8
X_2545__446 VPWR VGND net445 sg13g2_tiehi
XFILLER_2_161 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_decap_4
X_2160_ _0770_ net120 state\[52\] VPWR VGND sg13g2_nand2_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_596 VPWR VGND sg13g2_decap_8
XFILLER_34_544 VPWR VGND sg13g2_fill_1
XFILLER_34_577 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
X_2091_ VGND VPWR _0919_ _0735_ _0273_ net71 sg13g2_a21oi_1
XFILLER_21_227 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_457 VPWR VGND uio_oe[2] sg13g2_tiehi
X_1944_ net186 VPWR _0629_ VGND daisychain\[105\] net31 sg13g2_o21ai_1
X_1875_ VGND VPWR _0571_ _0572_ _0219_ _0573_ sg13g2_a21oi_1
X_2427_ net352 VGND VPWR _0243_ daisychain\[115\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_29_327 VPWR VGND sg13g2_decap_4
XFILLER_44_308 VPWR VGND sg13g2_decap_8
X_1309_ VPWR _0004_ state\[103\] VGND sg13g2_inv_1
X_2358_ net234 VGND VPWR _0174_ daisychain\[46\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2289_ VGND VPWR _0671_ _0834_ _0372_ net69 sg13g2_a21oi_1
XFILLER_25_511 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_4_437 VPWR VGND sg13g2_decap_8
XFILLER_16_511 VPWR VGND sg13g2_fill_1
XFILLER_16_555 VPWR VGND sg13g2_fill_1
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_36_809 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_11_271 VPWR VGND sg13g2_decap_8
XFILLER_12_750 VPWR VGND sg13g2_decap_8
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_8_765 VPWR VGND sg13g2_fill_1
XFILLER_7_242 VPWR VGND sg13g2_decap_8
X_1660_ VGND VPWR _0399_ _0400_ _0176_ _0401_ sg13g2_a21oi_1
X_1591_ state\[35\] daisychain\[35\] net144 _0990_ VPWR VGND sg13g2_mux2_1
XFILLER_38_168 VPWR VGND sg13g2_decap_8
X_2212_ _0796_ net130 state\[78\] VPWR VGND sg13g2_nand2_1
X_2143_ VGND VPWR _1023_ _0761_ _0299_ net79 sg13g2_a21oi_1
XFILLER_19_360 VPWR VGND sg13g2_fill_2
XFILLER_19_371 VPWR VGND sg13g2_fill_2
XFILLER_22_514 VPWR VGND sg13g2_decap_4
XFILLER_34_341 VPWR VGND sg13g2_decap_8
X_2074_ _0727_ net91 state\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_30_39 VPWR VGND sg13g2_decap_8
X_1927_ _0615_ net165 _0614_ VPWR VGND sg13g2_nand2_1
X_1858_ VGND VPWR net111 daisychain\[87\] _0560_ net54 sg13g2_a21oi_1
XFILLER_39_37 VPWR VGND sg13g2_decap_8
X_1789_ net194 VPWR _0505_ VGND daisychain\[74\] net39 sg13g2_o21ai_1
XFILLER_25_330 VPWR VGND sg13g2_fill_1
XFILLER_29_157 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_9_518 VPWR VGND sg13g2_decap_4
XFILLER_4_234 VPWR VGND sg13g2_decap_8
X_2499__348 VPWR VGND net347 sg13g2_tiehi
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_16_374 VPWR VGND sg13g2_fill_1
XFILLER_17_820 VPWR VGND sg13g2_fill_2
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND state\[123\] sg13g2_antennanp
X_1712_ _0443_ net171 _0442_ VPWR VGND sg13g2_nand2_1
X_1643_ VGND VPWR net115 daisychain\[44\] _0388_ net57 sg13g2_a21oi_1
XFILLER_4_790 VPWR VGND sg13g2_fill_1
X_1574_ net184 VPWR _0977_ VGND daisychain\[31\] net29 sg13g2_o21ai_1
XFILLER_19_190 VPWR VGND sg13g2_decap_8
XFILLER_26_127 VPWR VGND sg13g2_decap_8
X_2126_ _0753_ net115 state\[35\] VPWR VGND sg13g2_nand2_1
X_2057_ VGND VPWR _0849_ _0718_ _0256_ net68 sg13g2_a21oi_1
XFILLER_22_311 VPWR VGND sg13g2_fill_2
XFILLER_22_344 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_34_182 VPWR VGND sg13g2_decap_8
XFILLER_35_672 VPWR VGND sg13g2_fill_2
XFILLER_35_694 VPWR VGND sg13g2_decap_8
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_13_333 VPWR VGND sg13g2_decap_4
XFILLER_17_127 VPWR VGND sg13g2_decap_8
XFILLER_18_628 VPWR VGND sg13g2_fill_2
XFILLER_45_469 VPWR VGND sg13g2_decap_8
X_2351__249 VPWR VGND net248 sg13g2_tiehi
XFILLER_15_72 VPWR VGND sg13g2_decap_8
XFILLER_31_60 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_9_337 VPWR VGND sg13g2_decap_8
XFILLER_1_760 VPWR VGND sg13g2_fill_1
XFILLER_5_554 VPWR VGND sg13g2_fill_1
XFILLER_1_793 VPWR VGND sg13g2_fill_2
XFILLER_48_252 VPWR VGND sg13g2_decap_8
X_1290_ VPWR _0025_ state\[122\] VGND sg13g2_inv_1
XFILLER_17_672 VPWR VGND sg13g2_fill_1
XFILLER_17_683 VPWR VGND sg13g2_decap_8
XFILLER_31_130 VPWR VGND sg13g2_decap_8
X_1626_ state\[42\] daisychain\[42\] net144 _1018_ VPWR VGND sg13g2_mux2_1
X_1488_ VGND VPWR net91 daisychain\[13\] _0908_ net45 sg13g2_a21oi_1
X_1557_ _0963_ net160 _0962_ VPWR VGND sg13g2_nand2_1
XFILLER_14_119 VPWR VGND sg13g2_decap_8
XFILLER_27_414 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_39_296 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
X_2109_ VGND VPWR _0955_ _0744_ _0282_ net71 sg13g2_a21oi_1
XFILLER_10_314 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_decap_4
X_2461__244 VPWR VGND net243 sg13g2_tiehi
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_14_620 VPWR VGND sg13g2_decap_8
XFILLER_14_664 VPWR VGND sg13g2_decap_4
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_9_134 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
X_2460_ net247 VGND VPWR _0276_ state\[20\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_3_31 VPWR VGND sg13g2_fill_2
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_5_384 VPWR VGND sg13g2_decap_8
X_1342_ VPWR _0095_ state\[70\] VGND sg13g2_inv_1
X_1411_ VPWR _0039_ state\[1\] VGND sg13g2_inv_1
X_2391_ net424 VGND VPWR _0207_ daisychain\[79\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_20_601 VPWR VGND sg13g2_fill_2
XFILLER_20_623 VPWR VGND sg13g2_fill_1
XFILLER_20_656 VPWR VGND sg13g2_fill_1
XFILLER_20_689 VPWR VGND sg13g2_fill_2
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_32_483 VPWR VGND sg13g2_decap_4
Xfanout102 net103 net102 VPWR VGND sg13g2_buf_1
Xfanout113 net114 net113 VPWR VGND sg13g2_buf_1
X_1609_ net184 VPWR _1005_ VGND daisychain\[38\] net29 sg13g2_o21ai_1
Xfanout124 net131 net124 VPWR VGND sg13g2_buf_1
Xfanout135 net153 net135 VPWR VGND sg13g2_buf_1
Xfanout146 net147 net146 VPWR VGND sg13g2_buf_1
Xfanout157 net158 net157 VPWR VGND sg13g2_buf_1
Xfanout168 net176 net168 VPWR VGND sg13g2_buf_1
Xfanout179 net181 net179 VPWR VGND sg13g2_buf_1
XFILLER_27_299 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_43_704 VPWR VGND sg13g2_decap_4
XFILLER_10_111 VPWR VGND sg13g2_decap_8
XFILLER_10_188 VPWR VGND sg13g2_decap_8
XFILLER_11_678 VPWR VGND sg13g2_decap_4
XFILLER_6_148 VPWR VGND sg13g2_decap_8
XFILLER_7_605 VPWR VGND sg13g2_fill_2
XFILLER_2_343 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_19_778 VPWR VGND sg13g2_decap_8
XFILLER_33_214 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_46_575 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
X_1960_ VGND VPWR _0639_ _0640_ _0236_ _0641_ sg13g2_a21oi_1
X_1891_ state\[95\] daisychain\[95\] net142 _0586_ VPWR VGND sg13g2_mux2_1
XFILLER_5_181 VPWR VGND sg13g2_decap_8
X_2512_ net265 VGND VPWR _0328_ state\[72\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2443_ net315 VGND VPWR _0259_ state\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1325_ VPWR _0113_ state\[87\] VGND sg13g2_inv_1
X_2374_ net202 VGND VPWR _0190_ daisychain\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_12_409 VPWR VGND sg13g2_fill_1
XFILLER_24_258 VPWR VGND sg13g2_decap_8
XFILLER_24_269 VPWR VGND sg13g2_fill_1
XFILLER_33_39 VPWR VGND sg13g2_decap_8
XFILLER_37_586 VPWR VGND sg13g2_decap_8
XFILLER_20_486 VPWR VGND sg13g2_decap_8
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_16_715 VPWR VGND sg13g2_decap_8
XFILLER_15_247 VPWR VGND sg13g2_decap_8
XFILLER_30_228 VPWR VGND sg13g2_decap_8
XFILLER_7_424 VPWR VGND sg13g2_decap_4
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_3_630 VPWR VGND sg13g2_decap_8
XFILLER_19_531 VPWR VGND sg13g2_fill_1
XFILLER_48_91 VPWR VGND sg13g2_decap_8
X_2090_ _0735_ net99 state\[17\] VPWR VGND sg13g2_nand2_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_19_564 VPWR VGND sg13g2_fill_2
XFILLER_21_206 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_458 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_14_280 VPWR VGND sg13g2_decap_8
XFILLER_30_751 VPWR VGND sg13g2_fill_1
XFILLER_9_85 VPWR VGND sg13g2_decap_8
X_1943_ VGND VPWR net108 daisychain\[104\] _0628_ net53 sg13g2_a21oi_1
X_1874_ net194 VPWR _0573_ VGND daisychain\[91\] net39 sg13g2_o21ai_1
X_2426_ net354 VGND VPWR _0242_ daisychain\[114\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
X_1308_ VPWR _0005_ state\[104\] VGND sg13g2_inv_1
X_2492__376 VPWR VGND net375 sg13g2_tiehi
X_2357_ net236 VGND VPWR _0173_ daisychain\[45\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2288_ _0834_ net95 state\[116\] VPWR VGND sg13g2_nand2_1
XFILLER_12_239 VPWR VGND sg13g2_decap_8
XFILLER_20_250 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_20_261 VPWR VGND sg13g2_fill_2
XFILLER_4_416 VPWR VGND sg13g2_decap_8
XFILLER_0_600 VPWR VGND sg13g2_decap_8
XFILLER_0_622 VPWR VGND sg13g2_decap_8
XFILLER_0_666 VPWR VGND sg13g2_fill_2
XFILLER_48_637 VPWR VGND sg13g2_fill_2
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_44_810 VPWR VGND sg13g2_decap_8
XFILLER_44_821 VPWR VGND sg13g2_fill_2
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_11_250 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_fill_1
XFILLER_31_559 VPWR VGND sg13g2_decap_8
XFILLER_7_221 VPWR VGND sg13g2_decap_8
XFILLER_8_733 VPWR VGND sg13g2_fill_2
X_2330__291 VPWR VGND net290 sg13g2_tiehi
XFILLER_7_298 VPWR VGND sg13g2_decap_8
X_2406__395 VPWR VGND net394 sg13g2_tiehi
X_2361__229 VPWR VGND net228 sg13g2_tiehi
X_1590_ VGND VPWR _0987_ _0988_ _0162_ _0989_ sg13g2_a21oi_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_38_147 VPWR VGND sg13g2_decap_8
X_2211_ VGND VPWR _0515_ _0795_ _0333_ net85 sg13g2_a21oi_1
X_2142_ _0761_ net116 state\[43\] VPWR VGND sg13g2_nand2_1
X_2073_ VGND VPWR _0883_ _0726_ _0264_ net67 sg13g2_a21oi_1
XFILLER_30_18 VPWR VGND sg13g2_decap_8
X_1926_ state\[102\] daisychain\[102\] net142 _0614_ VPWR VGND sg13g2_mux2_1
X_1857_ _0559_ net172 _0558_ VPWR VGND sg13g2_nand2_1
X_1788_ VGND VPWR net124 daisychain\[73\] _0504_ net61 sg13g2_a21oi_1
XFILLER_29_136 VPWR VGND sg13g2_decap_8
X_2409_ net388 VGND VPWR _0225_ daisychain\[97\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_38_681 VPWR VGND sg13g2_fill_2
XFILLER_40_301 VPWR VGND sg13g2_decap_8
X_2457__260 VPWR VGND net259 sg13g2_tiehi
XFILLER_25_386 VPWR VGND sg13g2_decap_8
XFILLER_25_397 VPWR VGND sg13g2_fill_1
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_5_703 VPWR VGND sg13g2_fill_1
XFILLER_4_213 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_16_353 VPWR VGND sg13g2_decap_8
XFILLER_16_364 VPWR VGND sg13g2_fill_1
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_44_673 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_6_75 VPWR VGND sg13g2_decap_8
X_1711_ state\[59\] daisychain\[59\] net147 _0442_ VPWR VGND sg13g2_mux2_1
X_1642_ _0387_ net169 _0386_ VPWR VGND sg13g2_nand2_1
XFILLER_39_401 VPWR VGND sg13g2_decap_4
X_1573_ VGND VPWR net106 daisychain\[30\] _0976_ net51 sg13g2_a21oi_1
XFILLER_13_0 VPWR VGND sg13g2_fill_2
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_34_161 VPWR VGND sg13g2_decap_8
XFILLER_35_651 VPWR VGND sg13g2_fill_2
X_2125_ VGND VPWR _0987_ _0752_ _0290_ net72 sg13g2_a21oi_1
X_2056_ _0718_ net93 state\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_10_529 VPWR VGND sg13g2_fill_1
XFILLER_41_28 VPWR VGND sg13g2_decap_8
X_1909_ net187 VPWR _0601_ VGND daisychain\[98\] net32 sg13g2_o21ai_1
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_17_106 VPWR VGND sg13g2_decap_8
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_15_40 VPWR VGND sg13g2_fill_1
XFILLER_25_194 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_9_316 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_fill_1
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_41_687 VPWR VGND sg13g2_fill_1
XFILLER_49_743 VPWR VGND sg13g2_decap_8
XFILLER_5_566 VPWR VGND sg13g2_decap_4
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
X_2553__310 VPWR VGND net309 sg13g2_tiehi
XFILLER_31_186 VPWR VGND sg13g2_decap_8
XFILLER_32_621 VPWR VGND sg13g2_fill_2
XFILLER_8_382 VPWR VGND sg13g2_decap_8
X_1556_ state\[28\] daisychain\[28\] net138 _0962_ VPWR VGND sg13g2_mux2_1
X_1625_ VGND VPWR _1015_ _1016_ _0169_ _1017_ sg13g2_a21oi_1
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_39_275 VPWR VGND sg13g2_decap_8
X_1487_ _0907_ net156 _0906_ VPWR VGND sg13g2_nand2_1
XFILLER_27_448 VPWR VGND sg13g2_fill_2
XFILLER_27_459 VPWR VGND sg13g2_fill_2
X_2108_ _0744_ net102 state\[26\] VPWR VGND sg13g2_nand2_1
X_2039_ net178 VPWR _0705_ VGND daisychain\[124\] net26 sg13g2_o21ai_1
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_7_809 VPWR VGND sg13g2_decap_8
XFILLER_2_503 VPWR VGND sg13g2_fill_1
XFILLER_18_437 VPWR VGND sg13g2_fill_2
XFILLER_18_459 VPWR VGND sg13g2_fill_1
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_46_702 VPWR VGND sg13g2_fill_2
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_14_610 VPWR VGND sg13g2_fill_1
XFILLER_26_83 VPWR VGND sg13g2_fill_1
XFILLER_41_473 VPWR VGND sg13g2_decap_8
XFILLER_41_495 VPWR VGND sg13g2_fill_2
XFILLER_9_113 VPWR VGND sg13g2_decap_8
XFILLER_5_363 VPWR VGND sg13g2_decap_8
X_1410_ VPWR _0050_ state\[2\] VGND sg13g2_inv_1
XFILLER_3_98 VPWR VGND sg13g2_decap_8
X_1341_ VPWR _0096_ state\[71\] VGND sg13g2_inv_1
X_2390_ net426 VGND VPWR _0206_ daisychain\[78\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_20_635 VPWR VGND sg13g2_fill_1
XFILLER_20_668 VPWR VGND sg13g2_fill_2
X_2488__392 VPWR VGND net391 sg13g2_tiehi
X_1539_ net183 VPWR _0949_ VGND daisychain\[24\] net28 sg13g2_o21ai_1
Xfanout103 net132 net103 VPWR VGND sg13g2_buf_1
Xfanout114 net132 net114 VPWR VGND sg13g2_buf_1
Xfanout125 net126 net125 VPWR VGND sg13g2_buf_1
Xfanout136 net153 net136 VPWR VGND sg13g2_buf_1
Xfanout147 net152 net147 VPWR VGND sg13g2_buf_1
X_1608_ VGND VPWR net105 daisychain\[37\] _1004_ net51 sg13g2_a21oi_1
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
Xfanout158 net177 net158 VPWR VGND sg13g2_buf_1
Xfanout169 net176 net169 VPWR VGND sg13g2_buf_1
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_43_749 VPWR VGND sg13g2_fill_1
XFILLER_10_167 VPWR VGND sg13g2_decap_8
XFILLER_12_85 VPWR VGND sg13g2_decap_8
XFILLER_2_322 VPWR VGND sg13g2_decap_8
XFILLER_6_127 VPWR VGND sg13g2_decap_8
XFILLER_2_399 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_18_267 VPWR VGND sg13g2_fill_1
XFILLER_18_278 VPWR VGND sg13g2_decap_8
XFILLER_19_746 VPWR VGND sg13g2_decap_8
XFILLER_46_521 VPWR VGND sg13g2_fill_2
XFILLER_14_462 VPWR VGND sg13g2_decap_4
X_1890_ VGND VPWR _0583_ _0584_ _0222_ _0585_ sg13g2_a21oi_1
XFILLER_5_160 VPWR VGND sg13g2_decap_8
X_2511_ net273 VGND VPWR _0327_ state\[71\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2442_ net319 VGND VPWR _0258_ state\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2373_ net204 VGND VPWR _0189_ daisychain\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_17_19 VPWR VGND sg13g2_fill_2
XFILLER_37_532 VPWR VGND sg13g2_fill_1
X_1324_ VPWR _0114_ state\[88\] VGND sg13g2_inv_1
X_2555__246 VPWR VGND net245 sg13g2_tiehi
X_2371__209 VPWR VGND net208 sg13g2_tiehi
X_2340__271 VPWR VGND net270 sg13g2_tiehi
XFILLER_24_237 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_33_771 VPWR VGND sg13g2_fill_2
XFILLER_33_793 VPWR VGND sg13g2_fill_2
X_2416__375 VPWR VGND net374 sg13g2_tiehi
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_15_226 VPWR VGND sg13g2_decap_8
XFILLER_43_513 VPWR VGND sg13g2_decap_4
XFILLER_11_476 VPWR VGND sg13g2_fill_2
XFILLER_23_270 VPWR VGND sg13g2_fill_2
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_30_207 VPWR VGND sg13g2_decap_8
XFILLER_7_403 VPWR VGND sg13g2_decap_8
XFILLER_7_458 VPWR VGND sg13g2_fill_1
XFILLER_24_8 VPWR VGND sg13g2_fill_1
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_459 VPWR VGND uio_oe[4] sg13g2_tiehi
X_1942_ _0627_ net164 _0626_ VPWR VGND sg13g2_nand2_1
XFILLER_30_785 VPWR VGND sg13g2_fill_1
X_1873_ VGND VPWR net126 daisychain\[90\] _0572_ net61 sg13g2_a21oi_1
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_6_491 VPWR VGND sg13g2_decap_8
X_2561__294 VPWR VGND net293 sg13g2_tiehi
X_2425_ net356 VGND VPWR _0241_ daisychain\[113\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2356_ net238 VGND VPWR _0172_ daisychain\[44\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_44_28 VPWR VGND sg13g2_decap_8
X_1307_ VPWR _0006_ state\[105\] VGND sg13g2_inv_1
X_2287_ VGND VPWR _0667_ _0833_ _0371_ net69 sg13g2_a21oi_1
XFILLER_12_218 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
X_2319__313 VPWR VGND net312 sg13g2_tiehi
XFILLER_16_546 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_31_516 VPWR VGND sg13g2_fill_2
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_7_200 VPWR VGND sg13g2_decap_8
XFILLER_7_277 VPWR VGND sg13g2_decap_8
XFILLER_8_701 VPWR VGND sg13g2_fill_1
XFILLER_8_756 VPWR VGND sg13g2_decap_8
XFILLER_39_605 VPWR VGND sg13g2_decap_8
XFILLER_39_627 VPWR VGND sg13g2_fill_1
X_2210_ _0795_ net127 state\[77\] VPWR VGND sg13g2_nand2_1
XFILLER_15_4 VPWR VGND sg13g2_fill_1
XFILLER_35_800 VPWR VGND sg13g2_fill_1
XFILLER_38_126 VPWR VGND sg13g2_decap_8
X_2141_ VGND VPWR _1019_ _0760_ _0298_ net79 sg13g2_a21oi_1
X_2072_ _0726_ net92 state\[8\] VPWR VGND sg13g2_nand2_1
X_1925_ VGND VPWR _0611_ _0612_ _0229_ _0613_ sg13g2_a21oi_1
XFILLER_30_593 VPWR VGND sg13g2_fill_1
X_1856_ state\[88\] daisychain\[88\] net142 _0558_ VPWR VGND sg13g2_mux2_1
X_1787_ _0503_ net172 _0502_ VPWR VGND sg13g2_nand2_1
XFILLER_29_115 VPWR VGND sg13g2_decap_8
XFILLER_39_28 VPWR VGND sg13g2_decap_4
X_2408_ net390 VGND VPWR _0224_ daisychain\[96\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2339_ net272 VGND VPWR _0155_ daisychain\[27\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_38_660 VPWR VGND sg13g2_fill_2
XFILLER_41_814 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_5_715 VPWR VGND sg13g2_decap_8
X_2464__232 VPWR VGND net231 sg13g2_tiehi
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_20_30 VPWR VGND sg13g2_fill_2
XFILLER_20_96 VPWR VGND sg13g2_decap_8
XFILLER_4_269 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_16_332 VPWR VGND sg13g2_fill_2
XFILLER_17_822 VPWR VGND sg13g2_fill_1
XFILLER_29_94 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_12_560 VPWR VGND sg13g2_fill_2
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_8_531 VPWR VGND sg13g2_decap_8
X_2512__266 VPWR VGND net265 sg13g2_tiehi
XFILLER_12_593 VPWR VGND sg13g2_fill_2
XFILLER_6_54 VPWR VGND sg13g2_decap_8
XFILLER_8_542 VPWR VGND sg13g2_fill_1
X_2443__316 VPWR VGND net315 sg13g2_tiehi
X_1710_ VGND VPWR _0439_ _0440_ _0186_ _0441_ sg13g2_a21oi_1
X_1641_ state\[45\] daisychain\[45\] net145 _0386_ VPWR VGND sg13g2_mux2_1
X_1572_ _0975_ net162 _0974_ VPWR VGND sg13g2_nand2_1
XFILLER_3_280 VPWR VGND sg13g2_decap_8
X_2124_ _0752_ net105 state\[34\] VPWR VGND sg13g2_nand2_1
XFILLER_26_118 VPWR VGND sg13g2_decap_4
XFILLER_34_140 VPWR VGND sg13g2_decap_8
XFILLER_35_674 VPWR VGND sg13g2_fill_1
XFILLER_47_490 VPWR VGND sg13g2_decap_8
X_2055_ VGND VPWR _0715_ _0716_ _0255_ _0717_ sg13g2_a21oi_1
X_1908_ VGND VPWR net112 daisychain\[97\] _0600_ net54 sg13g2_a21oi_1
X_1839_ net194 VPWR _0545_ VGND daisychain\[84\] net39 sg13g2_o21ai_1
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_25_173 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_decap_4
XFILLER_41_655 VPWR VGND sg13g2_fill_2
XFILLER_31_95 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_49_766 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_fill_1
XFILLER_16_184 VPWR VGND sg13g2_decap_8
XFILLER_36_449 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_31_165 VPWR VGND sg13g2_decap_8
XFILLER_8_361 VPWR VGND sg13g2_decap_8
X_1555_ VGND VPWR _0959_ _0960_ _0155_ _0961_ sg13g2_a21oi_1
X_2380__447 VPWR VGND net446 sg13g2_tiehi
X_1624_ net190 VPWR _1017_ VGND daisychain\[41\] net35 sg13g2_o21ai_1
XFILLER_27_427 VPWR VGND sg13g2_decap_8
XFILLER_39_254 VPWR VGND sg13g2_decap_8
X_1486_ state\[14\] daisychain\[14\] net134 _0906_ VPWR VGND sg13g2_mux2_1
X_2107_ VGND VPWR _0951_ _0743_ _0281_ net72 sg13g2_a21oi_1
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_35_460 VPWR VGND sg13g2_fill_2
X_2350__251 VPWR VGND net250 sg13g2_tiehi
X_2038_ VGND VPWR net89 daisychain\[123\] _0704_ net48 sg13g2_a21oi_1
XFILLER_10_349 VPWR VGND sg13g2_decap_8
XFILLER_6_309 VPWR VGND sg13g2_decap_8
X_2426__355 VPWR VGND net354 sg13g2_tiehi
XFILLER_18_416 VPWR VGND sg13g2_decap_4
XFILLER_26_482 VPWR VGND sg13g2_decap_4
XFILLER_26_62 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_decap_4
XFILLER_46_736 VPWR VGND sg13g2_fill_1
XFILLER_46_758 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_4
XFILLER_9_169 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_342 VPWR VGND sg13g2_decap_8
X_1340_ VPWR _0097_ state\[72\] VGND sg13g2_inv_1
X_2327__297 VPWR VGND net296 sg13g2_tiehi
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_20_603 VPWR VGND sg13g2_fill_1
XFILLER_32_441 VPWR VGND sg13g2_fill_1
XFILLER_37_769 VPWR VGND sg13g2_fill_2
XFILLER_9_681 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_8_clk clknet_2_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
X_1469_ net179 VPWR _0893_ VGND daisychain\[10\] net23 sg13g2_o21ai_1
X_1538_ VGND VPWR net104 daisychain\[23\] _0948_ net51 sg13g2_a21oi_1
Xfanout104 net106 net104 VPWR VGND sg13g2_buf_1
Xfanout115 net118 net115 VPWR VGND sg13g2_buf_1
Xfanout126 net131 net126 VPWR VGND sg13g2_buf_1
Xfanout137 net140 net137 VPWR VGND sg13g2_buf_1
Xfanout148 net152 net148 VPWR VGND sg13g2_buf_1
Xfanout159 net163 net159 VPWR VGND sg13g2_buf_1
X_1607_ _1003_ net161 _1002_ VPWR VGND sg13g2_nand2_1
XFILLER_15_408 VPWR VGND sg13g2_decap_8
XFILLER_27_224 VPWR VGND sg13g2_decap_8
XFILLER_36_791 VPWR VGND sg13g2_fill_2
X_2495__364 VPWR VGND net363 sg13g2_tiehi
XFILLER_10_146 VPWR VGND sg13g2_decap_8
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_6_106 VPWR VGND sg13g2_decap_8
XFILLER_2_301 VPWR VGND sg13g2_decap_8
XFILLER_2_378 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_4
X_2474__448 VPWR VGND net447 sg13g2_tiehi
XFILLER_18_235 VPWR VGND sg13g2_decap_8
XFILLER_33_249 VPWR VGND sg13g2_decap_8
XFILLER_10_691 VPWR VGND sg13g2_decap_8
X_2510_ net281 VGND VPWR _0326_ state\[70\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1323_ VPWR _0115_ state\[89\] VGND sg13g2_inv_1
X_2441_ net323 VGND VPWR _0257_ state\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2372_ net206 VGND VPWR _0188_ daisychain\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_24_216 VPWR VGND sg13g2_decap_8
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_33_783 VPWR VGND sg13g2_fill_2
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_15_205 VPWR VGND sg13g2_decap_8
XFILLER_16_739 VPWR VGND sg13g2_fill_2
XFILLER_31_709 VPWR VGND sg13g2_fill_1
XFILLER_11_433 VPWR VGND sg13g2_decap_8
XFILLER_11_444 VPWR VGND sg13g2_fill_1
XFILLER_23_74 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_fill_2
XFILLER_19_566 VPWR VGND sg13g2_fill_1
XFILLER_19_577 VPWR VGND sg13g2_decap_8
XFILLER_34_503 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
X_2515__242 VPWR VGND net241 sg13g2_tiehi
XFILLER_15_761 VPWR VGND sg13g2_decap_8
XFILLER_15_794 VPWR VGND sg13g2_fill_2
XFILLER_30_731 VPWR VGND sg13g2_fill_1
XFILLER_30_764 VPWR VGND sg13g2_fill_1
X_1941_ state\[105\] daisychain\[105\] net141 _0626_ VPWR VGND sg13g2_mux2_1
X_1872_ _0571_ net173 _0570_ VPWR VGND sg13g2_nand2_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_1306_ VPWR _0007_ state\[106\] VGND sg13g2_inv_1
X_2424_ net358 VGND VPWR _0240_ daisychain\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2355_ net240 VGND VPWR _0171_ daisychain\[43\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2286_ _0833_ net95 state\[115\] VPWR VGND sg13g2_nand2_1
XFILLER_25_525 VPWR VGND sg13g2_decap_4
XFILLER_37_385 VPWR VGND sg13g2_fill_2
XFILLER_20_285 VPWR VGND sg13g2_fill_2
XFILLER_0_668 VPWR VGND sg13g2_fill_1
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_12_764 VPWR VGND sg13g2_fill_2
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_11_285 VPWR VGND sg13g2_decap_8
XFILLER_7_256 VPWR VGND sg13g2_decap_8
X_2549__382 VPWR VGND net381 sg13g2_tiehi
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_39_639 VPWR VGND sg13g2_decap_4
XFILLER_3_462 VPWR VGND sg13g2_decap_8
X_2140_ _0760_ net116 state\[42\] VPWR VGND sg13g2_nand2_1
XFILLER_34_322 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
X_2071_ VGND VPWR _0879_ _0725_ _0263_ net67 sg13g2_a21oi_1
XFILLER_22_528 VPWR VGND sg13g2_fill_2
XFILLER_30_550 VPWR VGND sg13g2_fill_1
XFILLER_34_399 VPWR VGND sg13g2_fill_1
X_1924_ net188 VPWR _0613_ VGND daisychain\[101\] net33 sg13g2_o21ai_1
X_1855_ VGND VPWR _0555_ _0556_ _0215_ _0557_ sg13g2_a21oi_1
X_1786_ state\[74\] daisychain\[74\] net148 _0502_ VPWR VGND sg13g2_mux2_1
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_45_609 VPWR VGND sg13g2_decap_8
X_2407_ net392 VGND VPWR _0223_ daisychain\[95\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2338_ net274 VGND VPWR _0154_ daisychain\[26\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2269_ VGND VPWR _0631_ _0824_ _0362_ net75 sg13g2_a21oi_1
XFILLER_13_539 VPWR VGND sg13g2_fill_2
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_38_694 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
X_2390__427 VPWR VGND net426 sg13g2_tiehi
XFILLER_4_248 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_20_75 VPWR VGND sg13g2_decap_8
X_2360__231 VPWR VGND net230 sg13g2_tiehi
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_29_73 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_44_631 VPWR VGND sg13g2_fill_2
XFILLER_44_653 VPWR VGND sg13g2_fill_1
XFILLER_48_469 VPWR VGND sg13g2_decap_8
X_2471__204 VPWR VGND net203 sg13g2_tiehi
X_2436__335 VPWR VGND net334 sg13g2_tiehi
XFILLER_12_583 VPWR VGND sg13g2_decap_4
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_8_554 VPWR VGND sg13g2_decap_8
XFILLER_8_598 VPWR VGND sg13g2_decap_8
X_1640_ VGND VPWR _1027_ _0384_ _0172_ _0385_ sg13g2_a21oi_1
X_1571_ state\[31\] daisychain\[31\] net139 _0974_ VPWR VGND sg13g2_mux2_1
X_2123_ VGND VPWR _0983_ _0751_ _0289_ net73 sg13g2_a21oi_1
XFILLER_22_358 VPWR VGND sg13g2_fill_2
XFILLER_34_196 VPWR VGND sg13g2_decap_8
XFILLER_35_653 VPWR VGND sg13g2_fill_1
X_2530__378 VPWR VGND net377 sg13g2_tiehi
X_2337__277 VPWR VGND net276 sg13g2_tiehi
X_2054_ net178 VPWR _0717_ VGND daisychain\[127\] net26 sg13g2_o21ai_1
X_1907_ _0599_ net166 _0598_ VPWR VGND sg13g2_nand2_1
X_1838_ VGND VPWR net124 daisychain\[83\] _0544_ net61 sg13g2_a21oi_1
XFILLER_2_719 VPWR VGND sg13g2_decap_8
X_1769_ net196 VPWR _0489_ VGND daisychain\[70\] net41 sg13g2_o21ai_1
XFILLER_14_815 VPWR VGND sg13g2_decap_8
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_15_86 VPWR VGND sg13g2_decap_8
XFILLER_25_152 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_41_678 VPWR VGND sg13g2_decap_8
XFILLER_31_74 VPWR VGND sg13g2_decap_8
X_2542__238 VPWR VGND net237 sg13g2_tiehi
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_16_163 VPWR VGND sg13g2_decap_8
XFILLER_17_620 VPWR VGND sg13g2_decap_4
XFILLER_20_807 VPWR VGND sg13g2_fill_1
XFILLER_32_623 VPWR VGND sg13g2_fill_1
XFILLER_32_656 VPWR VGND sg13g2_fill_2
XFILLER_44_483 VPWR VGND sg13g2_decap_8
XFILLER_20_818 VPWR VGND sg13g2_fill_2
XFILLER_31_144 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
X_1485_ VGND VPWR _0903_ _0904_ _0141_ _0905_ sg13g2_a21oi_1
X_1554_ net182 VPWR _0961_ VGND daisychain\[27\] net27 sg13g2_o21ai_1
X_1623_ VGND VPWR net116 daisychain\[40\] _1016_ net57 sg13g2_a21oi_1
.ends

