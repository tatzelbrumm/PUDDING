VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO heichips25_pudding
  CLASS BLOCK ;
  FOREIGN heichips25_pudding ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 21.580 3.150 23.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 41.580 3.150 43.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 61.580 3.150 63.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 81.580 3.150 83.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 101.580 3.150 103.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 121.580 3.150 123.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 141.580 3.150 143.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 161.580 3.150 163.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 181.580 3.150 183.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 201.580 3.150 203.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 221.580 3.150 223.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 241.580 3.150 243.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 261.580 3.150 263.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 281.580 3.150 283.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 301.580 3.150 303.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 321.580 3.150 323.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 341.580 3.150 343.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 361.580 3.150 363.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 381.580 3.150 383.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 401.580 3.560 403.780 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 421.580 3.560 423.780 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 441.580 3.560 443.780 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 461.580 3.560 463.780 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 481.580 3.560 483.780 193.000 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 22.480 496.800 24.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 42.480 496.800 44.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 62.480 496.800 64.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 82.480 496.800 84.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 102.480 496.800 104.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 122.480 496.800 124.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 142.480 496.800 144.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 162.480 496.800 164.680 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 182.480 496.800 184.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 15.380 3.560 17.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 35.380 3.560 37.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 55.380 3.560 57.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 75.380 3.560 77.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 95.380 3.560 97.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 115.380 3.560 117.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 135.380 3.560 137.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 155.380 3.560 157.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 175.380 3.560 177.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 195.380 3.560 197.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 215.380 3.560 217.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 235.380 3.560 237.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 255.380 3.560 257.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 275.380 3.560 277.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 295.380 3.560 297.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 315.380 3.560 317.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 335.380 3.560 337.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 355.380 3.560 357.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 375.380 3.560 377.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 395.380 3.560 397.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 415.380 3.560 417.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 435.380 3.560 437.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 455.380 3.560 457.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 475.380 3.560 477.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 495.380 3.560 497.580 193.000 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 16.280 497.580 18.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 36.280 497.580 38.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 56.280 497.580 58.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 76.280 497.580 78.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 96.280 497.580 98.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 116.280 497.580 118.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 136.280 497.580 138.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 156.280 497.580 158.480 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 2.880 176.280 497.580 178.480 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.340 0.400 183.740 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.140 0.400 179.540 ;
    END
  END ena
  PIN i_in
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER Metal3 ;
        RECT 400.000 107.930 500.000 108.630 ;
    END
  END i_in
  PIN i_out
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 66.047997 ;
    PORT
      LAYER Metal3 ;
        RECT 400.000 99.745 500.000 100.445 ;
    END
  END i_out
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.540 0.400 187.940 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.940 0.400 112.340 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.140 0.400 116.540 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.340 0.400 120.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.540 0.400 124.940 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.740 0.400 129.140 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.940 0.400 133.340 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.140 0.400 137.540 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.340 0.400 141.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.540 0.400 145.940 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.740 0.400 150.140 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.940 0.400 154.340 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.140 0.400 158.540 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.340 0.400 162.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.540 0.400 166.940 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.740 0.400 171.140 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.940 0.400 175.340 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.340 0.400 78.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.540 0.400 82.940 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.400 87.140 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.940 0.400 91.340 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.140 0.400 95.540 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.340 0.400 99.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.540 0.400 103.940 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.740 0.400 108.140 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.740 0.400 45.140 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.140 0.400 53.540 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.540 0.400 61.940 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.740 0.400 66.140 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.940 0.400 70.340 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.140 0.400 74.540 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.140 0.400 11.540 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.540 0.400 19.940 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.940 0.400 28.340 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.340 0.400 36.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 400.000 192.930 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 403.000 193.000 ;
      LAYER Metal2 ;
        RECT 2.775 3.635 403.000 192.925 ;
      LAYER Metal3 ;
        RECT 0.400 188.150 403.000 192.880 ;
        RECT 0.610 187.330 403.000 188.150 ;
        RECT 0.400 183.950 403.000 187.330 ;
        RECT 0.610 183.130 403.000 183.950 ;
        RECT 0.400 179.750 403.000 183.130 ;
        RECT 0.610 178.930 403.000 179.750 ;
        RECT 0.400 175.550 403.000 178.930 ;
        RECT 0.610 174.730 403.000 175.550 ;
        RECT 0.400 171.350 403.000 174.730 ;
        RECT 0.610 170.530 403.000 171.350 ;
        RECT 0.400 167.150 403.000 170.530 ;
        RECT 0.610 166.330 403.000 167.150 ;
        RECT 0.400 162.950 403.000 166.330 ;
        RECT 0.610 162.130 403.000 162.950 ;
        RECT 0.400 158.750 403.000 162.130 ;
        RECT 0.610 157.930 403.000 158.750 ;
        RECT 0.400 154.550 403.000 157.930 ;
        RECT 0.610 153.730 403.000 154.550 ;
        RECT 0.400 150.350 403.000 153.730 ;
        RECT 0.610 149.530 403.000 150.350 ;
        RECT 0.400 146.150 403.000 149.530 ;
        RECT 0.610 145.330 403.000 146.150 ;
        RECT 0.400 141.950 403.000 145.330 ;
        RECT 0.610 141.130 403.000 141.950 ;
        RECT 0.400 137.750 403.000 141.130 ;
        RECT 0.610 136.930 403.000 137.750 ;
        RECT 0.400 133.550 403.000 136.930 ;
        RECT 0.610 132.730 403.000 133.550 ;
        RECT 0.400 129.350 403.000 132.730 ;
        RECT 0.610 128.530 403.000 129.350 ;
        RECT 0.400 125.150 403.000 128.530 ;
        RECT 0.610 124.330 403.000 125.150 ;
        RECT 0.400 120.950 403.000 124.330 ;
        RECT 0.610 120.130 403.000 120.950 ;
        RECT 0.400 116.750 403.000 120.130 ;
        RECT 0.610 115.930 403.000 116.750 ;
        RECT 0.400 112.550 403.000 115.930 ;
        RECT 0.610 111.730 403.000 112.550 ;
        RECT 0.400 108.840 403.000 111.730 ;
        RECT 0.400 108.350 399.790 108.840 ;
        RECT 0.610 107.720 399.790 108.350 ;
        RECT 0.610 107.530 403.000 107.720 ;
        RECT 0.400 104.150 403.000 107.530 ;
        RECT 0.610 103.330 403.000 104.150 ;
        RECT 0.400 100.655 403.000 103.330 ;
        RECT 0.400 99.950 399.790 100.655 ;
        RECT 0.610 99.535 399.790 99.950 ;
        RECT 0.610 99.130 403.000 99.535 ;
        RECT 0.400 95.750 403.000 99.130 ;
        RECT 0.610 94.930 403.000 95.750 ;
        RECT 0.400 91.550 403.000 94.930 ;
        RECT 0.610 90.730 403.000 91.550 ;
        RECT 0.400 87.350 403.000 90.730 ;
        RECT 0.610 86.530 403.000 87.350 ;
        RECT 0.400 83.150 403.000 86.530 ;
        RECT 0.610 82.330 403.000 83.150 ;
        RECT 0.400 78.950 403.000 82.330 ;
        RECT 0.610 78.130 403.000 78.950 ;
        RECT 0.400 74.750 403.000 78.130 ;
        RECT 0.610 73.930 403.000 74.750 ;
        RECT 0.400 70.550 403.000 73.930 ;
        RECT 0.610 69.730 403.000 70.550 ;
        RECT 0.400 66.350 403.000 69.730 ;
        RECT 0.610 65.530 403.000 66.350 ;
        RECT 0.400 62.150 403.000 65.530 ;
        RECT 0.610 61.330 403.000 62.150 ;
        RECT 0.400 57.950 403.000 61.330 ;
        RECT 0.610 57.130 403.000 57.950 ;
        RECT 0.400 53.750 403.000 57.130 ;
        RECT 0.610 52.930 403.000 53.750 ;
        RECT 0.400 49.550 403.000 52.930 ;
        RECT 0.610 48.730 403.000 49.550 ;
        RECT 0.400 45.350 403.000 48.730 ;
        RECT 0.610 44.530 403.000 45.350 ;
        RECT 0.400 41.150 403.000 44.530 ;
        RECT 0.610 40.330 403.000 41.150 ;
        RECT 0.400 36.950 403.000 40.330 ;
        RECT 0.610 36.130 403.000 36.950 ;
        RECT 0.400 32.750 403.000 36.130 ;
        RECT 0.610 31.930 403.000 32.750 ;
        RECT 0.400 28.550 403.000 31.930 ;
        RECT 0.610 27.730 403.000 28.550 ;
        RECT 0.400 24.350 403.000 27.730 ;
        RECT 0.610 23.530 403.000 24.350 ;
        RECT 0.400 20.150 403.000 23.530 ;
        RECT 0.610 19.330 403.000 20.150 ;
        RECT 0.400 15.950 403.000 19.330 ;
        RECT 0.610 15.130 403.000 15.950 ;
        RECT 0.400 11.750 403.000 15.130 ;
        RECT 0.610 10.930 403.000 11.750 ;
        RECT 0.400 3.680 403.000 10.930 ;
      LAYER Metal4 ;
        RECT 13.340 3.635 400.000 192.925 ;
      LAYER Metal5 ;
        RECT 15.515 3.470 400.000 193.090 ;
  END
END heichips25_pudding
END LIBRARY

