magic
tech ihp-sg13g2
timestamp 1771125512
use pmosHV  pmosHV_0
timestamp 1771125512
transform 1 0 0 0 1 0
box -62 -62 3330 3262
<< end >>
