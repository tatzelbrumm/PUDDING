module heichips25_pudding (clk,
    ena,
    i_in,
    i_out,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 inout i_in;
 inout i_out;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire \bias[0] ;
 wire \bias[1] ;
 wire dacout;
 wire \daisychain[0] ;
 wire \daisychain[100] ;
 wire \daisychain[101] ;
 wire \daisychain[102] ;
 wire \daisychain[103] ;
 wire \daisychain[104] ;
 wire \daisychain[105] ;
 wire \daisychain[106] ;
 wire \daisychain[107] ;
 wire \daisychain[108] ;
 wire \daisychain[109] ;
 wire \daisychain[10] ;
 wire \daisychain[110] ;
 wire \daisychain[111] ;
 wire \daisychain[112] ;
 wire \daisychain[113] ;
 wire \daisychain[114] ;
 wire \daisychain[115] ;
 wire \daisychain[116] ;
 wire \daisychain[117] ;
 wire \daisychain[118] ;
 wire \daisychain[119] ;
 wire \daisychain[11] ;
 wire \daisychain[120] ;
 wire \daisychain[121] ;
 wire \daisychain[122] ;
 wire \daisychain[123] ;
 wire \daisychain[124] ;
 wire \daisychain[125] ;
 wire \daisychain[126] ;
 wire \daisychain[127] ;
 wire \daisychain[12] ;
 wire \daisychain[13] ;
 wire \daisychain[14] ;
 wire \daisychain[15] ;
 wire \daisychain[16] ;
 wire \daisychain[17] ;
 wire \daisychain[18] ;
 wire \daisychain[19] ;
 wire \daisychain[1] ;
 wire \daisychain[20] ;
 wire \daisychain[21] ;
 wire \daisychain[22] ;
 wire \daisychain[23] ;
 wire \daisychain[24] ;
 wire \daisychain[25] ;
 wire \daisychain[26] ;
 wire \daisychain[27] ;
 wire \daisychain[28] ;
 wire \daisychain[29] ;
 wire \daisychain[2] ;
 wire \daisychain[30] ;
 wire \daisychain[31] ;
 wire \daisychain[32] ;
 wire \daisychain[33] ;
 wire \daisychain[34] ;
 wire \daisychain[35] ;
 wire \daisychain[36] ;
 wire \daisychain[37] ;
 wire \daisychain[38] ;
 wire \daisychain[39] ;
 wire \daisychain[3] ;
 wire \daisychain[40] ;
 wire \daisychain[41] ;
 wire \daisychain[42] ;
 wire \daisychain[43] ;
 wire \daisychain[44] ;
 wire \daisychain[45] ;
 wire \daisychain[46] ;
 wire \daisychain[47] ;
 wire \daisychain[48] ;
 wire \daisychain[49] ;
 wire \daisychain[4] ;
 wire \daisychain[50] ;
 wire \daisychain[51] ;
 wire \daisychain[52] ;
 wire \daisychain[53] ;
 wire \daisychain[54] ;
 wire \daisychain[55] ;
 wire \daisychain[56] ;
 wire \daisychain[57] ;
 wire \daisychain[58] ;
 wire \daisychain[59] ;
 wire \daisychain[5] ;
 wire \daisychain[60] ;
 wire \daisychain[61] ;
 wire \daisychain[62] ;
 wire \daisychain[63] ;
 wire \daisychain[64] ;
 wire \daisychain[65] ;
 wire \daisychain[66] ;
 wire \daisychain[67] ;
 wire \daisychain[68] ;
 wire \daisychain[69] ;
 wire \daisychain[6] ;
 wire \daisychain[70] ;
 wire \daisychain[71] ;
 wire \daisychain[72] ;
 wire \daisychain[73] ;
 wire \daisychain[74] ;
 wire \daisychain[75] ;
 wire \daisychain[76] ;
 wire \daisychain[77] ;
 wire \daisychain[78] ;
 wire \daisychain[79] ;
 wire \daisychain[7] ;
 wire \daisychain[80] ;
 wire \daisychain[81] ;
 wire \daisychain[82] ;
 wire \daisychain[83] ;
 wire \daisychain[84] ;
 wire \daisychain[85] ;
 wire \daisychain[86] ;
 wire \daisychain[87] ;
 wire \daisychain[88] ;
 wire \daisychain[89] ;
 wire \daisychain[8] ;
 wire \daisychain[90] ;
 wire \daisychain[91] ;
 wire \daisychain[92] ;
 wire \daisychain[93] ;
 wire \daisychain[94] ;
 wire \daisychain[95] ;
 wire \daisychain[96] ;
 wire \daisychain[97] ;
 wire \daisychain[98] ;
 wire \daisychain[99] ;
 wire \daisychain[9] ;
 wire \digitalen.g[0].u.OUTN ;
 wire \digitalen.g[0].u.OUTP ;
 wire \digitalen.g[1].u.OUTN ;
 wire \digitalen.g[1].u.OUTP ;
 wire \digitalen.g[2].u.OUTN ;
 wire \digitalen.g[2].u.OUTP ;
 wire \digitalen.g[3].u.OUTN ;
 wire \digitalen.g[3].u.OUTP ;
 wire \iref[0] ;
 wire \iref[1] ;
 wire net1;
 wire \state[0] ;
 wire \state[100] ;
 wire \state[101] ;
 wire \state[102] ;
 wire \state[103] ;
 wire \state[104] ;
 wire \state[105] ;
 wire \state[106] ;
 wire \state[107] ;
 wire \state[108] ;
 wire \state[109] ;
 wire \state[10] ;
 wire \state[110] ;
 wire \state[111] ;
 wire \state[112] ;
 wire \state[113] ;
 wire \state[114] ;
 wire \state[115] ;
 wire \state[116] ;
 wire \state[117] ;
 wire \state[118] ;
 wire \state[119] ;
 wire \state[11] ;
 wire \state[120] ;
 wire \state[121] ;
 wire \state[122] ;
 wire \state[123] ;
 wire \state[124] ;
 wire \state[125] ;
 wire \state[126] ;
 wire \state[127] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[16] ;
 wire \state[17] ;
 wire \state[18] ;
 wire \state[19] ;
 wire \state[1] ;
 wire \state[20] ;
 wire \state[21] ;
 wire \state[22] ;
 wire \state[23] ;
 wire \state[24] ;
 wire \state[25] ;
 wire \state[26] ;
 wire \state[27] ;
 wire \state[28] ;
 wire \state[29] ;
 wire \state[2] ;
 wire \state[30] ;
 wire \state[31] ;
 wire \state[32] ;
 wire \state[33] ;
 wire \state[34] ;
 wire \state[35] ;
 wire \state[36] ;
 wire \state[37] ;
 wire \state[38] ;
 wire \state[39] ;
 wire \state[3] ;
 wire \state[40] ;
 wire \state[41] ;
 wire \state[42] ;
 wire \state[43] ;
 wire \state[44] ;
 wire \state[45] ;
 wire \state[46] ;
 wire \state[47] ;
 wire \state[48] ;
 wire \state[49] ;
 wire \state[4] ;
 wire \state[50] ;
 wire \state[51] ;
 wire \state[52] ;
 wire \state[53] ;
 wire \state[54] ;
 wire \state[55] ;
 wire \state[56] ;
 wire \state[57] ;
 wire \state[58] ;
 wire \state[59] ;
 wire \state[5] ;
 wire \state[60] ;
 wire \state[61] ;
 wire \state[62] ;
 wire \state[63] ;
 wire \state[64] ;
 wire \state[65] ;
 wire \state[66] ;
 wire \state[67] ;
 wire \state[68] ;
 wire \state[69] ;
 wire \state[6] ;
 wire \state[70] ;
 wire \state[71] ;
 wire \state[72] ;
 wire \state[73] ;
 wire \state[74] ;
 wire \state[75] ;
 wire \state[76] ;
 wire \state[77] ;
 wire \state[78] ;
 wire \state[79] ;
 wire \state[7] ;
 wire \state[80] ;
 wire \state[81] ;
 wire \state[82] ;
 wire \state[83] ;
 wire \state[84] ;
 wire \state[85] ;
 wire \state[86] ;
 wire \state[87] ;
 wire \state[88] ;
 wire \state[89] ;
 wire \state[8] ;
 wire \state[90] ;
 wire \state[91] ;
 wire \state[92] ;
 wire \state[93] ;
 wire \state[94] ;
 wire \state[95] ;
 wire \state[96] ;
 wire \state[97] ;
 wire \state[98] ;
 wire \state[99] ;
 wire \state[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \vdda[0] ;
 wire \vdda[1] ;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _0898_ (.Y(_0695_),
    .A(\daisychain[123] ));
 sg13g2_inv_1 _0899_ (.Y(_0696_),
    .A(net138));
 sg13g2_inv_1 _0900_ (.Y(_0028_),
    .A(\state[125] ));
 sg13g2_inv_1 _0901_ (.Y(_0697_),
    .A(\daisychain[125] ));
 sg13g2_inv_1 _0902_ (.Y(_0698_),
    .A(\daisychain[124] ));
 sg13g2_inv_1 _0903_ (.Y(_0029_),
    .A(\state[126] ));
 sg13g2_inv_1 _0904_ (.Y(_0699_),
    .A(\daisychain[126] ));
 sg13g2_inv_1 _0905_ (.Y(_0030_),
    .A(\state[127] ));
 sg13g2_inv_1 _0906_ (.Y(_0700_),
    .A(\daisychain[127] ));
 sg13g2_inv_1 _0907_ (.Y(_0000_),
    .A(\state[0] ));
 sg13g2_inv_1 _0908_ (.Y(_0039_),
    .A(\state[1] ));
 sg13g2_inv_1 _0909_ (.Y(_0050_),
    .A(\state[2] ));
 sg13g2_inv_1 _0910_ (.Y(_0061_),
    .A(\state[3] ));
 sg13g2_inv_1 _0911_ (.Y(_0072_),
    .A(\state[4] ));
 sg13g2_inv_1 _0912_ (.Y(_0083_),
    .A(\state[5] ));
 sg13g2_inv_1 _0913_ (.Y(_0094_),
    .A(\state[6] ));
 sg13g2_inv_1 _0914_ (.Y(_0105_),
    .A(\state[7] ));
 sg13g2_inv_1 _0915_ (.Y(_0116_),
    .A(\state[8] ));
 sg13g2_inv_1 _0916_ (.Y(_0127_),
    .A(\state[9] ));
 sg13g2_inv_1 _0917_ (.Y(_0011_),
    .A(\state[10] ));
 sg13g2_inv_1 _0918_ (.Y(_0022_),
    .A(\state[11] ));
 sg13g2_inv_1 _0919_ (.Y(_0031_),
    .A(\state[12] ));
 sg13g2_inv_1 _0920_ (.Y(_0032_),
    .A(\state[13] ));
 sg13g2_inv_1 _0921_ (.Y(_0033_),
    .A(\state[14] ));
 sg13g2_inv_1 _0922_ (.Y(_0034_),
    .A(\state[15] ));
 sg13g2_inv_1 _0923_ (.Y(_0035_),
    .A(\state[16] ));
 sg13g2_inv_1 _0924_ (.Y(_0036_),
    .A(\state[17] ));
 sg13g2_inv_1 _0925_ (.Y(_0037_),
    .A(\state[18] ));
 sg13g2_inv_1 _0926_ (.Y(_0038_),
    .A(\state[19] ));
 sg13g2_inv_1 _0927_ (.Y(_0040_),
    .A(\state[20] ));
 sg13g2_inv_1 _0928_ (.Y(_0041_),
    .A(\state[21] ));
 sg13g2_inv_1 _0929_ (.Y(_0042_),
    .A(\state[22] ));
 sg13g2_inv_1 _0930_ (.Y(_0043_),
    .A(\state[23] ));
 sg13g2_inv_1 _0931_ (.Y(_0044_),
    .A(\state[24] ));
 sg13g2_inv_1 _0932_ (.Y(_0045_),
    .A(\state[25] ));
 sg13g2_inv_1 _0933_ (.Y(_0046_),
    .A(\state[26] ));
 sg13g2_inv_1 _0934_ (.Y(_0047_),
    .A(\state[27] ));
 sg13g2_inv_1 _0935_ (.Y(_0048_),
    .A(\state[28] ));
 sg13g2_inv_1 _0936_ (.Y(_0049_),
    .A(\state[29] ));
 sg13g2_inv_1 _0937_ (.Y(_0051_),
    .A(\state[30] ));
 sg13g2_inv_1 _0938_ (.Y(_0052_),
    .A(\state[31] ));
 sg13g2_inv_1 _0939_ (.Y(_0053_),
    .A(\state[32] ));
 sg13g2_inv_1 _0940_ (.Y(_0054_),
    .A(\state[33] ));
 sg13g2_inv_1 _0941_ (.Y(_0055_),
    .A(\state[34] ));
 sg13g2_inv_1 _0942_ (.Y(_0056_),
    .A(\state[35] ));
 sg13g2_inv_1 _0943_ (.Y(_0057_),
    .A(\state[36] ));
 sg13g2_inv_1 _0944_ (.Y(_0058_),
    .A(\state[37] ));
 sg13g2_inv_1 _0945_ (.Y(_0059_),
    .A(\state[38] ));
 sg13g2_inv_1 _0946_ (.Y(_0060_),
    .A(\state[39] ));
 sg13g2_inv_1 _0947_ (.Y(_0062_),
    .A(\state[40] ));
 sg13g2_inv_1 _0948_ (.Y(_0063_),
    .A(\state[41] ));
 sg13g2_inv_1 _0949_ (.Y(_0064_),
    .A(\state[42] ));
 sg13g2_inv_1 _0950_ (.Y(_0065_),
    .A(\state[43] ));
 sg13g2_inv_1 _0951_ (.Y(_0066_),
    .A(\state[44] ));
 sg13g2_inv_1 _0952_ (.Y(_0067_),
    .A(\state[45] ));
 sg13g2_inv_1 _0953_ (.Y(_0068_),
    .A(\state[46] ));
 sg13g2_inv_1 _0954_ (.Y(_0069_),
    .A(\state[47] ));
 sg13g2_inv_1 _0955_ (.Y(_0070_),
    .A(\state[48] ));
 sg13g2_inv_1 _0956_ (.Y(_0071_),
    .A(\state[49] ));
 sg13g2_inv_1 _0957_ (.Y(_0073_),
    .A(\state[50] ));
 sg13g2_inv_1 _0958_ (.Y(_0074_),
    .A(\state[51] ));
 sg13g2_inv_1 _0959_ (.Y(_0075_),
    .A(\state[52] ));
 sg13g2_inv_1 _0960_ (.Y(_0076_),
    .A(\state[53] ));
 sg13g2_inv_1 _0961_ (.Y(_0077_),
    .A(\state[54] ));
 sg13g2_inv_1 _0962_ (.Y(_0078_),
    .A(\state[55] ));
 sg13g2_inv_1 _0963_ (.Y(_0079_),
    .A(\state[56] ));
 sg13g2_inv_1 _0964_ (.Y(_0080_),
    .A(\state[57] ));
 sg13g2_inv_1 _0965_ (.Y(_0081_),
    .A(\state[58] ));
 sg13g2_inv_1 _0966_ (.Y(_0082_),
    .A(\state[59] ));
 sg13g2_inv_1 _0967_ (.Y(_0084_),
    .A(\state[60] ));
 sg13g2_inv_1 _0968_ (.Y(_0085_),
    .A(\state[61] ));
 sg13g2_inv_1 _0969_ (.Y(_0086_),
    .A(\state[62] ));
 sg13g2_inv_1 _0970_ (.Y(_0087_),
    .A(\state[63] ));
 sg13g2_inv_1 _0971_ (.Y(_0088_),
    .A(\state[64] ));
 sg13g2_inv_1 _0972_ (.Y(_0089_),
    .A(\state[65] ));
 sg13g2_inv_1 _0973_ (.Y(_0090_),
    .A(\state[66] ));
 sg13g2_inv_1 _0974_ (.Y(_0091_),
    .A(\state[67] ));
 sg13g2_inv_1 _0975_ (.Y(_0092_),
    .A(\state[68] ));
 sg13g2_inv_1 _0976_ (.Y(_0093_),
    .A(\state[69] ));
 sg13g2_inv_1 _0977_ (.Y(_0095_),
    .A(\state[70] ));
 sg13g2_inv_1 _0978_ (.Y(_0096_),
    .A(\state[71] ));
 sg13g2_inv_1 _0979_ (.Y(_0097_),
    .A(\state[72] ));
 sg13g2_inv_1 _0980_ (.Y(_0098_),
    .A(\state[73] ));
 sg13g2_inv_1 _0981_ (.Y(_0099_),
    .A(\state[74] ));
 sg13g2_inv_1 _0982_ (.Y(_0100_),
    .A(\state[75] ));
 sg13g2_inv_1 _0983_ (.Y(_0101_),
    .A(\state[76] ));
 sg13g2_inv_1 _0984_ (.Y(_0102_),
    .A(\state[77] ));
 sg13g2_inv_1 _0985_ (.Y(_0103_),
    .A(\state[78] ));
 sg13g2_inv_1 _0986_ (.Y(_0104_),
    .A(\state[79] ));
 sg13g2_inv_1 _0987_ (.Y(_0106_),
    .A(\state[80] ));
 sg13g2_inv_1 _0988_ (.Y(_0107_),
    .A(\state[81] ));
 sg13g2_inv_1 _0989_ (.Y(_0108_),
    .A(\state[82] ));
 sg13g2_inv_1 _0990_ (.Y(_0109_),
    .A(\state[83] ));
 sg13g2_inv_1 _0991_ (.Y(_0110_),
    .A(\state[84] ));
 sg13g2_inv_1 _0992_ (.Y(_0111_),
    .A(\state[85] ));
 sg13g2_inv_1 _0993_ (.Y(_0112_),
    .A(\state[86] ));
 sg13g2_inv_1 _0994_ (.Y(_0113_),
    .A(\state[87] ));
 sg13g2_inv_1 _0995_ (.Y(_0114_),
    .A(\state[88] ));
 sg13g2_inv_1 _0996_ (.Y(_0115_),
    .A(\state[89] ));
 sg13g2_inv_1 _0997_ (.Y(_0117_),
    .A(\state[90] ));
 sg13g2_inv_1 _0998_ (.Y(_0118_),
    .A(\state[91] ));
 sg13g2_inv_1 _0999_ (.Y(_0119_),
    .A(\state[92] ));
 sg13g2_inv_1 _1000_ (.Y(_0120_),
    .A(\state[93] ));
 sg13g2_inv_1 _1001_ (.Y(_0121_),
    .A(\state[94] ));
 sg13g2_inv_1 _1002_ (.Y(_0122_),
    .A(\state[95] ));
 sg13g2_inv_1 _1003_ (.Y(_0123_),
    .A(\state[96] ));
 sg13g2_inv_1 _1004_ (.Y(_0124_),
    .A(\state[97] ));
 sg13g2_inv_1 _1005_ (.Y(_0125_),
    .A(\state[98] ));
 sg13g2_inv_1 _1006_ (.Y(_0126_),
    .A(\state[99] ));
 sg13g2_inv_1 _1007_ (.Y(_0001_),
    .A(\state[100] ));
 sg13g2_inv_1 _1008_ (.Y(_0002_),
    .A(\state[101] ));
 sg13g2_inv_1 _1009_ (.Y(_0003_),
    .A(\state[102] ));
 sg13g2_inv_1 _1010_ (.Y(_0004_),
    .A(\state[103] ));
 sg13g2_inv_1 _1011_ (.Y(_0005_),
    .A(\state[104] ));
 sg13g2_inv_1 _1012_ (.Y(_0006_),
    .A(\state[105] ));
 sg13g2_inv_1 _1013_ (.Y(_0007_),
    .A(\state[106] ));
 sg13g2_inv_1 _1014_ (.Y(_0008_),
    .A(\state[107] ));
 sg13g2_inv_1 _1015_ (.Y(_0009_),
    .A(\state[108] ));
 sg13g2_inv_1 _1016_ (.Y(_0010_),
    .A(\state[109] ));
 sg13g2_inv_1 _1017_ (.Y(_0012_),
    .A(\state[110] ));
 sg13g2_inv_1 _1018_ (.Y(_0013_),
    .A(\state[111] ));
 sg13g2_inv_1 _1019_ (.Y(_0014_),
    .A(\state[112] ));
 sg13g2_inv_1 _1020_ (.Y(_0015_),
    .A(\state[113] ));
 sg13g2_inv_1 _1021_ (.Y(_0016_),
    .A(\state[114] ));
 sg13g2_inv_1 _1022_ (.Y(_0017_),
    .A(\state[115] ));
 sg13g2_inv_1 _1023_ (.Y(_0018_),
    .A(\state[116] ));
 sg13g2_inv_1 _1024_ (.Y(_0019_),
    .A(\state[117] ));
 sg13g2_inv_1 _1025_ (.Y(_0020_),
    .A(\state[118] ));
 sg13g2_inv_1 _1026_ (.Y(_0021_),
    .A(\state[119] ));
 sg13g2_inv_1 _1027_ (.Y(_0023_),
    .A(\state[120] ));
 sg13g2_inv_1 _1028_ (.Y(_0024_),
    .A(\state[121] ));
 sg13g2_inv_1 _1029_ (.Y(_0025_),
    .A(\state[122] ));
 sg13g2_inv_1 _1030_ (.Y(_0026_),
    .A(\state[123] ));
 sg13g2_inv_1 _1031_ (.Y(_0027_),
    .A(\state[124] ));
 sg13g2_inv_1 _1032_ (.Y(_0701_),
    .A(\daisychain[0] ));
 sg13g2_inv_1 _1033_ (.Y(_0702_),
    .A(\daisychain[1] ));
 sg13g2_inv_1 _1034_ (.Y(_0703_),
    .A(\daisychain[2] ));
 sg13g2_inv_1 _1035_ (.Y(_0704_),
    .A(\daisychain[3] ));
 sg13g2_inv_1 _1036_ (.Y(_0705_),
    .A(\daisychain[4] ));
 sg13g2_inv_1 _1037_ (.Y(_0706_),
    .A(\daisychain[5] ));
 sg13g2_inv_1 _1038_ (.Y(_0707_),
    .A(\daisychain[6] ));
 sg13g2_inv_1 _1039_ (.Y(_0708_),
    .A(\daisychain[7] ));
 sg13g2_inv_1 _1040_ (.Y(_0709_),
    .A(\daisychain[8] ));
 sg13g2_inv_1 _1041_ (.Y(_0710_),
    .A(\daisychain[9] ));
 sg13g2_inv_1 _1042_ (.Y(_0711_),
    .A(\daisychain[10] ));
 sg13g2_inv_1 _1043_ (.Y(_0712_),
    .A(\daisychain[11] ));
 sg13g2_inv_1 _1044_ (.Y(_0713_),
    .A(\daisychain[12] ));
 sg13g2_inv_1 _1045_ (.Y(_0714_),
    .A(\daisychain[13] ));
 sg13g2_inv_1 _1046_ (.Y(_0715_),
    .A(\daisychain[14] ));
 sg13g2_inv_1 _1047_ (.Y(_0716_),
    .A(\daisychain[15] ));
 sg13g2_inv_1 _1048_ (.Y(_0717_),
    .A(\daisychain[16] ));
 sg13g2_inv_1 _1049_ (.Y(_0718_),
    .A(\daisychain[17] ));
 sg13g2_inv_1 _1050_ (.Y(_0719_),
    .A(\daisychain[18] ));
 sg13g2_inv_1 _1051_ (.Y(_0720_),
    .A(\daisychain[19] ));
 sg13g2_inv_1 _1052_ (.Y(_0721_),
    .A(\daisychain[20] ));
 sg13g2_inv_1 _1053_ (.Y(_0722_),
    .A(\daisychain[21] ));
 sg13g2_inv_1 _1054_ (.Y(_0723_),
    .A(\daisychain[22] ));
 sg13g2_inv_1 _1055_ (.Y(_0724_),
    .A(\daisychain[23] ));
 sg13g2_inv_1 _1056_ (.Y(_0725_),
    .A(\daisychain[24] ));
 sg13g2_inv_1 _1057_ (.Y(_0726_),
    .A(\daisychain[25] ));
 sg13g2_inv_1 _1058_ (.Y(_0727_),
    .A(\daisychain[26] ));
 sg13g2_inv_1 _1059_ (.Y(_0728_),
    .A(\daisychain[27] ));
 sg13g2_inv_1 _1060_ (.Y(_0729_),
    .A(\daisychain[28] ));
 sg13g2_inv_1 _1061_ (.Y(_0730_),
    .A(\daisychain[29] ));
 sg13g2_inv_1 _1062_ (.Y(_0731_),
    .A(\daisychain[30] ));
 sg13g2_inv_1 _1063_ (.Y(_0732_),
    .A(\daisychain[31] ));
 sg13g2_inv_1 _1064_ (.Y(_0733_),
    .A(\daisychain[32] ));
 sg13g2_inv_1 _1065_ (.Y(_0734_),
    .A(\daisychain[33] ));
 sg13g2_inv_1 _1066_ (.Y(_0735_),
    .A(\daisychain[34] ));
 sg13g2_inv_1 _1067_ (.Y(_0736_),
    .A(\daisychain[35] ));
 sg13g2_inv_1 _1068_ (.Y(_0737_),
    .A(\daisychain[36] ));
 sg13g2_inv_1 _1069_ (.Y(_0738_),
    .A(\daisychain[37] ));
 sg13g2_inv_1 _1070_ (.Y(_0739_),
    .A(\daisychain[38] ));
 sg13g2_inv_1 _1071_ (.Y(_0740_),
    .A(\daisychain[39] ));
 sg13g2_inv_1 _1072_ (.Y(_0741_),
    .A(\daisychain[40] ));
 sg13g2_inv_1 _1073_ (.Y(_0742_),
    .A(\daisychain[41] ));
 sg13g2_inv_1 _1074_ (.Y(_0743_),
    .A(\daisychain[42] ));
 sg13g2_inv_1 _1075_ (.Y(_0744_),
    .A(\daisychain[43] ));
 sg13g2_inv_1 _1076_ (.Y(_0745_),
    .A(\daisychain[44] ));
 sg13g2_inv_1 _1077_ (.Y(_0746_),
    .A(\daisychain[45] ));
 sg13g2_inv_1 _1078_ (.Y(_0747_),
    .A(\daisychain[46] ));
 sg13g2_inv_1 _1079_ (.Y(_0748_),
    .A(\daisychain[47] ));
 sg13g2_inv_1 _1080_ (.Y(_0749_),
    .A(\daisychain[48] ));
 sg13g2_inv_1 _1081_ (.Y(_0750_),
    .A(\daisychain[49] ));
 sg13g2_inv_1 _1082_ (.Y(_0751_),
    .A(\daisychain[50] ));
 sg13g2_inv_1 _1083_ (.Y(_0752_),
    .A(\daisychain[51] ));
 sg13g2_inv_1 _1084_ (.Y(_0753_),
    .A(\daisychain[52] ));
 sg13g2_inv_1 _1085_ (.Y(_0754_),
    .A(\daisychain[53] ));
 sg13g2_inv_1 _1086_ (.Y(_0755_),
    .A(\daisychain[54] ));
 sg13g2_inv_1 _1087_ (.Y(_0756_),
    .A(\daisychain[55] ));
 sg13g2_inv_1 _1088_ (.Y(_0757_),
    .A(\daisychain[56] ));
 sg13g2_inv_1 _1089_ (.Y(_0758_),
    .A(\daisychain[57] ));
 sg13g2_inv_1 _1090_ (.Y(_0759_),
    .A(\daisychain[58] ));
 sg13g2_inv_1 _1091_ (.Y(_0760_),
    .A(\daisychain[59] ));
 sg13g2_inv_1 _1092_ (.Y(_0761_),
    .A(\daisychain[60] ));
 sg13g2_inv_1 _1093_ (.Y(_0762_),
    .A(\daisychain[61] ));
 sg13g2_inv_1 _1094_ (.Y(_0763_),
    .A(\daisychain[62] ));
 sg13g2_inv_1 _1095_ (.Y(_0764_),
    .A(\daisychain[63] ));
 sg13g2_inv_1 _1096_ (.Y(_0765_),
    .A(\daisychain[64] ));
 sg13g2_inv_1 _1097_ (.Y(_0766_),
    .A(\daisychain[65] ));
 sg13g2_inv_1 _1098_ (.Y(_0767_),
    .A(\daisychain[66] ));
 sg13g2_inv_1 _1099_ (.Y(_0768_),
    .A(\daisychain[67] ));
 sg13g2_inv_1 _1100_ (.Y(_0769_),
    .A(\daisychain[68] ));
 sg13g2_inv_1 _1101_ (.Y(_0770_),
    .A(\daisychain[69] ));
 sg13g2_inv_1 _1102_ (.Y(_0771_),
    .A(\daisychain[70] ));
 sg13g2_inv_1 _1103_ (.Y(_0772_),
    .A(\daisychain[71] ));
 sg13g2_inv_1 _1104_ (.Y(_0773_),
    .A(\daisychain[72] ));
 sg13g2_inv_1 _1105_ (.Y(_0774_),
    .A(\daisychain[73] ));
 sg13g2_inv_1 _1106_ (.Y(_0775_),
    .A(\daisychain[74] ));
 sg13g2_inv_1 _1107_ (.Y(_0776_),
    .A(\daisychain[75] ));
 sg13g2_inv_1 _1108_ (.Y(_0777_),
    .A(\daisychain[76] ));
 sg13g2_inv_1 _1109_ (.Y(_0778_),
    .A(\daisychain[77] ));
 sg13g2_inv_1 _1110_ (.Y(_0779_),
    .A(\daisychain[78] ));
 sg13g2_inv_1 _1111_ (.Y(_0780_),
    .A(\daisychain[79] ));
 sg13g2_inv_1 _1112_ (.Y(_0781_),
    .A(\daisychain[80] ));
 sg13g2_inv_1 _1113_ (.Y(_0782_),
    .A(\daisychain[81] ));
 sg13g2_inv_1 _1114_ (.Y(_0783_),
    .A(\daisychain[82] ));
 sg13g2_inv_1 _1115_ (.Y(_0784_),
    .A(\daisychain[83] ));
 sg13g2_inv_1 _1116_ (.Y(_0785_),
    .A(\daisychain[84] ));
 sg13g2_inv_1 _1117_ (.Y(_0786_),
    .A(\daisychain[85] ));
 sg13g2_inv_1 _1118_ (.Y(_0787_),
    .A(\daisychain[86] ));
 sg13g2_inv_1 _1119_ (.Y(_0788_),
    .A(\daisychain[87] ));
 sg13g2_inv_1 _1120_ (.Y(_0789_),
    .A(\daisychain[88] ));
 sg13g2_inv_1 _1121_ (.Y(_0790_),
    .A(\daisychain[89] ));
 sg13g2_inv_1 _1122_ (.Y(_0791_),
    .A(\daisychain[90] ));
 sg13g2_inv_1 _1123_ (.Y(_0792_),
    .A(\daisychain[91] ));
 sg13g2_inv_1 _1124_ (.Y(_0793_),
    .A(\daisychain[92] ));
 sg13g2_inv_1 _1125_ (.Y(_0794_),
    .A(\daisychain[93] ));
 sg13g2_inv_1 _1126_ (.Y(_0795_),
    .A(\daisychain[94] ));
 sg13g2_inv_1 _1127_ (.Y(_0796_),
    .A(\daisychain[95] ));
 sg13g2_inv_1 _1128_ (.Y(_0797_),
    .A(\daisychain[96] ));
 sg13g2_inv_1 _1129_ (.Y(_0798_),
    .A(\daisychain[97] ));
 sg13g2_inv_1 _1130_ (.Y(_0799_),
    .A(\daisychain[98] ));
 sg13g2_inv_1 _1131_ (.Y(_0800_),
    .A(\daisychain[99] ));
 sg13g2_inv_1 _1132_ (.Y(_0801_),
    .A(\daisychain[100] ));
 sg13g2_inv_1 _1133_ (.Y(_0802_),
    .A(\daisychain[101] ));
 sg13g2_inv_1 _1134_ (.Y(_0803_),
    .A(\daisychain[102] ));
 sg13g2_inv_1 _1135_ (.Y(_0804_),
    .A(\daisychain[103] ));
 sg13g2_inv_1 _1136_ (.Y(_0805_),
    .A(\daisychain[104] ));
 sg13g2_inv_1 _1137_ (.Y(_0806_),
    .A(\daisychain[105] ));
 sg13g2_inv_1 _1138_ (.Y(_0807_),
    .A(\daisychain[106] ));
 sg13g2_inv_1 _1139_ (.Y(_0808_),
    .A(\daisychain[107] ));
 sg13g2_inv_1 _1140_ (.Y(_0809_),
    .A(\daisychain[108] ));
 sg13g2_inv_1 _1141_ (.Y(_0810_),
    .A(\daisychain[109] ));
 sg13g2_inv_1 _1142_ (.Y(_0811_),
    .A(\daisychain[110] ));
 sg13g2_inv_1 _1143_ (.Y(_0812_),
    .A(\daisychain[111] ));
 sg13g2_inv_1 _1144_ (.Y(_0813_),
    .A(\daisychain[112] ));
 sg13g2_inv_1 _1145_ (.Y(_0814_),
    .A(\daisychain[113] ));
 sg13g2_inv_1 _1146_ (.Y(_0815_),
    .A(\daisychain[114] ));
 sg13g2_inv_1 _1147_ (.Y(_0816_),
    .A(\daisychain[115] ));
 sg13g2_inv_1 _1148_ (.Y(_0817_),
    .A(\daisychain[116] ));
 sg13g2_inv_1 _1149_ (.Y(_0818_),
    .A(\daisychain[117] ));
 sg13g2_inv_1 _1150_ (.Y(_0819_),
    .A(\daisychain[118] ));
 sg13g2_inv_1 _1151_ (.Y(_0820_),
    .A(\daisychain[119] ));
 sg13g2_inv_1 _1152_ (.Y(_0821_),
    .A(\daisychain[120] ));
 sg13g2_inv_1 _1153_ (.Y(_0822_),
    .A(\daisychain[121] ));
 sg13g2_inv_1 _1154_ (.Y(_0823_),
    .A(\daisychain[122] ));
 sg13g2_o21ai_1 _1155_ (.B1(net150),
    .Y(_0824_),
    .A1(net104),
    .A2(\state[0] ));
 sg13g2_a21o_1 _1156_ (.A2(_0701_),
    .A1(net104),
    .B1(_0824_),
    .X(_0825_));
 sg13g2_nor2_1 _1157_ (.A(net137),
    .B(net3),
    .Y(_0826_));
 sg13g2_a21oi_1 _1158_ (.A1(net68),
    .A2(net2),
    .Y(_0827_),
    .B1(net27));
 sg13g2_a22oi_1 _1159_ (.Y(_0128_),
    .B1(_0827_),
    .B2(_0825_),
    .A2(net37),
    .A1(_0701_));
 sg13g2_o21ai_1 _1160_ (.B1(net143),
    .Y(_0828_),
    .A1(net97),
    .A2(\state[1] ));
 sg13g2_a21o_1 _1161_ (.A2(_0702_),
    .A1(net97),
    .B1(_0828_),
    .X(_0829_));
 sg13g2_a21oi_1 _1162_ (.A1(net75),
    .A2(\daisychain[0] ),
    .Y(_0830_),
    .B1(net37));
 sg13g2_a22oi_1 _1163_ (.Y(_0129_),
    .B1(_0829_),
    .B2(_0830_),
    .A2(net38),
    .A1(_0702_));
 sg13g2_o21ai_1 _1164_ (.B1(net147),
    .Y(_0831_),
    .A1(net101),
    .A2(\state[2] ));
 sg13g2_a21o_1 _1165_ (.A2(_0703_),
    .A1(net101),
    .B1(_0831_),
    .X(_0832_));
 sg13g2_a21oi_1 _1166_ (.A1(net75),
    .A2(\daisychain[1] ),
    .Y(_0833_),
    .B1(net38));
 sg13g2_a22oi_1 _1167_ (.Y(_0130_),
    .B1(_0832_),
    .B2(_0833_),
    .A2(net38),
    .A1(_0703_));
 sg13g2_o21ai_1 _1168_ (.B1(net147),
    .Y(_0834_),
    .A1(net101),
    .A2(\state[3] ));
 sg13g2_a21o_1 _1169_ (.A2(_0704_),
    .A1(net102),
    .B1(_0834_),
    .X(_0835_));
 sg13g2_a21oi_1 _1170_ (.A1(net71),
    .A2(\daisychain[2] ),
    .Y(_0836_),
    .B1(net35));
 sg13g2_a22oi_1 _1171_ (.Y(_0131_),
    .B1(_0835_),
    .B2(_0836_),
    .A2(net35),
    .A1(_0704_));
 sg13g2_o21ai_1 _1172_ (.B1(net143),
    .Y(_0837_),
    .A1(net97),
    .A2(\state[4] ));
 sg13g2_a21o_1 _1173_ (.A2(_0705_),
    .A1(net97),
    .B1(_0837_),
    .X(_0838_));
 sg13g2_a21oi_1 _1174_ (.A1(net71),
    .A2(\daisychain[3] ),
    .Y(_0839_),
    .B1(net31));
 sg13g2_a22oi_1 _1175_ (.Y(_0132_),
    .B1(_0838_),
    .B2(_0839_),
    .A2(net31),
    .A1(_0705_));
 sg13g2_o21ai_1 _1176_ (.B1(net142),
    .Y(_0840_),
    .A1(net96),
    .A2(\state[5] ));
 sg13g2_a21o_1 _1177_ (.A2(_0706_),
    .A1(net96),
    .B1(_0840_),
    .X(_0841_));
 sg13g2_a21oi_1 _1178_ (.A1(net71),
    .A2(\daisychain[4] ),
    .Y(_0842_),
    .B1(net30));
 sg13g2_a22oi_1 _1179_ (.Y(_0133_),
    .B1(_0841_),
    .B2(_0842_),
    .A2(net30),
    .A1(_0706_));
 sg13g2_o21ai_1 _1180_ (.B1(net142),
    .Y(_0843_),
    .A1(net96),
    .A2(\state[6] ));
 sg13g2_a21o_1 _1181_ (.A2(_0707_),
    .A1(net96),
    .B1(_0843_),
    .X(_0844_));
 sg13g2_a21oi_1 _1182_ (.A1(net71),
    .A2(\daisychain[5] ),
    .Y(_0845_),
    .B1(net30));
 sg13g2_a22oi_1 _1183_ (.Y(_0134_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(net25),
    .A1(_0707_));
 sg13g2_o21ai_1 _1184_ (.B1(net139),
    .Y(_0846_),
    .A1(net92),
    .A2(\state[7] ));
 sg13g2_a21o_1 _1185_ (.A2(_0708_),
    .A1(net92),
    .B1(_0846_),
    .X(_0847_));
 sg13g2_a21oi_1 _1186_ (.A1(net68),
    .A2(\daisychain[6] ),
    .Y(_0848_),
    .B1(net25));
 sg13g2_a22oi_1 _1187_ (.Y(_0135_),
    .B1(_0847_),
    .B2(_0848_),
    .A2(net26),
    .A1(_0708_));
 sg13g2_o21ai_1 _1188_ (.B1(net139),
    .Y(_0849_),
    .A1(net92),
    .A2(\state[8] ));
 sg13g2_a21o_1 _1189_ (.A2(_0709_),
    .A1(net92),
    .B1(_0849_),
    .X(_0850_));
 sg13g2_a21oi_1 _1190_ (.A1(net68),
    .A2(\daisychain[7] ),
    .Y(_0851_),
    .B1(net25));
 sg13g2_a22oi_1 _1191_ (.Y(_0136_),
    .B1(_0850_),
    .B2(_0851_),
    .A2(net25),
    .A1(_0709_));
 sg13g2_o21ai_1 _1192_ (.B1(net139),
    .Y(_0852_),
    .A1(net92),
    .A2(\state[9] ));
 sg13g2_a21o_1 _1193_ (.A2(_0710_),
    .A1(net92),
    .B1(_0852_),
    .X(_0853_));
 sg13g2_a21oi_1 _1194_ (.A1(net68),
    .A2(\daisychain[8] ),
    .Y(_0854_),
    .B1(net25));
 sg13g2_a22oi_1 _1195_ (.Y(_0137_),
    .B1(_0853_),
    .B2(_0854_),
    .A2(net25),
    .A1(_0710_));
 sg13g2_o21ai_1 _1196_ (.B1(net139),
    .Y(_0855_),
    .A1(net92),
    .A2(\state[10] ));
 sg13g2_a21o_1 _1197_ (.A2(_0711_),
    .A1(net92),
    .B1(_0855_),
    .X(_0856_));
 sg13g2_a21oi_1 _1198_ (.A1(net68),
    .A2(\daisychain[9] ),
    .Y(_0857_),
    .B1(net25));
 sg13g2_a22oi_1 _1199_ (.Y(_0138_),
    .B1(_0856_),
    .B2(_0857_),
    .A2(net25),
    .A1(_0711_));
 sg13g2_o21ai_1 _1200_ (.B1(net139),
    .Y(_0858_),
    .A1(net93),
    .A2(\state[11] ));
 sg13g2_a21o_1 _1201_ (.A2(_0712_),
    .A1(net93),
    .B1(_0858_),
    .X(_0859_));
 sg13g2_a21oi_1 _1202_ (.A1(net68),
    .A2(\daisychain[10] ),
    .Y(_0860_),
    .B1(net26));
 sg13g2_a22oi_1 _1203_ (.Y(_0139_),
    .B1(_0859_),
    .B2(_0860_),
    .A2(net26),
    .A1(_0712_));
 sg13g2_o21ai_1 _1204_ (.B1(net142),
    .Y(_0861_),
    .A1(net96),
    .A2(\state[12] ));
 sg13g2_a21o_1 _1205_ (.A2(_0713_),
    .A1(net93),
    .B1(_0861_),
    .X(_0862_));
 sg13g2_a21oi_1 _1206_ (.A1(net68),
    .A2(\daisychain[11] ),
    .Y(_0863_),
    .B1(net26));
 sg13g2_a22oi_1 _1207_ (.Y(_0140_),
    .B1(_0862_),
    .B2(_0863_),
    .A2(net26),
    .A1(_0713_));
 sg13g2_o21ai_1 _1208_ (.B1(net142),
    .Y(_0864_),
    .A1(net96),
    .A2(\state[13] ));
 sg13g2_a21o_1 _1209_ (.A2(_0714_),
    .A1(net96),
    .B1(_0864_),
    .X(_0865_));
 sg13g2_a21oi_1 _1210_ (.A1(net71),
    .A2(\daisychain[12] ),
    .Y(_0866_),
    .B1(net30));
 sg13g2_a22oi_1 _1211_ (.Y(_0141_),
    .B1(_0865_),
    .B2(_0866_),
    .A2(net30),
    .A1(_0714_));
 sg13g2_o21ai_1 _1212_ (.B1(net143),
    .Y(_0867_),
    .A1(net97),
    .A2(\state[14] ));
 sg13g2_a21o_1 _1213_ (.A2(_0715_),
    .A1(net97),
    .B1(_0867_),
    .X(_0868_));
 sg13g2_a21oi_1 _1214_ (.A1(net74),
    .A2(\daisychain[13] ),
    .Y(_0869_),
    .B1(net30));
 sg13g2_a22oi_1 _1215_ (.Y(_0142_),
    .B1(_0868_),
    .B2(_0869_),
    .A2(net30),
    .A1(_0715_));
 sg13g2_o21ai_1 _1216_ (.B1(net143),
    .Y(_0870_),
    .A1(net97),
    .A2(\state[15] ));
 sg13g2_a21o_1 _1217_ (.A2(_0716_),
    .A1(net97),
    .B1(_0870_),
    .X(_0871_));
 sg13g2_a21oi_1 _1218_ (.A1(net74),
    .A2(\daisychain[14] ),
    .Y(_0872_),
    .B1(net31));
 sg13g2_a22oi_1 _1219_ (.Y(_0143_),
    .B1(_0871_),
    .B2(_0872_),
    .A2(net31),
    .A1(_0716_));
 sg13g2_o21ai_1 _1220_ (.B1(net142),
    .Y(_0873_),
    .A1(net96),
    .A2(\state[16] ));
 sg13g2_a21o_1 _1221_ (.A2(_0717_),
    .A1(net98),
    .B1(_0873_),
    .X(_0874_));
 sg13g2_a21oi_1 _1222_ (.A1(net71),
    .A2(\daisychain[15] ),
    .Y(_0875_),
    .B1(net30));
 sg13g2_a22oi_1 _1223_ (.Y(_0144_),
    .B1(_0874_),
    .B2(_0875_),
    .A2(net32),
    .A1(_0717_));
 sg13g2_o21ai_1 _1224_ (.B1(net145),
    .Y(_0876_),
    .A1(net98),
    .A2(\state[17] ));
 sg13g2_a21o_1 _1225_ (.A2(_0718_),
    .A1(net98),
    .B1(_0876_),
    .X(_0877_));
 sg13g2_a21oi_1 _1226_ (.A1(net71),
    .A2(\daisychain[16] ),
    .Y(_0878_),
    .B1(net32));
 sg13g2_a22oi_1 _1227_ (.Y(_0145_),
    .B1(_0877_),
    .B2(_0878_),
    .A2(net32),
    .A1(_0718_));
 sg13g2_o21ai_1 _1228_ (.B1(net145),
    .Y(_0879_),
    .A1(net98),
    .A2(\state[18] ));
 sg13g2_a21o_1 _1229_ (.A2(_0719_),
    .A1(net98),
    .B1(_0879_),
    .X(_0880_));
 sg13g2_a21oi_1 _1230_ (.A1(net71),
    .A2(\daisychain[17] ),
    .Y(_0881_),
    .B1(net32));
 sg13g2_a22oi_1 _1231_ (.Y(_0146_),
    .B1(_0880_),
    .B2(_0881_),
    .A2(net32),
    .A1(_0719_));
 sg13g2_o21ai_1 _1232_ (.B1(net146),
    .Y(_0882_),
    .A1(net99),
    .A2(\state[19] ));
 sg13g2_a21o_1 _1233_ (.A2(_0720_),
    .A1(net99),
    .B1(_0882_),
    .X(_0883_));
 sg13g2_a21oi_1 _1234_ (.A1(net72),
    .A2(\daisychain[18] ),
    .Y(_0884_),
    .B1(net34));
 sg13g2_a22oi_1 _1235_ (.Y(_0147_),
    .B1(_0883_),
    .B2(_0884_),
    .A2(net34),
    .A1(_0720_));
 sg13g2_o21ai_1 _1236_ (.B1(net147),
    .Y(_0885_),
    .A1(net101),
    .A2(\state[20] ));
 sg13g2_a21o_1 _1237_ (.A2(_0721_),
    .A1(net101),
    .B1(_0885_),
    .X(_0886_));
 sg13g2_a21oi_1 _1238_ (.A1(net72),
    .A2(\daisychain[19] ),
    .Y(_0887_),
    .B1(net34));
 sg13g2_a22oi_1 _1239_ (.Y(_0148_),
    .B1(_0886_),
    .B2(_0887_),
    .A2(net35),
    .A1(_0721_));
 sg13g2_o21ai_1 _1240_ (.B1(net147),
    .Y(_0888_),
    .A1(net101),
    .A2(\state[21] ));
 sg13g2_a21o_1 _1241_ (.A2(_0722_),
    .A1(net101),
    .B1(_0888_),
    .X(_0889_));
 sg13g2_a21oi_1 _1242_ (.A1(net74),
    .A2(\daisychain[20] ),
    .Y(_0890_),
    .B1(net31));
 sg13g2_a22oi_1 _1243_ (.Y(_0149_),
    .B1(_0889_),
    .B2(_0890_),
    .A2(net31),
    .A1(_0722_));
 sg13g2_o21ai_1 _1244_ (.B1(net147),
    .Y(_0891_),
    .A1(net102),
    .A2(\state[22] ));
 sg13g2_a21o_1 _1245_ (.A2(_0723_),
    .A1(net101),
    .B1(_0891_),
    .X(_0892_));
 sg13g2_a21oi_1 _1246_ (.A1(net73),
    .A2(\daisychain[21] ),
    .Y(_0893_),
    .B1(net35));
 sg13g2_a22oi_1 _1247_ (.Y(_0150_),
    .B1(_0892_),
    .B2(_0893_),
    .A2(net35),
    .A1(_0723_));
 sg13g2_o21ai_1 _1248_ (.B1(net148),
    .Y(_0894_),
    .A1(net102),
    .A2(\state[23] ));
 sg13g2_a21o_1 _1249_ (.A2(_0724_),
    .A1(net102),
    .B1(_0894_),
    .X(_0895_));
 sg13g2_a21oi_1 _1250_ (.A1(net73),
    .A2(\daisychain[22] ),
    .Y(_0896_),
    .B1(net35));
 sg13g2_a22oi_1 _1251_ (.Y(_0151_),
    .B1(_0895_),
    .B2(_0896_),
    .A2(net35),
    .A1(_0724_));
 sg13g2_o21ai_1 _1252_ (.B1(net148),
    .Y(_0897_),
    .A1(net102),
    .A2(\state[24] ));
 sg13g2_a21o_1 _1253_ (.A2(_0725_),
    .A1(net102),
    .B1(_0897_),
    .X(_0384_));
 sg13g2_a21oi_1 _1254_ (.A1(net73),
    .A2(\daisychain[23] ),
    .Y(_0385_),
    .B1(net35));
 sg13g2_a22oi_1 _1255_ (.Y(_0152_),
    .B1(_0384_),
    .B2(_0385_),
    .A2(net36),
    .A1(_0725_));
 sg13g2_o21ai_1 _1256_ (.B1(net146),
    .Y(_0386_),
    .A1(net99),
    .A2(\state[25] ));
 sg13g2_a21o_1 _1257_ (.A2(_0726_),
    .A1(net99),
    .B1(_0386_),
    .X(_0387_));
 sg13g2_a21oi_1 _1258_ (.A1(net72),
    .A2(\daisychain[24] ),
    .Y(_0388_),
    .B1(net36));
 sg13g2_a22oi_1 _1259_ (.Y(_0153_),
    .B1(_0387_),
    .B2(_0388_),
    .A2(net33),
    .A1(_0726_));
 sg13g2_o21ai_1 _1260_ (.B1(net146),
    .Y(_0389_),
    .A1(net99),
    .A2(\state[26] ));
 sg13g2_a21o_1 _1261_ (.A2(_0727_),
    .A1(net99),
    .B1(_0389_),
    .X(_0390_));
 sg13g2_a21oi_1 _1262_ (.A1(net72),
    .A2(\daisychain[25] ),
    .Y(_0391_),
    .B1(net33));
 sg13g2_a22oi_1 _1263_ (.Y(_0154_),
    .B1(_0390_),
    .B2(_0391_),
    .A2(net33),
    .A1(_0727_));
 sg13g2_o21ai_1 _1264_ (.B1(net146),
    .Y(_0392_),
    .A1(net99),
    .A2(\state[27] ));
 sg13g2_a21o_1 _1265_ (.A2(_0728_),
    .A1(net99),
    .B1(_0392_),
    .X(_0393_));
 sg13g2_a21oi_1 _1266_ (.A1(net72),
    .A2(\daisychain[26] ),
    .Y(_0394_),
    .B1(net34));
 sg13g2_a22oi_1 _1267_ (.Y(_0155_),
    .B1(_0393_),
    .B2(_0394_),
    .A2(net34),
    .A1(_0728_));
 sg13g2_o21ai_1 _1268_ (.B1(net146),
    .Y(_0395_),
    .A1(net100),
    .A2(\state[28] ));
 sg13g2_a21o_1 _1269_ (.A2(_0729_),
    .A1(net100),
    .B1(_0395_),
    .X(_0396_));
 sg13g2_a21oi_1 _1270_ (.A1(net72),
    .A2(\daisychain[27] ),
    .Y(_0397_),
    .B1(net34));
 sg13g2_a22oi_1 _1271_ (.Y(_0156_),
    .B1(_0396_),
    .B2(_0397_),
    .A2(net33),
    .A1(_0729_));
 sg13g2_o21ai_1 _1272_ (.B1(net146),
    .Y(_0398_),
    .A1(net100),
    .A2(\state[29] ));
 sg13g2_a21o_1 _1273_ (.A2(_0730_),
    .A1(net100),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_a21oi_1 _1274_ (.A1(net72),
    .A2(\daisychain[28] ),
    .Y(_0400_),
    .B1(net33));
 sg13g2_a22oi_1 _1275_ (.Y(_0157_),
    .B1(_0399_),
    .B2(_0400_),
    .A2(net33),
    .A1(_0730_));
 sg13g2_o21ai_1 _1276_ (.B1(net158),
    .Y(_0401_),
    .A1(net112),
    .A2(\state[30] ));
 sg13g2_a21o_1 _1277_ (.A2(_0731_),
    .A1(net112),
    .B1(_0401_),
    .X(_0402_));
 sg13g2_a21oi_1 _1278_ (.A1(net72),
    .A2(\daisychain[29] ),
    .Y(_0403_),
    .B1(net33));
 sg13g2_a22oi_1 _1279_ (.Y(_0158_),
    .B1(_0402_),
    .B2(_0403_),
    .A2(net45),
    .A1(_0731_));
 sg13g2_o21ai_1 _1280_ (.B1(net158),
    .Y(_0404_),
    .A1(net112),
    .A2(\state[31] ));
 sg13g2_a21o_1 _1281_ (.A2(_0732_),
    .A1(net112),
    .B1(_0404_),
    .X(_0405_));
 sg13g2_a21oi_1 _1282_ (.A1(net79),
    .A2(\daisychain[30] ),
    .Y(_0406_),
    .B1(net45));
 sg13g2_a22oi_1 _1283_ (.Y(_0159_),
    .B1(_0405_),
    .B2(_0406_),
    .A2(net45),
    .A1(_0732_));
 sg13g2_o21ai_1 _1284_ (.B1(net158),
    .Y(_0407_),
    .A1(net112),
    .A2(\state[32] ));
 sg13g2_a21o_1 _1285_ (.A2(_0733_),
    .A1(net112),
    .B1(_0407_),
    .X(_0408_));
 sg13g2_a21oi_1 _1286_ (.A1(net79),
    .A2(\daisychain[31] ),
    .Y(_0409_),
    .B1(net45));
 sg13g2_a22oi_1 _1287_ (.Y(_0160_),
    .B1(_0408_),
    .B2(_0409_),
    .A2(net45),
    .A1(_0733_));
 sg13g2_o21ai_1 _1288_ (.B1(net158),
    .Y(_0410_),
    .A1(net112),
    .A2(\state[33] ));
 sg13g2_a21o_1 _1289_ (.A2(_0734_),
    .A1(net112),
    .B1(_0410_),
    .X(_0411_));
 sg13g2_a21oi_1 _1290_ (.A1(net79),
    .A2(\daisychain[32] ),
    .Y(_0412_),
    .B1(net45));
 sg13g2_a22oi_1 _1291_ (.Y(_0161_),
    .B1(_0411_),
    .B2(_0412_),
    .A2(net45),
    .A1(_0734_));
 sg13g2_o21ai_1 _1292_ (.B1(net158),
    .Y(_0413_),
    .A1(net113),
    .A2(\state[34] ));
 sg13g2_a21o_1 _1293_ (.A2(_0735_),
    .A1(net113),
    .B1(_0413_),
    .X(_0414_));
 sg13g2_a21oi_1 _1294_ (.A1(net73),
    .A2(\daisychain[33] ),
    .Y(_0415_),
    .B1(net33));
 sg13g2_a22oi_1 _1295_ (.Y(_0162_),
    .B1(_0414_),
    .B2(_0415_),
    .A2(net36),
    .A1(_0735_));
 sg13g2_o21ai_1 _1296_ (.B1(net161),
    .Y(_0416_),
    .A1(net102),
    .A2(\state[35] ));
 sg13g2_a21o_1 _1297_ (.A2(_0736_),
    .A1(net103),
    .B1(_0416_),
    .X(_0417_));
 sg13g2_a21oi_1 _1298_ (.A1(net73),
    .A2(\daisychain[34] ),
    .Y(_0418_),
    .B1(net34));
 sg13g2_a22oi_1 _1299_ (.Y(_0163_),
    .B1(_0417_),
    .B2(_0418_),
    .A2(net36),
    .A1(_0736_));
 sg13g2_o21ai_1 _1300_ (.B1(net161),
    .Y(_0419_),
    .A1(net115),
    .A2(\state[36] ));
 sg13g2_a21o_1 _1301_ (.A2(_0737_),
    .A1(net115),
    .B1(_0419_),
    .X(_0420_));
 sg13g2_a21oi_1 _1302_ (.A1(net80),
    .A2(\daisychain[35] ),
    .Y(_0421_),
    .B1(net48));
 sg13g2_a22oi_1 _1303_ (.Y(_0164_),
    .B1(_0420_),
    .B2(_0421_),
    .A2(net48),
    .A1(_0737_));
 sg13g2_o21ai_1 _1304_ (.B1(net161),
    .Y(_0422_),
    .A1(net115),
    .A2(\state[37] ));
 sg13g2_a21o_1 _1305_ (.A2(_0738_),
    .A1(net115),
    .B1(_0422_),
    .X(_0423_));
 sg13g2_a21oi_1 _1306_ (.A1(net80),
    .A2(\daisychain[36] ),
    .Y(_0424_),
    .B1(net48));
 sg13g2_a22oi_1 _1307_ (.Y(_0165_),
    .B1(_0423_),
    .B2(_0424_),
    .A2(net48),
    .A1(_0738_));
 sg13g2_o21ai_1 _1308_ (.B1(net161),
    .Y(_0425_),
    .A1(net115),
    .A2(\state[38] ));
 sg13g2_a21o_1 _1309_ (.A2(_0739_),
    .A1(net113),
    .B1(_0425_),
    .X(_0426_));
 sg13g2_a21oi_1 _1310_ (.A1(net80),
    .A2(\daisychain[37] ),
    .Y(_0427_),
    .B1(net48));
 sg13g2_a22oi_1 _1311_ (.Y(_0166_),
    .B1(_0426_),
    .B2(_0427_),
    .A2(net48),
    .A1(_0739_));
 sg13g2_o21ai_1 _1312_ (.B1(net159),
    .Y(_0428_),
    .A1(net113),
    .A2(\state[39] ));
 sg13g2_a21o_1 _1313_ (.A2(_0740_),
    .A1(net113),
    .B1(_0428_),
    .X(_0429_));
 sg13g2_a21oi_1 _1314_ (.A1(net79),
    .A2(\daisychain[38] ),
    .Y(_0430_),
    .B1(net45));
 sg13g2_a22oi_1 _1315_ (.Y(_0167_),
    .B1(_0429_),
    .B2(_0430_),
    .A2(net47),
    .A1(_0740_));
 sg13g2_o21ai_1 _1316_ (.B1(net159),
    .Y(_0431_),
    .A1(net113),
    .A2(\state[40] ));
 sg13g2_a21o_1 _1317_ (.A2(_0741_),
    .A1(net113),
    .B1(_0431_),
    .X(_0432_));
 sg13g2_a21oi_1 _1318_ (.A1(net79),
    .A2(\daisychain[39] ),
    .Y(_0433_),
    .B1(net46));
 sg13g2_a22oi_1 _1319_ (.Y(_0168_),
    .B1(_0432_),
    .B2(_0433_),
    .A2(net46),
    .A1(_0741_));
 sg13g2_o21ai_1 _1320_ (.B1(net159),
    .Y(_0434_),
    .A1(net114),
    .A2(\state[41] ));
 sg13g2_a21o_1 _1321_ (.A2(_0742_),
    .A1(net114),
    .B1(_0434_),
    .X(_0435_));
 sg13g2_a21oi_1 _1322_ (.A1(net79),
    .A2(\daisychain[40] ),
    .Y(_0436_),
    .B1(net46));
 sg13g2_a22oi_1 _1323_ (.Y(_0169_),
    .B1(_0435_),
    .B2(_0436_),
    .A2(net46),
    .A1(_0742_));
 sg13g2_o21ai_1 _1324_ (.B1(net159),
    .Y(_0437_),
    .A1(net114),
    .A2(\state[42] ));
 sg13g2_a21o_1 _1325_ (.A2(_0743_),
    .A1(net114),
    .B1(_0437_),
    .X(_0438_));
 sg13g2_a21oi_1 _1326_ (.A1(net79),
    .A2(\daisychain[41] ),
    .Y(_0439_),
    .B1(net46));
 sg13g2_a22oi_1 _1327_ (.Y(_0170_),
    .B1(_0438_),
    .B2(_0439_),
    .A2(net46),
    .A1(_0743_));
 sg13g2_o21ai_1 _1328_ (.B1(net163),
    .Y(_0440_),
    .A1(net119),
    .A2(\state[43] ));
 sg13g2_a21o_1 _1329_ (.A2(_0744_),
    .A1(net119),
    .B1(_0440_),
    .X(_0441_));
 sg13g2_a21oi_1 _1330_ (.A1(net79),
    .A2(\daisychain[42] ),
    .Y(_0442_),
    .B1(net46));
 sg13g2_a22oi_1 _1331_ (.Y(_0171_),
    .B1(_0441_),
    .B2(_0442_),
    .A2(net46),
    .A1(_0744_));
 sg13g2_o21ai_1 _1332_ (.B1(net163),
    .Y(_0443_),
    .A1(net119),
    .A2(\state[44] ));
 sg13g2_a21o_1 _1333_ (.A2(_0745_),
    .A1(net119),
    .B1(_0443_),
    .X(_0444_));
 sg13g2_a21oi_1 _1334_ (.A1(net81),
    .A2(\daisychain[43] ),
    .Y(_0445_),
    .B1(net50));
 sg13g2_a22oi_1 _1335_ (.Y(_0172_),
    .B1(_0444_),
    .B2(_0445_),
    .A2(net50),
    .A1(_0745_));
 sg13g2_o21ai_1 _1336_ (.B1(net163),
    .Y(_0446_),
    .A1(net119),
    .A2(\state[45] ));
 sg13g2_a21o_1 _1337_ (.A2(_0746_),
    .A1(net119),
    .B1(_0446_),
    .X(_0447_));
 sg13g2_a21oi_1 _1338_ (.A1(net81),
    .A2(\daisychain[44] ),
    .Y(_0448_),
    .B1(net50));
 sg13g2_a22oi_1 _1339_ (.Y(_0173_),
    .B1(_0447_),
    .B2(_0448_),
    .A2(net51),
    .A1(_0746_));
 sg13g2_o21ai_1 _1340_ (.B1(net162),
    .Y(_0449_),
    .A1(net115),
    .A2(\state[46] ));
 sg13g2_a21o_1 _1341_ (.A2(_0747_),
    .A1(net115),
    .B1(_0449_),
    .X(_0450_));
 sg13g2_a21oi_1 _1342_ (.A1(net80),
    .A2(\daisychain[45] ),
    .Y(_0451_),
    .B1(net47));
 sg13g2_a22oi_1 _1343_ (.Y(_0174_),
    .B1(_0450_),
    .B2(_0451_),
    .A2(net48),
    .A1(_0747_));
 sg13g2_o21ai_1 _1344_ (.B1(net162),
    .Y(_0452_),
    .A1(net115),
    .A2(\state[47] ));
 sg13g2_a21o_1 _1345_ (.A2(_0748_),
    .A1(net116),
    .B1(_0452_),
    .X(_0453_));
 sg13g2_a21oi_1 _1346_ (.A1(net80),
    .A2(\daisychain[46] ),
    .Y(_0454_),
    .B1(net48));
 sg13g2_a22oi_1 _1347_ (.Y(_0175_),
    .B1(_0453_),
    .B2(_0454_),
    .A2(net49),
    .A1(_0748_));
 sg13g2_o21ai_1 _1348_ (.B1(net162),
    .Y(_0455_),
    .A1(net116),
    .A2(\state[48] ));
 sg13g2_a21o_1 _1349_ (.A2(_0749_),
    .A1(net116),
    .B1(_0455_),
    .X(_0456_));
 sg13g2_a21oi_1 _1350_ (.A1(net80),
    .A2(\daisychain[47] ),
    .Y(_0457_),
    .B1(net49));
 sg13g2_a22oi_1 _1351_ (.Y(_0176_),
    .B1(_0456_),
    .B2(_0457_),
    .A2(net49),
    .A1(_0749_));
 sg13g2_o21ai_1 _1352_ (.B1(net167),
    .Y(_0458_),
    .A1(net120),
    .A2(\state[49] ));
 sg13g2_a21o_1 _1353_ (.A2(_0750_),
    .A1(net120),
    .B1(_0458_),
    .X(_0459_));
 sg13g2_a21oi_1 _1354_ (.A1(net83),
    .A2(\daisychain[48] ),
    .Y(_0460_),
    .B1(net54));
 sg13g2_a22oi_1 _1355_ (.Y(_0177_),
    .B1(_0459_),
    .B2(_0460_),
    .A2(net54),
    .A1(_0750_));
 sg13g2_o21ai_1 _1356_ (.B1(net167),
    .Y(_0461_),
    .A1(net120),
    .A2(\state[50] ));
 sg13g2_a21o_1 _1357_ (.A2(_0751_),
    .A1(net120),
    .B1(_0461_),
    .X(_0462_));
 sg13g2_a21oi_1 _1358_ (.A1(net83),
    .A2(\daisychain[49] ),
    .Y(_0463_),
    .B1(net54));
 sg13g2_a22oi_1 _1359_ (.Y(_0178_),
    .B1(_0462_),
    .B2(_0463_),
    .A2(net54),
    .A1(_0751_));
 sg13g2_o21ai_1 _1360_ (.B1(net167),
    .Y(_0464_),
    .A1(net120),
    .A2(\state[51] ));
 sg13g2_a21o_1 _1361_ (.A2(_0752_),
    .A1(net120),
    .B1(_0464_),
    .X(_0465_));
 sg13g2_a21oi_1 _1362_ (.A1(net83),
    .A2(\daisychain[50] ),
    .Y(_0466_),
    .B1(net54));
 sg13g2_a22oi_1 _1363_ (.Y(_0179_),
    .B1(_0465_),
    .B2(_0466_),
    .A2(net54),
    .A1(_0752_));
 sg13g2_o21ai_1 _1364_ (.B1(net164),
    .Y(_0467_),
    .A1(net118),
    .A2(\state[52] ));
 sg13g2_a21o_1 _1365_ (.A2(_0753_),
    .A1(net118),
    .B1(_0467_),
    .X(_0468_));
 sg13g2_a21oi_1 _1366_ (.A1(net81),
    .A2(\daisychain[51] ),
    .Y(_0469_),
    .B1(net51));
 sg13g2_a22oi_1 _1367_ (.Y(_0180_),
    .B1(_0468_),
    .B2(_0469_),
    .A2(net51),
    .A1(_0753_));
 sg13g2_o21ai_1 _1368_ (.B1(net165),
    .Y(_0470_),
    .A1(net118),
    .A2(\state[53] ));
 sg13g2_a21o_1 _1369_ (.A2(_0754_),
    .A1(net119),
    .B1(_0470_),
    .X(_0471_));
 sg13g2_a21oi_1 _1370_ (.A1(net81),
    .A2(\daisychain[52] ),
    .Y(_0472_),
    .B1(net51));
 sg13g2_a22oi_1 _1371_ (.Y(_0181_),
    .B1(_0471_),
    .B2(_0472_),
    .A2(net51),
    .A1(_0754_));
 sg13g2_o21ai_1 _1372_ (.B1(net164),
    .Y(_0473_),
    .A1(net117),
    .A2(\state[54] ));
 sg13g2_a21o_1 _1373_ (.A2(_0755_),
    .A1(net117),
    .B1(_0473_),
    .X(_0474_));
 sg13g2_a21oi_1 _1374_ (.A1(net81),
    .A2(\daisychain[53] ),
    .Y(_0475_),
    .B1(net51));
 sg13g2_a22oi_1 _1375_ (.Y(_0182_),
    .B1(_0474_),
    .B2(_0475_),
    .A2(net50),
    .A1(_0755_));
 sg13g2_o21ai_1 _1376_ (.B1(net164),
    .Y(_0476_),
    .A1(net117),
    .A2(\state[55] ));
 sg13g2_a21o_1 _1377_ (.A2(_0756_),
    .A1(net119),
    .B1(_0476_),
    .X(_0477_));
 sg13g2_a21oi_1 _1378_ (.A1(net81),
    .A2(\daisychain[54] ),
    .Y(_0478_),
    .B1(net50));
 sg13g2_a22oi_1 _1379_ (.Y(_0183_),
    .B1(_0477_),
    .B2(_0478_),
    .A2(net50),
    .A1(_0756_));
 sg13g2_o21ai_1 _1380_ (.B1(net164),
    .Y(_0479_),
    .A1(net117),
    .A2(\state[56] ));
 sg13g2_a21o_1 _1381_ (.A2(_0757_),
    .A1(net117),
    .B1(_0479_),
    .X(_0480_));
 sg13g2_a21oi_1 _1382_ (.A1(net81),
    .A2(\daisychain[55] ),
    .Y(_0481_),
    .B1(net50));
 sg13g2_a22oi_1 _1383_ (.Y(_0184_),
    .B1(_0480_),
    .B2(_0481_),
    .A2(net50),
    .A1(_0757_));
 sg13g2_o21ai_1 _1384_ (.B1(net164),
    .Y(_0482_),
    .A1(net117),
    .A2(\state[57] ));
 sg13g2_a21o_1 _1385_ (.A2(_0758_),
    .A1(net117),
    .B1(_0482_),
    .X(_0483_));
 sg13g2_a21oi_1 _1386_ (.A1(net81),
    .A2(\daisychain[56] ),
    .Y(_0484_),
    .B1(net52));
 sg13g2_a22oi_1 _1387_ (.Y(_0185_),
    .B1(_0483_),
    .B2(_0484_),
    .A2(net52),
    .A1(_0758_));
 sg13g2_o21ai_1 _1388_ (.B1(net164),
    .Y(_0485_),
    .A1(net117),
    .A2(\state[58] ));
 sg13g2_a21o_1 _1389_ (.A2(_0759_),
    .A1(net118),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_a21oi_1 _1390_ (.A1(net82),
    .A2(\daisychain[57] ),
    .Y(_0487_),
    .B1(net52));
 sg13g2_a22oi_1 _1391_ (.Y(_0186_),
    .B1(_0486_),
    .B2(_0487_),
    .A2(net52),
    .A1(_0759_));
 sg13g2_o21ai_1 _1392_ (.B1(net165),
    .Y(_0488_),
    .A1(net118),
    .A2(\state[59] ));
 sg13g2_a21o_1 _1393_ (.A2(_0760_),
    .A1(net118),
    .B1(_0488_),
    .X(_0489_));
 sg13g2_a21oi_1 _1394_ (.A1(net82),
    .A2(\daisychain[58] ),
    .Y(_0490_),
    .B1(net52));
 sg13g2_a22oi_1 _1395_ (.Y(_0187_),
    .B1(_0489_),
    .B2(_0490_),
    .A2(net52),
    .A1(_0760_));
 sg13g2_o21ai_1 _1396_ (.B1(net165),
    .Y(_0491_),
    .A1(net118),
    .A2(\state[60] ));
 sg13g2_a21o_1 _1397_ (.A2(_0761_),
    .A1(net122),
    .B1(_0491_),
    .X(_0492_));
 sg13g2_a21oi_1 _1398_ (.A1(net82),
    .A2(\daisychain[59] ),
    .Y(_0493_),
    .B1(net52));
 sg13g2_a22oi_1 _1399_ (.Y(_0188_),
    .B1(_0492_),
    .B2(_0493_),
    .A2(net52),
    .A1(_0761_));
 sg13g2_o21ai_1 _1400_ (.B1(net167),
    .Y(_0494_),
    .A1(net120),
    .A2(\state[61] ));
 sg13g2_a21o_1 _1401_ (.A2(_0762_),
    .A1(net120),
    .B1(_0494_),
    .X(_0495_));
 sg13g2_a21oi_1 _1402_ (.A1(net82),
    .A2(\daisychain[60] ),
    .Y(_0496_),
    .B1(net53));
 sg13g2_a22oi_1 _1403_ (.Y(_0189_),
    .B1(_0495_),
    .B2(_0496_),
    .A2(net54),
    .A1(_0762_));
 sg13g2_o21ai_1 _1404_ (.B1(net167),
    .Y(_0497_),
    .A1(net121),
    .A2(\state[62] ));
 sg13g2_a21o_1 _1405_ (.A2(_0763_),
    .A1(net121),
    .B1(_0497_),
    .X(_0498_));
 sg13g2_a21oi_1 _1406_ (.A1(net83),
    .A2(\daisychain[61] ),
    .Y(_0499_),
    .B1(net54));
 sg13g2_a22oi_1 _1407_ (.Y(_0190_),
    .B1(_0498_),
    .B2(_0499_),
    .A2(net55),
    .A1(_0763_));
 sg13g2_o21ai_1 _1408_ (.B1(net168),
    .Y(_0500_),
    .A1(net121),
    .A2(\state[63] ));
 sg13g2_a21o_1 _1409_ (.A2(_0764_),
    .A1(net121),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_a21oi_1 _1410_ (.A1(net83),
    .A2(\daisychain[62] ),
    .Y(_0502_),
    .B1(net55));
 sg13g2_a22oi_1 _1411_ (.Y(_0191_),
    .B1(_0501_),
    .B2(_0502_),
    .A2(net55),
    .A1(_0764_));
 sg13g2_o21ai_1 _1412_ (.B1(net175),
    .Y(_0503_),
    .A1(net128),
    .A2(\state[64] ));
 sg13g2_a21o_1 _1413_ (.A2(_0765_),
    .A1(net128),
    .B1(_0503_),
    .X(_0504_));
 sg13g2_a21oi_1 _1414_ (.A1(net87),
    .A2(\daisychain[63] ),
    .Y(_0505_),
    .B1(net61));
 sg13g2_a22oi_1 _1415_ (.Y(_0192_),
    .B1(_0504_),
    .B2(_0505_),
    .A2(net61),
    .A1(_0765_));
 sg13g2_o21ai_1 _1416_ (.B1(net175),
    .Y(_0506_),
    .A1(net129),
    .A2(\state[65] ));
 sg13g2_a21o_1 _1417_ (.A2(_0766_),
    .A1(net129),
    .B1(_0506_),
    .X(_0507_));
 sg13g2_a21oi_1 _1418_ (.A1(net87),
    .A2(\daisychain[64] ),
    .Y(_0508_),
    .B1(net62));
 sg13g2_a22oi_1 _1419_ (.Y(_0193_),
    .B1(_0507_),
    .B2(_0508_),
    .A2(net62),
    .A1(_0766_));
 sg13g2_o21ai_1 _1420_ (.B1(net176),
    .Y(_0509_),
    .A1(net129),
    .A2(\state[66] ));
 sg13g2_a21o_1 _1421_ (.A2(_0767_),
    .A1(net129),
    .B1(_0509_),
    .X(_0510_));
 sg13g2_a21oi_1 _1422_ (.A1(net87),
    .A2(\daisychain[65] ),
    .Y(_0511_),
    .B1(net62));
 sg13g2_a22oi_1 _1423_ (.Y(_0194_),
    .B1(_0510_),
    .B2(_0511_),
    .A2(net62),
    .A1(_0767_));
 sg13g2_o21ai_1 _1424_ (.B1(net178),
    .Y(_0512_),
    .A1(net131),
    .A2(\state[67] ));
 sg13g2_a21o_1 _1425_ (.A2(_0768_),
    .A1(net131),
    .B1(_0512_),
    .X(_0513_));
 sg13g2_a21oi_1 _1426_ (.A1(net86),
    .A2(\daisychain[66] ),
    .Y(_0514_),
    .B1(net64));
 sg13g2_a22oi_1 _1427_ (.Y(_0195_),
    .B1(_0513_),
    .B2(_0514_),
    .A2(net64),
    .A1(_0768_));
 sg13g2_o21ai_1 _1428_ (.B1(net178),
    .Y(_0515_),
    .A1(net131),
    .A2(\state[68] ));
 sg13g2_a21o_1 _1429_ (.A2(_0769_),
    .A1(net131),
    .B1(_0515_),
    .X(_0516_));
 sg13g2_a21oi_1 _1430_ (.A1(net86),
    .A2(\daisychain[67] ),
    .Y(_0517_),
    .B1(net64));
 sg13g2_a22oi_1 _1431_ (.Y(_0196_),
    .B1(_0516_),
    .B2(_0517_),
    .A2(net64),
    .A1(_0769_));
 sg13g2_o21ai_1 _1432_ (.B1(net178),
    .Y(_0518_),
    .A1(net131),
    .A2(\state[69] ));
 sg13g2_a21o_1 _1433_ (.A2(_0770_),
    .A1(net131),
    .B1(_0518_),
    .X(_0519_));
 sg13g2_a21oi_1 _1434_ (.A1(net86),
    .A2(\daisychain[68] ),
    .Y(_0520_),
    .B1(net64));
 sg13g2_a22oi_1 _1435_ (.Y(_0197_),
    .B1(_0519_),
    .B2(_0520_),
    .A2(net64),
    .A1(_0770_));
 sg13g2_o21ai_1 _1436_ (.B1(net178),
    .Y(_0521_),
    .A1(net132),
    .A2(\state[70] ));
 sg13g2_a21o_1 _1437_ (.A2(_0771_),
    .A1(net132),
    .B1(_0521_),
    .X(_0522_));
 sg13g2_a21oi_1 _1438_ (.A1(net88),
    .A2(\daisychain[69] ),
    .Y(_0523_),
    .B1(net64));
 sg13g2_a22oi_1 _1439_ (.Y(_0198_),
    .B1(_0522_),
    .B2(_0523_),
    .A2(net64),
    .A1(_0771_));
 sg13g2_o21ai_1 _1440_ (.B1(net179),
    .Y(_0524_),
    .A1(net132),
    .A2(\state[71] ));
 sg13g2_a21o_1 _1441_ (.A2(_0772_),
    .A1(net132),
    .B1(_0524_),
    .X(_0525_));
 sg13g2_a21oi_1 _1442_ (.A1(net87),
    .A2(\daisychain[70] ),
    .Y(_0526_),
    .B1(net65));
 sg13g2_a22oi_1 _1443_ (.Y(_0199_),
    .B1(_0525_),
    .B2(_0526_),
    .A2(net65),
    .A1(_0772_));
 sg13g2_o21ai_1 _1444_ (.B1(net179),
    .Y(_0527_),
    .A1(net132),
    .A2(\state[72] ));
 sg13g2_a21o_1 _1445_ (.A2(_0773_),
    .A1(net130),
    .B1(_0527_),
    .X(_0528_));
 sg13g2_a21oi_1 _1446_ (.A1(net86),
    .A2(\daisychain[71] ),
    .Y(_0529_),
    .B1(net63));
 sg13g2_a22oi_1 _1447_ (.Y(_0200_),
    .B1(_0528_),
    .B2(_0529_),
    .A2(net63),
    .A1(_0773_));
 sg13g2_o21ai_1 _1448_ (.B1(net177),
    .Y(_0530_),
    .A1(net130),
    .A2(\state[73] ));
 sg13g2_a21o_1 _1449_ (.A2(_0774_),
    .A1(net130),
    .B1(_0530_),
    .X(_0531_));
 sg13g2_a21oi_1 _1450_ (.A1(net86),
    .A2(\daisychain[72] ),
    .Y(_0532_),
    .B1(net63));
 sg13g2_a22oi_1 _1451_ (.Y(_0201_),
    .B1(_0531_),
    .B2(_0532_),
    .A2(net65),
    .A1(_0774_));
 sg13g2_o21ai_1 _1452_ (.B1(net178),
    .Y(_0533_),
    .A1(net131),
    .A2(\state[74] ));
 sg13g2_a21o_1 _1453_ (.A2(_0775_),
    .A1(net130),
    .B1(_0533_),
    .X(_0534_));
 sg13g2_a21oi_1 _1454_ (.A1(net86),
    .A2(\daisychain[73] ),
    .Y(_0535_),
    .B1(net65));
 sg13g2_a22oi_1 _1455_ (.Y(_0202_),
    .B1(_0534_),
    .B2(_0535_),
    .A2(net63),
    .A1(_0775_));
 sg13g2_o21ai_1 _1456_ (.B1(net178),
    .Y(_0536_),
    .A1(net131),
    .A2(\state[75] ));
 sg13g2_a21o_1 _1457_ (.A2(_0776_),
    .A1(net130),
    .B1(_0536_),
    .X(_0537_));
 sg13g2_a21oi_1 _1458_ (.A1(net86),
    .A2(\daisychain[74] ),
    .Y(_0538_),
    .B1(net63));
 sg13g2_a22oi_1 _1459_ (.Y(_0203_),
    .B1(_0537_),
    .B2(_0538_),
    .A2(net63),
    .A1(_0776_));
 sg13g2_o21ai_1 _1460_ (.B1(net177),
    .Y(_0539_),
    .A1(net130),
    .A2(\state[76] ));
 sg13g2_a21o_1 _1461_ (.A2(_0777_),
    .A1(net130),
    .B1(_0539_),
    .X(_0540_));
 sg13g2_a21oi_1 _1462_ (.A1(net86),
    .A2(\daisychain[75] ),
    .Y(_0541_),
    .B1(net63));
 sg13g2_a22oi_1 _1463_ (.Y(_0204_),
    .B1(_0540_),
    .B2(_0541_),
    .A2(net63),
    .A1(_0777_));
 sg13g2_o21ai_1 _1464_ (.B1(net175),
    .Y(_0542_),
    .A1(net128),
    .A2(\state[77] ));
 sg13g2_a21o_1 _1465_ (.A2(_0778_),
    .A1(net128),
    .B1(_0542_),
    .X(_0543_));
 sg13g2_a21oi_1 _1466_ (.A1(net87),
    .A2(\daisychain[76] ),
    .Y(_0544_),
    .B1(net61));
 sg13g2_a22oi_1 _1467_ (.Y(_0205_),
    .B1(_0543_),
    .B2(_0544_),
    .A2(net61),
    .A1(_0778_));
 sg13g2_o21ai_1 _1468_ (.B1(net175),
    .Y(_0545_),
    .A1(net128),
    .A2(\state[78] ));
 sg13g2_a21o_1 _1469_ (.A2(_0779_),
    .A1(net128),
    .B1(_0545_),
    .X(_0546_));
 sg13g2_a21oi_1 _1470_ (.A1(net87),
    .A2(\daisychain[77] ),
    .Y(_0547_),
    .B1(net61));
 sg13g2_a22oi_1 _1471_ (.Y(_0206_),
    .B1(_0546_),
    .B2(_0547_),
    .A2(net61),
    .A1(_0779_));
 sg13g2_o21ai_1 _1472_ (.B1(net175),
    .Y(_0548_),
    .A1(net128),
    .A2(\state[79] ));
 sg13g2_a21o_1 _1473_ (.A2(_0780_),
    .A1(net128),
    .B1(_0548_),
    .X(_0549_));
 sg13g2_a21oi_1 _1474_ (.A1(net87),
    .A2(\daisychain[78] ),
    .Y(_0550_),
    .B1(net61));
 sg13g2_a22oi_1 _1475_ (.Y(_0207_),
    .B1(_0549_),
    .B2(_0550_),
    .A2(net61),
    .A1(_0780_));
 sg13g2_o21ai_1 _1476_ (.B1(net170),
    .Y(_0551_),
    .A1(net123),
    .A2(\state[80] ));
 sg13g2_a21o_1 _1477_ (.A2(_0781_),
    .A1(net123),
    .B1(_0551_),
    .X(_0552_));
 sg13g2_a21oi_1 _1478_ (.A1(net85),
    .A2(\daisychain[79] ),
    .Y(_0553_),
    .B1(net56));
 sg13g2_a22oi_1 _1479_ (.Y(_0208_),
    .B1(_0552_),
    .B2(_0553_),
    .A2(net56),
    .A1(_0781_));
 sg13g2_o21ai_1 _1480_ (.B1(net170),
    .Y(_0554_),
    .A1(net123),
    .A2(\state[81] ));
 sg13g2_a21o_1 _1481_ (.A2(_0782_),
    .A1(net123),
    .B1(_0554_),
    .X(_0555_));
 sg13g2_a21oi_1 _1482_ (.A1(net85),
    .A2(\daisychain[80] ),
    .Y(_0556_),
    .B1(net56));
 sg13g2_a22oi_1 _1483_ (.Y(_0209_),
    .B1(_0555_),
    .B2(_0556_),
    .A2(net56),
    .A1(_0782_));
 sg13g2_o21ai_1 _1484_ (.B1(net170),
    .Y(_0557_),
    .A1(net127),
    .A2(\state[82] ));
 sg13g2_a21o_1 _1485_ (.A2(_0783_),
    .A1(net127),
    .B1(_0557_),
    .X(_0558_));
 sg13g2_a21oi_1 _1486_ (.A1(net85),
    .A2(\daisychain[81] ),
    .Y(_0559_),
    .B1(net60));
 sg13g2_a22oi_1 _1487_ (.Y(_0210_),
    .B1(_0558_),
    .B2(_0559_),
    .A2(net60),
    .A1(_0783_));
 sg13g2_o21ai_1 _1488_ (.B1(net172),
    .Y(_0560_),
    .A1(net125),
    .A2(\state[83] ));
 sg13g2_a21o_1 _1489_ (.A2(_0784_),
    .A1(net125),
    .B1(_0560_),
    .X(_0561_));
 sg13g2_a21oi_1 _1490_ (.A1(net84),
    .A2(\daisychain[82] ),
    .Y(_0562_),
    .B1(net58));
 sg13g2_a22oi_1 _1491_ (.Y(_0211_),
    .B1(_0561_),
    .B2(_0562_),
    .A2(net58),
    .A1(_0784_));
 sg13g2_o21ai_1 _1492_ (.B1(net177),
    .Y(_0563_),
    .A1(net125),
    .A2(\state[84] ));
 sg13g2_a21o_1 _1493_ (.A2(_0785_),
    .A1(net125),
    .B1(_0563_),
    .X(_0564_));
 sg13g2_a21oi_1 _1494_ (.A1(net84),
    .A2(\daisychain[83] ),
    .Y(_0565_),
    .B1(net58));
 sg13g2_a22oi_1 _1495_ (.Y(_0212_),
    .B1(_0564_),
    .B2(_0565_),
    .A2(net58),
    .A1(_0785_));
 sg13g2_o21ai_1 _1496_ (.B1(net177),
    .Y(_0566_),
    .A1(net130),
    .A2(\state[85] ));
 sg13g2_a21o_1 _1497_ (.A2(_0786_),
    .A1(net125),
    .B1(_0566_),
    .X(_0567_));
 sg13g2_a21oi_1 _1498_ (.A1(net84),
    .A2(\daisychain[84] ),
    .Y(_0568_),
    .B1(net58));
 sg13g2_a22oi_1 _1499_ (.Y(_0213_),
    .B1(_0567_),
    .B2(_0568_),
    .A2(net58),
    .A1(_0786_));
 sg13g2_o21ai_1 _1500_ (.B1(net177),
    .Y(_0569_),
    .A1(net133),
    .A2(\state[86] ));
 sg13g2_a21o_1 _1501_ (.A2(_0787_),
    .A1(net125),
    .B1(_0569_),
    .X(_0570_));
 sg13g2_a21oi_1 _1502_ (.A1(net84),
    .A2(\daisychain[85] ),
    .Y(_0571_),
    .B1(net58));
 sg13g2_a22oi_1 _1503_ (.Y(_0214_),
    .B1(_0570_),
    .B2(_0571_),
    .A2(net58),
    .A1(_0787_));
 sg13g2_o21ai_1 _1504_ (.B1(net172),
    .Y(_0572_),
    .A1(net125),
    .A2(\state[87] ));
 sg13g2_a21o_1 _1505_ (.A2(_0788_),
    .A1(net126),
    .B1(_0572_),
    .X(_0573_));
 sg13g2_a21oi_1 _1506_ (.A1(net85),
    .A2(\daisychain[86] ),
    .Y(_0574_),
    .B1(net59));
 sg13g2_a22oi_1 _1507_ (.Y(_0215_),
    .B1(_0573_),
    .B2(_0574_),
    .A2(net59),
    .A1(_0788_));
 sg13g2_o21ai_1 _1508_ (.B1(net171),
    .Y(_0575_),
    .A1(net124),
    .A2(\state[88] ));
 sg13g2_a21o_1 _1509_ (.A2(_0789_),
    .A1(net124),
    .B1(_0575_),
    .X(_0576_));
 sg13g2_a21oi_1 _1510_ (.A1(net84),
    .A2(\daisychain[87] ),
    .Y(_0577_),
    .B1(net57));
 sg13g2_a22oi_1 _1511_ (.Y(_0216_),
    .B1(_0576_),
    .B2(_0577_),
    .A2(net57),
    .A1(_0789_));
 sg13g2_o21ai_1 _1512_ (.B1(net154),
    .Y(_0578_),
    .A1(net108),
    .A2(\state[89] ));
 sg13g2_a21o_1 _1513_ (.A2(_0790_),
    .A1(net108),
    .B1(_0578_),
    .X(_0579_));
 sg13g2_a21oi_1 _1514_ (.A1(net76),
    .A2(\daisychain[88] ),
    .Y(_0580_),
    .B1(net41));
 sg13g2_a22oi_1 _1515_ (.Y(_0217_),
    .B1(_0579_),
    .B2(_0580_),
    .A2(net41),
    .A1(_0790_));
 sg13g2_o21ai_1 _1516_ (.B1(net171),
    .Y(_0581_),
    .A1(net124),
    .A2(\state[90] ));
 sg13g2_a21o_1 _1517_ (.A2(_0791_),
    .A1(net126),
    .B1(_0581_),
    .X(_0582_));
 sg13g2_a21oi_1 _1518_ (.A1(net76),
    .A2(\daisychain[89] ),
    .Y(_0583_),
    .B1(net41));
 sg13g2_a22oi_1 _1519_ (.Y(_0218_),
    .B1(_0582_),
    .B2(_0583_),
    .A2(net43),
    .A1(_0791_));
 sg13g2_o21ai_1 _1520_ (.B1(net172),
    .Y(_0584_),
    .A1(net126),
    .A2(\state[91] ));
 sg13g2_a21o_1 _1521_ (.A2(_0792_),
    .A1(net126),
    .B1(_0584_),
    .X(_0585_));
 sg13g2_a21oi_1 _1522_ (.A1(net84),
    .A2(\daisychain[90] ),
    .Y(_0586_),
    .B1(net57));
 sg13g2_a22oi_1 _1523_ (.Y(_0219_),
    .B1(_0585_),
    .B2(_0586_),
    .A2(net59),
    .A1(_0792_));
 sg13g2_o21ai_1 _1524_ (.B1(net172),
    .Y(_0587_),
    .A1(net125),
    .A2(\state[92] ));
 sg13g2_a21o_1 _1525_ (.A2(_0793_),
    .A1(net124),
    .B1(_0587_),
    .X(_0588_));
 sg13g2_a21oi_1 _1526_ (.A1(net84),
    .A2(\daisychain[91] ),
    .Y(_0589_),
    .B1(net59));
 sg13g2_a22oi_1 _1527_ (.Y(_0220_),
    .B1(_0588_),
    .B2(_0589_),
    .A2(net57),
    .A1(_0793_));
 sg13g2_o21ai_1 _1528_ (.B1(net171),
    .Y(_0590_),
    .A1(net124),
    .A2(\state[93] ));
 sg13g2_a21o_1 _1529_ (.A2(_0794_),
    .A1(net124),
    .B1(_0590_),
    .X(_0591_));
 sg13g2_a21oi_1 _1530_ (.A1(net84),
    .A2(\daisychain[92] ),
    .Y(_0592_),
    .B1(net57));
 sg13g2_a22oi_1 _1531_ (.Y(_0221_),
    .B1(_0591_),
    .B2(_0592_),
    .A2(net57),
    .A1(_0794_));
 sg13g2_o21ai_1 _1532_ (.B1(net154),
    .Y(_0593_),
    .A1(net108),
    .A2(\state[94] ));
 sg13g2_a21o_1 _1533_ (.A2(_0795_),
    .A1(net108),
    .B1(_0593_),
    .X(_0594_));
 sg13g2_a21oi_1 _1534_ (.A1(net76),
    .A2(\daisychain[93] ),
    .Y(_0595_),
    .B1(net41));
 sg13g2_a22oi_1 _1535_ (.Y(_0222_),
    .B1(_0594_),
    .B2(_0595_),
    .A2(net41),
    .A1(_0795_));
 sg13g2_o21ai_1 _1536_ (.B1(net154),
    .Y(_0596_),
    .A1(net108),
    .A2(\state[95] ));
 sg13g2_a21o_1 _1537_ (.A2(_0796_),
    .A1(net109),
    .B1(_0596_),
    .X(_0597_));
 sg13g2_a21oi_1 _1538_ (.A1(net76),
    .A2(\daisychain[94] ),
    .Y(_0598_),
    .B1(net41));
 sg13g2_a22oi_1 _1539_ (.Y(_0223_),
    .B1(_0597_),
    .B2(_0598_),
    .A2(net43),
    .A1(_0796_));
 sg13g2_o21ai_1 _1540_ (.B1(net154),
    .Y(_0599_),
    .A1(net109),
    .A2(\state[96] ));
 sg13g2_a21o_1 _1541_ (.A2(_0797_),
    .A1(net109),
    .B1(_0599_),
    .X(_0600_));
 sg13g2_a21oi_1 _1542_ (.A1(net76),
    .A2(\daisychain[95] ),
    .Y(_0601_),
    .B1(net42));
 sg13g2_a22oi_1 _1543_ (.Y(_0224_),
    .B1(_0600_),
    .B2(_0601_),
    .A2(net42),
    .A1(_0797_));
 sg13g2_o21ai_1 _1544_ (.B1(net154),
    .Y(_0602_),
    .A1(net109),
    .A2(\state[97] ));
 sg13g2_a21o_1 _1545_ (.A2(_0798_),
    .A1(net109),
    .B1(_0602_),
    .X(_0603_));
 sg13g2_a21oi_1 _1546_ (.A1(net76),
    .A2(\daisychain[96] ),
    .Y(_0604_),
    .B1(net42));
 sg13g2_a22oi_1 _1547_ (.Y(_0225_),
    .B1(_0603_),
    .B2(_0604_),
    .A2(net42),
    .A1(_0798_));
 sg13g2_o21ai_1 _1548_ (.B1(net155),
    .Y(_0605_),
    .A1(net108),
    .A2(\state[98] ));
 sg13g2_a21o_1 _1549_ (.A2(_0799_),
    .A1(net108),
    .B1(_0605_),
    .X(_0606_));
 sg13g2_a21oi_1 _1550_ (.A1(net76),
    .A2(\daisychain[97] ),
    .Y(_0607_),
    .B1(net42));
 sg13g2_a22oi_1 _1551_ (.Y(_0226_),
    .B1(_0606_),
    .B2(_0607_),
    .A2(net42),
    .A1(_0799_));
 sg13g2_o21ai_1 _1552_ (.B1(net155),
    .Y(_0608_),
    .A1(net110),
    .A2(\state[99] ));
 sg13g2_a21o_1 _1553_ (.A2(_0800_),
    .A1(net108),
    .B1(_0608_),
    .X(_0609_));
 sg13g2_a21oi_1 _1554_ (.A1(net77),
    .A2(\daisychain[98] ),
    .Y(_0610_),
    .B1(net41));
 sg13g2_a22oi_1 _1555_ (.Y(_0227_),
    .B1(_0609_),
    .B2(_0610_),
    .A2(net41),
    .A1(_0800_));
 sg13g2_o21ai_1 _1556_ (.B1(net171),
    .Y(_0611_),
    .A1(net124),
    .A2(\state[100] ));
 sg13g2_a21o_1 _1557_ (.A2(_0801_),
    .A1(net124),
    .B1(_0611_),
    .X(_0612_));
 sg13g2_a21oi_1 _1558_ (.A1(net77),
    .A2(\daisychain[99] ),
    .Y(_0613_),
    .B1(net57));
 sg13g2_a22oi_1 _1559_ (.Y(_0228_),
    .B1(_0612_),
    .B2(_0613_),
    .A2(net57),
    .A1(_0801_));
 sg13g2_o21ai_1 _1560_ (.B1(net170),
    .Y(_0614_),
    .A1(net123),
    .A2(\state[101] ));
 sg13g2_a21o_1 _1561_ (.A2(_0802_),
    .A1(net123),
    .B1(_0614_),
    .X(_0615_));
 sg13g2_a21oi_1 _1562_ (.A1(net85),
    .A2(\daisychain[100] ),
    .Y(_0616_),
    .B1(net56));
 sg13g2_a22oi_1 _1563_ (.Y(_0229_),
    .B1(_0615_),
    .B2(_0616_),
    .A2(net56),
    .A1(_0802_));
 sg13g2_o21ai_1 _1564_ (.B1(net170),
    .Y(_0617_),
    .A1(net123),
    .A2(\state[102] ));
 sg13g2_a21o_1 _1565_ (.A2(_0803_),
    .A1(net123),
    .B1(_0617_),
    .X(_0618_));
 sg13g2_a21oi_1 _1566_ (.A1(net85),
    .A2(\daisychain[101] ),
    .Y(_0619_),
    .B1(net56));
 sg13g2_a22oi_1 _1567_ (.Y(_0230_),
    .B1(_0618_),
    .B2(_0619_),
    .A2(net56),
    .A1(_0803_));
 sg13g2_o21ai_1 _1568_ (.B1(net153),
    .Y(_0620_),
    .A1(net110),
    .A2(\state[103] ));
 sg13g2_a21o_1 _1569_ (.A2(_0804_),
    .A1(net110),
    .B1(_0620_),
    .X(_0621_));
 sg13g2_a21oi_1 _1570_ (.A1(net77),
    .A2(\daisychain[102] ),
    .Y(_0622_),
    .B1(net40));
 sg13g2_a22oi_1 _1571_ (.Y(_0231_),
    .B1(_0621_),
    .B2(_0622_),
    .A2(net43),
    .A1(_0804_));
 sg13g2_o21ai_1 _1572_ (.B1(net156),
    .Y(_0623_),
    .A1(net107),
    .A2(\state[104] ));
 sg13g2_a21o_1 _1573_ (.A2(_0805_),
    .A1(net107),
    .B1(_0623_),
    .X(_0624_));
 sg13g2_a21oi_1 _1574_ (.A1(net77),
    .A2(\daisychain[103] ),
    .Y(_0625_),
    .B1(net43));
 sg13g2_a22oi_1 _1575_ (.Y(_0232_),
    .B1(_0624_),
    .B2(_0625_),
    .A2(net40),
    .A1(_0805_));
 sg13g2_o21ai_1 _1576_ (.B1(net153),
    .Y(_0626_),
    .A1(net107),
    .A2(\state[105] ));
 sg13g2_a21o_1 _1577_ (.A2(_0806_),
    .A1(net107),
    .B1(_0626_),
    .X(_0627_));
 sg13g2_a21oi_1 _1578_ (.A1(net77),
    .A2(\daisychain[104] ),
    .Y(_0628_),
    .B1(net40));
 sg13g2_a22oi_1 _1579_ (.Y(_0233_),
    .B1(_0627_),
    .B2(_0628_),
    .A2(net40),
    .A1(_0806_));
 sg13g2_o21ai_1 _1580_ (.B1(net152),
    .Y(_0629_),
    .A1(net106),
    .A2(\state[106] ));
 sg13g2_a21o_1 _1581_ (.A2(_0807_),
    .A1(net106),
    .B1(_0629_),
    .X(_0630_));
 sg13g2_a21oi_1 _1582_ (.A1(net76),
    .A2(\daisychain[105] ),
    .Y(_0631_),
    .B1(net42));
 sg13g2_a22oi_1 _1583_ (.Y(_0234_),
    .B1(_0630_),
    .B2(_0631_),
    .A2(net39),
    .A1(_0807_));
 sg13g2_o21ai_1 _1584_ (.B1(net151),
    .Y(_0632_),
    .A1(net105),
    .A2(\state[107] ));
 sg13g2_a21o_1 _1585_ (.A2(_0808_),
    .A1(net105),
    .B1(_0632_),
    .X(_0633_));
 sg13g2_a21oi_1 _1586_ (.A1(net78),
    .A2(\daisychain[106] ),
    .Y(_0634_),
    .B1(net39));
 sg13g2_a22oi_1 _1587_ (.Y(_0235_),
    .B1(_0633_),
    .B2(_0634_),
    .A2(net38),
    .A1(_0808_));
 sg13g2_o21ai_1 _1588_ (.B1(net151),
    .Y(_0635_),
    .A1(net105),
    .A2(\state[108] ));
 sg13g2_a21o_1 _1589_ (.A2(_0809_),
    .A1(net105),
    .B1(_0635_),
    .X(_0636_));
 sg13g2_a21oi_1 _1590_ (.A1(net75),
    .A2(\daisychain[107] ),
    .Y(_0637_),
    .B1(net38));
 sg13g2_a22oi_1 _1591_ (.Y(_0236_),
    .B1(_0636_),
    .B2(_0637_),
    .A2(net39),
    .A1(_0809_));
 sg13g2_o21ai_1 _1592_ (.B1(net153),
    .Y(_0638_),
    .A1(net107),
    .A2(\state[109] ));
 sg13g2_a21o_1 _1593_ (.A2(_0810_),
    .A1(net107),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_a21oi_1 _1594_ (.A1(net77),
    .A2(\daisychain[108] ),
    .Y(_0640_),
    .B1(net40));
 sg13g2_a22oi_1 _1595_ (.Y(_0237_),
    .B1(_0639_),
    .B2(_0640_),
    .A2(net40),
    .A1(_0810_));
 sg13g2_o21ai_1 _1596_ (.B1(net153),
    .Y(_0641_),
    .A1(net107),
    .A2(\state[110] ));
 sg13g2_a21o_1 _1597_ (.A2(_0811_),
    .A1(net107),
    .B1(_0641_),
    .X(_0642_));
 sg13g2_a21oi_1 _1598_ (.A1(net77),
    .A2(\daisychain[109] ),
    .Y(_0643_),
    .B1(net40));
 sg13g2_a22oi_1 _1599_ (.Y(_0238_),
    .B1(_0642_),
    .B2(_0643_),
    .A2(net40),
    .A1(_0811_));
 sg13g2_o21ai_1 _1600_ (.B1(net151),
    .Y(_0644_),
    .A1(net105),
    .A2(\state[111] ));
 sg13g2_a21o_1 _1601_ (.A2(_0812_),
    .A1(net106),
    .B1(_0644_),
    .X(_0645_));
 sg13g2_a21oi_1 _1602_ (.A1(net75),
    .A2(\daisychain[110] ),
    .Y(_0646_),
    .B1(net39));
 sg13g2_a22oi_1 _1603_ (.Y(_0239_),
    .B1(_0645_),
    .B2(_0646_),
    .A2(net39),
    .A1(_0812_));
 sg13g2_o21ai_1 _1604_ (.B1(net150),
    .Y(_0647_),
    .A1(net104),
    .A2(\state[112] ));
 sg13g2_a21o_1 _1605_ (.A2(_0813_),
    .A1(net104),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_a21oi_1 _1606_ (.A1(net75),
    .A2(\daisychain[111] ),
    .Y(_0649_),
    .B1(net37));
 sg13g2_a22oi_1 _1607_ (.Y(_0240_),
    .B1(_0648_),
    .B2(_0649_),
    .A2(net37),
    .A1(_0813_));
 sg13g2_o21ai_1 _1608_ (.B1(net150),
    .Y(_0650_),
    .A1(net104),
    .A2(\state[113] ));
 sg13g2_a21o_1 _1609_ (.A2(_0814_),
    .A1(net104),
    .B1(_0650_),
    .X(_0651_));
 sg13g2_a21oi_1 _1610_ (.A1(net75),
    .A2(\daisychain[112] ),
    .Y(_0652_),
    .B1(net37));
 sg13g2_a22oi_1 _1611_ (.Y(_0241_),
    .B1(_0651_),
    .B2(_0652_),
    .A2(net37),
    .A1(_0814_));
 sg13g2_o21ai_1 _1612_ (.B1(net151),
    .Y(_0653_),
    .A1(net104),
    .A2(\state[114] ));
 sg13g2_a21o_1 _1613_ (.A2(_0815_),
    .A1(net104),
    .B1(_0653_),
    .X(_0654_));
 sg13g2_a21oi_1 _1614_ (.A1(net75),
    .A2(\daisychain[113] ),
    .Y(_0655_),
    .B1(net37));
 sg13g2_a22oi_1 _1615_ (.Y(_0242_),
    .B1(_0654_),
    .B2(_0655_),
    .A2(net37),
    .A1(_0815_));
 sg13g2_o21ai_1 _1616_ (.B1(net152),
    .Y(_0656_),
    .A1(net105),
    .A2(\state[115] ));
 sg13g2_a21o_1 _1617_ (.A2(_0816_),
    .A1(net105),
    .B1(_0656_),
    .X(_0657_));
 sg13g2_a21oi_1 _1618_ (.A1(net75),
    .A2(\daisychain[114] ),
    .Y(_0658_),
    .B1(net38));
 sg13g2_a22oi_1 _1619_ (.Y(_0243_),
    .B1(_0657_),
    .B2(_0658_),
    .A2(net38),
    .A1(_0816_));
 sg13g2_o21ai_1 _1620_ (.B1(net150),
    .Y(_0659_),
    .A1(net94),
    .A2(\state[116] ));
 sg13g2_a21o_1 _1621_ (.A2(_0817_),
    .A1(net94),
    .B1(_0659_),
    .X(_0660_));
 sg13g2_a21oi_1 _1622_ (.A1(net68),
    .A2(\daisychain[115] ),
    .Y(_0661_),
    .B1(net27));
 sg13g2_a22oi_1 _1623_ (.Y(_0244_),
    .B1(_0660_),
    .B2(_0661_),
    .A2(net27),
    .A1(_0817_));
 sg13g2_o21ai_1 _1624_ (.B1(net140),
    .Y(_0662_),
    .A1(net94),
    .A2(\state[117] ));
 sg13g2_a21o_1 _1625_ (.A2(_0818_),
    .A1(net94),
    .B1(_0662_),
    .X(_0663_));
 sg13g2_a21oi_1 _1626_ (.A1(net69),
    .A2(\daisychain[116] ),
    .Y(_0664_),
    .B1(net27));
 sg13g2_a22oi_1 _1627_ (.Y(_0245_),
    .B1(_0663_),
    .B2(_0664_),
    .A2(net28),
    .A1(_0818_));
 sg13g2_o21ai_1 _1628_ (.B1(net140),
    .Y(_0665_),
    .A1(net94),
    .A2(\state[118] ));
 sg13g2_a21o_1 _1629_ (.A2(_0819_),
    .A1(net94),
    .B1(_0665_),
    .X(_0666_));
 sg13g2_a21oi_1 _1630_ (.A1(net69),
    .A2(\daisychain[117] ),
    .Y(_0667_),
    .B1(net28));
 sg13g2_a22oi_1 _1631_ (.Y(_0246_),
    .B1(_0666_),
    .B2(_0667_),
    .A2(net28),
    .A1(_0819_));
 sg13g2_o21ai_1 _1632_ (.B1(net140),
    .Y(_0668_),
    .A1(net95),
    .A2(\state[119] ));
 sg13g2_a21o_1 _1633_ (.A2(_0820_),
    .A1(net95),
    .B1(_0668_),
    .X(_0669_));
 sg13g2_a21oi_1 _1634_ (.A1(net69),
    .A2(\daisychain[118] ),
    .Y(_0670_),
    .B1(net27));
 sg13g2_a22oi_1 _1635_ (.Y(_0247_),
    .B1(_0669_),
    .B2(_0670_),
    .A2(net27),
    .A1(_0820_));
 sg13g2_o21ai_1 _1636_ (.B1(net140),
    .Y(_0671_),
    .A1(net94),
    .A2(\state[120] ));
 sg13g2_a21o_1 _1637_ (.A2(_0821_),
    .A1(net94),
    .B1(_0671_),
    .X(_0672_));
 sg13g2_a21oi_1 _1638_ (.A1(net69),
    .A2(\daisychain[119] ),
    .Y(_0673_),
    .B1(net27));
 sg13g2_a22oi_1 _1639_ (.Y(_0248_),
    .B1(_0672_),
    .B2(_0673_),
    .A2(net27),
    .A1(_0821_));
 sg13g2_o21ai_1 _1640_ (.B1(net138),
    .Y(_0674_),
    .A1(net90),
    .A2(\state[121] ));
 sg13g2_a21o_1 _1641_ (.A2(_0822_),
    .A1(net90),
    .B1(_0674_),
    .X(_0675_));
 sg13g2_a21oi_1 _1642_ (.A1(net70),
    .A2(\daisychain[120] ),
    .Y(_0676_),
    .B1(net23));
 sg13g2_a22oi_1 _1643_ (.Y(_0249_),
    .B1(_0675_),
    .B2(_0676_),
    .A2(net23),
    .A1(_0822_));
 sg13g2_o21ai_1 _1644_ (.B1(net138),
    .Y(_0677_),
    .A1(net90),
    .A2(\state[122] ));
 sg13g2_a21o_1 _1645_ (.A2(_0823_),
    .A1(net90),
    .B1(_0677_),
    .X(_0678_));
 sg13g2_a21oi_1 _1646_ (.A1(net70),
    .A2(\daisychain[121] ),
    .Y(_0679_),
    .B1(net23));
 sg13g2_a22oi_1 _1647_ (.Y(_0250_),
    .B1(_0678_),
    .B2(_0679_),
    .A2(net23),
    .A1(_0823_));
 sg13g2_o21ai_1 _1648_ (.B1(net138),
    .Y(_0680_),
    .A1(net90),
    .A2(\state[123] ));
 sg13g2_a21o_1 _1649_ (.A2(net90),
    .A1(_0695_),
    .B1(_0680_),
    .X(_0681_));
 sg13g2_a21oi_1 _1650_ (.A1(net70),
    .A2(\daisychain[122] ),
    .Y(_0682_),
    .B1(net23));
 sg13g2_a22oi_1 _1651_ (.Y(_0251_),
    .B1(_0681_),
    .B2(_0682_),
    .A2(net23),
    .A1(_0695_));
 sg13g2_o21ai_1 _1652_ (.B1(net138),
    .Y(_0683_),
    .A1(net90),
    .A2(\state[124] ));
 sg13g2_a21o_1 _1653_ (.A2(_0698_),
    .A1(net90),
    .B1(_0683_),
    .X(_0684_));
 sg13g2_a21oi_1 _1654_ (.A1(\daisychain[123] ),
    .A2(net70),
    .Y(_0685_),
    .B1(net23));
 sg13g2_a22oi_1 _1655_ (.Y(_0252_),
    .B1(_0684_),
    .B2(_0685_),
    .A2(net24),
    .A1(_0698_));
 sg13g2_o21ai_1 _1656_ (.B1(net137),
    .Y(_0686_),
    .A1(\state[125] ),
    .A2(net91));
 sg13g2_a21o_1 _1657_ (.A2(net91),
    .A1(_0697_),
    .B1(_0686_),
    .X(_0687_));
 sg13g2_a21oi_1 _1658_ (.A1(net70),
    .A2(\daisychain[124] ),
    .Y(_0688_),
    .B1(net23));
 sg13g2_a22oi_1 _1659_ (.Y(_0253_),
    .B1(_0687_),
    .B2(_0688_),
    .A2(net24),
    .A1(_0697_));
 sg13g2_o21ai_1 _1660_ (.B1(net137),
    .Y(_0689_),
    .A1(net91),
    .A2(\state[126] ));
 sg13g2_a21o_1 _1661_ (.A2(_0699_),
    .A1(net91),
    .B1(_0689_),
    .X(_0690_));
 sg13g2_a21oi_1 _1662_ (.A1(net70),
    .A2(\daisychain[125] ),
    .Y(_0691_),
    .B1(net24));
 sg13g2_a22oi_1 _1663_ (.Y(_0254_),
    .B1(_0690_),
    .B2(_0691_),
    .A2(net24),
    .A1(_0699_));
 sg13g2_o21ai_1 _1664_ (.B1(net137),
    .Y(_0692_),
    .A1(net91),
    .A2(\state[127] ));
 sg13g2_a21o_1 _1665_ (.A2(_0700_),
    .A1(net91),
    .B1(_0692_),
    .X(_0693_));
 sg13g2_a21oi_1 _1666_ (.A1(net70),
    .A2(\daisychain[126] ),
    .Y(_0694_),
    .B1(net24));
 sg13g2_a22oi_1 _1667_ (.Y(_0255_),
    .B1(_0693_),
    .B2(_0694_),
    .A2(net24),
    .A1(_0700_));
 sg13g2_o21ai_1 _1668_ (.B1(_0825_),
    .Y(_0256_),
    .A1(net150),
    .A2(_0000_));
 sg13g2_o21ai_1 _1669_ (.B1(_0829_),
    .Y(_0257_),
    .A1(net143),
    .A2(_0039_));
 sg13g2_o21ai_1 _1670_ (.B1(_0832_),
    .Y(_0258_),
    .A1(net147),
    .A2(_0050_));
 sg13g2_o21ai_1 _1671_ (.B1(_0835_),
    .Y(_0259_),
    .A1(net147),
    .A2(_0061_));
 sg13g2_o21ai_1 _1672_ (.B1(_0838_),
    .Y(_0260_),
    .A1(net144),
    .A2(_0072_));
 sg13g2_o21ai_1 _1673_ (.B1(_0841_),
    .Y(_0261_),
    .A1(net142),
    .A2(_0083_));
 sg13g2_o21ai_1 _1674_ (.B1(_0844_),
    .Y(_0262_),
    .A1(net144),
    .A2(_0094_));
 sg13g2_o21ai_1 _1675_ (.B1(_0847_),
    .Y(_0263_),
    .A1(net139),
    .A2(_0105_));
 sg13g2_o21ai_1 _1676_ (.B1(_0850_),
    .Y(_0264_),
    .A1(net139),
    .A2(_0116_));
 sg13g2_o21ai_1 _1677_ (.B1(_0853_),
    .Y(_0265_),
    .A1(net139),
    .A2(_0127_));
 sg13g2_o21ai_1 _1678_ (.B1(_0856_),
    .Y(_0266_),
    .A1(net140),
    .A2(_0011_));
 sg13g2_o21ai_1 _1679_ (.B1(_0859_),
    .Y(_0267_),
    .A1(net140),
    .A2(_0022_));
 sg13g2_o21ai_1 _1680_ (.B1(_0862_),
    .Y(_0268_),
    .A1(net144),
    .A2(_0031_));
 sg13g2_o21ai_1 _1681_ (.B1(_0865_),
    .Y(_0269_),
    .A1(net142),
    .A2(_0032_));
 sg13g2_o21ai_1 _1682_ (.B1(_0868_),
    .Y(_0270_),
    .A1(net143),
    .A2(_0033_));
 sg13g2_o21ai_1 _1683_ (.B1(_0871_),
    .Y(_0271_),
    .A1(net143),
    .A2(_0034_));
 sg13g2_o21ai_1 _1684_ (.B1(_0874_),
    .Y(_0272_),
    .A1(net142),
    .A2(_0035_));
 sg13g2_o21ai_1 _1685_ (.B1(_0877_),
    .Y(_0273_),
    .A1(net145),
    .A2(_0036_));
 sg13g2_o21ai_1 _1686_ (.B1(_0880_),
    .Y(_0274_),
    .A1(net145),
    .A2(_0037_));
 sg13g2_o21ai_1 _1687_ (.B1(_0883_),
    .Y(_0275_),
    .A1(net146),
    .A2(_0038_));
 sg13g2_o21ai_1 _1688_ (.B1(_0886_),
    .Y(_0276_),
    .A1(net147),
    .A2(_0040_));
 sg13g2_o21ai_1 _1689_ (.B1(_0889_),
    .Y(_0277_),
    .A1(net143),
    .A2(_0041_));
 sg13g2_o21ai_1 _1690_ (.B1(_0892_),
    .Y(_0278_),
    .A1(net148),
    .A2(_0042_));
 sg13g2_o21ai_1 _1691_ (.B1(_0895_),
    .Y(_0279_),
    .A1(net148),
    .A2(_0043_));
 sg13g2_o21ai_1 _1692_ (.B1(_0384_),
    .Y(_0280_),
    .A1(net148),
    .A2(_0044_));
 sg13g2_o21ai_1 _1693_ (.B1(_0387_),
    .Y(_0281_),
    .A1(net148),
    .A2(_0045_));
 sg13g2_o21ai_1 _1694_ (.B1(_0390_),
    .Y(_0282_),
    .A1(net149),
    .A2(_0046_));
 sg13g2_o21ai_1 _1695_ (.B1(_0393_),
    .Y(_0283_),
    .A1(net146),
    .A2(_0047_));
 sg13g2_o21ai_1 _1696_ (.B1(_0396_),
    .Y(_0284_),
    .A1(net149),
    .A2(_0048_));
 sg13g2_o21ai_1 _1697_ (.B1(_0399_),
    .Y(_0285_),
    .A1(net149),
    .A2(_0049_));
 sg13g2_o21ai_1 _1698_ (.B1(_0402_),
    .Y(_0286_),
    .A1(net158),
    .A2(_0051_));
 sg13g2_o21ai_1 _1699_ (.B1(_0405_),
    .Y(_0287_),
    .A1(net158),
    .A2(_0052_));
 sg13g2_o21ai_1 _1700_ (.B1(_0408_),
    .Y(_0288_),
    .A1(net158),
    .A2(_0053_));
 sg13g2_o21ai_1 _1701_ (.B1(_0411_),
    .Y(_0289_),
    .A1(net160),
    .A2(_0054_));
 sg13g2_o21ai_1 _1702_ (.B1(_0414_),
    .Y(_0290_),
    .A1(net161),
    .A2(_0055_));
 sg13g2_o21ai_1 _1703_ (.B1(_0417_),
    .Y(_0291_),
    .A1(net148),
    .A2(_0056_));
 sg13g2_o21ai_1 _1704_ (.B1(_0420_),
    .Y(_0292_),
    .A1(net161),
    .A2(_0057_));
 sg13g2_o21ai_1 _1705_ (.B1(_0423_),
    .Y(_0293_),
    .A1(net161),
    .A2(_0058_));
 sg13g2_o21ai_1 _1706_ (.B1(_0426_),
    .Y(_0294_),
    .A1(net161),
    .A2(_0059_));
 sg13g2_o21ai_1 _1707_ (.B1(_0429_),
    .Y(_0295_),
    .A1(net159),
    .A2(_0060_));
 sg13g2_o21ai_1 _1708_ (.B1(_0432_),
    .Y(_0296_),
    .A1(net159),
    .A2(_0062_));
 sg13g2_o21ai_1 _1709_ (.B1(_0435_),
    .Y(_0297_),
    .A1(net159),
    .A2(_0063_));
 sg13g2_o21ai_1 _1710_ (.B1(_0438_),
    .Y(_0298_),
    .A1(net159),
    .A2(_0064_));
 sg13g2_o21ai_1 _1711_ (.B1(_0441_),
    .Y(_0299_),
    .A1(net163),
    .A2(_0065_));
 sg13g2_o21ai_1 _1712_ (.B1(_0444_),
    .Y(_0300_),
    .A1(net163),
    .A2(_0066_));
 sg13g2_o21ai_1 _1713_ (.B1(_0447_),
    .Y(_0301_),
    .A1(net160),
    .A2(_0067_));
 sg13g2_o21ai_1 _1714_ (.B1(_0450_),
    .Y(_0302_),
    .A1(net162),
    .A2(_0068_));
 sg13g2_o21ai_1 _1715_ (.B1(_0453_),
    .Y(_0303_),
    .A1(net162),
    .A2(_0069_));
 sg13g2_o21ai_1 _1716_ (.B1(_0456_),
    .Y(_0304_),
    .A1(net162),
    .A2(_0070_));
 sg13g2_o21ai_1 _1717_ (.B1(_0459_),
    .Y(_0305_),
    .A1(net167),
    .A2(_0071_));
 sg13g2_o21ai_1 _1718_ (.B1(_0462_),
    .Y(_0306_),
    .A1(net167),
    .A2(_0073_));
 sg13g2_o21ai_1 _1719_ (.B1(_0465_),
    .Y(_0307_),
    .A1(net167),
    .A2(_0074_));
 sg13g2_o21ai_1 _1720_ (.B1(_0468_),
    .Y(_0308_),
    .A1(net163),
    .A2(_0075_));
 sg13g2_o21ai_1 _1721_ (.B1(_0471_),
    .Y(_0309_),
    .A1(net166),
    .A2(_0076_));
 sg13g2_o21ai_1 _1722_ (.B1(_0474_),
    .Y(_0310_),
    .A1(net165),
    .A2(_0077_));
 sg13g2_o21ai_1 _1723_ (.B1(_0477_),
    .Y(_0311_),
    .A1(net163),
    .A2(_0078_));
 sg13g2_o21ai_1 _1724_ (.B1(_0480_),
    .Y(_0312_),
    .A1(net163),
    .A2(_0079_));
 sg13g2_o21ai_1 _1725_ (.B1(_0483_),
    .Y(_0313_),
    .A1(net164),
    .A2(_0080_));
 sg13g2_o21ai_1 _1726_ (.B1(_0486_),
    .Y(_0314_),
    .A1(net164),
    .A2(_0081_));
 sg13g2_o21ai_1 _1727_ (.B1(_0489_),
    .Y(_0315_),
    .A1(net165),
    .A2(_0082_));
 sg13g2_o21ai_1 _1728_ (.B1(_0492_),
    .Y(_0316_),
    .A1(net165),
    .A2(_0084_));
 sg13g2_o21ai_1 _1729_ (.B1(_0495_),
    .Y(_0317_),
    .A1(net168),
    .A2(_0085_));
 sg13g2_o21ai_1 _1730_ (.B1(_0498_),
    .Y(_0318_),
    .A1(net168),
    .A2(_0086_));
 sg13g2_o21ai_1 _1731_ (.B1(_0501_),
    .Y(_0319_),
    .A1(net168),
    .A2(_0087_));
 sg13g2_o21ai_1 _1732_ (.B1(_0504_),
    .Y(_0320_),
    .A1(net176),
    .A2(_0088_));
 sg13g2_o21ai_1 _1733_ (.B1(_0507_),
    .Y(_0321_),
    .A1(net176),
    .A2(_0089_));
 sg13g2_o21ai_1 _1734_ (.B1(_0510_),
    .Y(_0322_),
    .A1(net176),
    .A2(_0090_));
 sg13g2_o21ai_1 _1735_ (.B1(_0513_),
    .Y(_0323_),
    .A1(net178),
    .A2(_0091_));
 sg13g2_o21ai_1 _1736_ (.B1(_0516_),
    .Y(_0324_),
    .A1(net178),
    .A2(_0092_));
 sg13g2_o21ai_1 _1737_ (.B1(_0519_),
    .Y(_0325_),
    .A1(net179),
    .A2(_0093_));
 sg13g2_o21ai_1 _1738_ (.B1(_0522_),
    .Y(_0326_),
    .A1(net179),
    .A2(_0095_));
 sg13g2_o21ai_1 _1739_ (.B1(_0525_),
    .Y(_0327_),
    .A1(net179),
    .A2(_0096_));
 sg13g2_o21ai_1 _1740_ (.B1(_0528_),
    .Y(_0328_),
    .A1(net180),
    .A2(_0097_));
 sg13g2_o21ai_1 _1741_ (.B1(_0531_),
    .Y(_0329_),
    .A1(net180),
    .A2(_0098_));
 sg13g2_o21ai_1 _1742_ (.B1(_0534_),
    .Y(_0330_),
    .A1(net177),
    .A2(_0099_));
 sg13g2_o21ai_1 _1743_ (.B1(_0537_),
    .Y(_0331_),
    .A1(net177),
    .A2(_0100_));
 sg13g2_o21ai_1 _1744_ (.B1(_0540_),
    .Y(_0332_),
    .A1(net177),
    .A2(_0101_));
 sg13g2_o21ai_1 _1745_ (.B1(_0543_),
    .Y(_0333_),
    .A1(net175),
    .A2(_0102_));
 sg13g2_o21ai_1 _1746_ (.B1(_0546_),
    .Y(_0334_),
    .A1(net175),
    .A2(_0103_));
 sg13g2_o21ai_1 _1747_ (.B1(_0549_),
    .Y(_0335_),
    .A1(net175),
    .A2(_0104_));
 sg13g2_o21ai_1 _1748_ (.B1(_0552_),
    .Y(_0336_),
    .A1(net170),
    .A2(_0106_));
 sg13g2_o21ai_1 _1749_ (.B1(_0555_),
    .Y(_0337_),
    .A1(net174),
    .A2(_0107_));
 sg13g2_o21ai_1 _1750_ (.B1(_0558_),
    .Y(_0338_),
    .A1(net174),
    .A2(_0108_));
 sg13g2_o21ai_1 _1751_ (.B1(_0561_),
    .Y(_0339_),
    .A1(net172),
    .A2(_0109_));
 sg13g2_o21ai_1 _1752_ (.B1(_0564_),
    .Y(_0340_),
    .A1(net172),
    .A2(_0110_));
 sg13g2_o21ai_1 _1753_ (.B1(_0567_),
    .Y(_0341_),
    .A1(net172),
    .A2(_0111_));
 sg13g2_o21ai_1 _1754_ (.B1(_0570_),
    .Y(_0342_),
    .A1(net172),
    .A2(_0112_));
 sg13g2_o21ai_1 _1755_ (.B1(_0573_),
    .Y(_0343_),
    .A1(net173),
    .A2(_0113_));
 sg13g2_o21ai_1 _1756_ (.B1(_0576_),
    .Y(_0344_),
    .A1(net171),
    .A2(_0114_));
 sg13g2_o21ai_1 _1757_ (.B1(_0579_),
    .Y(_0345_),
    .A1(net155),
    .A2(_0115_));
 sg13g2_o21ai_1 _1758_ (.B1(_0582_),
    .Y(_0346_),
    .A1(net173),
    .A2(_0117_));
 sg13g2_o21ai_1 _1759_ (.B1(_0585_),
    .Y(_0347_),
    .A1(net173),
    .A2(_0118_));
 sg13g2_o21ai_1 _1760_ (.B1(_0588_),
    .Y(_0348_),
    .A1(net171),
    .A2(_0119_));
 sg13g2_o21ai_1 _1761_ (.B1(_0591_),
    .Y(_0349_),
    .A1(net171),
    .A2(_0120_));
 sg13g2_o21ai_1 _1762_ (.B1(_0594_),
    .Y(_0350_),
    .A1(net155),
    .A2(_0121_));
 sg13g2_o21ai_1 _1763_ (.B1(_0597_),
    .Y(_0351_),
    .A1(net155),
    .A2(_0122_));
 sg13g2_o21ai_1 _1764_ (.B1(_0600_),
    .Y(_0352_),
    .A1(net154),
    .A2(_0123_));
 sg13g2_o21ai_1 _1765_ (.B1(_0603_),
    .Y(_0353_),
    .A1(net154),
    .A2(_0124_));
 sg13g2_o21ai_1 _1766_ (.B1(_0606_),
    .Y(_0354_),
    .A1(net154),
    .A2(_0125_));
 sg13g2_o21ai_1 _1767_ (.B1(_0609_),
    .Y(_0355_),
    .A1(net156),
    .A2(_0126_));
 sg13g2_o21ai_1 _1768_ (.B1(_0612_),
    .Y(_0356_),
    .A1(net171),
    .A2(_0001_));
 sg13g2_o21ai_1 _1769_ (.B1(_0615_),
    .Y(_0357_),
    .A1(net170),
    .A2(_0002_));
 sg13g2_o21ai_1 _1770_ (.B1(_0618_),
    .Y(_0358_),
    .A1(net170),
    .A2(_0003_));
 sg13g2_o21ai_1 _1771_ (.B1(_0621_),
    .Y(_0359_),
    .A1(net156),
    .A2(_0004_));
 sg13g2_o21ai_1 _1772_ (.B1(_0624_),
    .Y(_0360_),
    .A1(net153),
    .A2(_0005_));
 sg13g2_o21ai_1 _1773_ (.B1(_0627_),
    .Y(_0361_),
    .A1(net153),
    .A2(_0006_));
 sg13g2_o21ai_1 _1774_ (.B1(_0630_),
    .Y(_0362_),
    .A1(net152),
    .A2(_0007_));
 sg13g2_o21ai_1 _1775_ (.B1(_0633_),
    .Y(_0363_),
    .A1(net151),
    .A2(_0008_));
 sg13g2_o21ai_1 _1776_ (.B1(_0636_),
    .Y(_0364_),
    .A1(net151),
    .A2(_0009_));
 sg13g2_o21ai_1 _1777_ (.B1(_0639_),
    .Y(_0365_),
    .A1(net153),
    .A2(_0010_));
 sg13g2_o21ai_1 _1778_ (.B1(_0642_),
    .Y(_0366_),
    .A1(net153),
    .A2(_0012_));
 sg13g2_o21ai_1 _1779_ (.B1(_0645_),
    .Y(_0367_),
    .A1(net152),
    .A2(_0013_));
 sg13g2_o21ai_1 _1780_ (.B1(_0648_),
    .Y(_0368_),
    .A1(net150),
    .A2(_0014_));
 sg13g2_o21ai_1 _1781_ (.B1(_0651_),
    .Y(_0369_),
    .A1(net150),
    .A2(_0015_));
 sg13g2_o21ai_1 _1782_ (.B1(_0654_),
    .Y(_0370_),
    .A1(net152),
    .A2(_0016_));
 sg13g2_o21ai_1 _1783_ (.B1(_0657_),
    .Y(_0371_),
    .A1(net150),
    .A2(_0017_));
 sg13g2_o21ai_1 _1784_ (.B1(_0660_),
    .Y(_0372_),
    .A1(net151),
    .A2(_0018_));
 sg13g2_o21ai_1 _1785_ (.B1(_0663_),
    .Y(_0373_),
    .A1(net140),
    .A2(_0019_));
 sg13g2_o21ai_1 _1786_ (.B1(_0666_),
    .Y(_0374_),
    .A1(net141),
    .A2(_0020_));
 sg13g2_o21ai_1 _1787_ (.B1(_0669_),
    .Y(_0375_),
    .A1(net141),
    .A2(_0021_));
 sg13g2_o21ai_1 _1788_ (.B1(_0672_),
    .Y(_0376_),
    .A1(net141),
    .A2(_0023_));
 sg13g2_o21ai_1 _1789_ (.B1(_0675_),
    .Y(_0377_),
    .A1(net137),
    .A2(_0024_));
 sg13g2_o21ai_1 _1790_ (.B1(_0678_),
    .Y(_0378_),
    .A1(net138),
    .A2(_0025_));
 sg13g2_o21ai_1 _1791_ (.B1(_0681_),
    .Y(_0379_),
    .A1(net138),
    .A2(_0026_));
 sg13g2_o21ai_1 _1792_ (.B1(_0684_),
    .Y(_0380_),
    .A1(net141),
    .A2(_0027_));
 sg13g2_o21ai_1 _1793_ (.B1(_0687_),
    .Y(_0381_),
    .A1(net137),
    .A2(_0028_));
 sg13g2_o21ai_1 _1794_ (.B1(_0690_),
    .Y(_0382_),
    .A1(net137),
    .A2(_0029_));
 sg13g2_o21ai_1 _1795_ (.B1(_0693_),
    .Y(_0383_),
    .A1(net137),
    .A2(_0030_));
 sg13g2_dfrbpq_1 _1796_ (.RESET_B(net196),
    .D(_0128_),
    .Q(\daisychain[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1797_ (.RESET_B(net197),
    .D(_0129_),
    .Q(\daisychain[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1798_ (.RESET_B(net197),
    .D(_0130_),
    .Q(\daisychain[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1799_ (.RESET_B(net188),
    .D(_0131_),
    .Q(\daisychain[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1800_ (.RESET_B(net189),
    .D(_0132_),
    .Q(\daisychain[4] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1801_ (.RESET_B(net189),
    .D(_0133_),
    .Q(\daisychain[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1802_ (.RESET_B(net186),
    .D(_0134_),
    .Q(\daisychain[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1803_ (.RESET_B(net185),
    .D(_0135_),
    .Q(\daisychain[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1804_ (.RESET_B(net185),
    .D(_0136_),
    .Q(\daisychain[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1805_ (.RESET_B(net185),
    .D(_0137_),
    .Q(\daisychain[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1806_ (.RESET_B(net185),
    .D(_0138_),
    .Q(\daisychain[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1807_ (.RESET_B(net185),
    .D(_0139_),
    .Q(\daisychain[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1808_ (.RESET_B(net189),
    .D(_0140_),
    .Q(\daisychain[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1809_ (.RESET_B(net189),
    .D(_0141_),
    .Q(\daisychain[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1810_ (.RESET_B(net188),
    .D(_0142_),
    .Q(\daisychain[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1811_ (.RESET_B(net188),
    .D(_0143_),
    .Q(\daisychain[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1812_ (.RESET_B(net190),
    .D(_0144_),
    .Q(\daisychain[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1813_ (.RESET_B(net190),
    .D(_0145_),
    .Q(\daisychain[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1814_ (.RESET_B(net190),
    .D(_0146_),
    .Q(\daisychain[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1815_ (.RESET_B(net191),
    .D(_0147_),
    .Q(\daisychain[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1816_ (.RESET_B(net188),
    .D(_0148_),
    .Q(\daisychain[20] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1817_ (.RESET_B(net193),
    .D(_0149_),
    .Q(\daisychain[21] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1818_ (.RESET_B(net193),
    .D(_0150_),
    .Q(\daisychain[22] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1819_ (.RESET_B(net193),
    .D(_0151_),
    .Q(\daisychain[23] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1820_ (.RESET_B(net194),
    .D(_0152_),
    .Q(\daisychain[24] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1821_ (.RESET_B(net191),
    .D(_0153_),
    .Q(\daisychain[25] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1822_ (.RESET_B(net191),
    .D(_0154_),
    .Q(\daisychain[26] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1823_ (.RESET_B(net191),
    .D(_0155_),
    .Q(\daisychain[27] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1824_ (.RESET_B(net191),
    .D(_0156_),
    .Q(\daisychain[28] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1825_ (.RESET_B(net191),
    .D(_0157_),
    .Q(\daisychain[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1826_ (.RESET_B(net204),
    .D(_0158_),
    .Q(\daisychain[30] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1827_ (.RESET_B(net204),
    .D(_0159_),
    .Q(\daisychain[31] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1828_ (.RESET_B(net204),
    .D(_0160_),
    .Q(\daisychain[32] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1829_ (.RESET_B(net192),
    .D(_0161_),
    .Q(\daisychain[33] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1830_ (.RESET_B(net192),
    .D(_0162_),
    .Q(\daisychain[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1831_ (.RESET_B(net194),
    .D(_0163_),
    .Q(\daisychain[35] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1832_ (.RESET_B(net207),
    .D(_0164_),
    .Q(\daisychain[36] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1833_ (.RESET_B(net207),
    .D(_0165_),
    .Q(\daisychain[37] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1834_ (.RESET_B(net204),
    .D(_0166_),
    .Q(\daisychain[38] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1835_ (.RESET_B(net204),
    .D(_0167_),
    .Q(\daisychain[39] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1836_ (.RESET_B(net205),
    .D(_0168_),
    .Q(\daisychain[40] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1837_ (.RESET_B(net204),
    .D(_0169_),
    .Q(\daisychain[41] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1838_ (.RESET_B(net205),
    .D(_0170_),
    .Q(\daisychain[42] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1839_ (.RESET_B(net205),
    .D(_0171_),
    .Q(\daisychain[43] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1840_ (.RESET_B(net205),
    .D(_0172_),
    .Q(\daisychain[44] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1841_ (.RESET_B(net205),
    .D(_0173_),
    .Q(\daisychain[45] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1842_ (.RESET_B(net207),
    .D(_0174_),
    .Q(\daisychain[46] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1843_ (.RESET_B(net207),
    .D(_0175_),
    .Q(\daisychain[47] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1844_ (.RESET_B(net207),
    .D(_0176_),
    .Q(\daisychain[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1845_ (.RESET_B(net212),
    .D(_0177_),
    .Q(\daisychain[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1846_ (.RESET_B(net212),
    .D(_0178_),
    .Q(\daisychain[50] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1847_ (.RESET_B(net212),
    .D(_0179_),
    .Q(\daisychain[51] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1848_ (.RESET_B(net211),
    .D(_0180_),
    .Q(\daisychain[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1849_ (.RESET_B(net211),
    .D(_0181_),
    .Q(\daisychain[53] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1850_ (.RESET_B(net211),
    .D(_0182_),
    .Q(\daisychain[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1851_ (.RESET_B(net211),
    .D(_0183_),
    .Q(\daisychain[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1852_ (.RESET_B(net211),
    .D(_0184_),
    .Q(\daisychain[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1853_ (.RESET_B(net209),
    .D(_0185_),
    .Q(\daisychain[57] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1854_ (.RESET_B(net209),
    .D(_0186_),
    .Q(\daisychain[58] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1855_ (.RESET_B(net209),
    .D(_0187_),
    .Q(\daisychain[59] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1856_ (.RESET_B(net209),
    .D(_0188_),
    .Q(\daisychain[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1857_ (.RESET_B(net212),
    .D(_0189_),
    .Q(\daisychain[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1858_ (.RESET_B(net212),
    .D(_0190_),
    .Q(\daisychain[62] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1859_ (.RESET_B(net213),
    .D(_0191_),
    .Q(\daisychain[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1860_ (.RESET_B(net219),
    .D(_0192_),
    .Q(\daisychain[64] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1861_ (.RESET_B(net219),
    .D(_0193_),
    .Q(\daisychain[65] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1862_ (.RESET_B(net219),
    .D(_0194_),
    .Q(\daisychain[66] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1863_ (.RESET_B(net221),
    .D(_0195_),
    .Q(\daisychain[67] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1864_ (.RESET_B(net221),
    .D(_0196_),
    .Q(\daisychain[68] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1865_ (.RESET_B(net221),
    .D(_0197_),
    .Q(\daisychain[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1866_ (.RESET_B(net221),
    .D(_0198_),
    .Q(\daisychain[70] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1867_ (.RESET_B(net220),
    .D(_0199_),
    .Q(\daisychain[71] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1868_ (.RESET_B(net220),
    .D(_0200_),
    .Q(\daisychain[72] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1869_ (.RESET_B(net220),
    .D(_0201_),
    .Q(\daisychain[73] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1870_ (.RESET_B(net220),
    .D(_0202_),
    .Q(\daisychain[74] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1871_ (.RESET_B(net220),
    .D(_0203_),
    .Q(\daisychain[75] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1872_ (.RESET_B(net220),
    .D(_0204_),
    .Q(\daisychain[76] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1873_ (.RESET_B(net219),
    .D(_0205_),
    .Q(\daisychain[77] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1874_ (.RESET_B(net219),
    .D(_0206_),
    .Q(\daisychain[78] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1875_ (.RESET_B(net215),
    .D(_0207_),
    .Q(\daisychain[79] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1876_ (.RESET_B(net215),
    .D(_0208_),
    .Q(\daisychain[80] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1877_ (.RESET_B(net215),
    .D(_0209_),
    .Q(\daisychain[81] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1878_ (.RESET_B(net217),
    .D(_0210_),
    .Q(\daisychain[82] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1879_ (.RESET_B(net217),
    .D(_0211_),
    .Q(\daisychain[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1880_ (.RESET_B(net217),
    .D(_0212_),
    .Q(\daisychain[84] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1881_ (.RESET_B(net217),
    .D(_0213_),
    .Q(\daisychain[85] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1882_ (.RESET_B(net217),
    .D(_0214_),
    .Q(\daisychain[86] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1883_ (.RESET_B(net216),
    .D(_0215_),
    .Q(\daisychain[87] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1884_ (.RESET_B(net201),
    .D(_0216_),
    .Q(\daisychain[88] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1885_ (.RESET_B(net201),
    .D(_0217_),
    .Q(\daisychain[89] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1886_ (.RESET_B(net216),
    .D(_0218_),
    .Q(\daisychain[90] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1887_ (.RESET_B(net216),
    .D(_0219_),
    .Q(\daisychain[91] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1888_ (.RESET_B(net216),
    .D(_0220_),
    .Q(\daisychain[92] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1889_ (.RESET_B(net201),
    .D(_0221_),
    .Q(\daisychain[93] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1890_ (.RESET_B(net201),
    .D(_0222_),
    .Q(\daisychain[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1891_ (.RESET_B(net202),
    .D(_0223_),
    .Q(\daisychain[95] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1892_ (.RESET_B(net202),
    .D(_0224_),
    .Q(\daisychain[96] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1893_ (.RESET_B(net202),
    .D(_0225_),
    .Q(\daisychain[97] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1894_ (.RESET_B(net201),
    .D(_0226_),
    .Q(\daisychain[98] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1895_ (.RESET_B(net201),
    .D(_0227_),
    .Q(\daisychain[99] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1896_ (.RESET_B(net216),
    .D(_0228_),
    .Q(\daisychain[100] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1897_ (.RESET_B(net215),
    .D(_0229_),
    .Q(\daisychain[101] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1898_ (.RESET_B(net199),
    .D(_0230_),
    .Q(\daisychain[102] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1899_ (.RESET_B(net200),
    .D(_0231_),
    .Q(\daisychain[103] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1900_ (.RESET_B(net199),
    .D(_0232_),
    .Q(\daisychain[104] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1901_ (.RESET_B(net199),
    .D(_0233_),
    .Q(\daisychain[105] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1902_ (.RESET_B(net203),
    .D(_0234_),
    .Q(\daisychain[106] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1903_ (.RESET_B(net197),
    .D(_0235_),
    .Q(\daisychain[107] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1904_ (.RESET_B(net197),
    .D(_0236_),
    .Q(\daisychain[108] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1905_ (.RESET_B(net199),
    .D(_0237_),
    .Q(\daisychain[109] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1906_ (.RESET_B(net197),
    .D(_0238_),
    .Q(\daisychain[110] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1907_ (.RESET_B(net197),
    .D(_0239_),
    .Q(\daisychain[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1908_ (.RESET_B(net196),
    .D(_0240_),
    .Q(\daisychain[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1909_ (.RESET_B(net196),
    .D(_0241_),
    .Q(\daisychain[113] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1910_ (.RESET_B(net196),
    .D(_0242_),
    .Q(\daisychain[114] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1911_ (.RESET_B(net196),
    .D(_0243_),
    .Q(\daisychain[115] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1912_ (.RESET_B(net186),
    .D(_0244_),
    .Q(\daisychain[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1913_ (.RESET_B(net186),
    .D(_0245_),
    .Q(\daisychain[117] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1914_ (.RESET_B(net186),
    .D(_0246_),
    .Q(\daisychain[118] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1915_ (.RESET_B(net186),
    .D(_0247_),
    .Q(\daisychain[119] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1916_ (.RESET_B(net186),
    .D(_0248_),
    .Q(\daisychain[120] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1917_ (.RESET_B(net183),
    .D(_0249_),
    .Q(\daisychain[121] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1918_ (.RESET_B(net183),
    .D(_0250_),
    .Q(\daisychain[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1919_ (.RESET_B(net183),
    .D(_0251_),
    .Q(\daisychain[123] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1920_ (.RESET_B(net183),
    .D(_0252_),
    .Q(\daisychain[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1921_ (.RESET_B(net183),
    .D(_0253_),
    .Q(\daisychain[125] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1922_ (.RESET_B(net183),
    .D(_0254_),
    .Q(\daisychain[126] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1923_ (.RESET_B(net184),
    .D(_0255_),
    .Q(\daisychain[127] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1924_ (.RESET_B(net196),
    .D(_0256_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1925_ (.RESET_B(net188),
    .D(_0257_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1926_ (.RESET_B(net193),
    .D(_0258_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1927_ (.RESET_B(net193),
    .D(_0259_),
    .Q(\state[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1928_ (.RESET_B(net188),
    .D(_0260_),
    .Q(\state[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1929_ (.RESET_B(net190),
    .D(_0261_),
    .Q(\state[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1930_ (.RESET_B(net189),
    .D(_0262_),
    .Q(\state[6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1931_ (.RESET_B(net185),
    .D(_0263_),
    .Q(\state[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1932_ (.RESET_B(net185),
    .D(_0264_),
    .Q(\state[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1933_ (.RESET_B(net185),
    .D(_0265_),
    .Q(\state[9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1934_ (.RESET_B(net187),
    .D(_0266_),
    .Q(\state[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1935_ (.RESET_B(net187),
    .D(_0267_),
    .Q(\state[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1936_ (.RESET_B(net189),
    .D(_0268_),
    .Q(\state[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1937_ (.RESET_B(net189),
    .D(_0269_),
    .Q(\state[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1938_ (.RESET_B(net188),
    .D(_0270_),
    .Q(\state[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1939_ (.RESET_B(net188),
    .D(_0271_),
    .Q(\state[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1940_ (.RESET_B(net189),
    .D(_0272_),
    .Q(\state[16] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1941_ (.RESET_B(net190),
    .D(_0273_),
    .Q(\state[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1942_ (.RESET_B(net190),
    .D(_0274_),
    .Q(\state[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1943_ (.RESET_B(net191),
    .D(_0275_),
    .Q(\state[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1944_ (.RESET_B(net193),
    .D(_0276_),
    .Q(\state[20] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1945_ (.RESET_B(net193),
    .D(_0277_),
    .Q(\state[21] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1946_ (.RESET_B(net193),
    .D(_0278_),
    .Q(\state[22] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1947_ (.RESET_B(net194),
    .D(_0279_),
    .Q(\state[23] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1948_ (.RESET_B(net194),
    .D(_0280_),
    .Q(\state[24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1949_ (.RESET_B(net194),
    .D(_0281_),
    .Q(\state[25] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1950_ (.RESET_B(net192),
    .D(_0282_),
    .Q(\state[26] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1951_ (.RESET_B(net191),
    .D(_0283_),
    .Q(\state[27] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1952_ (.RESET_B(net192),
    .D(_0284_),
    .Q(\state[28] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1953_ (.RESET_B(net192),
    .D(_0285_),
    .Q(\state[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1954_ (.RESET_B(net204),
    .D(_0286_),
    .Q(\state[30] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1955_ (.RESET_B(net204),
    .D(_0287_),
    .Q(\state[31] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1956_ (.RESET_B(net206),
    .D(_0288_),
    .Q(\state[32] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1957_ (.RESET_B(net206),
    .D(_0289_),
    .Q(\state[33] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1958_ (.RESET_B(net207),
    .D(_0290_),
    .Q(\state[34] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1959_ (.RESET_B(net194),
    .D(_0291_),
    .Q(\state[35] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1960_ (.RESET_B(net207),
    .D(_0292_),
    .Q(\state[36] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1961_ (.RESET_B(net207),
    .D(_0293_),
    .Q(\state[37] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1962_ (.RESET_B(net208),
    .D(_0294_),
    .Q(\state[38] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1963_ (.RESET_B(net205),
    .D(_0295_),
    .Q(\state[39] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1964_ (.RESET_B(net206),
    .D(_0296_),
    .Q(\state[40] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1965_ (.RESET_B(net205),
    .D(_0297_),
    .Q(\state[41] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1966_ (.RESET_B(net205),
    .D(_0298_),
    .Q(\state[42] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1967_ (.RESET_B(net211),
    .D(_0299_),
    .Q(\state[43] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1968_ (.RESET_B(net211),
    .D(_0300_),
    .Q(\state[44] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1969_ (.RESET_B(net211),
    .D(_0301_),
    .Q(\state[45] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1970_ (.RESET_B(net212),
    .D(_0302_),
    .Q(\state[46] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1971_ (.RESET_B(net208),
    .D(_0303_),
    .Q(\state[47] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1972_ (.RESET_B(net208),
    .D(_0304_),
    .Q(\state[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1973_ (.RESET_B(net212),
    .D(_0305_),
    .Q(\state[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1974_ (.RESET_B(net212),
    .D(_0306_),
    .Q(\state[50] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1975_ (.RESET_B(net213),
    .D(_0307_),
    .Q(\state[51] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1976_ (.RESET_B(net210),
    .D(_0308_),
    .Q(\state[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1977_ (.RESET_B(net210),
    .D(_0309_),
    .Q(\state[53] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1978_ (.RESET_B(net210),
    .D(_0310_),
    .Q(\state[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1979_ (.RESET_B(net209),
    .D(_0311_),
    .Q(\state[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1980_ (.RESET_B(net209),
    .D(_0312_),
    .Q(\state[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1981_ (.RESET_B(net209),
    .D(_0313_),
    .Q(\state[57] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1982_ (.RESET_B(net209),
    .D(_0314_),
    .Q(\state[58] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1983_ (.RESET_B(net210),
    .D(_0315_),
    .Q(\state[59] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1984_ (.RESET_B(net210),
    .D(_0316_),
    .Q(\state[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1985_ (.RESET_B(net213),
    .D(_0317_),
    .Q(\state[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1986_ (.RESET_B(net213),
    .D(_0318_),
    .Q(\state[62] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1987_ (.RESET_B(net213),
    .D(_0319_),
    .Q(\state[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1988_ (.RESET_B(net224),
    .D(_0320_),
    .Q(\state[64] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1989_ (.RESET_B(net224),
    .D(_0321_),
    .Q(\state[65] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1990_ (.RESET_B(net224),
    .D(_0322_),
    .Q(\state[66] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1991_ (.RESET_B(net221),
    .D(_0323_),
    .Q(\state[67] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1992_ (.RESET_B(net221),
    .D(_0324_),
    .Q(\state[68] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1993_ (.RESET_B(net222),
    .D(_0325_),
    .Q(\state[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1994_ (.RESET_B(net222),
    .D(_0326_),
    .Q(\state[70] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1995_ (.RESET_B(net222),
    .D(_0327_),
    .Q(\state[71] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1996_ (.RESET_B(net222),
    .D(_0328_),
    .Q(\state[72] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1997_ (.RESET_B(net222),
    .D(_0329_),
    .Q(\state[73] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1998_ (.RESET_B(net221),
    .D(_0330_),
    .Q(\state[74] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1999_ (.RESET_B(net221),
    .D(_0331_),
    .Q(\state[75] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2000_ (.RESET_B(net220),
    .D(_0332_),
    .Q(\state[76] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2001_ (.RESET_B(net219),
    .D(_0333_),
    .Q(\state[77] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2002_ (.RESET_B(net219),
    .D(_0334_),
    .Q(\state[78] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2003_ (.RESET_B(net219),
    .D(_0335_),
    .Q(\state[79] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2004_ (.RESET_B(net215),
    .D(_0336_),
    .Q(\state[80] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2005_ (.RESET_B(net215),
    .D(_0337_),
    .Q(\state[81] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2006_ (.RESET_B(net225),
    .D(_0338_),
    .Q(\state[82] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2007_ (.RESET_B(net217),
    .D(_0339_),
    .Q(\state[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2008_ (.RESET_B(net220),
    .D(_0340_),
    .Q(\state[84] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2009_ (.RESET_B(net223),
    .D(_0341_),
    .Q(\state[85] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2010_ (.RESET_B(net223),
    .D(_0342_),
    .Q(\state[86] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2011_ (.RESET_B(net217),
    .D(_0343_),
    .Q(\state[87] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2012_ (.RESET_B(net216),
    .D(_0344_),
    .Q(\state[88] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2013_ (.RESET_B(net202),
    .D(_0345_),
    .Q(\state[89] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2014_ (.RESET_B(net218),
    .D(_0346_),
    .Q(\state[90] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2015_ (.RESET_B(net218),
    .D(_0347_),
    .Q(\state[91] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2016_ (.RESET_B(net217),
    .D(_0348_),
    .Q(\state[92] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2017_ (.RESET_B(net216),
    .D(_0349_),
    .Q(\state[93] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2018_ (.RESET_B(net201),
    .D(_0350_),
    .Q(\state[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2019_ (.RESET_B(net202),
    .D(_0351_),
    .Q(\state[95] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2020_ (.RESET_B(net202),
    .D(_0352_),
    .Q(\state[96] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2021_ (.RESET_B(net202),
    .D(_0353_),
    .Q(\state[97] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2022_ (.RESET_B(net201),
    .D(_0354_),
    .Q(\state[98] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2023_ (.RESET_B(net200),
    .D(_0355_),
    .Q(\state[99] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2024_ (.RESET_B(net216),
    .D(_0356_),
    .Q(\state[100] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2025_ (.RESET_B(net215),
    .D(_0357_),
    .Q(\state[101] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2026_ (.RESET_B(net215),
    .D(_0358_),
    .Q(\state[102] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2027_ (.RESET_B(net200),
    .D(_0359_),
    .Q(\state[103] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2028_ (.RESET_B(net200),
    .D(_0360_),
    .Q(\state[104] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2029_ (.RESET_B(net199),
    .D(_0361_),
    .Q(\state[105] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2030_ (.RESET_B(net203),
    .D(_0362_),
    .Q(\state[106] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2031_ (.RESET_B(net199),
    .D(_0363_),
    .Q(\state[107] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2032_ (.RESET_B(net197),
    .D(_0364_),
    .Q(\state[108] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2033_ (.RESET_B(net199),
    .D(_0365_),
    .Q(\state[109] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2034_ (.RESET_B(net199),
    .D(_0366_),
    .Q(\state[110] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2035_ (.RESET_B(net197),
    .D(_0367_),
    .Q(\state[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2036_ (.RESET_B(net196),
    .D(_0368_),
    .Q(\state[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2037_ (.RESET_B(net198),
    .D(_0369_),
    .Q(\state[113] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2038_ (.RESET_B(net198),
    .D(_0370_),
    .Q(\state[114] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2039_ (.RESET_B(net196),
    .D(_0371_),
    .Q(\state[115] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2040_ (.RESET_B(net198),
    .D(_0372_),
    .Q(\state[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2041_ (.RESET_B(net186),
    .D(_0373_),
    .Q(\state[117] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2042_ (.RESET_B(net187),
    .D(_0374_),
    .Q(\state[118] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2043_ (.RESET_B(net187),
    .D(_0375_),
    .Q(\state[119] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2044_ (.RESET_B(net186),
    .D(_0376_),
    .Q(\state[120] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2045_ (.RESET_B(net184),
    .D(_0377_),
    .Q(\state[121] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2046_ (.RESET_B(net183),
    .D(_0378_),
    .Q(\state[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2047_ (.RESET_B(net183),
    .D(_0379_),
    .Q(\state[123] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2048_ (.RESET_B(net184),
    .D(_0380_),
    .Q(\state[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2049_ (.RESET_B(net184),
    .D(_0381_),
    .Q(\state[125] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2050_ (.RESET_B(net184),
    .D(_0382_),
    .Q(\state[126] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2051_ (.RESET_B(net184),
    .D(_0383_),
    .Q(\state[127] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_tiehi heichips25_pudding_228 (.L_HI(net228));
 sg13g2_tiehi heichips25_pudding_229 (.L_HI(net229));
 sg13g2_tiehi heichips25_pudding_230 (.L_HI(net230));
 sg13g2_tiehi heichips25_pudding_231 (.L_HI(net231));
 sg13g2_tiehi heichips25_pudding_232 (.L_HI(net232));
 sg13g2_tiehi heichips25_pudding_233 (.L_HI(net233));
 sg13g2_tiehi heichips25_pudding_234 (.L_HI(net234));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _2060_ (.A(\state[120] ),
    .X(net7));
 sg13g2_buf_1 _2061_ (.A(\state[121] ),
    .X(net8));
 sg13g2_buf_1 _2062_ (.A(\state[122] ),
    .X(net9));
 sg13g2_buf_1 _2063_ (.A(\state[123] ),
    .X(net10));
 sg13g2_buf_1 _2064_ (.A(\state[124] ),
    .X(net11));
 sg13g2_buf_1 _2065_ (.A(\state[125] ),
    .X(net12));
 sg13g2_buf_1 _2066_ (.A(\state[126] ),
    .X(net13));
 sg13g2_buf_1 _2067_ (.A(\state[127] ),
    .X(net14));
 sg13g2_buf_1 _2068_ (.A(\daisychain[120] ),
    .X(net15));
 sg13g2_buf_1 _2069_ (.A(\daisychain[121] ),
    .X(net16));
 sg13g2_buf_1 _2070_ (.A(\daisychain[122] ),
    .X(net17));
 sg13g2_buf_1 _2071_ (.A(\daisychain[123] ),
    .X(net18));
 sg13g2_buf_1 _2072_ (.A(\daisychain[124] ),
    .X(net19));
 sg13g2_buf_1 _2073_ (.A(\daisychain[125] ),
    .X(net20));
 sg13g2_buf_1 _2074_ (.A(\daisychain[126] ),
    .X(net21));
 sg13g2_buf_1 _2075_ (.A(\daisychain[127] ),
    .X(net22));
 dac128module dac (.Iout(dacout),
    .EN({\digitalen.g[3].u.OUTP ,
    \digitalen.g[2].u.OUTP ,
    \digitalen.g[1].u.OUTP ,
    \digitalen.g[0].u.OUTP }),
    .ENB({\digitalen.g[3].u.OUTN ,
    \digitalen.g[2].u.OUTN ,
    \digitalen.g[1].u.OUTN ,
    \digitalen.g[0].u.OUTN }),
    .ON({\state[127] ,
    \state[126] ,
    \state[125] ,
    \state[124] ,
    \state[123] ,
    \state[122] ,
    \state[121] ,
    \state[120] ,
    \state[119] ,
    \state[118] ,
    \state[117] ,
    \state[116] ,
    \state[115] ,
    \state[114] ,
    \state[113] ,
    \state[112] ,
    \state[111] ,
    \state[110] ,
    \state[109] ,
    \state[108] ,
    \state[107] ,
    \state[106] ,
    \state[105] ,
    \state[104] ,
    \state[103] ,
    \state[102] ,
    \state[101] ,
    \state[100] ,
    \state[99] ,
    \state[98] ,
    \state[97] ,
    \state[96] ,
    \state[95] ,
    \state[94] ,
    \state[93] ,
    \state[92] ,
    \state[91] ,
    \state[90] ,
    \state[89] ,
    \state[88] ,
    \state[87] ,
    \state[86] ,
    \state[85] ,
    \state[84] ,
    \state[83] ,
    \state[82] ,
    \state[81] ,
    \state[80] ,
    \state[79] ,
    \state[78] ,
    \state[77] ,
    \state[76] ,
    \state[75] ,
    \state[74] ,
    \state[73] ,
    \state[72] ,
    \state[71] ,
    \state[70] ,
    \state[69] ,
    \state[68] ,
    \state[67] ,
    \state[66] ,
    \state[65] ,
    \state[64] ,
    \state[63] ,
    \state[62] ,
    \state[61] ,
    \state[60] ,
    \state[59] ,
    \state[58] ,
    \state[57] ,
    \state[56] ,
    \state[55] ,
    \state[54] ,
    \state[53] ,
    \state[52] ,
    \state[51] ,
    \state[50] ,
    \state[49] ,
    \state[48] ,
    \state[47] ,
    \state[46] ,
    \state[45] ,
    \state[44] ,
    \state[43] ,
    \state[42] ,
    \state[41] ,
    \state[40] ,
    \state[39] ,
    \state[38] ,
    \state[37] ,
    \state[36] ,
    \state[35] ,
    \state[34] ,
    \state[33] ,
    \state[32] ,
    \state[31] ,
    \state[30] ,
    \state[29] ,
    \state[28] ,
    \state[27] ,
    \state[26] ,
    \state[25] ,
    \state[24] ,
    \state[23] ,
    \state[22] ,
    \state[21] ,
    \state[20] ,
    \state[19] ,
    \state[18] ,
    \state[17] ,
    \state[16] ,
    \state[15] ,
    \state[14] ,
    \state[13] ,
    \state[12] ,
    \state[11] ,
    \state[10] ,
    \state[9] ,
    \state[8] ,
    \state[7] ,
    \state[6] ,
    \state[5] ,
    \state[4] ,
    \state[3] ,
    \state[2] ,
    \state[1] ,
    \state[0] }),
    .ONB({_0030_,
    _0029_,
    _0028_,
    _0027_,
    _0026_,
    _0025_,
    _0024_,
    _0023_,
    _0021_,
    _0020_,
    _0019_,
    _0018_,
    _0017_,
    _0016_,
    _0015_,
    _0014_,
    _0013_,
    _0012_,
    _0010_,
    _0009_,
    _0008_,
    _0007_,
    _0006_,
    _0005_,
    _0004_,
    _0003_,
    _0002_,
    _0001_,
    _0126_,
    _0125_,
    _0124_,
    _0123_,
    _0122_,
    _0121_,
    _0120_,
    _0119_,
    _0118_,
    _0117_,
    _0115_,
    _0114_,
    _0113_,
    _0112_,
    _0111_,
    _0110_,
    _0109_,
    _0108_,
    _0107_,
    _0106_,
    _0104_,
    _0103_,
    _0102_,
    _0101_,
    _0100_,
    _0099_,
    _0098_,
    _0097_,
    _0096_,
    _0095_,
    _0093_,
    _0092_,
    _0091_,
    _0090_,
    _0089_,
    _0088_,
    _0087_,
    _0086_,
    _0085_,
    _0084_,
    _0082_,
    _0081_,
    _0080_,
    _0079_,
    _0078_,
    _0077_,
    _0076_,
    _0075_,
    _0074_,
    _0073_,
    _0071_,
    _0070_,
    _0069_,
    _0068_,
    _0067_,
    _0066_,
    _0065_,
    _0064_,
    _0063_,
    _0062_,
    _0060_,
    _0059_,
    _0058_,
    _0057_,
    _0056_,
    _0055_,
    _0054_,
    _0053_,
    _0052_,
    _0051_,
    _0049_,
    _0048_,
    _0047_,
    _0046_,
    _0045_,
    _0044_,
    _0043_,
    _0042_,
    _0041_,
    _0040_,
    _0038_,
    _0037_,
    _0036_,
    _0035_,
    _0034_,
    _0033_,
    _0032_,
    _0031_,
    _0022_,
    _0011_,
    _0127_,
    _0116_,
    _0105_,
    _0094_,
    _0083_,
    _0072_,
    _0061_,
    _0050_,
    _0039_,
    _0000_}),
    .VbiasP({\bias[1] ,
    \bias[0] }),
    .VcascP({\iref[1] ,
    \iref[0] }));
 sg13g2_inv_1 \digitalen.g[0].u.inv1  (.Y(\digitalen.g[0].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[0].u.inv2  (.Y(\digitalen.g[0].u.OUTP ),
    .A(\digitalen.g[0].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[1].u.inv1  (.Y(\digitalen.g[1].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[1].u.inv2  (.Y(\digitalen.g[1].u.OUTP ),
    .A(\digitalen.g[1].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[2].u.inv1  (.Y(\digitalen.g[2].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[2].u.inv2  (.Y(\digitalen.g[2].u.OUTP ),
    .A(\digitalen.g[2].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[3].u.inv1  (.Y(\digitalen.g[3].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[3].u.inv2  (.Y(\digitalen.g[3].u.OUTP ),
    .A(\digitalen.g[3].u.OUTN ));
 analog_wires wires (.Iout(dacout),
    .i_in(i_in),
    .i_out(i_out),
    .VDDA({\vdda[1] ,
    \vdda[0] }),
    .VbiasP({\bias[1] ,
    \bias[0] }),
    .VcascP({\iref[1] ,
    \iref[0] }));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]));
 sg13g2_buf_1 fanout23 (.A(net24),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net29),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(net29),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net29),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(net29),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(_0826_),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net32),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net44),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net34),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net36),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net36),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net44),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net38),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net44),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net43),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net42),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(net67),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net47),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(net49),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(net49),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net67),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net53),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net53),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(net55),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net67),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(net60),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net59),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(net59),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net66),
    .X(net60));
 sg13g2_buf_1 fanout61 (.A(net66),
    .X(net61));
 sg13g2_buf_1 fanout62 (.A(net66),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(net65),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(net65),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(net67),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(_0826_),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(net89),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net89),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(net74),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(net78),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(net78),
    .X(net75));
 sg13g2_buf_1 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net78),
    .X(net77));
 sg13g2_buf_1 fanout78 (.A(net89),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(net88),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net83),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_1 fanout83 (.A(net88),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(net85),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net88),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(_0696_),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net136),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(net136),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net95),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net136),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net98),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(net111),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net103),
    .X(net99));
 sg13g2_buf_1 fanout100 (.A(net103),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(net111),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_1 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net111),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net110),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_1 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(net135),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net116),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(net116),
    .X(net114));
 sg13g2_buf_1 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net135),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(net122),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net122),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(net122),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(net135),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(net127),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(net126),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net134),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net134),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(net134),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net133),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net133),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net5),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net141),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net182),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(net157),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(net149),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(net157),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net157),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net156),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net156),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(net182),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_1 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(net169),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net169),
    .X(net161));
 sg13g2_buf_1 fanout162 (.A(net169),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net166),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(net166),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(net169),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_1 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net182),
    .X(net169));
 sg13g2_buf_1 fanout170 (.A(net174),
    .X(net170));
 sg13g2_buf_1 fanout171 (.A(net173),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net181),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net181),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net181),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net180),
    .X(net177));
 sg13g2_buf_1 fanout178 (.A(net180),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_1 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net4),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net227),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net227),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net187),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net227),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net190),
    .X(net188));
 sg13g2_buf_1 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net226),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net195),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(net195),
    .X(net192));
 sg13g2_buf_1 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_1 fanout195 (.A(net226),
    .X(net195));
 sg13g2_buf_1 fanout196 (.A(net198),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_1 fanout198 (.A(net203),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net203),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(net203),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_1 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_1 fanout203 (.A(net226),
    .X(net203));
 sg13g2_buf_1 fanout204 (.A(net206),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_1 fanout206 (.A(net208),
    .X(net206));
 sg13g2_buf_1 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_1 fanout208 (.A(net226),
    .X(net208));
 sg13g2_buf_1 fanout209 (.A(net214),
    .X(net209));
 sg13g2_buf_1 fanout210 (.A(net214),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(net214),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net214),
    .X(net212));
 sg13g2_buf_1 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_1 fanout214 (.A(net226),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net225),
    .X(net215));
 sg13g2_buf_1 fanout216 (.A(net218),
    .X(net216));
 sg13g2_buf_1 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_1 fanout218 (.A(net225),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(net224),
    .X(net219));
 sg13g2_buf_1 fanout220 (.A(net223),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(net223),
    .X(net221));
 sg13g2_buf_1 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_1 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_1 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_1 fanout225 (.A(net226),
    .X(net225));
 sg13g2_buf_1 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_1 fanout227 (.A(net1),
    .X(net227));
 sg13g2_tiehi heichips25_pudding (.L_HI(net));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_16 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_0_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_6_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0007_));
 sg13g2_antennanp ANTENNA_2 (.A(_0012_));
 sg13g2_antennanp ANTENNA_3 (.A(_0047_));
 sg13g2_antennanp ANTENNA_4 (.A(_0112_));
 sg13g2_antennanp ANTENNA_5 (.A(\state[56] ));
 sg13g2_antennanp ANTENNA_6 (.A(\state[83] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_4 FILLER_0_609 ();
 sg13g2_fill_1 FILLER_0_613 ();
 sg13g2_fill_1 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_4 FILLER_0_678 ();
 sg13g2_decap_4 FILLER_0_685 ();
 sg13g2_fill_1 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_783 ();
 sg13g2_fill_1 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_4 FILLER_1_595 ();
 sg13g2_fill_2 FILLER_1_599 ();
 sg13g2_fill_2 FILLER_1_628 ();
 sg13g2_decap_4 FILLER_1_774 ();
 sg13g2_fill_1 FILLER_1_778 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_4 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_fill_2 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_586 ();
 sg13g2_fill_2 FILLER_2_593 ();
 sg13g2_fill_1 FILLER_2_595 ();
 sg13g2_fill_2 FILLER_2_599 ();
 sg13g2_fill_1 FILLER_2_601 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_fill_2 FILLER_2_634 ();
 sg13g2_fill_1 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_fill_2 FILLER_2_662 ();
 sg13g2_fill_1 FILLER_2_675 ();
 sg13g2_decap_4 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_692 ();
 sg13g2_decap_4 FILLER_2_699 ();
 sg13g2_decap_8 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_723 ();
 sg13g2_decap_4 FILLER_2_730 ();
 sg13g2_fill_2 FILLER_2_734 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_fill_2 FILLER_2_784 ();
 sg13g2_fill_1 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_807 ();
 sg13g2_decap_8 FILLER_2_814 ();
 sg13g2_fill_2 FILLER_2_821 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_fill_2 FILLER_3_574 ();
 sg13g2_fill_1 FILLER_3_576 ();
 sg13g2_decap_8 FILLER_3_604 ();
 sg13g2_decap_4 FILLER_3_611 ();
 sg13g2_fill_1 FILLER_3_615 ();
 sg13g2_fill_1 FILLER_3_623 ();
 sg13g2_fill_2 FILLER_3_629 ();
 sg13g2_fill_1 FILLER_3_631 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_fill_1 FILLER_3_662 ();
 sg13g2_fill_2 FILLER_3_672 ();
 sg13g2_fill_1 FILLER_3_674 ();
 sg13g2_fill_2 FILLER_3_716 ();
 sg13g2_fill_1 FILLER_3_718 ();
 sg13g2_fill_2 FILLER_3_746 ();
 sg13g2_fill_2 FILLER_3_756 ();
 sg13g2_fill_2 FILLER_3_761 ();
 sg13g2_fill_1 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_769 ();
 sg13g2_decap_8 FILLER_3_776 ();
 sg13g2_decap_8 FILLER_3_783 ();
 sg13g2_fill_2 FILLER_3_790 ();
 sg13g2_fill_1 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_decap_8 FILLER_4_473 ();
 sg13g2_decap_8 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_8 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_501 ();
 sg13g2_decap_8 FILLER_4_508 ();
 sg13g2_decap_8 FILLER_4_515 ();
 sg13g2_decap_8 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_4_529 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_4 FILLER_4_550 ();
 sg13g2_fill_1 FILLER_4_586 ();
 sg13g2_decap_8 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_fill_1 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_fill_1 FILLER_4_732 ();
 sg13g2_decap_4 FILLER_4_778 ();
 sg13g2_fill_1 FILLER_4_782 ();
 sg13g2_fill_1 FILLER_4_822 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_fill_1 FILLER_5_536 ();
 sg13g2_decap_4 FILLER_5_543 ();
 sg13g2_fill_2 FILLER_5_547 ();
 sg13g2_fill_2 FILLER_5_552 ();
 sg13g2_fill_1 FILLER_5_554 ();
 sg13g2_decap_8 FILLER_5_566 ();
 sg13g2_fill_1 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_577 ();
 sg13g2_fill_2 FILLER_5_584 ();
 sg13g2_decap_4 FILLER_5_618 ();
 sg13g2_fill_1 FILLER_5_622 ();
 sg13g2_fill_1 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_fill_2 FILLER_5_658 ();
 sg13g2_fill_1 FILLER_5_660 ();
 sg13g2_fill_1 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_fill_2 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_fill_2 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_fill_2 FILLER_6_529 ();
 sg13g2_fill_1 FILLER_6_531 ();
 sg13g2_decap_8 FILLER_6_559 ();
 sg13g2_fill_2 FILLER_6_566 ();
 sg13g2_fill_1 FILLER_6_575 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_fill_2 FILLER_6_595 ();
 sg13g2_fill_1 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_fill_2 FILLER_6_663 ();
 sg13g2_decap_8 FILLER_6_681 ();
 sg13g2_decap_8 FILLER_6_688 ();
 sg13g2_decap_8 FILLER_6_695 ();
 sg13g2_fill_1 FILLER_6_702 ();
 sg13g2_fill_1 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_4 FILLER_6_742 ();
 sg13g2_fill_1 FILLER_6_752 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_772 ();
 sg13g2_decap_8 FILLER_6_779 ();
 sg13g2_decap_8 FILLER_6_786 ();
 sg13g2_fill_1 FILLER_6_793 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_4 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_4 FILLER_7_532 ();
 sg13g2_fill_2 FILLER_7_536 ();
 sg13g2_decap_8 FILLER_7_555 ();
 sg13g2_decap_4 FILLER_7_562 ();
 sg13g2_fill_1 FILLER_7_566 ();
 sg13g2_decap_8 FILLER_7_599 ();
 sg13g2_decap_8 FILLER_7_606 ();
 sg13g2_fill_2 FILLER_7_613 ();
 sg13g2_fill_1 FILLER_7_615 ();
 sg13g2_decap_4 FILLER_7_621 ();
 sg13g2_decap_8 FILLER_7_684 ();
 sg13g2_decap_8 FILLER_7_691 ();
 sg13g2_fill_2 FILLER_7_698 ();
 sg13g2_fill_1 FILLER_7_700 ();
 sg13g2_decap_4 FILLER_7_733 ();
 sg13g2_fill_1 FILLER_7_737 ();
 sg13g2_fill_2 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_484 ();
 sg13g2_fill_1 FILLER_8_491 ();
 sg13g2_decap_8 FILLER_8_498 ();
 sg13g2_decap_8 FILLER_8_505 ();
 sg13g2_fill_2 FILLER_8_512 ();
 sg13g2_fill_1 FILLER_8_514 ();
 sg13g2_decap_8 FILLER_8_520 ();
 sg13g2_decap_4 FILLER_8_527 ();
 sg13g2_fill_1 FILLER_8_531 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_4 FILLER_8_571 ();
 sg13g2_fill_2 FILLER_8_575 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_2 FILLER_8_586 ();
 sg13g2_decap_8 FILLER_8_621 ();
 sg13g2_decap_4 FILLER_8_628 ();
 sg13g2_fill_2 FILLER_8_632 ();
 sg13g2_fill_1 FILLER_8_639 ();
 sg13g2_decap_8 FILLER_8_643 ();
 sg13g2_decap_8 FILLER_8_650 ();
 sg13g2_fill_2 FILLER_8_657 ();
 sg13g2_fill_1 FILLER_8_659 ();
 sg13g2_fill_1 FILLER_8_668 ();
 sg13g2_fill_2 FILLER_8_679 ();
 sg13g2_fill_1 FILLER_8_681 ();
 sg13g2_decap_8 FILLER_8_713 ();
 sg13g2_fill_2 FILLER_8_720 ();
 sg13g2_fill_1 FILLER_8_722 ();
 sg13g2_decap_4 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_fill_1 FILLER_8_773 ();
 sg13g2_decap_4 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_4 FILLER_9_459 ();
 sg13g2_fill_1 FILLER_9_463 ();
 sg13g2_fill_1 FILLER_9_491 ();
 sg13g2_fill_2 FILLER_9_519 ();
 sg13g2_fill_1 FILLER_9_548 ();
 sg13g2_fill_2 FILLER_9_552 ();
 sg13g2_decap_8 FILLER_9_580 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_8 FILLER_9_594 ();
 sg13g2_decap_8 FILLER_9_629 ();
 sg13g2_decap_4 FILLER_9_636 ();
 sg13g2_fill_1 FILLER_9_640 ();
 sg13g2_decap_4 FILLER_9_672 ();
 sg13g2_fill_2 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_691 ();
 sg13g2_fill_2 FILLER_9_698 ();
 sg13g2_fill_1 FILLER_9_700 ();
 sg13g2_fill_2 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_4 FILLER_9_784 ();
 sg13g2_fill_2 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_4 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_478 ();
 sg13g2_fill_2 FILLER_10_485 ();
 sg13g2_fill_1 FILLER_10_487 ();
 sg13g2_decap_4 FILLER_10_493 ();
 sg13g2_fill_2 FILLER_10_509 ();
 sg13g2_fill_2 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_551 ();
 sg13g2_decap_8 FILLER_10_558 ();
 sg13g2_fill_2 FILLER_10_600 ();
 sg13g2_fill_1 FILLER_10_602 ();
 sg13g2_fill_2 FILLER_10_614 ();
 sg13g2_decap_4 FILLER_10_643 ();
 sg13g2_fill_1 FILLER_10_647 ();
 sg13g2_fill_1 FILLER_10_654 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_4 FILLER_10_674 ();
 sg13g2_fill_2 FILLER_10_678 ();
 sg13g2_fill_1 FILLER_10_718 ();
 sg13g2_fill_1 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_fill_2 FILLER_10_762 ();
 sg13g2_fill_1 FILLER_10_768 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_fill_2 FILLER_10_786 ();
 sg13g2_fill_2 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_4 FILLER_11_431 ();
 sg13g2_fill_2 FILLER_11_435 ();
 sg13g2_fill_1 FILLER_11_464 ();
 sg13g2_fill_2 FILLER_11_469 ();
 sg13g2_fill_1 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_499 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_fill_1 FILLER_11_577 ();
 sg13g2_decap_4 FILLER_11_582 ();
 sg13g2_fill_2 FILLER_11_586 ();
 sg13g2_decap_4 FILLER_11_615 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_4 FILLER_11_641 ();
 sg13g2_fill_1 FILLER_11_645 ();
 sg13g2_decap_8 FILLER_11_687 ();
 sg13g2_fill_2 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_4 FILLER_11_738 ();
 sg13g2_fill_1 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_765 ();
 sg13g2_decap_4 FILLER_11_772 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_fill_2 FILLER_11_821 ();
 sg13g2_decap_4 FILLER_12_4 ();
 sg13g2_fill_1 FILLER_12_8 ();
 sg13g2_decap_8 FILLER_12_13 ();
 sg13g2_decap_8 FILLER_12_20 ();
 sg13g2_decap_8 FILLER_12_27 ();
 sg13g2_decap_8 FILLER_12_34 ();
 sg13g2_decap_8 FILLER_12_41 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_decap_8 FILLER_12_55 ();
 sg13g2_decap_8 FILLER_12_62 ();
 sg13g2_decap_8 FILLER_12_69 ();
 sg13g2_decap_8 FILLER_12_76 ();
 sg13g2_decap_8 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_90 ();
 sg13g2_decap_8 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_104 ();
 sg13g2_decap_8 FILLER_12_111 ();
 sg13g2_decap_8 FILLER_12_118 ();
 sg13g2_decap_8 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_decap_8 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_decap_8 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_251 ();
 sg13g2_decap_8 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_265 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_12_419 ();
 sg13g2_decap_8 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_12_433 ();
 sg13g2_fill_2 FILLER_12_440 ();
 sg13g2_decap_4 FILLER_12_448 ();
 sg13g2_fill_1 FILLER_12_452 ();
 sg13g2_fill_1 FILLER_12_456 ();
 sg13g2_fill_2 FILLER_12_520 ();
 sg13g2_fill_1 FILLER_12_531 ();
 sg13g2_decap_4 FILLER_12_559 ();
 sg13g2_fill_1 FILLER_12_563 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_4 FILLER_12_595 ();
 sg13g2_fill_2 FILLER_12_622 ();
 sg13g2_fill_1 FILLER_12_624 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_fill_2 FILLER_12_662 ();
 sg13g2_fill_1 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_4 FILLER_12_686 ();
 sg13g2_fill_1 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_fill_2 FILLER_12_709 ();
 sg13g2_fill_1 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_4 FILLER_12_735 ();
 sg13g2_fill_1 FILLER_12_739 ();
 sg13g2_fill_1 FILLER_12_751 ();
 sg13g2_decap_8 FILLER_12_779 ();
 sg13g2_decap_4 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_4 FILLER_13_431 ();
 sg13g2_fill_1 FILLER_13_435 ();
 sg13g2_decap_8 FILLER_13_458 ();
 sg13g2_decap_4 FILLER_13_465 ();
 sg13g2_decap_8 FILLER_13_478 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_decap_8 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_499 ();
 sg13g2_fill_1 FILLER_13_506 ();
 sg13g2_decap_8 FILLER_13_510 ();
 sg13g2_fill_2 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_fill_1 FILLER_13_567 ();
 sg13g2_fill_1 FILLER_13_573 ();
 sg13g2_fill_1 FILLER_13_606 ();
 sg13g2_fill_2 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_659 ();
 sg13g2_fill_2 FILLER_13_666 ();
 sg13g2_decap_8 FILLER_13_702 ();
 sg13g2_decap_8 FILLER_13_713 ();
 sg13g2_fill_2 FILLER_13_720 ();
 sg13g2_fill_2 FILLER_13_749 ();
 sg13g2_fill_1 FILLER_13_756 ();
 sg13g2_fill_2 FILLER_13_761 ();
 sg13g2_decap_4 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_808 ();
 sg13g2_decap_8 FILLER_13_815 ();
 sg13g2_fill_1 FILLER_13_822 ();
 sg13g2_decap_4 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_8 ();
 sg13g2_decap_8 FILLER_14_13 ();
 sg13g2_decap_8 FILLER_14_20 ();
 sg13g2_decap_8 FILLER_14_27 ();
 sg13g2_decap_8 FILLER_14_34 ();
 sg13g2_decap_8 FILLER_14_41 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_decap_8 FILLER_14_55 ();
 sg13g2_decap_8 FILLER_14_62 ();
 sg13g2_decap_8 FILLER_14_69 ();
 sg13g2_decap_8 FILLER_14_76 ();
 sg13g2_decap_8 FILLER_14_83 ();
 sg13g2_decap_8 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_97 ();
 sg13g2_decap_8 FILLER_14_104 ();
 sg13g2_decap_8 FILLER_14_111 ();
 sg13g2_decap_8 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_decap_8 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_decap_8 FILLER_14_174 ();
 sg13g2_decap_8 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_decap_8 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_4 FILLER_14_419 ();
 sg13g2_decap_8 FILLER_14_484 ();
 sg13g2_decap_4 FILLER_14_491 ();
 sg13g2_fill_1 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_535 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_fill_2 FILLER_14_605 ();
 sg13g2_fill_1 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_622 ();
 sg13g2_fill_2 FILLER_14_629 ();
 sg13g2_decap_4 FILLER_14_635 ();
 sg13g2_fill_2 FILLER_14_639 ();
 sg13g2_fill_1 FILLER_14_646 ();
 sg13g2_decap_4 FILLER_14_685 ();
 sg13g2_fill_1 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_764 ();
 sg13g2_decap_8 FILLER_14_771 ();
 sg13g2_decap_8 FILLER_14_778 ();
 sg13g2_decap_4 FILLER_14_785 ();
 sg13g2_fill_1 FILLER_14_789 ();
 sg13g2_fill_1 FILLER_14_822 ();
 sg13g2_decap_4 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_8 ();
 sg13g2_decap_8 FILLER_15_13 ();
 sg13g2_decap_8 FILLER_15_20 ();
 sg13g2_decap_8 FILLER_15_27 ();
 sg13g2_decap_8 FILLER_15_34 ();
 sg13g2_decap_8 FILLER_15_41 ();
 sg13g2_decap_8 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_62 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_139 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_decap_8 FILLER_15_160 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_230 ();
 sg13g2_decap_8 FILLER_15_237 ();
 sg13g2_decap_8 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_4 FILLER_15_419 ();
 sg13g2_decap_8 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_15_435 ();
 sg13g2_fill_1 FILLER_15_442 ();
 sg13g2_fill_2 FILLER_15_454 ();
 sg13g2_decap_4 FILLER_15_462 ();
 sg13g2_fill_2 FILLER_15_466 ();
 sg13g2_fill_2 FILLER_15_508 ();
 sg13g2_fill_1 FILLER_15_510 ();
 sg13g2_decap_4 FILLER_15_516 ();
 sg13g2_decap_8 FILLER_15_555 ();
 sg13g2_decap_4 FILLER_15_562 ();
 sg13g2_fill_2 FILLER_15_566 ();
 sg13g2_decap_8 FILLER_15_586 ();
 sg13g2_fill_1 FILLER_15_593 ();
 sg13g2_decap_4 FILLER_15_651 ();
 sg13g2_fill_1 FILLER_15_655 ();
 sg13g2_decap_4 FILLER_15_659 ();
 sg13g2_fill_1 FILLER_15_663 ();
 sg13g2_decap_8 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_698 ();
 sg13g2_decap_8 FILLER_15_705 ();
 sg13g2_decap_4 FILLER_15_712 ();
 sg13g2_fill_1 FILLER_15_716 ();
 sg13g2_fill_2 FILLER_15_747 ();
 sg13g2_fill_1 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_4 FILLER_15_784 ();
 sg13g2_fill_1 FILLER_15_788 ();
 sg13g2_fill_2 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_810 ();
 sg13g2_decap_4 FILLER_15_817 ();
 sg13g2_fill_2 FILLER_15_821 ();
 sg13g2_decap_4 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_8 ();
 sg13g2_decap_8 FILLER_16_13 ();
 sg13g2_decap_8 FILLER_16_20 ();
 sg13g2_decap_8 FILLER_16_27 ();
 sg13g2_decap_8 FILLER_16_34 ();
 sg13g2_decap_8 FILLER_16_41 ();
 sg13g2_decap_8 FILLER_16_48 ();
 sg13g2_decap_8 FILLER_16_55 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_decap_8 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_83 ();
 sg13g2_decap_8 FILLER_16_90 ();
 sg13g2_decap_8 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_195 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_4 FILLER_16_391 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_451 ();
 sg13g2_decap_4 FILLER_16_484 ();
 sg13g2_fill_2 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_493 ();
 sg13g2_decap_8 FILLER_16_500 ();
 sg13g2_fill_2 FILLER_16_514 ();
 sg13g2_fill_1 FILLER_16_516 ();
 sg13g2_decap_4 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_524 ();
 sg13g2_decap_8 FILLER_16_544 ();
 sg13g2_decap_8 FILLER_16_551 ();
 sg13g2_fill_1 FILLER_16_558 ();
 sg13g2_fill_2 FILLER_16_565 ();
 sg13g2_fill_1 FILLER_16_567 ();
 sg13g2_fill_2 FILLER_16_576 ();
 sg13g2_fill_1 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_4 FILLER_16_628 ();
 sg13g2_fill_2 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_8 FILLER_16_666 ();
 sg13g2_decap_4 FILLER_16_699 ();
 sg13g2_fill_2 FILLER_16_706 ();
 sg13g2_fill_2 FILLER_16_747 ();
 sg13g2_fill_1 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_755 ();
 sg13g2_fill_1 FILLER_16_762 ();
 sg13g2_fill_1 FILLER_16_800 ();
 sg13g2_fill_2 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_4 FILLER_16_818 ();
 sg13g2_fill_1 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_13 ();
 sg13g2_decap_8 FILLER_17_20 ();
 sg13g2_decap_8 FILLER_17_27 ();
 sg13g2_decap_8 FILLER_17_34 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_48 ();
 sg13g2_decap_8 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_62 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_decap_8 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_90 ();
 sg13g2_decap_8 FILLER_17_97 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_125 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_decap_8 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_decap_8 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_4 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_1 FILLER_17_402 ();
 sg13g2_fill_2 FILLER_17_424 ();
 sg13g2_fill_1 FILLER_17_426 ();
 sg13g2_fill_2 FILLER_17_433 ();
 sg13g2_decap_8 FILLER_17_442 ();
 sg13g2_decap_8 FILLER_17_449 ();
 sg13g2_decap_4 FILLER_17_456 ();
 sg13g2_decap_8 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_492 ();
 sg13g2_fill_2 FILLER_17_527 ();
 sg13g2_fill_1 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_decap_4 FILLER_17_604 ();
 sg13g2_fill_2 FILLER_17_608 ();
 sg13g2_fill_2 FILLER_17_648 ();
 sg13g2_fill_1 FILLER_17_650 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_fill_2 FILLER_17_663 ();
 sg13g2_fill_1 FILLER_17_665 ();
 sg13g2_fill_2 FILLER_17_726 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_decap_4 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_769 ();
 sg13g2_decap_4 FILLER_17_776 ();
 sg13g2_fill_2 FILLER_17_780 ();
 sg13g2_fill_1 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_4 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_433 ();
 sg13g2_fill_1 FILLER_18_440 ();
 sg13g2_decap_8 FILLER_18_446 ();
 sg13g2_decap_8 FILLER_18_453 ();
 sg13g2_decap_4 FILLER_18_460 ();
 sg13g2_fill_2 FILLER_18_464 ();
 sg13g2_fill_2 FILLER_18_498 ();
 sg13g2_fill_1 FILLER_18_500 ();
 sg13g2_fill_2 FILLER_18_553 ();
 sg13g2_decap_4 FILLER_18_563 ();
 sg13g2_decap_8 FILLER_18_579 ();
 sg13g2_decap_8 FILLER_18_586 ();
 sg13g2_decap_8 FILLER_18_593 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_decap_4 FILLER_18_624 ();
 sg13g2_fill_1 FILLER_18_628 ();
 sg13g2_fill_2 FILLER_18_636 ();
 sg13g2_fill_1 FILLER_18_642 ();
 sg13g2_decap_8 FILLER_18_680 ();
 sg13g2_decap_4 FILLER_18_687 ();
 sg13g2_fill_2 FILLER_18_691 ();
 sg13g2_decap_4 FILLER_18_700 ();
 sg13g2_fill_2 FILLER_18_704 ();
 sg13g2_decap_4 FILLER_18_719 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_4 FILLER_18_753 ();
 sg13g2_fill_1 FILLER_18_757 ();
 sg13g2_decap_8 FILLER_18_762 ();
 sg13g2_decap_8 FILLER_18_769 ();
 sg13g2_fill_1 FILLER_18_776 ();
 sg13g2_fill_1 FILLER_18_783 ();
 sg13g2_fill_2 FILLER_18_789 ();
 sg13g2_fill_1 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_797 ();
 sg13g2_decap_8 FILLER_18_804 ();
 sg13g2_decap_8 FILLER_18_811 ();
 sg13g2_decap_4 FILLER_18_818 ();
 sg13g2_fill_1 FILLER_18_822 ();
 sg13g2_decap_4 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_8 ();
 sg13g2_decap_8 FILLER_19_13 ();
 sg13g2_decap_8 FILLER_19_20 ();
 sg13g2_decap_8 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_34 ();
 sg13g2_decap_8 FILLER_19_41 ();
 sg13g2_decap_8 FILLER_19_48 ();
 sg13g2_decap_8 FILLER_19_55 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_decap_8 FILLER_19_83 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_decap_8 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_decap_8 FILLER_19_132 ();
 sg13g2_decap_8 FILLER_19_139 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_4 FILLER_19_272 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_decap_4 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_fill_2 FILLER_19_464 ();
 sg13g2_fill_1 FILLER_19_466 ();
 sg13g2_decap_8 FILLER_19_494 ();
 sg13g2_fill_2 FILLER_19_501 ();
 sg13g2_fill_1 FILLER_19_503 ();
 sg13g2_fill_2 FILLER_19_509 ();
 sg13g2_decap_8 FILLER_19_516 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_8 FILLER_19_530 ();
 sg13g2_fill_1 FILLER_19_537 ();
 sg13g2_fill_1 FILLER_19_543 ();
 sg13g2_fill_1 FILLER_19_569 ();
 sg13g2_decap_4 FILLER_19_624 ();
 sg13g2_decap_8 FILLER_19_646 ();
 sg13g2_decap_8 FILLER_19_653 ();
 sg13g2_decap_8 FILLER_19_660 ();
 sg13g2_decap_4 FILLER_19_667 ();
 sg13g2_decap_8 FILLER_19_675 ();
 sg13g2_decap_8 FILLER_19_682 ();
 sg13g2_fill_1 FILLER_19_689 ();
 sg13g2_fill_1 FILLER_19_695 ();
 sg13g2_fill_2 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_709 ();
 sg13g2_fill_1 FILLER_19_716 ();
 sg13g2_fill_2 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_4 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_8 ();
 sg13g2_decap_8 FILLER_20_13 ();
 sg13g2_decap_8 FILLER_20_20 ();
 sg13g2_decap_8 FILLER_20_27 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_decap_8 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_decap_4 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_decap_4 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_4 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_decap_4 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_4 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_decap_4 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_fill_1 FILLER_20_438 ();
 sg13g2_fill_2 FILLER_20_469 ();
 sg13g2_decap_4 FILLER_20_505 ();
 sg13g2_fill_1 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_528 ();
 sg13g2_fill_2 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_572 ();
 sg13g2_fill_1 FILLER_20_574 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_decap_4 FILLER_20_592 ();
 sg13g2_fill_2 FILLER_20_596 ();
 sg13g2_fill_1 FILLER_20_603 ();
 sg13g2_fill_2 FILLER_20_616 ();
 sg13g2_fill_1 FILLER_20_618 ();
 sg13g2_fill_1 FILLER_20_622 ();
 sg13g2_fill_1 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_661 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_fill_2 FILLER_20_675 ();
 sg13g2_fill_1 FILLER_20_680 ();
 sg13g2_fill_1 FILLER_20_717 ();
 sg13g2_decap_4 FILLER_20_736 ();
 sg13g2_fill_2 FILLER_20_743 ();
 sg13g2_decap_4 FILLER_20_751 ();
 sg13g2_fill_2 FILLER_20_755 ();
 sg13g2_decap_4 FILLER_20_760 ();
 sg13g2_fill_1 FILLER_20_764 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_fill_2 FILLER_20_775 ();
 sg13g2_fill_1 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_4 FILLER_20_799 ();
 sg13g2_decap_4 FILLER_20_806 ();
 sg13g2_fill_1 FILLER_20_810 ();
 sg13g2_decap_4 FILLER_20_814 ();
 sg13g2_fill_2 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_21_8 ();
 sg13g2_decap_4 FILLER_21_15 ();
 sg13g2_decap_8 FILLER_21_23 ();
 sg13g2_decap_8 FILLER_21_30 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_8 FILLER_21_44 ();
 sg13g2_decap_4 FILLER_21_51 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_131 ();
 sg13g2_decap_8 FILLER_21_138 ();
 sg13g2_decap_8 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_152 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_decap_8 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_decap_8 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_fill_2 FILLER_21_398 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_4 FILLER_21_410 ();
 sg13g2_fill_1 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_425 ();
 sg13g2_decap_8 FILLER_21_432 ();
 sg13g2_decap_4 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_443 ();
 sg13g2_fill_2 FILLER_21_450 ();
 sg13g2_fill_1 FILLER_21_452 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_465 ();
 sg13g2_fill_2 FILLER_21_484 ();
 sg13g2_fill_1 FILLER_21_489 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_13 ();
 sg13g2_decap_8 FILLER_22_20 ();
 sg13g2_decap_4 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_decap_8 FILLER_22_250 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_4 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_4 FILLER_22_401 ();
 sg13g2_fill_2 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_465 ();
 sg13g2_fill_2 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_479 ();
 sg13g2_fill_1 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_fill_2 FILLER_22_497 ();
 sg13g2_fill_2 FILLER_22_517 ();
 sg13g2_decap_8 FILLER_22_530 ();
 sg13g2_fill_1 FILLER_22_537 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_13 ();
 sg13g2_decap_8 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_27 ();
 sg13g2_decap_8 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_fill_1 FILLER_23_68 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_191 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_decap_8 FILLER_23_219 ();
 sg13g2_decap_8 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_decap_8 FILLER_23_240 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_8 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_282 ();
 sg13g2_decap_8 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_503 ();
 sg13g2_fill_2 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_fill_1 FILLER_23_543 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_4 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_decap_8 FILLER_24_43 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_fill_2 FILLER_24_57 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_4 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_325 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_395 ();
 sg13g2_decap_4 FILLER_24_457 ();
 sg13g2_fill_2 FILLER_24_461 ();
 sg13g2_fill_1 FILLER_24_473 ();
 sg13g2_fill_1 FILLER_24_490 ();
 sg13g2_fill_2 FILLER_24_515 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_decap_8 FILLER_25_117 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_decap_8 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_243 ();
 sg13g2_decap_8 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_257 ();
 sg13g2_decap_8 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_4 FILLER_25_349 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_410 ();
 sg13g2_fill_2 FILLER_25_437 ();
 sg13g2_decap_4 FILLER_25_493 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_fill_1 FILLER_25_543 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_6 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_4 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_4 FILLER_26_442 ();
 sg13g2_fill_2 FILLER_26_446 ();
 sg13g2_decap_8 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_decap_8 FILLER_26_466 ();
 sg13g2_decap_4 FILLER_26_473 ();
 sg13g2_fill_2 FILLER_26_477 ();
 sg13g2_fill_1 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_487 ();
 sg13g2_decap_8 FILLER_26_494 ();
 sg13g2_fill_1 FILLER_26_501 ();
 sg13g2_fill_1 FILLER_26_508 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_4 FILLER_26_531 ();
 sg13g2_fill_2 FILLER_26_535 ();
 sg13g2_fill_1 FILLER_26_543 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_decap_4 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_2 FILLER_27_429 ();
 sg13g2_fill_1 FILLER_27_431 ();
 sg13g2_decap_8 FILLER_27_464 ();
 sg13g2_fill_2 FILLER_27_485 ();
 sg13g2_fill_2 FILLER_27_524 ();
 sg13g2_fill_1 FILLER_27_529 ();
 sg13g2_fill_1 FILLER_27_536 ();
 sg13g2_fill_1 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_4 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_4 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_4 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_4 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_438 ();
 sg13g2_fill_2 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_492 ();
 sg13g2_decap_8 FILLER_28_499 ();
 sg13g2_fill_1 FILLER_28_506 ();
 sg13g2_decap_4 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_8 ();
 sg13g2_decap_8 FILLER_29_13 ();
 sg13g2_decap_8 FILLER_29_20 ();
 sg13g2_decap_8 FILLER_29_27 ();
 sg13g2_decap_8 FILLER_29_34 ();
 sg13g2_decap_8 FILLER_29_41 ();
 sg13g2_decap_8 FILLER_29_48 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_decap_8 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_69 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_448 ();
 sg13g2_decap_4 FILLER_29_455 ();
 sg13g2_fill_2 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_471 ();
 sg13g2_fill_2 FILLER_29_504 ();
 sg13g2_fill_2 FILLER_29_509 ();
 sg13g2_fill_2 FILLER_29_525 ();
 sg13g2_fill_1 FILLER_29_527 ();
 sg13g2_fill_2 FILLER_29_532 ();
 sg13g2_fill_1 FILLER_29_534 ();
 sg13g2_decap_4 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_8 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_decap_8 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_39 ();
 sg13g2_decap_8 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_decap_8 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_decap_8 FILLER_30_109 ();
 sg13g2_decap_8 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_443 ();
 sg13g2_fill_1 FILLER_30_452 ();
 sg13g2_decap_8 FILLER_30_458 ();
 sg13g2_decap_8 FILLER_30_465 ();
 sg13g2_decap_8 FILLER_30_472 ();
 sg13g2_decap_8 FILLER_30_479 ();
 sg13g2_decap_4 FILLER_30_491 ();
 sg13g2_fill_1 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_fill_1 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_4 FILLER_30_549 ();
 sg13g2_fill_1 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_559 ();
 sg13g2_fill_2 FILLER_30_569 ();
 sg13g2_fill_1 FILLER_30_571 ();
 sg13g2_fill_1 FILLER_30_575 ();
 sg13g2_fill_1 FILLER_30_579 ();
 sg13g2_fill_2 FILLER_30_593 ();
 sg13g2_decap_8 FILLER_30_598 ();
 sg13g2_decap_4 FILLER_30_605 ();
 sg13g2_fill_2 FILLER_30_609 ();
 sg13g2_decap_4 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_633 ();
 sg13g2_fill_2 FILLER_30_643 ();
 sg13g2_fill_2 FILLER_30_648 ();
 sg13g2_fill_1 FILLER_30_650 ();
 sg13g2_decap_4 FILLER_30_654 ();
 sg13g2_fill_1 FILLER_30_658 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_fill_1 FILLER_30_671 ();
 sg13g2_fill_2 FILLER_30_678 ();
 sg13g2_fill_1 FILLER_30_712 ();
 sg13g2_decap_4 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_734 ();
 sg13g2_fill_2 FILLER_30_740 ();
 sg13g2_fill_1 FILLER_30_742 ();
 sg13g2_fill_1 FILLER_30_746 ();
 sg13g2_fill_1 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_754 ();
 sg13g2_decap_8 FILLER_30_761 ();
 sg13g2_decap_4 FILLER_30_768 ();
 sg13g2_fill_1 FILLER_30_772 ();
 sg13g2_fill_2 FILLER_30_778 ();
 sg13g2_fill_2 FILLER_30_783 ();
 sg13g2_fill_1 FILLER_30_785 ();
 sg13g2_fill_1 FILLER_30_796 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_4 FILLER_30_807 ();
 sg13g2_fill_2 FILLER_30_811 ();
 sg13g2_decap_4 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_20 ();
 sg13g2_decap_8 FILLER_31_27 ();
 sg13g2_decap_8 FILLER_31_34 ();
 sg13g2_decap_8 FILLER_31_41 ();
 sg13g2_decap_8 FILLER_31_48 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_69 ();
 sg13g2_decap_8 FILLER_31_76 ();
 sg13g2_decap_8 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_90 ();
 sg13g2_decap_8 FILLER_31_97 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_decap_8 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_230 ();
 sg13g2_decap_8 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_258 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_4 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_610 ();
 sg13g2_fill_1 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_640 ();
 sg13g2_fill_1 FILLER_31_647 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_decap_4 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_696 ();
 sg13g2_decap_4 FILLER_31_703 ();
 sg13g2_fill_2 FILLER_31_707 ();
 sg13g2_decap_4 FILLER_31_767 ();
 sg13g2_fill_2 FILLER_31_771 ();
 sg13g2_fill_1 FILLER_31_786 ();
 sg13g2_decap_4 FILLER_31_818 ();
 sg13g2_fill_1 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_4 FILLER_32_382 ();
 sg13g2_decap_4 FILLER_32_389 ();
 sg13g2_decap_4 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_32_402 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_decap_4 FILLER_32_423 ();
 sg13g2_fill_1 FILLER_32_427 ();
 sg13g2_fill_2 FILLER_32_440 ();
 sg13g2_fill_2 FILLER_32_454 ();
 sg13g2_fill_2 FILLER_32_466 ();
 sg13g2_decap_8 FILLER_32_471 ();
 sg13g2_decap_8 FILLER_32_478 ();
 sg13g2_decap_4 FILLER_32_485 ();
 sg13g2_fill_2 FILLER_32_489 ();
 sg13g2_decap_8 FILLER_32_498 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_540 ();
 sg13g2_decap_4 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_551 ();
 sg13g2_decap_8 FILLER_32_564 ();
 sg13g2_decap_8 FILLER_32_571 ();
 sg13g2_decap_4 FILLER_32_578 ();
 sg13g2_fill_2 FILLER_32_589 ();
 sg13g2_fill_1 FILLER_32_591 ();
 sg13g2_decap_4 FILLER_32_597 ();
 sg13g2_fill_1 FILLER_32_601 ();
 sg13g2_fill_2 FILLER_32_655 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_decap_4 FILLER_32_671 ();
 sg13g2_fill_2 FILLER_32_691 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_fill_2 FILLER_32_705 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_fill_1 FILLER_32_711 ();
 sg13g2_decap_4 FILLER_32_727 ();
 sg13g2_fill_2 FILLER_32_731 ();
 sg13g2_fill_2 FILLER_32_740 ();
 sg13g2_fill_1 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_fill_1 FILLER_32_755 ();
 sg13g2_decap_4 FILLER_32_788 ();
 sg13g2_fill_1 FILLER_32_792 ();
 sg13g2_fill_1 FILLER_32_798 ();
 sg13g2_fill_2 FILLER_32_804 ();
 sg13g2_fill_1 FILLER_32_806 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_decap_4 FILLER_32_817 ();
 sg13g2_fill_2 FILLER_32_821 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_81 ();
 sg13g2_decap_8 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_452 ();
 sg13g2_decap_4 FILLER_33_487 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_fill_2 FILLER_33_558 ();
 sg13g2_decap_4 FILLER_33_569 ();
 sg13g2_fill_2 FILLER_33_573 ();
 sg13g2_fill_1 FILLER_33_617 ();
 sg13g2_fill_1 FILLER_33_627 ();
 sg13g2_fill_1 FILLER_33_635 ();
 sg13g2_decap_8 FILLER_33_641 ();
 sg13g2_decap_4 FILLER_33_648 ();
 sg13g2_fill_2 FILLER_33_679 ();
 sg13g2_fill_1 FILLER_33_681 ();
 sg13g2_fill_1 FILLER_33_709 ();
 sg13g2_fill_1 FILLER_33_716 ();
 sg13g2_fill_2 FILLER_33_726 ();
 sg13g2_decap_4 FILLER_33_737 ();
 sg13g2_decap_4 FILLER_33_746 ();
 sg13g2_fill_2 FILLER_33_755 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_fill_2 FILLER_33_774 ();
 sg13g2_fill_1 FILLER_33_776 ();
 sg13g2_fill_2 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_4 FILLER_34_399 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_2 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_34_431 ();
 sg13g2_decap_8 FILLER_34_463 ();
 sg13g2_decap_8 FILLER_34_470 ();
 sg13g2_decap_8 FILLER_34_477 ();
 sg13g2_decap_4 FILLER_34_500 ();
 sg13g2_decap_8 FILLER_34_507 ();
 sg13g2_decap_8 FILLER_34_514 ();
 sg13g2_fill_2 FILLER_34_521 ();
 sg13g2_fill_1 FILLER_34_555 ();
 sg13g2_decap_8 FILLER_34_583 ();
 sg13g2_decap_8 FILLER_34_590 ();
 sg13g2_decap_4 FILLER_34_597 ();
 sg13g2_fill_1 FILLER_34_601 ();
 sg13g2_decap_8 FILLER_34_640 ();
 sg13g2_decap_8 FILLER_34_647 ();
 sg13g2_fill_2 FILLER_34_654 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_fill_1 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_fill_2 FILLER_34_700 ();
 sg13g2_fill_2 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_fill_2 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_4 FILLER_35_406 ();
 sg13g2_fill_2 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_decap_4 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_458 ();
 sg13g2_decap_4 FILLER_35_465 ();
 sg13g2_fill_2 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_475 ();
 sg13g2_decap_4 FILLER_35_482 ();
 sg13g2_decap_8 FILLER_35_528 ();
 sg13g2_fill_1 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_4 FILLER_35_588 ();
 sg13g2_fill_1 FILLER_35_597 ();
 sg13g2_decap_4 FILLER_35_601 ();
 sg13g2_fill_1 FILLER_35_605 ();
 sg13g2_fill_2 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_624 ();
 sg13g2_decap_8 FILLER_35_636 ();
 sg13g2_fill_1 FILLER_35_670 ();
 sg13g2_fill_2 FILLER_35_683 ();
 sg13g2_fill_1 FILLER_35_685 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_fill_2 FILLER_35_703 ();
 sg13g2_fill_1 FILLER_35_705 ();
 sg13g2_fill_1 FILLER_35_733 ();
 sg13g2_fill_1 FILLER_35_737 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_752 ();
 sg13g2_decap_8 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_fill_2 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_493 ();
 sg13g2_decap_8 FILLER_36_500 ();
 sg13g2_decap_4 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_550 ();
 sg13g2_decap_8 FILLER_36_557 ();
 sg13g2_fill_2 FILLER_36_564 ();
 sg13g2_fill_1 FILLER_36_566 ();
 sg13g2_decap_8 FILLER_36_570 ();
 sg13g2_fill_1 FILLER_36_577 ();
 sg13g2_decap_4 FILLER_36_610 ();
 sg13g2_fill_2 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_622 ();
 sg13g2_fill_2 FILLER_36_644 ();
 sg13g2_fill_1 FILLER_36_646 ();
 sg13g2_decap_4 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_decap_4 FILLER_36_722 ();
 sg13g2_fill_1 FILLER_36_726 ();
 sg13g2_fill_2 FILLER_36_738 ();
 sg13g2_fill_1 FILLER_36_740 ();
 sg13g2_fill_1 FILLER_36_750 ();
 sg13g2_decap_4 FILLER_36_756 ();
 sg13g2_decap_4 FILLER_36_763 ();
 sg13g2_fill_2 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_fill_2 FILLER_36_820 ();
 sg13g2_fill_1 FILLER_36_822 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_decap_8 FILLER_37_426 ();
 sg13g2_decap_4 FILLER_37_433 ();
 sg13g2_decap_8 FILLER_37_447 ();
 sg13g2_decap_8 FILLER_37_454 ();
 sg13g2_decap_8 FILLER_37_461 ();
 sg13g2_decap_8 FILLER_37_468 ();
 sg13g2_decap_4 FILLER_37_475 ();
 sg13g2_fill_2 FILLER_37_490 ();
 sg13g2_fill_1 FILLER_37_492 ();
 sg13g2_fill_2 FILLER_37_505 ();
 sg13g2_decap_8 FILLER_37_540 ();
 sg13g2_fill_2 FILLER_37_579 ();
 sg13g2_decap_4 FILLER_37_594 ();
 sg13g2_fill_1 FILLER_37_598 ();
 sg13g2_decap_4 FILLER_37_602 ();
 sg13g2_fill_2 FILLER_37_671 ();
 sg13g2_fill_2 FILLER_37_677 ();
 sg13g2_fill_2 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_698 ();
 sg13g2_fill_1 FILLER_37_705 ();
 sg13g2_fill_2 FILLER_37_743 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_4 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_fill_1 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_425 ();
 sg13g2_decap_8 FILLER_38_432 ();
 sg13g2_decap_8 FILLER_38_439 ();
 sg13g2_decap_8 FILLER_38_446 ();
 sg13g2_decap_8 FILLER_38_453 ();
 sg13g2_decap_4 FILLER_38_460 ();
 sg13g2_fill_2 FILLER_38_464 ();
 sg13g2_fill_1 FILLER_38_496 ();
 sg13g2_fill_1 FILLER_38_528 ();
 sg13g2_fill_2 FILLER_38_534 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_fill_2 FILLER_38_553 ();
 sg13g2_fill_2 FILLER_38_575 ();
 sg13g2_fill_1 FILLER_38_582 ();
 sg13g2_decap_8 FILLER_38_618 ();
 sg13g2_fill_1 FILLER_38_625 ();
 sg13g2_decap_8 FILLER_38_642 ();
 sg13g2_decap_8 FILLER_38_649 ();
 sg13g2_decap_8 FILLER_38_656 ();
 sg13g2_decap_4 FILLER_38_663 ();
 sg13g2_fill_1 FILLER_38_667 ();
 sg13g2_fill_1 FILLER_38_679 ();
 sg13g2_fill_1 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_722 ();
 sg13g2_fill_1 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_754 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_4 FILLER_38_774 ();
 sg13g2_fill_1 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_4 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_500 ();
 sg13g2_decap_8 FILLER_39_507 ();
 sg13g2_fill_2 FILLER_39_514 ();
 sg13g2_decap_4 FILLER_39_548 ();
 sg13g2_decap_8 FILLER_39_583 ();
 sg13g2_fill_1 FILLER_39_590 ();
 sg13g2_decap_4 FILLER_39_623 ();
 sg13g2_fill_1 FILLER_39_659 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_fill_1 FILLER_39_702 ();
 sg13g2_decap_4 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_4 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_fill_2 FILLER_40_511 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_fill_2 FILLER_40_531 ();
 sg13g2_decap_8 FILLER_40_572 ();
 sg13g2_decap_8 FILLER_40_579 ();
 sg13g2_fill_2 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_decap_8 FILLER_40_612 ();
 sg13g2_decap_8 FILLER_40_619 ();
 sg13g2_fill_1 FILLER_40_626 ();
 sg13g2_decap_8 FILLER_40_639 ();
 sg13g2_decap_4 FILLER_40_646 ();
 sg13g2_fill_2 FILLER_40_650 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_decap_8 FILLER_40_669 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_decap_4 FILLER_40_688 ();
 sg13g2_fill_2 FILLER_40_724 ();
 sg13g2_fill_1 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_765 ();
 sg13g2_fill_1 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_771 ();
 sg13g2_decap_8 FILLER_40_778 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_fill_2 FILLER_41_518 ();
 sg13g2_fill_1 FILLER_41_560 ();
 sg13g2_fill_1 FILLER_41_588 ();
 sg13g2_fill_1 FILLER_41_625 ();
 sg13g2_fill_2 FILLER_41_632 ();
 sg13g2_decap_8 FILLER_41_639 ();
 sg13g2_fill_1 FILLER_41_646 ();
 sg13g2_decap_4 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_fill_2 FILLER_41_691 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_fill_2 FILLER_41_704 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_fill_2 FILLER_41_735 ();
 sg13g2_fill_1 FILLER_41_737 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_fill_2 FILLER_41_786 ();
 sg13g2_fill_1 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_fill_1 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_516 ();
 sg13g2_fill_1 FILLER_42_518 ();
 sg13g2_fill_2 FILLER_42_559 ();
 sg13g2_fill_1 FILLER_42_561 ();
 sg13g2_fill_2 FILLER_42_573 ();
 sg13g2_decap_8 FILLER_42_580 ();
 sg13g2_decap_8 FILLER_42_587 ();
 sg13g2_decap_8 FILLER_42_594 ();
 sg13g2_decap_8 FILLER_42_601 ();
 sg13g2_decap_8 FILLER_42_608 ();
 sg13g2_decap_4 FILLER_42_615 ();
 sg13g2_fill_1 FILLER_42_619 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_4 FILLER_42_669 ();
 sg13g2_fill_2 FILLER_42_673 ();
 sg13g2_decap_8 FILLER_42_705 ();
 sg13g2_decap_8 FILLER_42_712 ();
 sg13g2_fill_1 FILLER_42_719 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_506 ();
 sg13g2_fill_1 FILLER_43_537 ();
 sg13g2_fill_1 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_4 FILLER_43_607 ();
 sg13g2_fill_1 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_627 ();
 sg13g2_fill_2 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_636 ();
 sg13g2_decap_8 FILLER_43_641 ();
 sg13g2_decap_8 FILLER_43_648 ();
 sg13g2_fill_2 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_4 FILLER_43_684 ();
 sg13g2_fill_1 FILLER_43_688 ();
 sg13g2_decap_8 FILLER_43_726 ();
 sg13g2_fill_2 FILLER_43_733 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_fill_2 FILLER_43_746 ();
 sg13g2_fill_1 FILLER_43_748 ();
 sg13g2_decap_8 FILLER_43_752 ();
 sg13g2_decap_8 FILLER_43_759 ();
 sg13g2_decap_4 FILLER_43_766 ();
 sg13g2_fill_2 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_4 FILLER_43_782 ();
 sg13g2_fill_2 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_4 FILLER_43_817 ();
 sg13g2_fill_2 FILLER_43_821 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_fill_2 FILLER_44_532 ();
 sg13g2_fill_1 FILLER_44_540 ();
 sg13g2_decap_4 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_580 ();
 sg13g2_fill_2 FILLER_44_587 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_fill_2 FILLER_44_599 ();
 sg13g2_fill_1 FILLER_44_601 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_fill_1 FILLER_44_641 ();
 sg13g2_fill_2 FILLER_44_648 ();
 sg13g2_fill_1 FILLER_44_662 ();
 sg13g2_fill_2 FILLER_44_690 ();
 sg13g2_fill_2 FILLER_44_705 ();
 sg13g2_fill_1 FILLER_44_707 ();
 sg13g2_decap_4 FILLER_44_713 ();
 sg13g2_fill_1 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_4 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_813 ();
 sg13g2_fill_2 FILLER_44_820 ();
 sg13g2_fill_1 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_594 ();
 sg13g2_decap_4 FILLER_45_614 ();
 sg13g2_fill_2 FILLER_45_618 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_decap_8 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_decap_4 FILLER_45_697 ();
 sg13g2_fill_2 FILLER_45_701 ();
 sg13g2_decap_8 FILLER_45_706 ();
 sg13g2_decap_4 FILLER_45_746 ();
 sg13g2_fill_2 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_fill_2 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_fill_2 FILLER_46_574 ();
 sg13g2_fill_1 FILLER_46_593 ();
 sg13g2_decap_8 FILLER_46_639 ();
 sg13g2_decap_8 FILLER_46_646 ();
 sg13g2_decap_4 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_657 ();
 sg13g2_decap_4 FILLER_46_681 ();
 sg13g2_decap_8 FILLER_46_712 ();
 sg13g2_decap_8 FILLER_46_719 ();
 sg13g2_decap_8 FILLER_46_726 ();
 sg13g2_fill_2 FILLER_46_733 ();
 sg13g2_fill_1 FILLER_46_735 ();
 sg13g2_fill_2 FILLER_46_741 ();
 sg13g2_fill_1 FILLER_46_743 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_decap_4 FILLER_46_782 ();
 sg13g2_fill_2 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_fill_1 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_4 FILLER_47_574 ();
 sg13g2_fill_1 FILLER_47_578 ();
 sg13g2_decap_4 FILLER_47_632 ();
 sg13g2_fill_2 FILLER_47_690 ();
 sg13g2_decap_4 FILLER_47_774 ();
 sg13g2_decap_4 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_fill_1 FILLER_48_581 ();
 sg13g2_fill_1 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_fill_2 FILLER_48_658 ();
 sg13g2_fill_1 FILLER_48_660 ();
 sg13g2_fill_1 FILLER_48_667 ();
 sg13g2_fill_2 FILLER_48_753 ();
 sg13g2_fill_1 FILLER_48_789 ();
 sg13g2_fill_2 FILLER_48_820 ();
 sg13g2_fill_1 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_decap_8 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_585 ();
 sg13g2_fill_1 FILLER_49_592 ();
 sg13g2_decap_8 FILLER_49_596 ();
 sg13g2_decap_8 FILLER_49_603 ();
 sg13g2_decap_8 FILLER_49_610 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_4 FILLER_49_627 ();
 sg13g2_decap_8 FILLER_49_636 ();
 sg13g2_decap_8 FILLER_49_643 ();
 sg13g2_decap_8 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_657 ();
 sg13g2_fill_1 FILLER_49_664 ();
 sg13g2_fill_2 FILLER_49_694 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_fill_1 FILLER_49_763 ();
 sg13g2_decap_4 FILLER_49_774 ();
 sg13g2_fill_2 FILLER_49_778 ();
 sg13g2_fill_2 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 assign uio_oe[0] = net;
 assign uio_oe[1] = net228;
 assign uio_oe[2] = net229;
 assign uio_oe[3] = net230;
 assign uio_oe[4] = net231;
 assign uio_oe[5] = net232;
 assign uio_oe[6] = net233;
 assign uio_oe[7] = net234;
endmodule
