** sch_path: /home/cmaier/EDA/PUDDING/xschem/dac2u64out2in.sch
.subckt dac2u64out2in Iout ON[63] ON[62] ON[61] ON[60] ON[59] ON[58] ON[57] ON[56] ON[55] ON[54] ON[53] ON[52] ON[51] ON[50]
+ ON[49] ON[48] ON[47] ON[46] ON[45] ON[44] ON[43] ON[42] ON[41] ON[40] ON[39] ON[38] ON[37] ON[36] ON[35] ON[34] ON[33] ON[32] ON[31]
+ ON[30] ON[29] ON[28] ON[27] ON[26] ON[25] ON[24] ON[23] ON[22] ON[21] ON[20] ON[19] ON[18] ON[17] ON[16] ON[15] ON[14] ON[13] ON[12]
+ ON[11] ON[10] ON[9] ON[8] ON[7] ON[6] ON[5] ON[4] ON[3] ON[2] ON[1] ON[0] ONB[63] ONB[62] ONB[61] ONB[60] ONB[59] ONB[58] ONB[57]
+ ONB[56] ONB[55] ONB[54] ONB[53] ONB[52] ONB[51] ONB[50] ONB[49] ONB[48] ONB[47] ONB[46] ONB[45] ONB[44] ONB[43] ONB[42] ONB[41] ONB[40]
+ ONB[39] ONB[38] ONB[37] ONB[36] ONB[35] ONB[34] ONB[33] ONB[32] ONB[31] ONB[30] ONB[29] ONB[28] ONB[27] ONB[26] ONB[25] ONB[24] ONB[23]
+ ONB[22] ONB[21] ONB[20] ONB[19] ONB[18] ONB[17] ONB[16] ONB[15] ONB[14] ONB[13] ONB[12] ONB[11] ONB[10] ONB[9] ONB[8] ONB[7] ONB[6]
+ ONB[5] ONB[4] ONB[3] ONB[2] ONB[1] ONB[0] VSS VDD Vpcbias EN[1] EN[0] ENB[1] ENB[0]
*.PININFO Iout:O ON[63:0]:I ONB[63:0]:I VSS:B VDD:B Vpcbias:B EN[1:0]:I ENB[1:0]:I
Mcbias Vpcbias Vpcbias Vpbias VDD sg13_lv_pmos w=5.85u l=0.15u ng=1 m=2
xref[1] VDD Vpbias EN[1] ENB[1] Vpbias Vpcbias VSS unitsource2u
xref[0] VDD Vpbias EN[0] ENB[0] Vpbias Vpcbias VSS unitsource2u
xsrc[63] VDD Vpbias ON[63] ONB[63] Iout Vpcbias VSS unitsource2u
xsrc[62] VDD Vpbias ON[62] ONB[62] Iout Vpcbias VSS unitsource2u
xsrc[61] VDD Vpbias ON[61] ONB[61] Iout Vpcbias VSS unitsource2u
xsrc[60] VDD Vpbias ON[60] ONB[60] Iout Vpcbias VSS unitsource2u
xsrc[59] VDD Vpbias ON[59] ONB[59] Iout Vpcbias VSS unitsource2u
xsrc[58] VDD Vpbias ON[58] ONB[58] Iout Vpcbias VSS unitsource2u
xsrc[57] VDD Vpbias ON[57] ONB[57] Iout Vpcbias VSS unitsource2u
xsrc[56] VDD Vpbias ON[56] ONB[56] Iout Vpcbias VSS unitsource2u
xsrc[55] VDD Vpbias ON[55] ONB[55] Iout Vpcbias VSS unitsource2u
xsrc[54] VDD Vpbias ON[54] ONB[54] Iout Vpcbias VSS unitsource2u
xsrc[53] VDD Vpbias ON[53] ONB[53] Iout Vpcbias VSS unitsource2u
xsrc[52] VDD Vpbias ON[52] ONB[52] Iout Vpcbias VSS unitsource2u
xsrc[51] VDD Vpbias ON[51] ONB[51] Iout Vpcbias VSS unitsource2u
xsrc[50] VDD Vpbias ON[50] ONB[50] Iout Vpcbias VSS unitsource2u
xsrc[49] VDD Vpbias ON[49] ONB[49] Iout Vpcbias VSS unitsource2u
xsrc[48] VDD Vpbias ON[48] ONB[48] Iout Vpcbias VSS unitsource2u
xsrc[47] VDD Vpbias ON[47] ONB[47] Iout Vpcbias VSS unitsource2u
xsrc[46] VDD Vpbias ON[46] ONB[46] Iout Vpcbias VSS unitsource2u
xsrc[45] VDD Vpbias ON[45] ONB[45] Iout Vpcbias VSS unitsource2u
xsrc[44] VDD Vpbias ON[44] ONB[44] Iout Vpcbias VSS unitsource2u
xsrc[43] VDD Vpbias ON[43] ONB[43] Iout Vpcbias VSS unitsource2u
xsrc[42] VDD Vpbias ON[42] ONB[42] Iout Vpcbias VSS unitsource2u
xsrc[41] VDD Vpbias ON[41] ONB[41] Iout Vpcbias VSS unitsource2u
xsrc[40] VDD Vpbias ON[40] ONB[40] Iout Vpcbias VSS unitsource2u
xsrc[39] VDD Vpbias ON[39] ONB[39] Iout Vpcbias VSS unitsource2u
xsrc[38] VDD Vpbias ON[38] ONB[38] Iout Vpcbias VSS unitsource2u
xsrc[37] VDD Vpbias ON[37] ONB[37] Iout Vpcbias VSS unitsource2u
xsrc[36] VDD Vpbias ON[36] ONB[36] Iout Vpcbias VSS unitsource2u
xsrc[35] VDD Vpbias ON[35] ONB[35] Iout Vpcbias VSS unitsource2u
xsrc[34] VDD Vpbias ON[34] ONB[34] Iout Vpcbias VSS unitsource2u
xsrc[33] VDD Vpbias ON[33] ONB[33] Iout Vpcbias VSS unitsource2u
xsrc[32] VDD Vpbias ON[32] ONB[32] Iout Vpcbias VSS unitsource2u
xsrc[31] VDD Vpbias ON[31] ONB[31] Iout Vpcbias VSS unitsource2u
xsrc[30] VDD Vpbias ON[30] ONB[30] Iout Vpcbias VSS unitsource2u
xsrc[29] VDD Vpbias ON[29] ONB[29] Iout Vpcbias VSS unitsource2u
xsrc[28] VDD Vpbias ON[28] ONB[28] Iout Vpcbias VSS unitsource2u
xsrc[27] VDD Vpbias ON[27] ONB[27] Iout Vpcbias VSS unitsource2u
xsrc[26] VDD Vpbias ON[26] ONB[26] Iout Vpcbias VSS unitsource2u
xsrc[25] VDD Vpbias ON[25] ONB[25] Iout Vpcbias VSS unitsource2u
xsrc[24] VDD Vpbias ON[24] ONB[24] Iout Vpcbias VSS unitsource2u
xsrc[23] VDD Vpbias ON[23] ONB[23] Iout Vpcbias VSS unitsource2u
xsrc[22] VDD Vpbias ON[22] ONB[22] Iout Vpcbias VSS unitsource2u
xsrc[21] VDD Vpbias ON[21] ONB[21] Iout Vpcbias VSS unitsource2u
xsrc[20] VDD Vpbias ON[20] ONB[20] Iout Vpcbias VSS unitsource2u
xsrc[19] VDD Vpbias ON[19] ONB[19] Iout Vpcbias VSS unitsource2u
xsrc[18] VDD Vpbias ON[18] ONB[18] Iout Vpcbias VSS unitsource2u
xsrc[17] VDD Vpbias ON[17] ONB[17] Iout Vpcbias VSS unitsource2u
xsrc[16] VDD Vpbias ON[16] ONB[16] Iout Vpcbias VSS unitsource2u
xsrc[15] VDD Vpbias ON[15] ONB[15] Iout Vpcbias VSS unitsource2u
xsrc[14] VDD Vpbias ON[14] ONB[14] Iout Vpcbias VSS unitsource2u
xsrc[13] VDD Vpbias ON[13] ONB[13] Iout Vpcbias VSS unitsource2u
xsrc[12] VDD Vpbias ON[12] ONB[12] Iout Vpcbias VSS unitsource2u
xsrc[11] VDD Vpbias ON[11] ONB[11] Iout Vpcbias VSS unitsource2u
xsrc[10] VDD Vpbias ON[10] ONB[10] Iout Vpcbias VSS unitsource2u
xsrc[9] VDD Vpbias ON[9] ONB[9] Iout Vpcbias VSS unitsource2u
xsrc[8] VDD Vpbias ON[8] ONB[8] Iout Vpcbias VSS unitsource2u
xsrc[7] VDD Vpbias ON[7] ONB[7] Iout Vpcbias VSS unitsource2u
xsrc[6] VDD Vpbias ON[6] ONB[6] Iout Vpcbias VSS unitsource2u
xsrc[5] VDD Vpbias ON[5] ONB[5] Iout Vpcbias VSS unitsource2u
xsrc[4] VDD Vpbias ON[4] ONB[4] Iout Vpcbias VSS unitsource2u
xsrc[3] VDD Vpbias ON[3] ONB[3] Iout Vpcbias VSS unitsource2u
xsrc[2] VDD Vpbias ON[2] ONB[2] Iout Vpcbias VSS unitsource2u
xsrc[1] VDD Vpbias ON[1] ONB[1] Iout Vpcbias VSS unitsource2u
xsrc[0] VDD Vpbias ON[0] ONB[0] Iout Vpcbias VSS unitsource2u
**** begin user architecture code

* device parameters
.param l      = 5u
.param w      = 1.45u
.param lc     = 0.6u
.param wc     = 1.2u
.param lb     = 0.15u
.param wb     = 5.85u
.param lplogic= 0.13u
.param wplogic= 0.5u
.param lnlogic= 0.13u
.param wnlogic= 0.15u


**** end user architecture code
.ends

* expanding   symbol:  unitsource2u.sym # of pins=7
** sym_path: /home/cmaier/EDA/PUDDING/xschem/unitsource2u.sym
** sch_path: /home/cmaier/EDA/PUDDING/xschem/unitsource2u.sch
.subckt unitsource2u VDD VbiasP ON ONB Iout VcascP VSS
*.PININFO VSS:B VDD:B VbiasP:B VcascP:B ON:I ONB:I Iout:B
xnonoverlap VDD VSS ON ONB on_n off_n nonoverlap
xsw VDD off_n Vcasc on_n VcascP cascodeswitch_pmos
xsrc VDD VbiasP Vcasc Iout pcsource2u
.ends


* expanding   symbol:  nonoverlap.sym # of pins=6
** sym_path: /home/cmaier/EDA/PUDDING/xschem/nonoverlap.sym
** sch_path: /home/cmaier/EDA/PUDDING/xschem/nonoverlap.sch
.subckt nonoverlap VDD VSS INP INN OUTN OUTP
*.PININFO VSS:B VDD:B INP:I INN:I OUTP:O OUTN:O
M1 OUTN INP VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M2 OUTP INN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M3 OUTN OUTP VSS VSS sg13_lv_nmos w=0.15u l=0.52u ng=1 m=1
M4 OUTP OUTN VSS VSS sg13_lv_nmos w=0.15u l=0.52u ng=1 m=1
.ends


* expanding   symbol:  cascodeswitch_pmos.sym # of pins=5
** sym_path: /home/cmaier/EDA/PUDDING/xschem/cascodeswitch_pmos.sym
** sch_path: /home/cmaier/EDA/PUDDING/xschem/cascodeswitch_pmos.sch
.subckt cascodeswitch_pmos VDD off_n Vcasc on_n Vbpcasc
*.PININFO off_n:I Vbpcasc:I Vcasc:O on_n:I VDD:I
Mpullup Vcasc off_n VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
Mbias Vbpcasc on_n Vcasc VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  pcsource2u.sym # of pins=4
** sym_path: /home/cmaier/EDA/PUDDING/xschem/pcsource2u.sym
** sch_path: /home/cmaier/EDA/PUDDING/xschem/pcsource2u.sch
.subckt pcsource2u VDD VbiasP VcascodeP Iout
*.PININFO VcascodeP:I VbiasP:I Iout:O VDD:I
Msrc drain VbiasP VDD VDD sg13_lv_pmos w=1.45u l=5u ng=1 m=1
Mcasc Iout VcascodeP drain VDD sg13_lv_pmos w=1.2u l=0.6u ng=1 m=1
.ends

