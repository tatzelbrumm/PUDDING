* Extracted by KLayout with SG13G2 LVS runset on : 18/08/2025 23:22

.SUBCKT PCASCSRC16
M$1 \$1 \$2 \$19 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$2 \$19 \$3 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$3 \$1 \$2 \$20 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$4 \$20 \$4 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$5 \$1 \$2 \$22 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$6 \$22 \$5 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$7 \$1 \$2 \$23 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$8 \$23 \$6 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$9 \$1 \$2 \$25 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$10 \$25 \$7 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$11 \$1 \$2 \$26 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$12 \$26 \$8 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$13 \$1 \$2 \$27 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$14 \$27 \$9 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p PS=1.04u
+ PD=1.46u
M$15 \$1 \$2 \$29 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$16 \$29 \$10 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$17 \$1 \$2 \$30 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$18 \$30 \$11 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$19 \$1 \$2 \$32 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$20 \$32 \$12 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$21 \$1 \$2 \$33 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$22 \$33 \$13 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$23 \$1 \$2 \$34 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$24 \$34 \$14 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$25 \$1 \$2 \$31 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$26 \$31 \$15 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$27 \$1 \$2 \$28 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$28 \$28 \$16 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$29 \$1 \$2 \$24 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$30 \$24 \$17 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
M$31 \$1 \$2 \$21 \$1 sg13_lv_pmos L=2u W=0.74u AS=0.2516p AD=0.0956p PS=2.16u
+ PD=1.04u
M$32 \$21 \$18 \$35 \$1 sg13_lv_pmos L=0.3u W=0.3u AS=0.0956p AD=0.129p
+ PS=1.04u PD=1.46u
.ENDS PCASCSRC16
