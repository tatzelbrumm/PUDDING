VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC2U128OUT4IN_PINS
  CLASS BLOCK ;
  FOREIGN DAC2U128OUT4IN_PINS ;
  ORIGIN 1.900 4.910 ;
  SIZE 133.800 BY 26.190 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT -1.900 15.150 131.900 15.820 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 17.200 131.900 17.700 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 0.550 131.900 1.220 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 -1.330 131.900 -0.830 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -1.900 20.780 131.900 21.280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 -4.910 131.900 -4.410 ;
    END
  END VSS
  PIN VbiasP[1]
    PORT
      LAYER Metal1 ;
        RECT -1.000 10.040 131.000 14.970 ;
    END
  END VbiasP[1]
  PIN Iout
    PORT
      LAYER Metal1 ;
        RECT -1.900 7.835 131.900 8.535 ;
    END
  END Iout
  PIN VbiasP[0]
    PORT
      LAYER Metal1 ;
        RECT -1.000 1.400 131.000 6.330 ;
    END
  END VbiasP[0]
  PIN ON[64]
    PORT
      LAYER Metal2 ;
        RECT 128.130 20.990 128.420 21.280 ;
    END
  END ON[64]
  PIN ONB[64]
    PORT
      LAYER Metal2 ;
        RECT 127.580 20.990 127.870 21.280 ;
    END
  END ONB[64]
  PIN ON[65]
    PORT
      LAYER Metal2 ;
        RECT 126.130 20.990 126.420 21.280 ;
    END
  END ON[65]
  PIN ONB[65]
    PORT
      LAYER Metal2 ;
        RECT 125.580 20.990 125.870 21.280 ;
    END
  END ONB[65]
  PIN ON[66]
    PORT
      LAYER Metal2 ;
        RECT 124.130 20.990 124.420 21.280 ;
    END
  END ON[66]
  PIN ONB[66]
    PORT
      LAYER Metal2 ;
        RECT 123.580 20.990 123.870 21.280 ;
    END
  END ONB[66]
  PIN ON[67]
    PORT
      LAYER Metal2 ;
        RECT 122.130 20.990 122.420 21.280 ;
    END
  END ON[67]
  PIN ONB[67]
    PORT
      LAYER Metal2 ;
        RECT 121.580 20.990 121.870 21.280 ;
    END
  END ONB[67]
  PIN ON[68]
    PORT
      LAYER Metal2 ;
        RECT 120.130 20.990 120.420 21.280 ;
    END
  END ON[68]
  PIN ONB[68]
    PORT
      LAYER Metal2 ;
        RECT 119.580 20.990 119.870 21.280 ;
    END
  END ONB[68]
  PIN ON[69]
    PORT
      LAYER Metal2 ;
        RECT 118.130 20.990 118.420 21.280 ;
    END
  END ON[69]
  PIN ONB[69]
    PORT
      LAYER Metal2 ;
        RECT 117.580 20.990 117.870 21.280 ;
    END
  END ONB[69]
  PIN ON[70]
    PORT
      LAYER Metal2 ;
        RECT 116.130 20.990 116.420 21.280 ;
    END
  END ON[70]
  PIN ONB[70]
    PORT
      LAYER Metal2 ;
        RECT 115.580 20.990 115.870 21.280 ;
    END
  END ONB[70]
  PIN ON[71]
    PORT
      LAYER Metal2 ;
        RECT 114.130 20.990 114.420 21.280 ;
    END
  END ON[71]
  PIN ONB[71]
    PORT
      LAYER Metal2 ;
        RECT 113.580 20.990 113.870 21.280 ;
    END
  END ONB[71]
  PIN ON[72]
    PORT
      LAYER Metal2 ;
        RECT 112.130 20.990 112.420 21.280 ;
    END
  END ON[72]
  PIN ONB[72]
    PORT
      LAYER Metal2 ;
        RECT 111.580 20.990 111.870 21.280 ;
    END
  END ONB[72]
  PIN ON[73]
    PORT
      LAYER Metal2 ;
        RECT 110.130 20.990 110.420 21.280 ;
    END
  END ON[73]
  PIN ONB[73]
    PORT
      LAYER Metal2 ;
        RECT 109.580 20.990 109.870 21.280 ;
    END
  END ONB[73]
  PIN ON[74]
    PORT
      LAYER Metal2 ;
        RECT 108.130 20.990 108.420 21.280 ;
    END
  END ON[74]
  PIN ONB[74]
    PORT
      LAYER Metal2 ;
        RECT 107.580 20.990 107.870 21.280 ;
    END
  END ONB[74]
  PIN ON[75]
    PORT
      LAYER Metal2 ;
        RECT 106.130 20.990 106.420 21.280 ;
    END
  END ON[75]
  PIN ONB[75]
    PORT
      LAYER Metal2 ;
        RECT 105.580 20.990 105.870 21.280 ;
    END
  END ONB[75]
  PIN ON[76]
    PORT
      LAYER Metal2 ;
        RECT 104.130 20.990 104.420 21.280 ;
    END
  END ON[76]
  PIN ONB[76]
    PORT
      LAYER Metal2 ;
        RECT 103.580 20.990 103.870 21.280 ;
    END
  END ONB[76]
  PIN ON[77]
    PORT
      LAYER Metal2 ;
        RECT 102.130 20.990 102.420 21.280 ;
    END
  END ON[77]
  PIN ONB[77]
    PORT
      LAYER Metal2 ;
        RECT 101.580 20.990 101.870 21.280 ;
    END
  END ONB[77]
  PIN ON[78]
    PORT
      LAYER Metal2 ;
        RECT 100.130 20.990 100.420 21.280 ;
    END
  END ON[78]
  PIN ONB[78]
    PORT
      LAYER Metal2 ;
        RECT 99.580 20.990 99.870 21.280 ;
    END
  END ONB[78]
  PIN ON[79]
    PORT
      LAYER Metal2 ;
        RECT 98.130 20.990 98.420 21.280 ;
    END
  END ON[79]
  PIN ONB[79]
    PORT
      LAYER Metal2 ;
        RECT 97.580 20.990 97.870 21.280 ;
    END
  END ONB[79]
  PIN ON[80]
    PORT
      LAYER Metal2 ;
        RECT 96.130 20.990 96.420 21.280 ;
    END
  END ON[80]
  PIN ONB[80]
    PORT
      LAYER Metal2 ;
        RECT 95.580 20.990 95.870 21.280 ;
    END
  END ONB[80]
  PIN ON[81]
    PORT
      LAYER Metal2 ;
        RECT 94.130 20.990 94.420 21.280 ;
    END
  END ON[81]
  PIN ONB[81]
    PORT
      LAYER Metal2 ;
        RECT 93.580 20.990 93.870 21.280 ;
    END
  END ONB[81]
  PIN ON[82]
    PORT
      LAYER Metal2 ;
        RECT 92.130 20.990 92.420 21.280 ;
    END
  END ON[82]
  PIN ONB[82]
    PORT
      LAYER Metal2 ;
        RECT 91.580 20.990 91.870 21.280 ;
    END
  END ONB[82]
  PIN ON[83]
    PORT
      LAYER Metal2 ;
        RECT 90.130 20.990 90.420 21.280 ;
    END
  END ON[83]
  PIN ONB[83]
    PORT
      LAYER Metal2 ;
        RECT 89.580 20.990 89.870 21.280 ;
    END
  END ONB[83]
  PIN ON[84]
    PORT
      LAYER Metal2 ;
        RECT 88.130 20.990 88.420 21.280 ;
    END
  END ON[84]
  PIN ONB[84]
    PORT
      LAYER Metal2 ;
        RECT 87.580 20.990 87.870 21.280 ;
    END
  END ONB[84]
  PIN ON[85]
    PORT
      LAYER Metal2 ;
        RECT 86.130 20.990 86.420 21.280 ;
    END
  END ON[85]
  PIN ONB[85]
    PORT
      LAYER Metal2 ;
        RECT 85.580 20.990 85.870 21.280 ;
    END
  END ONB[85]
  PIN ON[86]
    PORT
      LAYER Metal2 ;
        RECT 84.130 20.990 84.420 21.280 ;
    END
  END ON[86]
  PIN ONB[86]
    PORT
      LAYER Metal2 ;
        RECT 83.580 20.990 83.870 21.280 ;
    END
  END ONB[86]
  PIN ON[87]
    PORT
      LAYER Metal2 ;
        RECT 82.130 20.990 82.420 21.280 ;
    END
  END ON[87]
  PIN ONB[87]
    PORT
      LAYER Metal2 ;
        RECT 81.580 20.990 81.870 21.280 ;
    END
  END ONB[87]
  PIN ON[88]
    PORT
      LAYER Metal2 ;
        RECT 80.130 20.990 80.420 21.280 ;
    END
  END ON[88]
  PIN ONB[88]
    PORT
      LAYER Metal2 ;
        RECT 79.580 20.990 79.870 21.280 ;
    END
  END ONB[88]
  PIN ON[89]
    PORT
      LAYER Metal2 ;
        RECT 78.130 20.990 78.420 21.280 ;
    END
  END ON[89]
  PIN ONB[89]
    PORT
      LAYER Metal2 ;
        RECT 77.580 20.990 77.870 21.280 ;
    END
  END ONB[89]
  PIN ON[90]
    PORT
      LAYER Metal2 ;
        RECT 76.130 20.990 76.420 21.280 ;
    END
  END ON[90]
  PIN ONB[90]
    PORT
      LAYER Metal2 ;
        RECT 75.580 20.990 75.870 21.280 ;
    END
  END ONB[90]
  PIN ON[91]
    PORT
      LAYER Metal2 ;
        RECT 74.130 20.990 74.420 21.280 ;
    END
  END ON[91]
  PIN ONB[91]
    PORT
      LAYER Metal2 ;
        RECT 73.580 20.990 73.870 21.280 ;
    END
  END ONB[91]
  PIN ON[92]
    PORT
      LAYER Metal2 ;
        RECT 72.130 20.990 72.420 21.280 ;
    END
  END ON[92]
  PIN ONB[92]
    PORT
      LAYER Metal2 ;
        RECT 71.580 20.990 71.870 21.280 ;
    END
  END ONB[92]
  PIN ON[93]
    PORT
      LAYER Metal2 ;
        RECT 70.130 20.990 70.420 21.280 ;
    END
  END ON[93]
  PIN ONB[93]
    PORT
      LAYER Metal2 ;
        RECT 69.580 20.990 69.870 21.280 ;
    END
  END ONB[93]
  PIN ON[94]
    PORT
      LAYER Metal2 ;
        RECT 68.130 20.990 68.420 21.280 ;
    END
  END ON[94]
  PIN ONB[94]
    PORT
      LAYER Metal2 ;
        RECT 67.580 20.990 67.870 21.280 ;
    END
  END ONB[94]
  PIN ON[95]
    PORT
      LAYER Metal2 ;
        RECT 66.130 20.990 66.420 21.280 ;
    END
  END ON[95]
  PIN ONB[95]
    PORT
      LAYER Metal2 ;
        RECT 65.580 20.990 65.870 21.280 ;
    END
  END ONB[95]
  PIN EN[2]
    PORT
      LAYER Metal2 ;
        RECT 130.130 20.990 130.420 21.280 ;
    END
  END EN[2]
  PIN ENB[2]
    PORT
      LAYER Metal2 ;
        RECT 129.580 20.990 129.870 21.280 ;
    END
  END ENB[2]
  PIN ON[97]
    PORT
      LAYER Metal2 ;
        RECT 62.130 20.990 62.420 21.280 ;
    END
  END ON[97]
  PIN ONB[97]
    PORT
      LAYER Metal2 ;
        RECT 61.580 20.990 61.870 21.280 ;
    END
  END ONB[97]
  PIN ON[98]
    PORT
      LAYER Metal2 ;
        RECT 60.130 20.990 60.420 21.280 ;
    END
  END ON[98]
  PIN ONB[98]
    PORT
      LAYER Metal2 ;
        RECT 59.580 20.990 59.870 21.280 ;
    END
  END ONB[98]
  PIN ON[99]
    PORT
      LAYER Metal2 ;
        RECT 58.130 20.990 58.420 21.280 ;
    END
  END ON[99]
  PIN ONB[99]
    PORT
      LAYER Metal2 ;
        RECT 57.580 20.990 57.870 21.280 ;
    END
  END ONB[99]
  PIN ON[100]
    PORT
      LAYER Metal2 ;
        RECT 56.130 20.990 56.420 21.280 ;
    END
  END ON[100]
  PIN ONB[100]
    PORT
      LAYER Metal2 ;
        RECT 55.580 20.990 55.870 21.280 ;
    END
  END ONB[100]
  PIN ON[101]
    PORT
      LAYER Metal2 ;
        RECT 54.130 20.990 54.420 21.280 ;
    END
  END ON[101]
  PIN ONB[101]
    PORT
      LAYER Metal2 ;
        RECT 53.580 20.990 53.870 21.280 ;
    END
  END ONB[101]
  PIN ON[102]
    PORT
      LAYER Metal2 ;
        RECT 52.130 20.990 52.420 21.280 ;
    END
  END ON[102]
  PIN ONB[102]
    PORT
      LAYER Metal2 ;
        RECT 51.580 20.990 51.870 21.280 ;
    END
  END ONB[102]
  PIN ON[103]
    PORT
      LAYER Metal2 ;
        RECT 50.130 20.990 50.420 21.280 ;
    END
  END ON[103]
  PIN ONB[103]
    PORT
      LAYER Metal2 ;
        RECT 49.580 20.990 49.870 21.280 ;
    END
  END ONB[103]
  PIN ON[104]
    PORT
      LAYER Metal2 ;
        RECT 48.130 20.990 48.420 21.280 ;
    END
  END ON[104]
  PIN ONB[104]
    PORT
      LAYER Metal2 ;
        RECT 47.580 20.990 47.870 21.280 ;
    END
  END ONB[104]
  PIN ON[105]
    PORT
      LAYER Metal2 ;
        RECT 46.130 20.990 46.420 21.280 ;
    END
  END ON[105]
  PIN ONB[105]
    PORT
      LAYER Metal2 ;
        RECT 45.580 20.990 45.870 21.280 ;
    END
  END ONB[105]
  PIN ON[106]
    PORT
      LAYER Metal2 ;
        RECT 44.130 20.990 44.420 21.280 ;
    END
  END ON[106]
  PIN ONB[106]
    PORT
      LAYER Metal2 ;
        RECT 43.580 20.990 43.870 21.280 ;
    END
  END ONB[106]
  PIN ON[107]
    PORT
      LAYER Metal2 ;
        RECT 42.130 20.990 42.420 21.280 ;
    END
  END ON[107]
  PIN ONB[107]
    PORT
      LAYER Metal2 ;
        RECT 41.580 20.990 41.870 21.280 ;
    END
  END ONB[107]
  PIN ON[108]
    PORT
      LAYER Metal2 ;
        RECT 40.130 20.990 40.420 21.280 ;
    END
  END ON[108]
  PIN ONB[108]
    PORT
      LAYER Metal2 ;
        RECT 39.580 20.990 39.870 21.280 ;
    END
  END ONB[108]
  PIN ON[109]
    PORT
      LAYER Metal2 ;
        RECT 38.130 20.990 38.420 21.280 ;
    END
  END ON[109]
  PIN ONB[109]
    PORT
      LAYER Metal2 ;
        RECT 37.580 20.990 37.870 21.280 ;
    END
  END ONB[109]
  PIN ON[110]
    PORT
      LAYER Metal2 ;
        RECT 36.130 20.990 36.420 21.280 ;
    END
  END ON[110]
  PIN ONB[110]
    PORT
      LAYER Metal2 ;
        RECT 35.580 20.990 35.870 21.280 ;
    END
  END ONB[110]
  PIN ON[111]
    PORT
      LAYER Metal2 ;
        RECT 34.130 20.990 34.420 21.280 ;
    END
  END ON[111]
  PIN ONB[111]
    PORT
      LAYER Metal2 ;
        RECT 33.580 20.990 33.870 21.280 ;
    END
  END ONB[111]
  PIN ON[112]
    PORT
      LAYER Metal2 ;
        RECT 32.130 20.990 32.420 21.280 ;
    END
  END ON[112]
  PIN ONB[112]
    PORT
      LAYER Metal2 ;
        RECT 31.580 20.990 31.870 21.280 ;
    END
  END ONB[112]
  PIN ON[113]
    PORT
      LAYER Metal2 ;
        RECT 30.130 20.990 30.420 21.280 ;
    END
  END ON[113]
  PIN ONB[113]
    PORT
      LAYER Metal2 ;
        RECT 29.580 20.990 29.870 21.280 ;
    END
  END ONB[113]
  PIN ON[114]
    PORT
      LAYER Metal2 ;
        RECT 28.130 20.990 28.420 21.280 ;
    END
  END ON[114]
  PIN ONB[114]
    PORT
      LAYER Metal2 ;
        RECT 27.580 20.990 27.870 21.280 ;
    END
  END ONB[114]
  PIN ON[115]
    PORT
      LAYER Metal2 ;
        RECT 26.130 20.990 26.420 21.280 ;
    END
  END ON[115]
  PIN ONB[115]
    PORT
      LAYER Metal2 ;
        RECT 25.580 20.990 25.870 21.280 ;
    END
  END ONB[115]
  PIN ON[116]
    PORT
      LAYER Metal2 ;
        RECT 24.130 20.990 24.420 21.280 ;
    END
  END ON[116]
  PIN ONB[116]
    PORT
      LAYER Metal2 ;
        RECT 23.580 20.990 23.870 21.280 ;
    END
  END ONB[116]
  PIN ON[117]
    PORT
      LAYER Metal2 ;
        RECT 22.130 20.990 22.420 21.280 ;
    END
  END ON[117]
  PIN ONB[117]
    PORT
      LAYER Metal2 ;
        RECT 21.580 20.990 21.870 21.280 ;
    END
  END ONB[117]
  PIN ON[118]
    PORT
      LAYER Metal2 ;
        RECT 20.130 20.990 20.420 21.280 ;
    END
  END ON[118]
  PIN ONB[118]
    PORT
      LAYER Metal2 ;
        RECT 19.580 20.990 19.870 21.280 ;
    END
  END ONB[118]
  PIN ON[119]
    PORT
      LAYER Metal2 ;
        RECT 18.130 20.990 18.420 21.280 ;
    END
  END ON[119]
  PIN ONB[119]
    PORT
      LAYER Metal2 ;
        RECT 17.580 20.990 17.870 21.280 ;
    END
  END ONB[119]
  PIN ON[120]
    PORT
      LAYER Metal2 ;
        RECT 16.130 20.990 16.420 21.280 ;
    END
  END ON[120]
  PIN ONB[120]
    PORT
      LAYER Metal2 ;
        RECT 15.580 20.990 15.870 21.280 ;
    END
  END ONB[120]
  PIN ON[121]
    PORT
      LAYER Metal2 ;
        RECT 14.130 20.990 14.420 21.280 ;
    END
  END ON[121]
  PIN ONB[121]
    PORT
      LAYER Metal2 ;
        RECT 13.580 20.990 13.870 21.280 ;
    END
  END ONB[121]
  PIN ON[122]
    PORT
      LAYER Metal2 ;
        RECT 12.130 20.990 12.420 21.280 ;
    END
  END ON[122]
  PIN ONB[122]
    PORT
      LAYER Metal2 ;
        RECT 11.580 20.990 11.870 21.280 ;
    END
  END ONB[122]
  PIN ON[123]
    PORT
      LAYER Metal2 ;
        RECT 10.130 20.990 10.420 21.280 ;
    END
  END ON[123]
  PIN ONB[123]
    PORT
      LAYER Metal2 ;
        RECT 9.580 20.990 9.870 21.280 ;
    END
  END ONB[123]
  PIN ON[124]
    PORT
      LAYER Metal2 ;
        RECT 8.130 20.990 8.420 21.280 ;
    END
  END ON[124]
  PIN ONB[124]
    PORT
      LAYER Metal2 ;
        RECT 7.580 20.990 7.870 21.280 ;
    END
  END ONB[124]
  PIN ON[125]
    PORT
      LAYER Metal2 ;
        RECT 6.130 20.990 6.420 21.280 ;
    END
  END ON[125]
  PIN ONB[125]
    PORT
      LAYER Metal2 ;
        RECT 5.580 20.990 5.870 21.280 ;
    END
  END ONB[125]
  PIN ON[126]
    PORT
      LAYER Metal2 ;
        RECT 4.130 20.990 4.420 21.280 ;
    END
  END ON[126]
  PIN ONB[126]
    PORT
      LAYER Metal2 ;
        RECT 3.580 20.990 3.870 21.280 ;
    END
  END ONB[126]
  PIN ON[127]
    PORT
      LAYER Metal2 ;
        RECT 2.130 20.990 2.420 21.280 ;
    END
  END ON[127]
  PIN ONB[127]
    PORT
      LAYER Metal2 ;
        RECT 1.580 20.990 1.870 21.280 ;
    END
  END ONB[127]
  PIN ON[96]
    PORT
      LAYER Metal2 ;
        RECT 64.130 20.990 64.420 21.280 ;
    END
  END ON[96]
  PIN ONB[96]
    PORT
      LAYER Metal2 ;
        RECT 63.580 20.990 63.870 21.280 ;
    END
  END ONB[96]
  PIN EN[3]
    PORT
      LAYER Metal2 ;
        RECT 0.130 20.990 0.420 21.280 ;
    END
  END EN[3]
  PIN ENB[3]
    PORT
      LAYER Metal2 ;
        RECT -0.420 20.990 -0.130 21.280 ;
    END
  END ENB[3]
  PIN ON[0]
    PORT
      LAYER Metal2 ;
        RECT 1.580 -4.910 1.870 -4.620 ;
    END
  END ON[0]
  PIN ONB[0]
    PORT
      LAYER Metal2 ;
        RECT 2.130 -4.910 2.420 -4.620 ;
    END
  END ONB[0]
  PIN ON[1]
    PORT
      LAYER Metal2 ;
        RECT 3.580 -4.910 3.870 -4.620 ;
    END
  END ON[1]
  PIN ONB[1]
    PORT
      LAYER Metal2 ;
        RECT 4.130 -4.910 4.420 -4.620 ;
    END
  END ONB[1]
  PIN ON[2]
    PORT
      LAYER Metal2 ;
        RECT 5.580 -4.910 5.870 -4.620 ;
    END
  END ON[2]
  PIN ONB[2]
    PORT
      LAYER Metal2 ;
        RECT 6.130 -4.910 6.420 -4.620 ;
    END
  END ONB[2]
  PIN ON[3]
    PORT
      LAYER Metal2 ;
        RECT 7.580 -4.910 7.870 -4.620 ;
    END
  END ON[3]
  PIN ONB[3]
    PORT
      LAYER Metal2 ;
        RECT 8.130 -4.910 8.420 -4.620 ;
    END
  END ONB[3]
  PIN ON[4]
    PORT
      LAYER Metal2 ;
        RECT 9.580 -4.910 9.870 -4.620 ;
    END
  END ON[4]
  PIN ONB[4]
    PORT
      LAYER Metal2 ;
        RECT 10.130 -4.910 10.420 -4.620 ;
    END
  END ONB[4]
  PIN ON[5]
    PORT
      LAYER Metal2 ;
        RECT 11.580 -4.910 11.870 -4.620 ;
    END
  END ON[5]
  PIN ONB[5]
    PORT
      LAYER Metal2 ;
        RECT 12.130 -4.910 12.420 -4.620 ;
    END
  END ONB[5]
  PIN ON[6]
    PORT
      LAYER Metal2 ;
        RECT 13.580 -4.910 13.870 -4.620 ;
    END
  END ON[6]
  PIN ONB[6]
    PORT
      LAYER Metal2 ;
        RECT 14.130 -4.910 14.420 -4.620 ;
    END
  END ONB[6]
  PIN ON[7]
    PORT
      LAYER Metal2 ;
        RECT 15.580 -4.910 15.870 -4.620 ;
    END
  END ON[7]
  PIN ONB[7]
    PORT
      LAYER Metal2 ;
        RECT 16.130 -4.910 16.420 -4.620 ;
    END
  END ONB[7]
  PIN ON[8]
    PORT
      LAYER Metal2 ;
        RECT 17.580 -4.910 17.870 -4.620 ;
    END
  END ON[8]
  PIN ONB[8]
    PORT
      LAYER Metal2 ;
        RECT 18.130 -4.910 18.420 -4.620 ;
    END
  END ONB[8]
  PIN ON[9]
    PORT
      LAYER Metal2 ;
        RECT 19.580 -4.910 19.870 -4.620 ;
    END
  END ON[9]
  PIN ONB[9]
    PORT
      LAYER Metal2 ;
        RECT 20.130 -4.910 20.420 -4.620 ;
    END
  END ONB[9]
  PIN ON[10]
    PORT
      LAYER Metal2 ;
        RECT 21.580 -4.910 21.870 -4.620 ;
    END
  END ON[10]
  PIN ONB[10]
    PORT
      LAYER Metal2 ;
        RECT 22.130 -4.910 22.420 -4.620 ;
    END
  END ONB[10]
  PIN ON[11]
    PORT
      LAYER Metal2 ;
        RECT 23.580 -4.910 23.870 -4.620 ;
    END
  END ON[11]
  PIN ONB[11]
    PORT
      LAYER Metal2 ;
        RECT 24.130 -4.910 24.420 -4.620 ;
    END
  END ONB[11]
  PIN ON[12]
    PORT
      LAYER Metal2 ;
        RECT 25.580 -4.910 25.870 -4.620 ;
    END
  END ON[12]
  PIN ONB[12]
    PORT
      LAYER Metal2 ;
        RECT 26.130 -4.910 26.420 -4.620 ;
    END
  END ONB[12]
  PIN ON[13]
    PORT
      LAYER Metal2 ;
        RECT 27.580 -4.910 27.870 -4.620 ;
    END
  END ON[13]
  PIN ONB[13]
    PORT
      LAYER Metal2 ;
        RECT 28.130 -4.910 28.420 -4.620 ;
    END
  END ONB[13]
  PIN ON[14]
    PORT
      LAYER Metal2 ;
        RECT 29.580 -4.910 29.870 -4.620 ;
    END
  END ON[14]
  PIN ONB[14]
    PORT
      LAYER Metal2 ;
        RECT 30.130 -4.910 30.420 -4.620 ;
    END
  END ONB[14]
  PIN ON[15]
    PORT
      LAYER Metal2 ;
        RECT 31.580 -4.910 31.870 -4.620 ;
    END
  END ON[15]
  PIN ONB[15]
    PORT
      LAYER Metal2 ;
        RECT 32.130 -4.910 32.420 -4.620 ;
    END
  END ONB[15]
  PIN ON[16]
    PORT
      LAYER Metal2 ;
        RECT 33.580 -4.910 33.870 -4.620 ;
    END
  END ON[16]
  PIN ONB[16]
    PORT
      LAYER Metal2 ;
        RECT 34.130 -4.910 34.420 -4.620 ;
    END
  END ONB[16]
  PIN ON[17]
    PORT
      LAYER Metal2 ;
        RECT 35.580 -4.910 35.870 -4.620 ;
    END
  END ON[17]
  PIN ONB[17]
    PORT
      LAYER Metal2 ;
        RECT 36.130 -4.910 36.420 -4.620 ;
    END
  END ONB[17]
  PIN ON[18]
    PORT
      LAYER Metal2 ;
        RECT 37.580 -4.910 37.870 -4.620 ;
    END
  END ON[18]
  PIN ONB[18]
    PORT
      LAYER Metal2 ;
        RECT 38.130 -4.910 38.420 -4.620 ;
    END
  END ONB[18]
  PIN ON[19]
    PORT
      LAYER Metal2 ;
        RECT 39.580 -4.910 39.870 -4.620 ;
    END
  END ON[19]
  PIN ONB[19]
    PORT
      LAYER Metal2 ;
        RECT 40.130 -4.910 40.420 -4.620 ;
    END
  END ONB[19]
  PIN ON[20]
    PORT
      LAYER Metal2 ;
        RECT 41.580 -4.910 41.870 -4.620 ;
    END
  END ON[20]
  PIN ONB[20]
    PORT
      LAYER Metal2 ;
        RECT 42.130 -4.910 42.420 -4.620 ;
    END
  END ONB[20]
  PIN ON[21]
    PORT
      LAYER Metal2 ;
        RECT 43.580 -4.910 43.870 -4.620 ;
    END
  END ON[21]
  PIN ONB[21]
    PORT
      LAYER Metal2 ;
        RECT 44.130 -4.910 44.420 -4.620 ;
    END
  END ONB[21]
  PIN ON[22]
    PORT
      LAYER Metal2 ;
        RECT 45.580 -4.910 45.870 -4.620 ;
    END
  END ON[22]
  PIN ONB[22]
    PORT
      LAYER Metal2 ;
        RECT 46.130 -4.910 46.420 -4.620 ;
    END
  END ONB[22]
  PIN ON[23]
    PORT
      LAYER Metal2 ;
        RECT 47.580 -4.910 47.870 -4.620 ;
    END
  END ON[23]
  PIN ONB[23]
    PORT
      LAYER Metal2 ;
        RECT 48.130 -4.910 48.420 -4.620 ;
    END
  END ONB[23]
  PIN ON[24]
    PORT
      LAYER Metal2 ;
        RECT 49.580 -4.910 49.870 -4.620 ;
    END
  END ON[24]
  PIN ONB[24]
    PORT
      LAYER Metal2 ;
        RECT 50.130 -4.910 50.420 -4.620 ;
    END
  END ONB[24]
  PIN ON[25]
    PORT
      LAYER Metal2 ;
        RECT 51.580 -4.910 51.870 -4.620 ;
    END
  END ON[25]
  PIN ONB[25]
    PORT
      LAYER Metal2 ;
        RECT 52.130 -4.910 52.420 -4.620 ;
    END
  END ONB[25]
  PIN ON[26]
    PORT
      LAYER Metal2 ;
        RECT 53.580 -4.910 53.870 -4.620 ;
    END
  END ON[26]
  PIN ONB[26]
    PORT
      LAYER Metal2 ;
        RECT 54.130 -4.910 54.420 -4.620 ;
    END
  END ONB[26]
  PIN ON[27]
    PORT
      LAYER Metal2 ;
        RECT 55.580 -4.910 55.870 -4.620 ;
    END
  END ON[27]
  PIN ONB[27]
    PORT
      LAYER Metal2 ;
        RECT 56.130 -4.910 56.420 -4.620 ;
    END
  END ONB[27]
  PIN ON[28]
    PORT
      LAYER Metal2 ;
        RECT 57.580 -4.910 57.870 -4.620 ;
    END
  END ON[28]
  PIN ONB[28]
    PORT
      LAYER Metal2 ;
        RECT 58.130 -4.910 58.420 -4.620 ;
    END
  END ONB[28]
  PIN ON[29]
    PORT
      LAYER Metal2 ;
        RECT 59.580 -4.910 59.870 -4.620 ;
    END
  END ON[29]
  PIN ONB[29]
    PORT
      LAYER Metal2 ;
        RECT 60.130 -4.910 60.420 -4.620 ;
    END
  END ONB[29]
  PIN ON[30]
    PORT
      LAYER Metal2 ;
        RECT 61.580 -4.910 61.870 -4.620 ;
    END
  END ON[30]
  PIN ONB[30]
    PORT
      LAYER Metal2 ;
        RECT 62.130 -4.910 62.420 -4.620 ;
    END
  END ONB[30]
  PIN ON[31]
    PORT
      LAYER Metal2 ;
        RECT 63.580 -4.910 63.870 -4.620 ;
    END
  END ON[31]
  PIN ONB[31]
    PORT
      LAYER Metal2 ;
        RECT 64.130 -4.910 64.420 -4.620 ;
    END
  END ONB[31]
  PIN EN[0]
    PORT
      LAYER Metal2 ;
        RECT -0.420 -4.910 -0.130 -4.620 ;
    END
  END EN[0]
  PIN ENB[0]
    PORT
      LAYER Metal2 ;
        RECT 0.130 -4.910 0.420 -4.620 ;
    END
  END ENB[0]
  PIN ON[33]
    PORT
      LAYER Metal2 ;
        RECT 67.580 -4.910 67.870 -4.620 ;
    END
  END ON[33]
  PIN ONB[33]
    PORT
      LAYER Metal2 ;
        RECT 68.130 -4.910 68.420 -4.620 ;
    END
  END ONB[33]
  PIN ON[34]
    PORT
      LAYER Metal2 ;
        RECT 69.580 -4.910 69.870 -4.620 ;
    END
  END ON[34]
  PIN ONB[34]
    PORT
      LAYER Metal2 ;
        RECT 70.130 -4.910 70.420 -4.620 ;
    END
  END ONB[34]
  PIN ON[35]
    PORT
      LAYER Metal2 ;
        RECT 71.580 -4.910 71.870 -4.620 ;
    END
  END ON[35]
  PIN ONB[35]
    PORT
      LAYER Metal2 ;
        RECT 72.130 -4.910 72.420 -4.620 ;
    END
  END ONB[35]
  PIN ON[36]
    PORT
      LAYER Metal2 ;
        RECT 73.580 -4.910 73.870 -4.620 ;
    END
  END ON[36]
  PIN ONB[36]
    PORT
      LAYER Metal2 ;
        RECT 74.130 -4.910 74.420 -4.620 ;
    END
  END ONB[36]
  PIN ON[37]
    PORT
      LAYER Metal2 ;
        RECT 75.580 -4.910 75.870 -4.620 ;
    END
  END ON[37]
  PIN ONB[37]
    PORT
      LAYER Metal2 ;
        RECT 76.130 -4.910 76.420 -4.620 ;
    END
  END ONB[37]
  PIN ON[38]
    PORT
      LAYER Metal2 ;
        RECT 77.580 -4.910 77.870 -4.620 ;
    END
  END ON[38]
  PIN ONB[38]
    PORT
      LAYER Metal2 ;
        RECT 78.130 -4.910 78.420 -4.620 ;
    END
  END ONB[38]
  PIN ON[39]
    PORT
      LAYER Metal2 ;
        RECT 79.580 -4.910 79.870 -4.620 ;
    END
  END ON[39]
  PIN ONB[39]
    PORT
      LAYER Metal2 ;
        RECT 80.130 -4.910 80.420 -4.620 ;
    END
  END ONB[39]
  PIN ON[40]
    PORT
      LAYER Metal2 ;
        RECT 81.580 -4.910 81.870 -4.620 ;
    END
  END ON[40]
  PIN ONB[40]
    PORT
      LAYER Metal2 ;
        RECT 82.130 -4.910 82.420 -4.620 ;
    END
  END ONB[40]
  PIN ON[41]
    PORT
      LAYER Metal2 ;
        RECT 83.580 -4.910 83.870 -4.620 ;
    END
  END ON[41]
  PIN ONB[41]
    PORT
      LAYER Metal2 ;
        RECT 84.130 -4.910 84.420 -4.620 ;
    END
  END ONB[41]
  PIN ON[42]
    PORT
      LAYER Metal2 ;
        RECT 85.580 -4.910 85.870 -4.620 ;
    END
  END ON[42]
  PIN ONB[42]
    PORT
      LAYER Metal2 ;
        RECT 86.130 -4.910 86.420 -4.620 ;
    END
  END ONB[42]
  PIN ON[43]
    PORT
      LAYER Metal2 ;
        RECT 87.580 -4.910 87.870 -4.620 ;
    END
  END ON[43]
  PIN ONB[43]
    PORT
      LAYER Metal2 ;
        RECT 88.130 -4.910 88.420 -4.620 ;
    END
  END ONB[43]
  PIN ON[44]
    PORT
      LAYER Metal2 ;
        RECT 89.580 -4.910 89.870 -4.620 ;
    END
  END ON[44]
  PIN ONB[44]
    PORT
      LAYER Metal2 ;
        RECT 90.130 -4.910 90.420 -4.620 ;
    END
  END ONB[44]
  PIN ON[45]
    PORT
      LAYER Metal2 ;
        RECT 91.580 -4.910 91.870 -4.620 ;
    END
  END ON[45]
  PIN ONB[45]
    PORT
      LAYER Metal2 ;
        RECT 92.130 -4.910 92.420 -4.620 ;
    END
  END ONB[45]
  PIN ON[46]
    PORT
      LAYER Metal2 ;
        RECT 93.580 -4.910 93.870 -4.620 ;
    END
  END ON[46]
  PIN ONB[46]
    PORT
      LAYER Metal2 ;
        RECT 94.130 -4.910 94.420 -4.620 ;
    END
  END ONB[46]
  PIN ON[47]
    PORT
      LAYER Metal2 ;
        RECT 95.580 -4.910 95.870 -4.620 ;
    END
  END ON[47]
  PIN ONB[47]
    PORT
      LAYER Metal2 ;
        RECT 96.130 -4.910 96.420 -4.620 ;
    END
  END ONB[47]
  PIN ON[48]
    PORT
      LAYER Metal2 ;
        RECT 97.580 -4.910 97.870 -4.620 ;
    END
  END ON[48]
  PIN ONB[48]
    PORT
      LAYER Metal2 ;
        RECT 98.130 -4.910 98.420 -4.620 ;
    END
  END ONB[48]
  PIN ON[49]
    PORT
      LAYER Metal2 ;
        RECT 99.580 -4.910 99.870 -4.620 ;
    END
  END ON[49]
  PIN ONB[49]
    PORT
      LAYER Metal2 ;
        RECT 100.130 -4.910 100.420 -4.620 ;
    END
  END ONB[49]
  PIN ON[50]
    PORT
      LAYER Metal2 ;
        RECT 101.580 -4.910 101.870 -4.620 ;
    END
  END ON[50]
  PIN ONB[50]
    PORT
      LAYER Metal2 ;
        RECT 102.130 -4.910 102.420 -4.620 ;
    END
  END ONB[50]
  PIN ON[51]
    PORT
      LAYER Metal2 ;
        RECT 103.580 -4.910 103.870 -4.620 ;
    END
  END ON[51]
  PIN ONB[51]
    PORT
      LAYER Metal2 ;
        RECT 104.130 -4.910 104.420 -4.620 ;
    END
  END ONB[51]
  PIN ON[52]
    PORT
      LAYER Metal2 ;
        RECT 105.580 -4.910 105.870 -4.620 ;
    END
  END ON[52]
  PIN ONB[52]
    PORT
      LAYER Metal2 ;
        RECT 106.130 -4.910 106.420 -4.620 ;
    END
  END ONB[52]
  PIN ON[53]
    PORT
      LAYER Metal2 ;
        RECT 107.580 -4.910 107.870 -4.620 ;
    END
  END ON[53]
  PIN ONB[53]
    PORT
      LAYER Metal2 ;
        RECT 108.130 -4.910 108.420 -4.620 ;
    END
  END ONB[53]
  PIN ON[54]
    PORT
      LAYER Metal2 ;
        RECT 109.580 -4.910 109.870 -4.620 ;
    END
  END ON[54]
  PIN ONB[54]
    PORT
      LAYER Metal2 ;
        RECT 110.130 -4.910 110.420 -4.620 ;
    END
  END ONB[54]
  PIN ON[55]
    PORT
      LAYER Metal2 ;
        RECT 111.580 -4.910 111.870 -4.620 ;
    END
  END ON[55]
  PIN ONB[55]
    PORT
      LAYER Metal2 ;
        RECT 112.130 -4.910 112.420 -4.620 ;
    END
  END ONB[55]
  PIN ON[56]
    PORT
      LAYER Metal2 ;
        RECT 113.580 -4.910 113.870 -4.620 ;
    END
  END ON[56]
  PIN ONB[56]
    PORT
      LAYER Metal2 ;
        RECT 114.130 -4.910 114.420 -4.620 ;
    END
  END ONB[56]
  PIN ON[57]
    PORT
      LAYER Metal2 ;
        RECT 115.580 -4.910 115.870 -4.620 ;
    END
  END ON[57]
  PIN ONB[57]
    PORT
      LAYER Metal2 ;
        RECT 116.130 -4.910 116.420 -4.620 ;
    END
  END ONB[57]
  PIN ON[58]
    PORT
      LAYER Metal2 ;
        RECT 117.580 -4.910 117.870 -4.620 ;
    END
  END ON[58]
  PIN ONB[58]
    PORT
      LAYER Metal2 ;
        RECT 118.130 -4.910 118.420 -4.620 ;
    END
  END ONB[58]
  PIN ON[59]
    PORT
      LAYER Metal2 ;
        RECT 119.580 -4.910 119.870 -4.620 ;
    END
  END ON[59]
  PIN ONB[59]
    PORT
      LAYER Metal2 ;
        RECT 120.130 -4.910 120.420 -4.620 ;
    END
  END ONB[59]
  PIN ON[60]
    PORT
      LAYER Metal2 ;
        RECT 121.580 -4.910 121.870 -4.620 ;
    END
  END ON[60]
  PIN ONB[60]
    PORT
      LAYER Metal2 ;
        RECT 122.130 -4.910 122.420 -4.620 ;
    END
  END ONB[60]
  PIN ON[61]
    PORT
      LAYER Metal2 ;
        RECT 123.580 -4.910 123.870 -4.620 ;
    END
  END ON[61]
  PIN ONB[61]
    PORT
      LAYER Metal2 ;
        RECT 124.130 -4.910 124.420 -4.620 ;
    END
  END ONB[61]
  PIN ON[62]
    PORT
      LAYER Metal2 ;
        RECT 125.580 -4.910 125.870 -4.620 ;
    END
  END ON[62]
  PIN ONB[62]
    PORT
      LAYER Metal2 ;
        RECT 126.130 -4.910 126.420 -4.620 ;
    END
  END ONB[62]
  PIN ON[63]
    PORT
      LAYER Metal2 ;
        RECT 127.580 -4.910 127.870 -4.620 ;
    END
  END ON[63]
  PIN ONB[63]
    PORT
      LAYER Metal2 ;
        RECT 128.130 -4.910 128.420 -4.620 ;
    END
  END ONB[63]
  PIN ON[32]
    PORT
      LAYER Metal2 ;
        RECT 65.580 -4.910 65.870 -4.620 ;
    END
  END ON[32]
  PIN ONB[32]
    PORT
      LAYER Metal2 ;
        RECT 66.130 -4.910 66.420 -4.620 ;
    END
  END ONB[32]
  PIN EN[1]
    PORT
      LAYER Metal2 ;
        RECT 129.580 -4.910 129.870 -4.620 ;
    END
  END EN[1]
  PIN ENB[1]
    PORT
      LAYER Metal2 ;
        RECT 130.130 -4.910 130.420 -4.620 ;
    END
  END ENB[1]
  PIN VcascP[1]
    PORT
      LAYER Metal3 ;
        RECT -1.900 16.020 131.900 16.720 ;
    END
  END VcascP[1]
  PIN VcascP[0]
    PORT
      LAYER Metal3 ;
        RECT -1.900 -0.350 131.900 0.350 ;
    END
  END VcascP[0]
END DAC2U128OUT4IN_PINS
END LIBRARY

