module heichips25_pudding (clk,
    ena,
    i_in,
    i_out,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 inout i_in;
 inout i_out;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire \bias[0] ;
 wire \bias[1] ;
 wire dacout;
 wire \daisychain[0] ;
 wire \daisychain[100] ;
 wire \daisychain[101] ;
 wire \daisychain[102] ;
 wire \daisychain[103] ;
 wire \daisychain[104] ;
 wire \daisychain[105] ;
 wire \daisychain[106] ;
 wire \daisychain[107] ;
 wire \daisychain[108] ;
 wire \daisychain[109] ;
 wire \daisychain[10] ;
 wire \daisychain[110] ;
 wire \daisychain[111] ;
 wire \daisychain[112] ;
 wire \daisychain[113] ;
 wire \daisychain[114] ;
 wire \daisychain[115] ;
 wire \daisychain[116] ;
 wire \daisychain[117] ;
 wire \daisychain[118] ;
 wire \daisychain[119] ;
 wire \daisychain[11] ;
 wire \daisychain[120] ;
 wire \daisychain[121] ;
 wire \daisychain[122] ;
 wire \daisychain[123] ;
 wire \daisychain[124] ;
 wire \daisychain[125] ;
 wire \daisychain[126] ;
 wire \daisychain[127] ;
 wire \daisychain[12] ;
 wire \daisychain[13] ;
 wire \daisychain[14] ;
 wire \daisychain[15] ;
 wire \daisychain[16] ;
 wire \daisychain[17] ;
 wire \daisychain[18] ;
 wire \daisychain[19] ;
 wire \daisychain[1] ;
 wire \daisychain[20] ;
 wire \daisychain[21] ;
 wire \daisychain[22] ;
 wire \daisychain[23] ;
 wire \daisychain[24] ;
 wire \daisychain[25] ;
 wire \daisychain[26] ;
 wire \daisychain[27] ;
 wire \daisychain[28] ;
 wire \daisychain[29] ;
 wire \daisychain[2] ;
 wire \daisychain[30] ;
 wire \daisychain[31] ;
 wire \daisychain[32] ;
 wire \daisychain[33] ;
 wire \daisychain[34] ;
 wire \daisychain[35] ;
 wire \daisychain[36] ;
 wire \daisychain[37] ;
 wire \daisychain[38] ;
 wire \daisychain[39] ;
 wire \daisychain[3] ;
 wire \daisychain[40] ;
 wire \daisychain[41] ;
 wire \daisychain[42] ;
 wire \daisychain[43] ;
 wire \daisychain[44] ;
 wire \daisychain[45] ;
 wire \daisychain[46] ;
 wire \daisychain[47] ;
 wire \daisychain[48] ;
 wire \daisychain[49] ;
 wire \daisychain[4] ;
 wire \daisychain[50] ;
 wire \daisychain[51] ;
 wire \daisychain[52] ;
 wire \daisychain[53] ;
 wire \daisychain[54] ;
 wire \daisychain[55] ;
 wire \daisychain[56] ;
 wire \daisychain[57] ;
 wire \daisychain[58] ;
 wire \daisychain[59] ;
 wire \daisychain[5] ;
 wire \daisychain[60] ;
 wire \daisychain[61] ;
 wire \daisychain[62] ;
 wire \daisychain[63] ;
 wire \daisychain[64] ;
 wire \daisychain[65] ;
 wire \daisychain[66] ;
 wire \daisychain[67] ;
 wire \daisychain[68] ;
 wire \daisychain[69] ;
 wire \daisychain[6] ;
 wire \daisychain[70] ;
 wire \daisychain[71] ;
 wire \daisychain[72] ;
 wire \daisychain[73] ;
 wire \daisychain[74] ;
 wire \daisychain[75] ;
 wire \daisychain[76] ;
 wire \daisychain[77] ;
 wire \daisychain[78] ;
 wire \daisychain[79] ;
 wire \daisychain[7] ;
 wire \daisychain[80] ;
 wire \daisychain[81] ;
 wire \daisychain[82] ;
 wire \daisychain[83] ;
 wire \daisychain[84] ;
 wire \daisychain[85] ;
 wire \daisychain[86] ;
 wire \daisychain[87] ;
 wire \daisychain[88] ;
 wire \daisychain[89] ;
 wire \daisychain[8] ;
 wire \daisychain[90] ;
 wire \daisychain[91] ;
 wire \daisychain[92] ;
 wire \daisychain[93] ;
 wire \daisychain[94] ;
 wire \daisychain[95] ;
 wire \daisychain[96] ;
 wire \daisychain[97] ;
 wire \daisychain[98] ;
 wire \daisychain[99] ;
 wire \daisychain[9] ;
 wire \digitalen.g[0].u.OUTN ;
 wire \digitalen.g[0].u.OUTP ;
 wire \digitalen.g[1].u.OUTN ;
 wire \digitalen.g[1].u.OUTP ;
 wire \digitalen.g[2].u.OUTN ;
 wire \digitalen.g[2].u.OUTP ;
 wire \digitalen.g[3].u.OUTN ;
 wire \digitalen.g[3].u.OUTP ;
 wire \iref[0] ;
 wire \iref[1] ;
 wire net1;
 wire \state[0] ;
 wire \state[100] ;
 wire \state[101] ;
 wire \state[102] ;
 wire \state[103] ;
 wire \state[104] ;
 wire \state[105] ;
 wire \state[106] ;
 wire \state[107] ;
 wire \state[108] ;
 wire \state[109] ;
 wire \state[10] ;
 wire \state[110] ;
 wire \state[111] ;
 wire \state[112] ;
 wire \state[113] ;
 wire \state[114] ;
 wire \state[115] ;
 wire \state[116] ;
 wire \state[117] ;
 wire \state[118] ;
 wire \state[119] ;
 wire \state[11] ;
 wire \state[120] ;
 wire \state[121] ;
 wire \state[122] ;
 wire \state[123] ;
 wire \state[124] ;
 wire \state[125] ;
 wire \state[126] ;
 wire \state[127] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[16] ;
 wire \state[17] ;
 wire \state[18] ;
 wire \state[19] ;
 wire \state[1] ;
 wire \state[20] ;
 wire \state[21] ;
 wire \state[22] ;
 wire \state[23] ;
 wire \state[24] ;
 wire \state[25] ;
 wire \state[26] ;
 wire \state[27] ;
 wire \state[28] ;
 wire \state[29] ;
 wire \state[2] ;
 wire \state[30] ;
 wire \state[31] ;
 wire \state[32] ;
 wire \state[33] ;
 wire \state[34] ;
 wire \state[35] ;
 wire \state[36] ;
 wire \state[37] ;
 wire \state[38] ;
 wire \state[39] ;
 wire \state[3] ;
 wire \state[40] ;
 wire \state[41] ;
 wire \state[42] ;
 wire \state[43] ;
 wire \state[44] ;
 wire \state[45] ;
 wire \state[46] ;
 wire \state[47] ;
 wire \state[48] ;
 wire \state[49] ;
 wire \state[4] ;
 wire \state[50] ;
 wire \state[51] ;
 wire \state[52] ;
 wire \state[53] ;
 wire \state[54] ;
 wire \state[55] ;
 wire \state[56] ;
 wire \state[57] ;
 wire \state[58] ;
 wire \state[59] ;
 wire \state[5] ;
 wire \state[60] ;
 wire \state[61] ;
 wire \state[62] ;
 wire \state[63] ;
 wire \state[64] ;
 wire \state[65] ;
 wire \state[66] ;
 wire \state[67] ;
 wire \state[68] ;
 wire \state[69] ;
 wire \state[6] ;
 wire \state[70] ;
 wire \state[71] ;
 wire \state[72] ;
 wire \state[73] ;
 wire \state[74] ;
 wire \state[75] ;
 wire \state[76] ;
 wire \state[77] ;
 wire \state[78] ;
 wire \state[79] ;
 wire \state[7] ;
 wire \state[80] ;
 wire \state[81] ;
 wire \state[82] ;
 wire \state[83] ;
 wire \state[84] ;
 wire \state[85] ;
 wire \state[86] ;
 wire \state[87] ;
 wire \state[88] ;
 wire \state[89] ;
 wire \state[8] ;
 wire \state[90] ;
 wire \state[91] ;
 wire \state[92] ;
 wire \state[93] ;
 wire \state[94] ;
 wire \state[95] ;
 wire \state[96] ;
 wire \state[97] ;
 wire \state[98] ;
 wire \state[99] ;
 wire \state[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _1284_ (.Y(_0030_),
    .A(\state[127] ));
 sg13g2_inv_1 _1285_ (.Y(_0846_),
    .A(net158));
 sg13g2_inv_1 _1286_ (.Y(_0029_),
    .A(\state[126] ));
 sg13g2_inv_1 _1287_ (.Y(_0028_),
    .A(\state[125] ));
 sg13g2_inv_1 _1288_ (.Y(_0027_),
    .A(\state[124] ));
 sg13g2_inv_1 _1289_ (.Y(_0026_),
    .A(\state[123] ));
 sg13g2_inv_1 _1290_ (.Y(_0025_),
    .A(\state[122] ));
 sg13g2_inv_1 _1291_ (.Y(_0024_),
    .A(\state[121] ));
 sg13g2_inv_1 _1292_ (.Y(_0023_),
    .A(\state[120] ));
 sg13g2_inv_1 _1293_ (.Y(_0021_),
    .A(\state[119] ));
 sg13g2_inv_1 _1294_ (.Y(_0020_),
    .A(\state[118] ));
 sg13g2_inv_1 _1295_ (.Y(_0019_),
    .A(\state[117] ));
 sg13g2_inv_1 _1296_ (.Y(_0018_),
    .A(\state[116] ));
 sg13g2_inv_1 _1297_ (.Y(_0017_),
    .A(\state[115] ));
 sg13g2_inv_1 _1298_ (.Y(_0016_),
    .A(\state[114] ));
 sg13g2_inv_1 _1299_ (.Y(_0015_),
    .A(\state[113] ));
 sg13g2_inv_1 _1300_ (.Y(_0014_),
    .A(\state[112] ));
 sg13g2_inv_1 _1301_ (.Y(_0013_),
    .A(\state[111] ));
 sg13g2_inv_1 _1302_ (.Y(_0012_),
    .A(\state[110] ));
 sg13g2_inv_1 _1303_ (.Y(_0010_),
    .A(\state[109] ));
 sg13g2_inv_1 _1304_ (.Y(_0009_),
    .A(\state[108] ));
 sg13g2_inv_1 _1305_ (.Y(_0008_),
    .A(\state[107] ));
 sg13g2_inv_1 _1306_ (.Y(_0007_),
    .A(\state[106] ));
 sg13g2_inv_1 _1307_ (.Y(_0006_),
    .A(\state[105] ));
 sg13g2_inv_1 _1308_ (.Y(_0005_),
    .A(\state[104] ));
 sg13g2_inv_1 _1309_ (.Y(_0004_),
    .A(\state[103] ));
 sg13g2_inv_1 _1310_ (.Y(_0003_),
    .A(\state[102] ));
 sg13g2_inv_1 _1311_ (.Y(_0002_),
    .A(\state[101] ));
 sg13g2_inv_1 _1312_ (.Y(_0001_),
    .A(\state[100] ));
 sg13g2_inv_1 _1313_ (.Y(_0126_),
    .A(\state[99] ));
 sg13g2_inv_1 _1314_ (.Y(_0125_),
    .A(\state[98] ));
 sg13g2_inv_1 _1315_ (.Y(_0124_),
    .A(\state[97] ));
 sg13g2_inv_1 _1316_ (.Y(_0123_),
    .A(\state[96] ));
 sg13g2_inv_1 _1317_ (.Y(_0122_),
    .A(\state[95] ));
 sg13g2_inv_1 _1318_ (.Y(_0121_),
    .A(\state[94] ));
 sg13g2_inv_1 _1319_ (.Y(_0120_),
    .A(\state[93] ));
 sg13g2_inv_1 _1320_ (.Y(_0119_),
    .A(\state[92] ));
 sg13g2_inv_1 _1321_ (.Y(_0118_),
    .A(\state[91] ));
 sg13g2_inv_1 _1322_ (.Y(_0117_),
    .A(\state[90] ));
 sg13g2_inv_1 _1323_ (.Y(_0115_),
    .A(\state[89] ));
 sg13g2_inv_1 _1324_ (.Y(_0114_),
    .A(\state[88] ));
 sg13g2_inv_1 _1325_ (.Y(_0113_),
    .A(\state[87] ));
 sg13g2_inv_1 _1326_ (.Y(_0112_),
    .A(\state[86] ));
 sg13g2_inv_1 _1327_ (.Y(_0111_),
    .A(\state[85] ));
 sg13g2_inv_1 _1328_ (.Y(_0110_),
    .A(\state[84] ));
 sg13g2_inv_1 _1329_ (.Y(_0109_),
    .A(\state[83] ));
 sg13g2_inv_1 _1330_ (.Y(_0108_),
    .A(\state[82] ));
 sg13g2_inv_1 _1331_ (.Y(_0107_),
    .A(\state[81] ));
 sg13g2_inv_1 _1332_ (.Y(_0106_),
    .A(\state[80] ));
 sg13g2_inv_1 _1333_ (.Y(_0104_),
    .A(\state[79] ));
 sg13g2_inv_1 _1334_ (.Y(_0103_),
    .A(\state[78] ));
 sg13g2_inv_1 _1335_ (.Y(_0102_),
    .A(\state[77] ));
 sg13g2_inv_1 _1336_ (.Y(_0101_),
    .A(\state[76] ));
 sg13g2_inv_1 _1337_ (.Y(_0100_),
    .A(\state[75] ));
 sg13g2_inv_1 _1338_ (.Y(_0099_),
    .A(\state[74] ));
 sg13g2_inv_1 _1339_ (.Y(_0098_),
    .A(\state[73] ));
 sg13g2_inv_1 _1340_ (.Y(_0097_),
    .A(\state[72] ));
 sg13g2_inv_1 _1341_ (.Y(_0096_),
    .A(\state[71] ));
 sg13g2_inv_1 _1342_ (.Y(_0095_),
    .A(\state[70] ));
 sg13g2_inv_1 _1343_ (.Y(_0093_),
    .A(\state[69] ));
 sg13g2_inv_1 _1344_ (.Y(_0092_),
    .A(\state[68] ));
 sg13g2_inv_1 _1345_ (.Y(_0091_),
    .A(\state[67] ));
 sg13g2_inv_1 _1346_ (.Y(_0090_),
    .A(\state[66] ));
 sg13g2_inv_1 _1347_ (.Y(_0089_),
    .A(\state[65] ));
 sg13g2_inv_1 _1348_ (.Y(_0088_),
    .A(\state[64] ));
 sg13g2_inv_1 _1349_ (.Y(_0087_),
    .A(\state[63] ));
 sg13g2_inv_1 _1350_ (.Y(_0086_),
    .A(\state[62] ));
 sg13g2_inv_1 _1351_ (.Y(_0085_),
    .A(\state[61] ));
 sg13g2_inv_1 _1352_ (.Y(_0084_),
    .A(\state[60] ));
 sg13g2_inv_1 _1353_ (.Y(_0082_),
    .A(\state[59] ));
 sg13g2_inv_1 _1354_ (.Y(_0081_),
    .A(\state[58] ));
 sg13g2_inv_1 _1355_ (.Y(_0080_),
    .A(\state[57] ));
 sg13g2_inv_1 _1356_ (.Y(_0079_),
    .A(\state[56] ));
 sg13g2_inv_1 _1357_ (.Y(_0078_),
    .A(\state[55] ));
 sg13g2_inv_1 _1358_ (.Y(_0077_),
    .A(\state[54] ));
 sg13g2_inv_1 _1359_ (.Y(_0076_),
    .A(\state[53] ));
 sg13g2_inv_1 _1360_ (.Y(_0075_),
    .A(\state[52] ));
 sg13g2_inv_1 _1361_ (.Y(_0074_),
    .A(\state[51] ));
 sg13g2_inv_1 _1362_ (.Y(_0073_),
    .A(\state[50] ));
 sg13g2_inv_1 _1363_ (.Y(_0071_),
    .A(\state[49] ));
 sg13g2_inv_1 _1364_ (.Y(_0070_),
    .A(\state[48] ));
 sg13g2_inv_1 _1365_ (.Y(_0069_),
    .A(\state[47] ));
 sg13g2_inv_1 _1366_ (.Y(_0068_),
    .A(\state[46] ));
 sg13g2_inv_1 _1367_ (.Y(_0067_),
    .A(\state[45] ));
 sg13g2_inv_1 _1368_ (.Y(_0066_),
    .A(\state[44] ));
 sg13g2_inv_1 _1369_ (.Y(_0065_),
    .A(\state[43] ));
 sg13g2_inv_1 _1370_ (.Y(_0064_),
    .A(\state[42] ));
 sg13g2_inv_1 _1371_ (.Y(_0063_),
    .A(\state[41] ));
 sg13g2_inv_1 _1372_ (.Y(_0062_),
    .A(\state[40] ));
 sg13g2_inv_1 _1373_ (.Y(_0060_),
    .A(\state[39] ));
 sg13g2_inv_1 _1374_ (.Y(_0059_),
    .A(\state[38] ));
 sg13g2_inv_1 _1375_ (.Y(_0058_),
    .A(\state[37] ));
 sg13g2_inv_1 _1376_ (.Y(_0057_),
    .A(\state[36] ));
 sg13g2_inv_1 _1377_ (.Y(_0056_),
    .A(\state[35] ));
 sg13g2_inv_1 _1378_ (.Y(_0055_),
    .A(\state[34] ));
 sg13g2_inv_1 _1379_ (.Y(_0054_),
    .A(\state[33] ));
 sg13g2_inv_1 _1380_ (.Y(_0053_),
    .A(\state[32] ));
 sg13g2_inv_1 _1381_ (.Y(_0052_),
    .A(\state[31] ));
 sg13g2_inv_1 _1382_ (.Y(_0051_),
    .A(\state[30] ));
 sg13g2_inv_1 _1383_ (.Y(_0049_),
    .A(\state[29] ));
 sg13g2_inv_1 _1384_ (.Y(_0048_),
    .A(\state[28] ));
 sg13g2_inv_1 _1385_ (.Y(_0047_),
    .A(\state[27] ));
 sg13g2_inv_1 _1386_ (.Y(_0046_),
    .A(\state[26] ));
 sg13g2_inv_1 _1387_ (.Y(_0045_),
    .A(\state[25] ));
 sg13g2_inv_1 _1388_ (.Y(_0044_),
    .A(\state[24] ));
 sg13g2_inv_1 _1389_ (.Y(_0043_),
    .A(\state[23] ));
 sg13g2_inv_1 _1390_ (.Y(_0042_),
    .A(\state[22] ));
 sg13g2_inv_1 _1391_ (.Y(_0041_),
    .A(\state[21] ));
 sg13g2_inv_1 _1392_ (.Y(_0040_),
    .A(\state[20] ));
 sg13g2_inv_1 _1393_ (.Y(_0038_),
    .A(\state[19] ));
 sg13g2_inv_1 _1394_ (.Y(_0037_),
    .A(\state[18] ));
 sg13g2_inv_1 _1395_ (.Y(_0036_),
    .A(\state[17] ));
 sg13g2_inv_1 _1396_ (.Y(_0035_),
    .A(\state[16] ));
 sg13g2_inv_1 _1397_ (.Y(_0034_),
    .A(\state[15] ));
 sg13g2_inv_1 _1398_ (.Y(_0033_),
    .A(\state[14] ));
 sg13g2_inv_1 _1399_ (.Y(_0032_),
    .A(\state[13] ));
 sg13g2_inv_1 _1400_ (.Y(_0031_),
    .A(\state[12] ));
 sg13g2_inv_1 _1401_ (.Y(_0022_),
    .A(\state[11] ));
 sg13g2_inv_1 _1402_ (.Y(_0011_),
    .A(\state[10] ));
 sg13g2_inv_1 _1403_ (.Y(_0127_),
    .A(\state[9] ));
 sg13g2_inv_1 _1404_ (.Y(_0116_),
    .A(\state[8] ));
 sg13g2_inv_1 _1405_ (.Y(_0105_),
    .A(\state[7] ));
 sg13g2_inv_1 _1406_ (.Y(_0094_),
    .A(\state[6] ));
 sg13g2_inv_1 _1407_ (.Y(_0083_),
    .A(\state[5] ));
 sg13g2_inv_1 _1408_ (.Y(_0072_),
    .A(\state[4] ));
 sg13g2_inv_1 _1409_ (.Y(_0061_),
    .A(\state[3] ));
 sg13g2_inv_1 _1410_ (.Y(_0050_),
    .A(\state[2] ));
 sg13g2_inv_1 _1411_ (.Y(_0039_),
    .A(\state[1] ));
 sg13g2_inv_1 _1412_ (.Y(_0000_),
    .A(\state[0] ));
 sg13g2_inv_1 _1413_ (.Y(_0847_),
    .A(net177));
 sg13g2_mux2_1 _1414_ (.A0(\state[0] ),
    .A1(\daisychain[0] ),
    .S(net133),
    .X(_0848_));
 sg13g2_nand2_1 _1415_ (.Y(_0849_),
    .A(net156),
    .B(_0848_));
 sg13g2_nor2_1 _1416_ (.A(net158),
    .B(net3),
    .Y(_0850_));
 sg13g2_or2_1 _1417_ (.X(_0851_),
    .B(net3),
    .A(net158));
 sg13g2_a21oi_1 _1418_ (.A1(net98),
    .A2(net2),
    .Y(_0852_),
    .B1(net48));
 sg13g2_o21ai_1 _1419_ (.B1(net178),
    .Y(_0853_),
    .A1(\daisychain[0] ),
    .A2(net23));
 sg13g2_a21oi_1 _1420_ (.A1(_0849_),
    .A2(_0852_),
    .Y(_0128_),
    .B1(_0853_));
 sg13g2_mux2_1 _1421_ (.A0(\state[1] ),
    .A1(\daisychain[1] ),
    .S(net133),
    .X(_0854_));
 sg13g2_nand2_1 _1422_ (.Y(_0855_),
    .A(net156),
    .B(_0854_));
 sg13g2_a21oi_1 _1423_ (.A1(net94),
    .A2(\daisychain[0] ),
    .Y(_0856_),
    .B1(net45));
 sg13g2_o21ai_1 _1424_ (.B1(net178),
    .Y(_0857_),
    .A1(\daisychain[1] ),
    .A2(net23));
 sg13g2_a21oi_1 _1425_ (.A1(_0855_),
    .A2(_0856_),
    .Y(_0129_),
    .B1(_0857_));
 sg13g2_mux2_1 _1426_ (.A0(\state[2] ),
    .A1(\daisychain[2] ),
    .S(net133),
    .X(_0858_));
 sg13g2_nand2_1 _1427_ (.Y(_0859_),
    .A(net156),
    .B(_0858_));
 sg13g2_a21oi_1 _1428_ (.A1(net94),
    .A2(\daisychain[1] ),
    .Y(_0860_),
    .B1(net45));
 sg13g2_o21ai_1 _1429_ (.B1(net178),
    .Y(_0861_),
    .A1(\daisychain[2] ),
    .A2(net23));
 sg13g2_a21oi_1 _1430_ (.A1(_0859_),
    .A2(_0860_),
    .Y(_0130_),
    .B1(_0861_));
 sg13g2_mux2_1 _1431_ (.A0(\state[3] ),
    .A1(\daisychain[3] ),
    .S(net133),
    .X(_0862_));
 sg13g2_nand2_1 _1432_ (.Y(_0863_),
    .A(net156),
    .B(_0862_));
 sg13g2_a21oi_1 _1433_ (.A1(net95),
    .A2(\daisychain[2] ),
    .Y(_0864_),
    .B1(net45));
 sg13g2_o21ai_1 _1434_ (.B1(net179),
    .Y(_0865_),
    .A1(\daisychain[3] ),
    .A2(net24));
 sg13g2_a21oi_1 _1435_ (.A1(_0863_),
    .A2(_0864_),
    .Y(_0131_),
    .B1(_0865_));
 sg13g2_mux2_1 _1436_ (.A0(\state[4] ),
    .A1(\daisychain[4] ),
    .S(net133),
    .X(_0866_));
 sg13g2_nand2_1 _1437_ (.Y(_0867_),
    .A(net156),
    .B(_0866_));
 sg13g2_a21oi_1 _1438_ (.A1(net95),
    .A2(\daisychain[3] ),
    .Y(_0868_),
    .B1(net46));
 sg13g2_o21ai_1 _1439_ (.B1(net179),
    .Y(_0869_),
    .A1(\daisychain[4] ),
    .A2(net24));
 sg13g2_a21oi_1 _1440_ (.A1(_0867_),
    .A2(_0868_),
    .Y(_0132_),
    .B1(_0869_));
 sg13g2_mux2_1 _1441_ (.A0(\state[5] ),
    .A1(\daisychain[5] ),
    .S(net134),
    .X(_0870_));
 sg13g2_nand2_1 _1442_ (.Y(_0871_),
    .A(net163),
    .B(_0870_));
 sg13g2_a21oi_1 _1443_ (.A1(net95),
    .A2(\daisychain[4] ),
    .Y(_0872_),
    .B1(net46));
 sg13g2_o21ai_1 _1444_ (.B1(net185),
    .Y(_0873_),
    .A1(\daisychain[5] ),
    .A2(net30));
 sg13g2_a21oi_1 _1445_ (.A1(_0871_),
    .A2(_0872_),
    .Y(_0133_),
    .B1(_0873_));
 sg13g2_mux2_1 _1446_ (.A0(\state[6] ),
    .A1(\daisychain[6] ),
    .S(net137),
    .X(_0874_));
 sg13g2_nand2_1 _1447_ (.Y(_0875_),
    .A(net163),
    .B(_0874_));
 sg13g2_a21oi_1 _1448_ (.A1(net107),
    .A2(\daisychain[5] ),
    .Y(_0876_),
    .B1(net53));
 sg13g2_o21ai_1 _1449_ (.B1(net185),
    .Y(_0877_),
    .A1(\daisychain[6] ),
    .A2(net30));
 sg13g2_a21oi_1 _1450_ (.A1(_0875_),
    .A2(_0876_),
    .Y(_0134_),
    .B1(_0877_));
 sg13g2_mux2_1 _1451_ (.A0(\state[7] ),
    .A1(\daisychain[7] ),
    .S(net137),
    .X(_0878_));
 sg13g2_nand2_1 _1452_ (.Y(_0879_),
    .A(net159),
    .B(_0878_));
 sg13g2_a21oi_1 _1453_ (.A1(net101),
    .A2(\daisychain[6] ),
    .Y(_0880_),
    .B1(net49));
 sg13g2_o21ai_1 _1454_ (.B1(net181),
    .Y(_0881_),
    .A1(\daisychain[7] ),
    .A2(net26));
 sg13g2_a21oi_1 _1455_ (.A1(_0879_),
    .A2(_0880_),
    .Y(_0135_),
    .B1(_0881_));
 sg13g2_mux2_1 _1456_ (.A0(\state[8] ),
    .A1(\daisychain[8] ),
    .S(net137),
    .X(_0882_));
 sg13g2_nand2_1 _1457_ (.Y(_0883_),
    .A(net159),
    .B(_0882_));
 sg13g2_a21oi_1 _1458_ (.A1(net101),
    .A2(\daisychain[7] ),
    .Y(_0884_),
    .B1(net49));
 sg13g2_o21ai_1 _1459_ (.B1(net181),
    .Y(_0885_),
    .A1(\daisychain[8] ),
    .A2(net26));
 sg13g2_a21oi_1 _1460_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0136_),
    .B1(_0885_));
 sg13g2_mux2_1 _1461_ (.A0(\state[9] ),
    .A1(\daisychain[9] ),
    .S(net133),
    .X(_0886_));
 sg13g2_nand2_1 _1462_ (.Y(_0887_),
    .A(net159),
    .B(_0886_));
 sg13g2_a21oi_1 _1463_ (.A1(net101),
    .A2(\daisychain[8] ),
    .Y(_0888_),
    .B1(net49));
 sg13g2_o21ai_1 _1464_ (.B1(net181),
    .Y(_0889_),
    .A1(\daisychain[9] ),
    .A2(net26));
 sg13g2_a21oi_1 _1465_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0137_),
    .B1(_0889_));
 sg13g2_mux2_1 _1466_ (.A0(\state[10] ),
    .A1(\daisychain[10] ),
    .S(net133),
    .X(_0890_));
 sg13g2_nand2_1 _1467_ (.Y(_0891_),
    .A(net156),
    .B(_0890_));
 sg13g2_a21oi_1 _1468_ (.A1(net92),
    .A2(\daisychain[9] ),
    .Y(_0892_),
    .B1(net45));
 sg13g2_o21ai_1 _1469_ (.B1(net178),
    .Y(_0893_),
    .A1(\daisychain[10] ),
    .A2(net23));
 sg13g2_a21oi_1 _1470_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0138_),
    .B1(_0893_));
 sg13g2_mux2_1 _1471_ (.A0(\state[11] ),
    .A1(\daisychain[11] ),
    .S(net133),
    .X(_0894_));
 sg13g2_nand2_1 _1472_ (.Y(_0895_),
    .A(net156),
    .B(_0894_));
 sg13g2_a21oi_1 _1473_ (.A1(net92),
    .A2(\daisychain[10] ),
    .Y(_0896_),
    .B1(net45));
 sg13g2_o21ai_1 _1474_ (.B1(net178),
    .Y(_0897_),
    .A1(\daisychain[11] ),
    .A2(net23));
 sg13g2_a21oi_1 _1475_ (.A1(_0895_),
    .A2(_0896_),
    .Y(_0139_),
    .B1(_0897_));
 sg13g2_mux2_1 _1476_ (.A0(\state[12] ),
    .A1(\daisychain[12] ),
    .S(net134),
    .X(_0898_));
 sg13g2_nand2_1 _1477_ (.Y(_0899_),
    .A(net156),
    .B(_0898_));
 sg13g2_a21oi_1 _1478_ (.A1(net92),
    .A2(\daisychain[11] ),
    .Y(_0900_),
    .B1(net45));
 sg13g2_o21ai_1 _1479_ (.B1(net178),
    .Y(_0901_),
    .A1(\daisychain[12] ),
    .A2(net23));
 sg13g2_a21oi_1 _1480_ (.A1(_0899_),
    .A2(_0900_),
    .Y(_0140_),
    .B1(_0901_));
 sg13g2_mux2_1 _1481_ (.A0(\state[13] ),
    .A1(\daisychain[13] ),
    .S(net134),
    .X(_0902_));
 sg13g2_nand2_1 _1482_ (.Y(_0903_),
    .A(net157),
    .B(_0902_));
 sg13g2_a21oi_1 _1483_ (.A1(net92),
    .A2(\daisychain[12] ),
    .Y(_0904_),
    .B1(net45));
 sg13g2_o21ai_1 _1484_ (.B1(net178),
    .Y(_0905_),
    .A1(\daisychain[13] ),
    .A2(net23));
 sg13g2_a21oi_1 _1485_ (.A1(_0903_),
    .A2(_0904_),
    .Y(_0141_),
    .B1(_0905_));
 sg13g2_mux2_1 _1486_ (.A0(\state[14] ),
    .A1(\daisychain[14] ),
    .S(net134),
    .X(_0906_));
 sg13g2_nand2_1 _1487_ (.Y(_0907_),
    .A(net157),
    .B(_0906_));
 sg13g2_a21oi_1 _1488_ (.A1(net93),
    .A2(\daisychain[13] ),
    .Y(_0908_),
    .B1(net45));
 sg13g2_o21ai_1 _1489_ (.B1(net178),
    .Y(_0909_),
    .A1(\daisychain[14] ),
    .A2(net23));
 sg13g2_a21oi_1 _1490_ (.A1(_0907_),
    .A2(_0908_),
    .Y(_0142_),
    .B1(_0909_));
 sg13g2_mux2_1 _1491_ (.A0(\state[15] ),
    .A1(\daisychain[15] ),
    .S(net137),
    .X(_0910_));
 sg13g2_nand2_1 _1492_ (.Y(_0911_),
    .A(net159),
    .B(_0910_));
 sg13g2_a21oi_1 _1493_ (.A1(net94),
    .A2(\daisychain[14] ),
    .Y(_0912_),
    .B1(net47));
 sg13g2_o21ai_1 _1494_ (.B1(net181),
    .Y(_0913_),
    .A1(\daisychain[15] ),
    .A2(net26));
 sg13g2_a21oi_1 _1495_ (.A1(_0911_),
    .A2(_0912_),
    .Y(_0143_),
    .B1(_0913_));
 sg13g2_mux2_1 _1496_ (.A0(\state[16] ),
    .A1(\daisychain[16] ),
    .S(net137),
    .X(_0914_));
 sg13g2_nand2_1 _1497_ (.Y(_0915_),
    .A(net159),
    .B(_0914_));
 sg13g2_a21oi_1 _1498_ (.A1(net99),
    .A2(\daisychain[15] ),
    .Y(_0916_),
    .B1(net49));
 sg13g2_o21ai_1 _1499_ (.B1(net181),
    .Y(_0917_),
    .A1(\daisychain[16] ),
    .A2(net26));
 sg13g2_a21oi_1 _1500_ (.A1(_0915_),
    .A2(_0916_),
    .Y(_0144_),
    .B1(_0917_));
 sg13g2_mux2_1 _1501_ (.A0(\state[17] ),
    .A1(\daisychain[17] ),
    .S(net137),
    .X(_0918_));
 sg13g2_nand2_1 _1502_ (.Y(_0919_),
    .A(net159),
    .B(_0918_));
 sg13g2_a21oi_1 _1503_ (.A1(net99),
    .A2(\daisychain[16] ),
    .Y(_0920_),
    .B1(net49));
 sg13g2_o21ai_1 _1504_ (.B1(net181),
    .Y(_0921_),
    .A1(\daisychain[17] ),
    .A2(net26));
 sg13g2_a21oi_1 _1505_ (.A1(_0919_),
    .A2(_0920_),
    .Y(_0145_),
    .B1(_0921_));
 sg13g2_mux2_1 _1506_ (.A0(\state[18] ),
    .A1(\daisychain[18] ),
    .S(net137),
    .X(_0922_));
 sg13g2_nand2_1 _1507_ (.Y(_0923_),
    .A(net159),
    .B(_0922_));
 sg13g2_a21oi_1 _1508_ (.A1(net99),
    .A2(\daisychain[17] ),
    .Y(_0924_),
    .B1(net49));
 sg13g2_o21ai_1 _1509_ (.B1(net181),
    .Y(_0925_),
    .A1(\daisychain[18] ),
    .A2(net26));
 sg13g2_a21oi_1 _1510_ (.A1(_0923_),
    .A2(_0924_),
    .Y(_0146_),
    .B1(_0925_));
 sg13g2_mux2_1 _1511_ (.A0(\state[19] ),
    .A1(\daisychain[19] ),
    .S(net137),
    .X(_0926_));
 sg13g2_nand2_1 _1512_ (.Y(_0927_),
    .A(net159),
    .B(_0926_));
 sg13g2_a21oi_1 _1513_ (.A1(net99),
    .A2(\daisychain[18] ),
    .Y(_0928_),
    .B1(net49));
 sg13g2_o21ai_1 _1514_ (.B1(net181),
    .Y(_0929_),
    .A1(\daisychain[19] ),
    .A2(net26));
 sg13g2_a21oi_1 _1515_ (.A1(_0927_),
    .A2(_0928_),
    .Y(_0147_),
    .B1(_0929_));
 sg13g2_mux2_1 _1516_ (.A0(\state[20] ),
    .A1(\daisychain[20] ),
    .S(net139),
    .X(_0930_));
 sg13g2_nand2_1 _1517_ (.Y(_0931_),
    .A(net161),
    .B(_0930_));
 sg13g2_a21oi_1 _1518_ (.A1(net99),
    .A2(\daisychain[19] ),
    .Y(_0932_),
    .B1(net50));
 sg13g2_o21ai_1 _1519_ (.B1(net183),
    .Y(_0933_),
    .A1(\daisychain[20] ),
    .A2(net28));
 sg13g2_a21oi_1 _1520_ (.A1(_0931_),
    .A2(_0932_),
    .Y(_0148_),
    .B1(_0933_));
 sg13g2_mux2_1 _1521_ (.A0(\state[21] ),
    .A1(\daisychain[21] ),
    .S(net139),
    .X(_0934_));
 sg13g2_nand2_1 _1522_ (.Y(_0935_),
    .A(net161),
    .B(_0934_));
 sg13g2_a21oi_1 _1523_ (.A1(net104),
    .A2(\daisychain[20] ),
    .Y(_0936_),
    .B1(net50));
 sg13g2_o21ai_1 _1524_ (.B1(net183),
    .Y(_0937_),
    .A1(\daisychain[21] ),
    .A2(net28));
 sg13g2_a21oi_1 _1525_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_0149_),
    .B1(_0937_));
 sg13g2_mux2_1 _1526_ (.A0(\state[22] ),
    .A1(\daisychain[22] ),
    .S(net139),
    .X(_0938_));
 sg13g2_nand2_1 _1527_ (.Y(_0939_),
    .A(net161),
    .B(_0938_));
 sg13g2_a21oi_1 _1528_ (.A1(net104),
    .A2(\daisychain[21] ),
    .Y(_0940_),
    .B1(net50));
 sg13g2_o21ai_1 _1529_ (.B1(net183),
    .Y(_0941_),
    .A1(\daisychain[22] ),
    .A2(net28));
 sg13g2_a21oi_1 _1530_ (.A1(_0939_),
    .A2(_0940_),
    .Y(_0150_),
    .B1(_0941_));
 sg13g2_mux2_1 _1531_ (.A0(\state[23] ),
    .A1(\daisychain[23] ),
    .S(net139),
    .X(_0942_));
 sg13g2_nand2_1 _1532_ (.Y(_0943_),
    .A(net161),
    .B(_0942_));
 sg13g2_a21oi_1 _1533_ (.A1(net104),
    .A2(\daisychain[22] ),
    .Y(_0944_),
    .B1(net50));
 sg13g2_o21ai_1 _1534_ (.B1(net183),
    .Y(_0945_),
    .A1(\daisychain[23] ),
    .A2(net28));
 sg13g2_a21oi_1 _1535_ (.A1(_0943_),
    .A2(_0944_),
    .Y(_0151_),
    .B1(_0945_));
 sg13g2_mux2_1 _1536_ (.A0(\state[24] ),
    .A1(\daisychain[24] ),
    .S(net139),
    .X(_0946_));
 sg13g2_nand2_1 _1537_ (.Y(_0947_),
    .A(net161),
    .B(_0946_));
 sg13g2_a21oi_1 _1538_ (.A1(net104),
    .A2(\daisychain[23] ),
    .Y(_0948_),
    .B1(net50));
 sg13g2_o21ai_1 _1539_ (.B1(net183),
    .Y(_0949_),
    .A1(\daisychain[24] ),
    .A2(net28));
 sg13g2_a21oi_1 _1540_ (.A1(_0947_),
    .A2(_0948_),
    .Y(_0152_),
    .B1(_0949_));
 sg13g2_mux2_1 _1541_ (.A0(\state[25] ),
    .A1(\daisychain[25] ),
    .S(net138),
    .X(_0950_));
 sg13g2_nand2_1 _1542_ (.Y(_0951_),
    .A(net160),
    .B(_0950_));
 sg13g2_a21oi_1 _1543_ (.A1(net100),
    .A2(\daisychain[24] ),
    .Y(_0952_),
    .B1(net50));
 sg13g2_o21ai_1 _1544_ (.B1(net182),
    .Y(_0953_),
    .A1(\daisychain[25] ),
    .A2(net27));
 sg13g2_a21oi_1 _1545_ (.A1(_0951_),
    .A2(_0952_),
    .Y(_0153_),
    .B1(_0953_));
 sg13g2_mux2_1 _1546_ (.A0(\state[26] ),
    .A1(\daisychain[26] ),
    .S(net138),
    .X(_0954_));
 sg13g2_nand2_1 _1547_ (.Y(_0955_),
    .A(net160),
    .B(_0954_));
 sg13g2_a21oi_1 _1548_ (.A1(net100),
    .A2(\daisychain[25] ),
    .Y(_0956_),
    .B1(net49));
 sg13g2_o21ai_1 _1549_ (.B1(net182),
    .Y(_0957_),
    .A1(\daisychain[26] ),
    .A2(net27));
 sg13g2_a21oi_1 _1550_ (.A1(_0955_),
    .A2(_0956_),
    .Y(_0154_),
    .B1(_0957_));
 sg13g2_mux2_1 _1551_ (.A0(\state[27] ),
    .A1(\daisychain[27] ),
    .S(net138),
    .X(_0958_));
 sg13g2_nand2_1 _1552_ (.Y(_0959_),
    .A(net160),
    .B(_0958_));
 sg13g2_a21oi_1 _1553_ (.A1(net100),
    .A2(\daisychain[26] ),
    .Y(_0960_),
    .B1(net52));
 sg13g2_o21ai_1 _1554_ (.B1(net182),
    .Y(_0961_),
    .A1(\daisychain[27] ),
    .A2(net27));
 sg13g2_a21oi_1 _1555_ (.A1(_0959_),
    .A2(_0960_),
    .Y(_0155_),
    .B1(_0961_));
 sg13g2_mux2_1 _1556_ (.A0(\state[28] ),
    .A1(\daisychain[28] ),
    .S(net138),
    .X(_0962_));
 sg13g2_nand2_1 _1557_ (.Y(_0963_),
    .A(net160),
    .B(_0962_));
 sg13g2_a21oi_1 _1558_ (.A1(net100),
    .A2(\daisychain[27] ),
    .Y(_0964_),
    .B1(net52));
 sg13g2_o21ai_1 _1559_ (.B1(net182),
    .Y(_0965_),
    .A1(\daisychain[28] ),
    .A2(net27));
 sg13g2_a21oi_1 _1560_ (.A1(_0963_),
    .A2(_0964_),
    .Y(_0156_),
    .B1(_0965_));
 sg13g2_mux2_1 _1561_ (.A0(\state[29] ),
    .A1(\daisychain[29] ),
    .S(net139),
    .X(_0966_));
 sg13g2_nand2_1 _1562_ (.Y(_0967_),
    .A(net161),
    .B(_0966_));
 sg13g2_a21oi_1 _1563_ (.A1(net100),
    .A2(\daisychain[28] ),
    .Y(_0968_),
    .B1(net51));
 sg13g2_o21ai_1 _1564_ (.B1(net183),
    .Y(_0969_),
    .A1(\daisychain[29] ),
    .A2(net28));
 sg13g2_a21oi_1 _1565_ (.A1(_0967_),
    .A2(_0968_),
    .Y(_0157_),
    .B1(_0969_));
 sg13g2_mux2_1 _1566_ (.A0(\state[30] ),
    .A1(\daisychain[30] ),
    .S(net140),
    .X(_0970_));
 sg13g2_nand2_1 _1567_ (.Y(_0971_),
    .A(net162),
    .B(_0970_));
 sg13g2_a21oi_1 _1568_ (.A1(net105),
    .A2(\daisychain[29] ),
    .Y(_0972_),
    .B1(net51));
 sg13g2_o21ai_1 _1569_ (.B1(net184),
    .Y(_0973_),
    .A1(\daisychain[30] ),
    .A2(net29));
 sg13g2_a21oi_1 _1570_ (.A1(_0971_),
    .A2(_0972_),
    .Y(_0158_),
    .B1(_0973_));
 sg13g2_mux2_1 _1571_ (.A0(\state[31] ),
    .A1(\daisychain[31] ),
    .S(net140),
    .X(_0974_));
 sg13g2_nand2_1 _1572_ (.Y(_0975_),
    .A(net162),
    .B(_0974_));
 sg13g2_a21oi_1 _1573_ (.A1(net105),
    .A2(\daisychain[30] ),
    .Y(_0976_),
    .B1(net51));
 sg13g2_o21ai_1 _1574_ (.B1(net184),
    .Y(_0977_),
    .A1(\daisychain[31] ),
    .A2(net29));
 sg13g2_a21oi_1 _1575_ (.A1(_0975_),
    .A2(_0976_),
    .Y(_0159_),
    .B1(_0977_));
 sg13g2_mux2_1 _1576_ (.A0(\state[32] ),
    .A1(\daisychain[32] ),
    .S(net140),
    .X(_0978_));
 sg13g2_nand2_1 _1577_ (.Y(_0979_),
    .A(net162),
    .B(_0978_));
 sg13g2_a21oi_1 _1578_ (.A1(net105),
    .A2(\daisychain[31] ),
    .Y(_0980_),
    .B1(net51));
 sg13g2_o21ai_1 _1579_ (.B1(net184),
    .Y(_0981_),
    .A1(\daisychain[32] ),
    .A2(net29));
 sg13g2_a21oi_1 _1580_ (.A1(_0979_),
    .A2(_0980_),
    .Y(_0160_),
    .B1(_0981_));
 sg13g2_mux2_1 _1581_ (.A0(\state[33] ),
    .A1(\daisychain[33] ),
    .S(net146),
    .X(_0982_));
 sg13g2_nand2_1 _1582_ (.Y(_0983_),
    .A(net169),
    .B(_0982_));
 sg13g2_a21oi_1 _1583_ (.A1(net105),
    .A2(\daisychain[32] ),
    .Y(_0984_),
    .B1(net51));
 sg13g2_o21ai_1 _1584_ (.B1(net191),
    .Y(_0985_),
    .A1(\daisychain[33] ),
    .A2(net36));
 sg13g2_a21oi_1 _1585_ (.A1(_0983_),
    .A2(_0984_),
    .Y(_0161_),
    .B1(_0985_));
 sg13g2_mux2_1 _1586_ (.A0(\state[34] ),
    .A1(\daisychain[34] ),
    .S(net145),
    .X(_0986_));
 sg13g2_nand2_1 _1587_ (.Y(_0987_),
    .A(net168),
    .B(_0986_));
 sg13g2_a21oi_1 _1588_ (.A1(net103),
    .A2(\daisychain[33] ),
    .Y(_0988_),
    .B1(net57));
 sg13g2_o21ai_1 _1589_ (.B1(net190),
    .Y(_0989_),
    .A1(\daisychain[34] ),
    .A2(net35));
 sg13g2_a21oi_1 _1590_ (.A1(_0987_),
    .A2(_0988_),
    .Y(_0162_),
    .B1(_0989_));
 sg13g2_mux2_1 _1591_ (.A0(\state[35] ),
    .A1(\daisychain[35] ),
    .S(net145),
    .X(_0990_));
 sg13g2_nand2_1 _1592_ (.Y(_0991_),
    .A(net168),
    .B(_0990_));
 sg13g2_a21oi_1 _1593_ (.A1(net103),
    .A2(\daisychain[34] ),
    .Y(_0992_),
    .B1(net57));
 sg13g2_o21ai_1 _1594_ (.B1(net190),
    .Y(_0993_),
    .A1(\daisychain[35] ),
    .A2(net35));
 sg13g2_a21oi_1 _1595_ (.A1(_0991_),
    .A2(_0992_),
    .Y(_0163_),
    .B1(_0993_));
 sg13g2_mux2_1 _1596_ (.A0(\state[36] ),
    .A1(\daisychain[36] ),
    .S(net145),
    .X(_0994_));
 sg13g2_nand2_1 _1597_ (.Y(_0995_),
    .A(net168),
    .B(_0994_));
 sg13g2_a21oi_1 _1598_ (.A1(net116),
    .A2(\daisychain[35] ),
    .Y(_0996_),
    .B1(net57));
 sg13g2_o21ai_1 _1599_ (.B1(net190),
    .Y(_0997_),
    .A1(\daisychain[36] ),
    .A2(net35));
 sg13g2_a21oi_1 _1600_ (.A1(_0995_),
    .A2(_0996_),
    .Y(_0164_),
    .B1(_0997_));
 sg13g2_mux2_1 _1601_ (.A0(\state[37] ),
    .A1(\daisychain[37] ),
    .S(net139),
    .X(_0998_));
 sg13g2_nand2_1 _1602_ (.Y(_0999_),
    .A(net161),
    .B(_0998_));
 sg13g2_a21oi_1 _1603_ (.A1(net103),
    .A2(\daisychain[36] ),
    .Y(_1000_),
    .B1(net57));
 sg13g2_o21ai_1 _1604_ (.B1(net183),
    .Y(_1001_),
    .A1(\daisychain[37] ),
    .A2(net28));
 sg13g2_a21oi_1 _1605_ (.A1(_0999_),
    .A2(_1000_),
    .Y(_0165_),
    .B1(_1001_));
 sg13g2_mux2_1 _1606_ (.A0(\state[38] ),
    .A1(\daisychain[38] ),
    .S(net139),
    .X(_1002_));
 sg13g2_nand2_1 _1607_ (.Y(_1003_),
    .A(net161),
    .B(_1002_));
 sg13g2_a21oi_1 _1608_ (.A1(net103),
    .A2(\daisychain[37] ),
    .Y(_1004_),
    .B1(net50));
 sg13g2_o21ai_1 _1609_ (.B1(net183),
    .Y(_1005_),
    .A1(\daisychain[38] ),
    .A2(net28));
 sg13g2_a21oi_1 _1610_ (.A1(_1003_),
    .A2(_1004_),
    .Y(_0166_),
    .B1(_1005_));
 sg13g2_mux2_1 _1611_ (.A0(\state[39] ),
    .A1(\daisychain[39] ),
    .S(net145),
    .X(_1006_));
 sg13g2_nand2_1 _1612_ (.Y(_1007_),
    .A(net168),
    .B(_1006_));
 sg13g2_a21oi_1 _1613_ (.A1(net103),
    .A2(\daisychain[38] ),
    .Y(_1008_),
    .B1(net50));
 sg13g2_o21ai_1 _1614_ (.B1(net190),
    .Y(_1009_),
    .A1(\daisychain[39] ),
    .A2(net35));
 sg13g2_a21oi_1 _1615_ (.A1(_1007_),
    .A2(_1008_),
    .Y(_0167_),
    .B1(_1009_));
 sg13g2_mux2_1 _1616_ (.A0(\state[40] ),
    .A1(\daisychain[40] ),
    .S(net145),
    .X(_1010_));
 sg13g2_nand2_1 _1617_ (.Y(_1011_),
    .A(net168),
    .B(_1010_));
 sg13g2_a21oi_1 _1618_ (.A1(net116),
    .A2(\daisychain[39] ),
    .Y(_1012_),
    .B1(net57));
 sg13g2_o21ai_1 _1619_ (.B1(net190),
    .Y(_1013_),
    .A1(\daisychain[40] ),
    .A2(net35));
 sg13g2_a21oi_1 _1620_ (.A1(_1011_),
    .A2(_1012_),
    .Y(_0168_),
    .B1(_1013_));
 sg13g2_mux2_1 _1621_ (.A0(\state[41] ),
    .A1(\daisychain[41] ),
    .S(net145),
    .X(_1014_));
 sg13g2_nand2_1 _1622_ (.Y(_1015_),
    .A(net168),
    .B(_1014_));
 sg13g2_a21oi_1 _1623_ (.A1(net115),
    .A2(\daisychain[40] ),
    .Y(_1016_),
    .B1(net57));
 sg13g2_o21ai_1 _1624_ (.B1(net190),
    .Y(_1017_),
    .A1(\daisychain[41] ),
    .A2(net35));
 sg13g2_a21oi_1 _1625_ (.A1(_1015_),
    .A2(_1016_),
    .Y(_0169_),
    .B1(_1017_));
 sg13g2_mux2_1 _1626_ (.A0(\state[42] ),
    .A1(\daisychain[42] ),
    .S(net145),
    .X(_1018_));
 sg13g2_nand2_1 _1627_ (.Y(_1019_),
    .A(net168),
    .B(_1018_));
 sg13g2_a21oi_1 _1628_ (.A1(net115),
    .A2(\daisychain[41] ),
    .Y(_1020_),
    .B1(net57));
 sg13g2_o21ai_1 _1629_ (.B1(net190),
    .Y(_1021_),
    .A1(\daisychain[42] ),
    .A2(net35));
 sg13g2_a21oi_1 _1630_ (.A1(_1019_),
    .A2(_1020_),
    .Y(_0170_),
    .B1(_1021_));
 sg13g2_mux2_1 _1631_ (.A0(\state[43] ),
    .A1(\daisychain[43] ),
    .S(net145),
    .X(_1022_));
 sg13g2_nand2_1 _1632_ (.Y(_1023_),
    .A(net168),
    .B(_1022_));
 sg13g2_a21oi_1 _1633_ (.A1(net115),
    .A2(\daisychain[42] ),
    .Y(_1024_),
    .B1(net57));
 sg13g2_o21ai_1 _1634_ (.B1(net190),
    .Y(_1025_),
    .A1(\daisychain[43] ),
    .A2(net35));
 sg13g2_a21oi_1 _1635_ (.A1(_1023_),
    .A2(_1024_),
    .Y(_0171_),
    .B1(_1025_));
 sg13g2_mux2_1 _1636_ (.A0(\state[44] ),
    .A1(\daisychain[44] ),
    .S(net146),
    .X(_1026_));
 sg13g2_nand2_1 _1637_ (.Y(_1027_),
    .A(net169),
    .B(_1026_));
 sg13g2_a21oi_1 _1638_ (.A1(net115),
    .A2(\daisychain[43] ),
    .Y(_0384_),
    .B1(net58));
 sg13g2_o21ai_1 _1639_ (.B1(net191),
    .Y(_0385_),
    .A1(\daisychain[44] ),
    .A2(net36));
 sg13g2_a21oi_1 _1640_ (.A1(_1027_),
    .A2(_0384_),
    .Y(_0172_),
    .B1(_0385_));
 sg13g2_mux2_1 _1641_ (.A0(\state[45] ),
    .A1(\daisychain[45] ),
    .S(net146),
    .X(_0386_));
 sg13g2_nand2_1 _1642_ (.Y(_0387_),
    .A(net169),
    .B(_0386_));
 sg13g2_a21oi_1 _1643_ (.A1(net116),
    .A2(\daisychain[44] ),
    .Y(_0388_),
    .B1(net58));
 sg13g2_o21ai_1 _1644_ (.B1(net191),
    .Y(_0389_),
    .A1(\daisychain[45] ),
    .A2(net36));
 sg13g2_a21oi_1 _1645_ (.A1(_0387_),
    .A2(_0388_),
    .Y(_0173_),
    .B1(_0389_));
 sg13g2_mux2_1 _1646_ (.A0(\state[46] ),
    .A1(\daisychain[46] ),
    .S(net146),
    .X(_0390_));
 sg13g2_nand2_1 _1647_ (.Y(_0391_),
    .A(net169),
    .B(_0390_));
 sg13g2_a21oi_1 _1648_ (.A1(net117),
    .A2(\daisychain[45] ),
    .Y(_0392_),
    .B1(net58));
 sg13g2_o21ai_1 _1649_ (.B1(net191),
    .Y(_0393_),
    .A1(\daisychain[46] ),
    .A2(net36));
 sg13g2_a21oi_1 _1650_ (.A1(_0391_),
    .A2(_0392_),
    .Y(_0174_),
    .B1(_0393_));
 sg13g2_mux2_1 _1651_ (.A0(\state[47] ),
    .A1(\daisychain[47] ),
    .S(net146),
    .X(_0394_));
 sg13g2_nand2_1 _1652_ (.Y(_0395_),
    .A(net169),
    .B(_0394_));
 sg13g2_a21oi_1 _1653_ (.A1(net117),
    .A2(\daisychain[46] ),
    .Y(_0396_),
    .B1(net58));
 sg13g2_o21ai_1 _1654_ (.B1(net191),
    .Y(_0397_),
    .A1(\daisychain[47] ),
    .A2(net36));
 sg13g2_a21oi_1 _1655_ (.A1(_0395_),
    .A2(_0396_),
    .Y(_0175_),
    .B1(_0397_));
 sg13g2_mux2_1 _1656_ (.A0(\state[48] ),
    .A1(\daisychain[48] ),
    .S(net148),
    .X(_0398_));
 sg13g2_nand2_1 _1657_ (.Y(_0399_),
    .A(net171),
    .B(_0398_));
 sg13g2_a21oi_1 _1658_ (.A1(net117),
    .A2(\daisychain[47] ),
    .Y(_0400_),
    .B1(net60));
 sg13g2_o21ai_1 _1659_ (.B1(net193),
    .Y(_0401_),
    .A1(\daisychain[48] ),
    .A2(net38));
 sg13g2_a21oi_1 _1660_ (.A1(_0399_),
    .A2(_0400_),
    .Y(_0176_),
    .B1(_0401_));
 sg13g2_mux2_1 _1661_ (.A0(\state[49] ),
    .A1(\daisychain[49] ),
    .S(net148),
    .X(_0402_));
 sg13g2_nand2_1 _1662_ (.Y(_0403_),
    .A(net171),
    .B(_0402_));
 sg13g2_a21oi_1 _1663_ (.A1(net122),
    .A2(\daisychain[48] ),
    .Y(_0404_),
    .B1(net60));
 sg13g2_o21ai_1 _1664_ (.B1(net193),
    .Y(_0405_),
    .A1(\daisychain[49] ),
    .A2(net38));
 sg13g2_a21oi_1 _1665_ (.A1(_0403_),
    .A2(_0404_),
    .Y(_0177_),
    .B1(_0405_));
 sg13g2_mux2_1 _1666_ (.A0(\state[50] ),
    .A1(\daisychain[50] ),
    .S(net147),
    .X(_0406_));
 sg13g2_nand2_1 _1667_ (.Y(_0407_),
    .A(net170),
    .B(_0406_));
 sg13g2_a21oi_1 _1668_ (.A1(net122),
    .A2(\daisychain[49] ),
    .Y(_0408_),
    .B1(net60));
 sg13g2_o21ai_1 _1669_ (.B1(net192),
    .Y(_0409_),
    .A1(\daisychain[50] ),
    .A2(net37));
 sg13g2_a21oi_1 _1670_ (.A1(_0407_),
    .A2(_0408_),
    .Y(_0178_),
    .B1(_0409_));
 sg13g2_mux2_1 _1671_ (.A0(\state[51] ),
    .A1(\daisychain[51] ),
    .S(net147),
    .X(_0410_));
 sg13g2_nand2_1 _1672_ (.Y(_0411_),
    .A(net170),
    .B(_0410_));
 sg13g2_a21oi_1 _1673_ (.A1(net118),
    .A2(\daisychain[50] ),
    .Y(_0412_),
    .B1(net59));
 sg13g2_o21ai_1 _1674_ (.B1(net192),
    .Y(_0413_),
    .A1(\daisychain[51] ),
    .A2(net37));
 sg13g2_a21oi_1 _1675_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0179_),
    .B1(_0413_));
 sg13g2_mux2_1 _1676_ (.A0(\state[52] ),
    .A1(\daisychain[52] ),
    .S(net147),
    .X(_0414_));
 sg13g2_nand2_1 _1677_ (.Y(_0415_),
    .A(net170),
    .B(_0414_));
 sg13g2_a21oi_1 _1678_ (.A1(net118),
    .A2(\daisychain[51] ),
    .Y(_0416_),
    .B1(net59));
 sg13g2_o21ai_1 _1679_ (.B1(net192),
    .Y(_0417_),
    .A1(\daisychain[52] ),
    .A2(net37));
 sg13g2_a21oi_1 _1680_ (.A1(_0415_),
    .A2(_0416_),
    .Y(_0180_),
    .B1(_0417_));
 sg13g2_mux2_1 _1681_ (.A0(\state[53] ),
    .A1(\daisychain[53] ),
    .S(net147),
    .X(_0418_));
 sg13g2_nand2_1 _1682_ (.Y(_0419_),
    .A(net170),
    .B(_0418_));
 sg13g2_a21oi_1 _1683_ (.A1(net118),
    .A2(\daisychain[52] ),
    .Y(_0420_),
    .B1(net59));
 sg13g2_o21ai_1 _1684_ (.B1(net192),
    .Y(_0421_),
    .A1(\daisychain[53] ),
    .A2(net37));
 sg13g2_a21oi_1 _1685_ (.A1(_0419_),
    .A2(_0420_),
    .Y(_0181_),
    .B1(_0421_));
 sg13g2_mux2_1 _1686_ (.A0(\state[54] ),
    .A1(\daisychain[54] ),
    .S(net147),
    .X(_0422_));
 sg13g2_nand2_1 _1687_ (.Y(_0423_),
    .A(net170),
    .B(_0422_));
 sg13g2_a21oi_1 _1688_ (.A1(net118),
    .A2(\daisychain[53] ),
    .Y(_0424_),
    .B1(net59));
 sg13g2_o21ai_1 _1689_ (.B1(net192),
    .Y(_0425_),
    .A1(\daisychain[54] ),
    .A2(net37));
 sg13g2_a21oi_1 _1690_ (.A1(_0423_),
    .A2(_0424_),
    .Y(_0182_),
    .B1(_0425_));
 sg13g2_mux2_1 _1691_ (.A0(\state[55] ),
    .A1(\daisychain[55] ),
    .S(net147),
    .X(_0426_));
 sg13g2_nand2_1 _1692_ (.Y(_0427_),
    .A(net170),
    .B(_0426_));
 sg13g2_a21oi_1 _1693_ (.A1(net118),
    .A2(\daisychain[54] ),
    .Y(_0428_),
    .B1(net59));
 sg13g2_o21ai_1 _1694_ (.B1(net192),
    .Y(_0429_),
    .A1(\daisychain[55] ),
    .A2(net37));
 sg13g2_a21oi_1 _1695_ (.A1(_0427_),
    .A2(_0428_),
    .Y(_0183_),
    .B1(_0429_));
 sg13g2_mux2_1 _1696_ (.A0(\state[56] ),
    .A1(\daisychain[56] ),
    .S(net147),
    .X(_0430_));
 sg13g2_nand2_1 _1697_ (.Y(_0431_),
    .A(net170),
    .B(_0430_));
 sg13g2_a21oi_1 _1698_ (.A1(net119),
    .A2(\daisychain[55] ),
    .Y(_0432_),
    .B1(net59));
 sg13g2_o21ai_1 _1699_ (.B1(net192),
    .Y(_0433_),
    .A1(\daisychain[56] ),
    .A2(net37));
 sg13g2_a21oi_1 _1700_ (.A1(_0431_),
    .A2(_0432_),
    .Y(_0184_),
    .B1(_0433_));
 sg13g2_mux2_1 _1701_ (.A0(\state[57] ),
    .A1(\daisychain[57] ),
    .S(net147),
    .X(_0434_));
 sg13g2_nand2_1 _1702_ (.Y(_0435_),
    .A(net170),
    .B(_0434_));
 sg13g2_a21oi_1 _1703_ (.A1(net119),
    .A2(\daisychain[56] ),
    .Y(_0436_),
    .B1(net59));
 sg13g2_o21ai_1 _1704_ (.B1(net192),
    .Y(_0437_),
    .A1(\daisychain[57] ),
    .A2(net37));
 sg13g2_a21oi_1 _1705_ (.A1(_0435_),
    .A2(_0436_),
    .Y(_0185_),
    .B1(_0437_));
 sg13g2_mux2_1 _1706_ (.A0(\state[58] ),
    .A1(\daisychain[58] ),
    .S(net148),
    .X(_0438_));
 sg13g2_nand2_1 _1707_ (.Y(_0439_),
    .A(net171),
    .B(_0438_));
 sg13g2_a21oi_1 _1708_ (.A1(net119),
    .A2(\daisychain[57] ),
    .Y(_0440_),
    .B1(net59));
 sg13g2_o21ai_1 _1709_ (.B1(net193),
    .Y(_0441_),
    .A1(\daisychain[58] ),
    .A2(net38));
 sg13g2_a21oi_1 _1710_ (.A1(_0439_),
    .A2(_0440_),
    .Y(_0186_),
    .B1(_0441_));
 sg13g2_mux2_1 _1711_ (.A0(\state[59] ),
    .A1(\daisychain[59] ),
    .S(net148),
    .X(_0442_));
 sg13g2_nand2_1 _1712_ (.Y(_0443_),
    .A(net171),
    .B(_0442_));
 sg13g2_a21oi_1 _1713_ (.A1(net119),
    .A2(\daisychain[58] ),
    .Y(_0444_),
    .B1(net60));
 sg13g2_o21ai_1 _1714_ (.B1(net193),
    .Y(_0445_),
    .A1(\daisychain[59] ),
    .A2(net38));
 sg13g2_a21oi_1 _1715_ (.A1(_0443_),
    .A2(_0444_),
    .Y(_0187_),
    .B1(_0445_));
 sg13g2_mux2_1 _1716_ (.A0(\state[60] ),
    .A1(\daisychain[60] ),
    .S(net148),
    .X(_0446_));
 sg13g2_nand2_1 _1717_ (.Y(_0447_),
    .A(net171),
    .B(_0446_));
 sg13g2_a21oi_1 _1718_ (.A1(net119),
    .A2(\daisychain[59] ),
    .Y(_0448_),
    .B1(net60));
 sg13g2_o21ai_1 _1719_ (.B1(net193),
    .Y(_0449_),
    .A1(\daisychain[60] ),
    .A2(net38));
 sg13g2_a21oi_1 _1720_ (.A1(_0447_),
    .A2(_0448_),
    .Y(_0188_),
    .B1(_0449_));
 sg13g2_mux2_1 _1721_ (.A0(\state[61] ),
    .A1(\daisychain[61] ),
    .S(net148),
    .X(_0450_));
 sg13g2_nand2_1 _1722_ (.Y(_0451_),
    .A(net171),
    .B(_0450_));
 sg13g2_a21oi_1 _1723_ (.A1(net120),
    .A2(\daisychain[60] ),
    .Y(_0452_),
    .B1(net60));
 sg13g2_o21ai_1 _1724_ (.B1(net193),
    .Y(_0453_),
    .A1(\daisychain[61] ),
    .A2(net38));
 sg13g2_a21oi_1 _1725_ (.A1(_0451_),
    .A2(_0452_),
    .Y(_0189_),
    .B1(_0453_));
 sg13g2_mux2_1 _1726_ (.A0(\state[62] ),
    .A1(\daisychain[62] ),
    .S(net148),
    .X(_0454_));
 sg13g2_nand2_1 _1727_ (.Y(_0455_),
    .A(net171),
    .B(_0454_));
 sg13g2_a21oi_1 _1728_ (.A1(net122),
    .A2(\daisychain[61] ),
    .Y(_0456_),
    .B1(net60));
 sg13g2_o21ai_1 _1729_ (.B1(net193),
    .Y(_0457_),
    .A1(\daisychain[62] ),
    .A2(net38));
 sg13g2_a21oi_1 _1730_ (.A1(_0455_),
    .A2(_0456_),
    .Y(_0190_),
    .B1(_0457_));
 sg13g2_mux2_1 _1731_ (.A0(\state[63] ),
    .A1(\daisychain[63] ),
    .S(net153),
    .X(_0458_));
 sg13g2_nand2_1 _1732_ (.Y(_0459_),
    .A(net176),
    .B(_0458_));
 sg13g2_a21oi_1 _1733_ (.A1(net122),
    .A2(\daisychain[62] ),
    .Y(_0460_),
    .B1(net65));
 sg13g2_o21ai_1 _1734_ (.B1(net198),
    .Y(_0461_),
    .A1(\daisychain[63] ),
    .A2(net43));
 sg13g2_a21oi_1 _1735_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0191_),
    .B1(_0461_));
 sg13g2_mux2_1 _1736_ (.A0(\state[64] ),
    .A1(\daisychain[64] ),
    .S(net152),
    .X(_0462_));
 sg13g2_nand2_1 _1737_ (.Y(_0463_),
    .A(net175),
    .B(_0462_));
 sg13g2_a21oi_1 _1738_ (.A1(net127),
    .A2(\daisychain[63] ),
    .Y(_0464_),
    .B1(net63));
 sg13g2_o21ai_1 _1739_ (.B1(net197),
    .Y(_0465_),
    .A1(\daisychain[64] ),
    .A2(net42));
 sg13g2_a21oi_1 _1740_ (.A1(_0463_),
    .A2(_0464_),
    .Y(_0192_),
    .B1(_0465_));
 sg13g2_mux2_1 _1741_ (.A0(\state[65] ),
    .A1(\daisychain[65] ),
    .S(net152),
    .X(_0466_));
 sg13g2_nand2_1 _1742_ (.Y(_0467_),
    .A(net175),
    .B(_0466_));
 sg13g2_a21oi_1 _1743_ (.A1(net127),
    .A2(\daisychain[64] ),
    .Y(_0468_),
    .B1(net63));
 sg13g2_o21ai_1 _1744_ (.B1(net197),
    .Y(_0469_),
    .A1(\daisychain[65] ),
    .A2(net42));
 sg13g2_a21oi_1 _1745_ (.A1(_0467_),
    .A2(_0468_),
    .Y(_0193_),
    .B1(_0469_));
 sg13g2_mux2_1 _1746_ (.A0(\state[66] ),
    .A1(\daisychain[66] ),
    .S(net151),
    .X(_0470_));
 sg13g2_nand2_1 _1747_ (.Y(_0471_),
    .A(net174),
    .B(_0470_));
 sg13g2_a21oi_1 _1748_ (.A1(net127),
    .A2(\daisychain[65] ),
    .Y(_0472_),
    .B1(net63));
 sg13g2_o21ai_1 _1749_ (.B1(net196),
    .Y(_0473_),
    .A1(\daisychain[66] ),
    .A2(net41));
 sg13g2_a21oi_1 _1750_ (.A1(_0471_),
    .A2(_0472_),
    .Y(_0194_),
    .B1(_0473_));
 sg13g2_mux2_1 _1751_ (.A0(\state[67] ),
    .A1(\daisychain[67] ),
    .S(net151),
    .X(_0474_));
 sg13g2_nand2_1 _1752_ (.Y(_0475_),
    .A(net174),
    .B(_0474_));
 sg13g2_a21oi_1 _1753_ (.A1(net129),
    .A2(\daisychain[66] ),
    .Y(_0476_),
    .B1(net62));
 sg13g2_o21ai_1 _1754_ (.B1(net196),
    .Y(_0477_),
    .A1(\daisychain[67] ),
    .A2(net41));
 sg13g2_a21oi_1 _1755_ (.A1(_0475_),
    .A2(_0476_),
    .Y(_0195_),
    .B1(_0477_));
 sg13g2_mux2_1 _1756_ (.A0(\state[68] ),
    .A1(\daisychain[68] ),
    .S(net151),
    .X(_0478_));
 sg13g2_nand2_1 _1757_ (.Y(_0479_),
    .A(net174),
    .B(_0478_));
 sg13g2_a21oi_1 _1758_ (.A1(net129),
    .A2(\daisychain[67] ),
    .Y(_0480_),
    .B1(net62));
 sg13g2_o21ai_1 _1759_ (.B1(net196),
    .Y(_0481_),
    .A1(\daisychain[68] ),
    .A2(net41));
 sg13g2_a21oi_1 _1760_ (.A1(_0479_),
    .A2(_0480_),
    .Y(_0196_),
    .B1(_0481_));
 sg13g2_mux2_1 _1761_ (.A0(\state[69] ),
    .A1(\daisychain[69] ),
    .S(net152),
    .X(_0482_));
 sg13g2_nand2_1 _1762_ (.Y(_0483_),
    .A(net175),
    .B(_0482_));
 sg13g2_a21oi_1 _1763_ (.A1(net129),
    .A2(\daisychain[68] ),
    .Y(_0484_),
    .B1(net62));
 sg13g2_o21ai_1 _1764_ (.B1(net197),
    .Y(_0485_),
    .A1(\daisychain[69] ),
    .A2(net42));
 sg13g2_a21oi_1 _1765_ (.A1(_0483_),
    .A2(_0484_),
    .Y(_0197_),
    .B1(_0485_));
 sg13g2_mux2_1 _1766_ (.A0(\state[70] ),
    .A1(\daisychain[70] ),
    .S(net152),
    .X(_0486_));
 sg13g2_nand2_1 _1767_ (.Y(_0487_),
    .A(net175),
    .B(_0486_));
 sg13g2_a21oi_1 _1768_ (.A1(net129),
    .A2(\daisychain[69] ),
    .Y(_0488_),
    .B1(net64));
 sg13g2_o21ai_1 _1769_ (.B1(net197),
    .Y(_0489_),
    .A1(\daisychain[70] ),
    .A2(net42));
 sg13g2_a21oi_1 _1770_ (.A1(_0487_),
    .A2(_0488_),
    .Y(_0198_),
    .B1(_0489_));
 sg13g2_mux2_1 _1771_ (.A0(\state[71] ),
    .A1(\daisychain[71] ),
    .S(net152),
    .X(_0490_));
 sg13g2_nand2_1 _1772_ (.Y(_0491_),
    .A(net175),
    .B(_0490_));
 sg13g2_a21oi_1 _1773_ (.A1(net129),
    .A2(\daisychain[70] ),
    .Y(_0492_),
    .B1(net63));
 sg13g2_o21ai_1 _1774_ (.B1(net197),
    .Y(_0493_),
    .A1(\daisychain[71] ),
    .A2(net42));
 sg13g2_a21oi_1 _1775_ (.A1(_0491_),
    .A2(_0492_),
    .Y(_0199_),
    .B1(_0493_));
 sg13g2_mux2_1 _1776_ (.A0(\state[72] ),
    .A1(\daisychain[72] ),
    .S(net151),
    .X(_0494_));
 sg13g2_nand2_1 _1777_ (.Y(_0495_),
    .A(net174),
    .B(_0494_));
 sg13g2_a21oi_1 _1778_ (.A1(net128),
    .A2(\daisychain[71] ),
    .Y(_0496_),
    .B1(net63));
 sg13g2_o21ai_1 _1779_ (.B1(net196),
    .Y(_0497_),
    .A1(\daisychain[72] ),
    .A2(net41));
 sg13g2_a21oi_1 _1780_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0200_),
    .B1(_0497_));
 sg13g2_mux2_1 _1781_ (.A0(\state[73] ),
    .A1(\daisychain[73] ),
    .S(net151),
    .X(_0498_));
 sg13g2_nand2_1 _1782_ (.Y(_0499_),
    .A(net174),
    .B(_0498_));
 sg13g2_a21oi_1 _1783_ (.A1(net128),
    .A2(\daisychain[72] ),
    .Y(_0500_),
    .B1(net62));
 sg13g2_o21ai_1 _1784_ (.B1(net196),
    .Y(_0501_),
    .A1(\daisychain[73] ),
    .A2(net41));
 sg13g2_a21oi_1 _1785_ (.A1(_0499_),
    .A2(_0500_),
    .Y(_0201_),
    .B1(_0501_));
 sg13g2_mux2_1 _1786_ (.A0(\state[74] ),
    .A1(\daisychain[74] ),
    .S(net149),
    .X(_0502_));
 sg13g2_nand2_1 _1787_ (.Y(_0503_),
    .A(net172),
    .B(_0502_));
 sg13g2_a21oi_1 _1788_ (.A1(net125),
    .A2(\daisychain[73] ),
    .Y(_0504_),
    .B1(net62));
 sg13g2_o21ai_1 _1789_ (.B1(net194),
    .Y(_0505_),
    .A1(\daisychain[74] ),
    .A2(net39));
 sg13g2_a21oi_1 _1790_ (.A1(_0503_),
    .A2(_0504_),
    .Y(_0202_),
    .B1(_0505_));
 sg13g2_mux2_1 _1791_ (.A0(\state[75] ),
    .A1(\daisychain[75] ),
    .S(net149),
    .X(_0506_));
 sg13g2_nand2_1 _1792_ (.Y(_0507_),
    .A(net172),
    .B(_0506_));
 sg13g2_a21oi_1 _1793_ (.A1(net125),
    .A2(\daisychain[74] ),
    .Y(_0508_),
    .B1(net61));
 sg13g2_o21ai_1 _1794_ (.B1(net194),
    .Y(_0509_),
    .A1(\daisychain[75] ),
    .A2(net39));
 sg13g2_a21oi_1 _1795_ (.A1(_0507_),
    .A2(_0508_),
    .Y(_0203_),
    .B1(_0509_));
 sg13g2_mux2_1 _1796_ (.A0(\state[76] ),
    .A1(\daisychain[76] ),
    .S(net151),
    .X(_0510_));
 sg13g2_nand2_1 _1797_ (.Y(_0511_),
    .A(net174),
    .B(_0510_));
 sg13g2_a21oi_1 _1798_ (.A1(net128),
    .A2(\daisychain[75] ),
    .Y(_0512_),
    .B1(net62));
 sg13g2_o21ai_1 _1799_ (.B1(net196),
    .Y(_0513_),
    .A1(\daisychain[76] ),
    .A2(net41));
 sg13g2_a21oi_1 _1800_ (.A1(_0511_),
    .A2(_0512_),
    .Y(_0204_),
    .B1(_0513_));
 sg13g2_mux2_1 _1801_ (.A0(\state[77] ),
    .A1(\daisychain[77] ),
    .S(net151),
    .X(_0514_));
 sg13g2_nand2_1 _1802_ (.Y(_0515_),
    .A(net174),
    .B(_0514_));
 sg13g2_a21oi_1 _1803_ (.A1(net128),
    .A2(\daisychain[76] ),
    .Y(_0516_),
    .B1(net62));
 sg13g2_o21ai_1 _1804_ (.B1(net196),
    .Y(_0517_),
    .A1(\daisychain[77] ),
    .A2(net41));
 sg13g2_a21oi_1 _1805_ (.A1(_0515_),
    .A2(_0516_),
    .Y(_0205_),
    .B1(_0517_));
 sg13g2_mux2_1 _1806_ (.A0(\state[78] ),
    .A1(\daisychain[78] ),
    .S(net151),
    .X(_0518_));
 sg13g2_nand2_1 _1807_ (.Y(_0519_),
    .A(net174),
    .B(_0518_));
 sg13g2_a21oi_1 _1808_ (.A1(net128),
    .A2(\daisychain[77] ),
    .Y(_0520_),
    .B1(net62));
 sg13g2_o21ai_1 _1809_ (.B1(net196),
    .Y(_0521_),
    .A1(\daisychain[78] ),
    .A2(net41));
 sg13g2_a21oi_1 _1810_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0206_),
    .B1(_0521_));
 sg13g2_mux2_1 _1811_ (.A0(\state[79] ),
    .A1(\daisychain[79] ),
    .S(net152),
    .X(_0522_));
 sg13g2_nand2_1 _1812_ (.Y(_0523_),
    .A(net175),
    .B(_0522_));
 sg13g2_a21oi_1 _1813_ (.A1(net127),
    .A2(\daisychain[78] ),
    .Y(_0524_),
    .B1(net63));
 sg13g2_o21ai_1 _1814_ (.B1(net197),
    .Y(_0525_),
    .A1(\daisychain[79] ),
    .A2(net42));
 sg13g2_a21oi_1 _1815_ (.A1(_0523_),
    .A2(_0524_),
    .Y(_0207_),
    .B1(_0525_));
 sg13g2_mux2_1 _1816_ (.A0(\state[80] ),
    .A1(\daisychain[80] ),
    .S(net149),
    .X(_0526_));
 sg13g2_nand2_1 _1817_ (.Y(_0527_),
    .A(net173),
    .B(_0526_));
 sg13g2_a21oi_1 _1818_ (.A1(net127),
    .A2(\daisychain[79] ),
    .Y(_0528_),
    .B1(net63));
 sg13g2_o21ai_1 _1819_ (.B1(net197),
    .Y(_0529_),
    .A1(\daisychain[80] ),
    .A2(net42));
 sg13g2_a21oi_1 _1820_ (.A1(_0527_),
    .A2(_0528_),
    .Y(_0208_),
    .B1(_0529_));
 sg13g2_mux2_1 _1821_ (.A0(\state[81] ),
    .A1(\daisychain[81] ),
    .S(net149),
    .X(_0530_));
 sg13g2_nand2_1 _1822_ (.Y(_0531_),
    .A(net173),
    .B(_0530_));
 sg13g2_a21oi_1 _1823_ (.A1(net126),
    .A2(\daisychain[80] ),
    .Y(_0532_),
    .B1(net61));
 sg13g2_o21ai_1 _1824_ (.B1(net195),
    .Y(_0533_),
    .A1(\daisychain[81] ),
    .A2(net40));
 sg13g2_a21oi_1 _1825_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0209_),
    .B1(_0533_));
 sg13g2_mux2_1 _1826_ (.A0(\state[82] ),
    .A1(\daisychain[82] ),
    .S(net149),
    .X(_0534_));
 sg13g2_nand2_1 _1827_ (.Y(_0535_),
    .A(net173),
    .B(_0534_));
 sg13g2_a21oi_1 _1828_ (.A1(net126),
    .A2(\daisychain[81] ),
    .Y(_0536_),
    .B1(net61));
 sg13g2_o21ai_1 _1829_ (.B1(net195),
    .Y(_0537_),
    .A1(\daisychain[82] ),
    .A2(net40));
 sg13g2_a21oi_1 _1830_ (.A1(_0535_),
    .A2(_0536_),
    .Y(_0210_),
    .B1(_0537_));
 sg13g2_mux2_1 _1831_ (.A0(\state[83] ),
    .A1(\daisychain[83] ),
    .S(net149),
    .X(_0538_));
 sg13g2_nand2_1 _1832_ (.Y(_0539_),
    .A(net172),
    .B(_0538_));
 sg13g2_a21oi_1 _1833_ (.A1(net125),
    .A2(\daisychain[82] ),
    .Y(_0540_),
    .B1(net61));
 sg13g2_o21ai_1 _1834_ (.B1(net194),
    .Y(_0541_),
    .A1(\daisychain[83] ),
    .A2(net39));
 sg13g2_a21oi_1 _1835_ (.A1(_0539_),
    .A2(_0540_),
    .Y(_0211_),
    .B1(_0541_));
 sg13g2_mux2_1 _1836_ (.A0(\state[84] ),
    .A1(\daisychain[84] ),
    .S(net150),
    .X(_0542_));
 sg13g2_nand2_1 _1837_ (.Y(_0543_),
    .A(net172),
    .B(_0542_));
 sg13g2_a21oi_1 _1838_ (.A1(net124),
    .A2(\daisychain[83] ),
    .Y(_0544_),
    .B1(net61));
 sg13g2_o21ai_1 _1839_ (.B1(net195),
    .Y(_0545_),
    .A1(\daisychain[84] ),
    .A2(net40));
 sg13g2_a21oi_1 _1840_ (.A1(_0543_),
    .A2(_0544_),
    .Y(_0212_),
    .B1(_0545_));
 sg13g2_mux2_1 _1841_ (.A0(\state[85] ),
    .A1(\daisychain[85] ),
    .S(net150),
    .X(_0546_));
 sg13g2_nand2_1 _1842_ (.Y(_0547_),
    .A(net172),
    .B(_0546_));
 sg13g2_a21oi_1 _1843_ (.A1(net124),
    .A2(\daisychain[84] ),
    .Y(_0548_),
    .B1(net61));
 sg13g2_o21ai_1 _1844_ (.B1(net194),
    .Y(_0549_),
    .A1(\daisychain[85] ),
    .A2(net39));
 sg13g2_a21oi_1 _1845_ (.A1(_0547_),
    .A2(_0548_),
    .Y(_0213_),
    .B1(_0549_));
 sg13g2_mux2_1 _1846_ (.A0(\state[86] ),
    .A1(\daisychain[86] ),
    .S(net150),
    .X(_0550_));
 sg13g2_nand2_1 _1847_ (.Y(_0551_),
    .A(net173),
    .B(_0550_));
 sg13g2_a21oi_1 _1848_ (.A1(net124),
    .A2(\daisychain[85] ),
    .Y(_0552_),
    .B1(net61));
 sg13g2_o21ai_1 _1849_ (.B1(net194),
    .Y(_0553_),
    .A1(\daisychain[86] ),
    .A2(net39));
 sg13g2_a21oi_1 _1850_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0214_),
    .B1(_0553_));
 sg13g2_mux2_1 _1851_ (.A0(\state[87] ),
    .A1(\daisychain[87] ),
    .S(net150),
    .X(_0554_));
 sg13g2_nand2_1 _1852_ (.Y(_0555_),
    .A(net172),
    .B(_0554_));
 sg13g2_a21oi_1 _1853_ (.A1(net124),
    .A2(\daisychain[86] ),
    .Y(_0556_),
    .B1(net64));
 sg13g2_o21ai_1 _1854_ (.B1(net194),
    .Y(_0557_),
    .A1(\daisychain[87] ),
    .A2(net39));
 sg13g2_a21oi_1 _1855_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0215_),
    .B1(_0557_));
 sg13g2_mux2_1 _1856_ (.A0(\state[88] ),
    .A1(\daisychain[88] ),
    .S(net142),
    .X(_0558_));
 sg13g2_nand2_1 _1857_ (.Y(_0559_),
    .A(net165),
    .B(_0558_));
 sg13g2_a21oi_1 _1858_ (.A1(net111),
    .A2(\daisychain[87] ),
    .Y(_0560_),
    .B1(net54));
 sg13g2_o21ai_1 _1859_ (.B1(net187),
    .Y(_0561_),
    .A1(\daisychain[88] ),
    .A2(net32));
 sg13g2_a21oi_1 _1860_ (.A1(_0559_),
    .A2(_0560_),
    .Y(_0216_),
    .B1(_0561_));
 sg13g2_mux2_1 _1861_ (.A0(\state[89] ),
    .A1(\daisychain[89] ),
    .S(net142),
    .X(_0562_));
 sg13g2_nand2_1 _1862_ (.Y(_0563_),
    .A(net172),
    .B(_0562_));
 sg13g2_a21oi_1 _1863_ (.A1(net111),
    .A2(\daisychain[88] ),
    .Y(_0564_),
    .B1(net54));
 sg13g2_o21ai_1 _1864_ (.B1(net194),
    .Y(_0565_),
    .A1(\daisychain[89] ),
    .A2(net39));
 sg13g2_a21oi_1 _1865_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0217_),
    .B1(_0565_));
 sg13g2_mux2_1 _1866_ (.A0(\state[90] ),
    .A1(\daisychain[90] ),
    .S(net150),
    .X(_0566_));
 sg13g2_nand2_1 _1867_ (.Y(_0567_),
    .A(net172),
    .B(_0566_));
 sg13g2_a21oi_1 _1868_ (.A1(net124),
    .A2(\daisychain[89] ),
    .Y(_0568_),
    .B1(net64));
 sg13g2_o21ai_1 _1869_ (.B1(net194),
    .Y(_0569_),
    .A1(\daisychain[90] ),
    .A2(net39));
 sg13g2_a21oi_1 _1870_ (.A1(_0567_),
    .A2(_0568_),
    .Y(_0218_),
    .B1(_0569_));
 sg13g2_mux2_1 _1871_ (.A0(\state[91] ),
    .A1(\daisychain[91] ),
    .S(net149),
    .X(_0570_));
 sg13g2_nand2_1 _1872_ (.Y(_0571_),
    .A(net173),
    .B(_0570_));
 sg13g2_a21oi_1 _1873_ (.A1(net124),
    .A2(\daisychain[90] ),
    .Y(_0572_),
    .B1(net64));
 sg13g2_o21ai_1 _1874_ (.B1(net195),
    .Y(_0573_),
    .A1(\daisychain[91] ),
    .A2(net40));
 sg13g2_a21oi_1 _1875_ (.A1(_0571_),
    .A2(_0572_),
    .Y(_0219_),
    .B1(_0573_));
 sg13g2_mux2_1 _1876_ (.A0(\state[92] ),
    .A1(\daisychain[92] ),
    .S(net149),
    .X(_0574_));
 sg13g2_nand2_1 _1877_ (.Y(_0575_),
    .A(net173),
    .B(_0574_));
 sg13g2_a21oi_1 _1878_ (.A1(net110),
    .A2(\daisychain[91] ),
    .Y(_0576_),
    .B1(net61));
 sg13g2_o21ai_1 _1879_ (.B1(net195),
    .Y(_0577_),
    .A1(\daisychain[92] ),
    .A2(net40));
 sg13g2_a21oi_1 _1880_ (.A1(_0575_),
    .A2(_0576_),
    .Y(_0220_),
    .B1(_0577_));
 sg13g2_mux2_1 _1881_ (.A0(\state[93] ),
    .A1(\daisychain[93] ),
    .S(net142),
    .X(_0578_));
 sg13g2_nand2_1 _1882_ (.Y(_0579_),
    .A(net165),
    .B(_0578_));
 sg13g2_a21oi_1 _1883_ (.A1(net113),
    .A2(\daisychain[92] ),
    .Y(_0580_),
    .B1(net55));
 sg13g2_o21ai_1 _1884_ (.B1(net187),
    .Y(_0581_),
    .A1(\daisychain[93] ),
    .A2(net32));
 sg13g2_a21oi_1 _1885_ (.A1(_0579_),
    .A2(_0580_),
    .Y(_0221_),
    .B1(_0581_));
 sg13g2_mux2_1 _1886_ (.A0(\state[94] ),
    .A1(\daisychain[94] ),
    .S(net142),
    .X(_0582_));
 sg13g2_nand2_1 _1887_ (.Y(_0583_),
    .A(net165),
    .B(_0582_));
 sg13g2_a21oi_1 _1888_ (.A1(net113),
    .A2(\daisychain[93] ),
    .Y(_0584_),
    .B1(net55));
 sg13g2_o21ai_1 _1889_ (.B1(net187),
    .Y(_0585_),
    .A1(\daisychain[94] ),
    .A2(net32));
 sg13g2_a21oi_1 _1890_ (.A1(_0583_),
    .A2(_0584_),
    .Y(_0222_),
    .B1(_0585_));
 sg13g2_mux2_1 _1891_ (.A0(\state[95] ),
    .A1(\daisychain[95] ),
    .S(net143),
    .X(_0586_));
 sg13g2_nand2_1 _1892_ (.Y(_0587_),
    .A(net165),
    .B(_0586_));
 sg13g2_a21oi_1 _1893_ (.A1(net111),
    .A2(\daisychain[94] ),
    .Y(_0588_),
    .B1(net54));
 sg13g2_o21ai_1 _1894_ (.B1(net187),
    .Y(_0589_),
    .A1(\daisychain[95] ),
    .A2(net32));
 sg13g2_a21oi_1 _1895_ (.A1(_0587_),
    .A2(_0588_),
    .Y(_0223_),
    .B1(_0589_));
 sg13g2_mux2_1 _1896_ (.A0(\state[96] ),
    .A1(\daisychain[96] ),
    .S(net143),
    .X(_0590_));
 sg13g2_nand2_1 _1897_ (.Y(_0591_),
    .A(net166),
    .B(_0590_));
 sg13g2_a21oi_1 _1898_ (.A1(net111),
    .A2(\daisychain[95] ),
    .Y(_0592_),
    .B1(net55));
 sg13g2_o21ai_1 _1899_ (.B1(net188),
    .Y(_0593_),
    .A1(\daisychain[96] ),
    .A2(net33));
 sg13g2_a21oi_1 _1900_ (.A1(_0591_),
    .A2(_0592_),
    .Y(_0224_),
    .B1(_0593_));
 sg13g2_mux2_1 _1901_ (.A0(\state[97] ),
    .A1(\daisychain[97] ),
    .S(net143),
    .X(_0594_));
 sg13g2_nand2_1 _1902_ (.Y(_0595_),
    .A(net166),
    .B(_0594_));
 sg13g2_a21oi_1 _1903_ (.A1(net112),
    .A2(\daisychain[96] ),
    .Y(_0596_),
    .B1(net54));
 sg13g2_o21ai_1 _1904_ (.B1(net188),
    .Y(_0597_),
    .A1(\daisychain[97] ),
    .A2(net33));
 sg13g2_a21oi_1 _1905_ (.A1(_0595_),
    .A2(_0596_),
    .Y(_0225_),
    .B1(_0597_));
 sg13g2_mux2_1 _1906_ (.A0(\state[98] ),
    .A1(\daisychain[98] ),
    .S(net141),
    .X(_0598_));
 sg13g2_nand2_1 _1907_ (.Y(_0599_),
    .A(net164),
    .B(_0598_));
 sg13g2_a21oi_1 _1908_ (.A1(net109),
    .A2(\daisychain[97] ),
    .Y(_0600_),
    .B1(net54));
 sg13g2_o21ai_1 _1909_ (.B1(net186),
    .Y(_0601_),
    .A1(\daisychain[98] ),
    .A2(net31));
 sg13g2_a21oi_1 _1910_ (.A1(_0599_),
    .A2(_0600_),
    .Y(_0226_),
    .B1(_0601_));
 sg13g2_mux2_1 _1911_ (.A0(\state[99] ),
    .A1(\daisychain[99] ),
    .S(net143),
    .X(_0602_));
 sg13g2_nand2_1 _1912_ (.Y(_0603_),
    .A(net166),
    .B(_0602_));
 sg13g2_a21oi_1 _1913_ (.A1(net109),
    .A2(\daisychain[98] ),
    .Y(_0604_),
    .B1(net54));
 sg13g2_o21ai_1 _1914_ (.B1(net188),
    .Y(_0605_),
    .A1(\daisychain[99] ),
    .A2(net33));
 sg13g2_a21oi_1 _1915_ (.A1(_0603_),
    .A2(_0604_),
    .Y(_0227_),
    .B1(_0605_));
 sg13g2_mux2_1 _1916_ (.A0(\state[100] ),
    .A1(\daisychain[100] ),
    .S(net143),
    .X(_0606_));
 sg13g2_nand2_1 _1917_ (.Y(_0607_),
    .A(net166),
    .B(_0606_));
 sg13g2_a21oi_1 _1918_ (.A1(net112),
    .A2(\daisychain[99] ),
    .Y(_0608_),
    .B1(net54));
 sg13g2_o21ai_1 _1919_ (.B1(net188),
    .Y(_0609_),
    .A1(\daisychain[100] ),
    .A2(net33));
 sg13g2_a21oi_1 _1920_ (.A1(_0607_),
    .A2(_0608_),
    .Y(_0228_),
    .B1(_0609_));
 sg13g2_mux2_1 _1921_ (.A0(\state[101] ),
    .A1(\daisychain[101] ),
    .S(net142),
    .X(_0610_));
 sg13g2_nand2_1 _1922_ (.Y(_0611_),
    .A(net165),
    .B(_0610_));
 sg13g2_a21oi_1 _1923_ (.A1(net112),
    .A2(\daisychain[100] ),
    .Y(_0612_),
    .B1(net54));
 sg13g2_o21ai_1 _1924_ (.B1(net187),
    .Y(_0613_),
    .A1(\daisychain[101] ),
    .A2(net32));
 sg13g2_a21oi_1 _1925_ (.A1(_0611_),
    .A2(_0612_),
    .Y(_0229_),
    .B1(_0613_));
 sg13g2_mux2_1 _1926_ (.A0(\state[102] ),
    .A1(\daisychain[102] ),
    .S(net142),
    .X(_0614_));
 sg13g2_nand2_1 _1927_ (.Y(_0615_),
    .A(net165),
    .B(_0614_));
 sg13g2_a21oi_1 _1928_ (.A1(net110),
    .A2(\daisychain[101] ),
    .Y(_0616_),
    .B1(net55));
 sg13g2_o21ai_1 _1929_ (.B1(net187),
    .Y(_0617_),
    .A1(\daisychain[102] ),
    .A2(net32));
 sg13g2_a21oi_1 _1930_ (.A1(_0615_),
    .A2(_0616_),
    .Y(_0230_),
    .B1(_0617_));
 sg13g2_mux2_1 _1931_ (.A0(\state[103] ),
    .A1(\daisychain[103] ),
    .S(net142),
    .X(_0618_));
 sg13g2_nand2_1 _1932_ (.Y(_0619_),
    .A(net165),
    .B(_0618_));
 sg13g2_a21oi_1 _1933_ (.A1(net110),
    .A2(\daisychain[102] ),
    .Y(_0620_),
    .B1(net55));
 sg13g2_o21ai_1 _1934_ (.B1(net187),
    .Y(_0621_),
    .A1(\daisychain[103] ),
    .A2(net32));
 sg13g2_a21oi_1 _1935_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0231_),
    .B1(_0621_));
 sg13g2_mux2_1 _1936_ (.A0(\state[104] ),
    .A1(\daisychain[104] ),
    .S(net142),
    .X(_0622_));
 sg13g2_nand2_1 _1937_ (.Y(_0623_),
    .A(net165),
    .B(_0622_));
 sg13g2_a21oi_1 _1938_ (.A1(net110),
    .A2(\daisychain[103] ),
    .Y(_0624_),
    .B1(net55));
 sg13g2_o21ai_1 _1939_ (.B1(net187),
    .Y(_0625_),
    .A1(\daisychain[104] ),
    .A2(net32));
 sg13g2_a21oi_1 _1940_ (.A1(_0623_),
    .A2(_0624_),
    .Y(_0232_),
    .B1(_0625_));
 sg13g2_mux2_1 _1941_ (.A0(\state[105] ),
    .A1(\daisychain[105] ),
    .S(net141),
    .X(_0626_));
 sg13g2_nand2_1 _1942_ (.Y(_0627_),
    .A(net163),
    .B(_0626_));
 sg13g2_a21oi_1 _1943_ (.A1(net107),
    .A2(\daisychain[104] ),
    .Y(_0628_),
    .B1(net53));
 sg13g2_o21ai_1 _1944_ (.B1(net185),
    .Y(_0629_),
    .A1(\daisychain[105] ),
    .A2(net30));
 sg13g2_a21oi_1 _1945_ (.A1(_0627_),
    .A2(_0628_),
    .Y(_0233_),
    .B1(_0629_));
 sg13g2_mux2_1 _1946_ (.A0(\state[106] ),
    .A1(\daisychain[106] ),
    .S(net141),
    .X(_0630_));
 sg13g2_nand2_1 _1947_ (.Y(_0631_),
    .A(net163),
    .B(_0630_));
 sg13g2_a21oi_1 _1948_ (.A1(net107),
    .A2(\daisychain[105] ),
    .Y(_0632_),
    .B1(net53));
 sg13g2_o21ai_1 _1949_ (.B1(net185),
    .Y(_0633_),
    .A1(\daisychain[106] ),
    .A2(net30));
 sg13g2_a21oi_1 _1950_ (.A1(_0631_),
    .A2(_0632_),
    .Y(_0234_),
    .B1(_0633_));
 sg13g2_mux2_1 _1951_ (.A0(\state[107] ),
    .A1(\daisychain[107] ),
    .S(net141),
    .X(_0634_));
 sg13g2_nand2_1 _1952_ (.Y(_0635_),
    .A(net163),
    .B(_0634_));
 sg13g2_a21oi_1 _1953_ (.A1(net107),
    .A2(\daisychain[106] ),
    .Y(_0636_),
    .B1(net53));
 sg13g2_o21ai_1 _1954_ (.B1(net185),
    .Y(_0637_),
    .A1(\daisychain[107] ),
    .A2(net30));
 sg13g2_a21oi_1 _1955_ (.A1(_0635_),
    .A2(_0636_),
    .Y(_0235_),
    .B1(_0637_));
 sg13g2_mux2_1 _1956_ (.A0(\state[108] ),
    .A1(\daisychain[108] ),
    .S(net141),
    .X(_0638_));
 sg13g2_nand2_1 _1957_ (.Y(_0639_),
    .A(net164),
    .B(_0638_));
 sg13g2_a21oi_1 _1958_ (.A1(net108),
    .A2(\daisychain[107] ),
    .Y(_0640_),
    .B1(net53));
 sg13g2_o21ai_1 _1959_ (.B1(net185),
    .Y(_0641_),
    .A1(\daisychain[108] ),
    .A2(net30));
 sg13g2_a21oi_1 _1960_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0236_),
    .B1(_0641_));
 sg13g2_mux2_1 _1961_ (.A0(\state[109] ),
    .A1(\daisychain[109] ),
    .S(net141),
    .X(_0642_));
 sg13g2_nand2_1 _1962_ (.Y(_0643_),
    .A(net164),
    .B(_0642_));
 sg13g2_a21oi_1 _1963_ (.A1(net108),
    .A2(\daisychain[108] ),
    .Y(_0644_),
    .B1(net53));
 sg13g2_o21ai_1 _1964_ (.B1(net186),
    .Y(_0645_),
    .A1(\daisychain[109] ),
    .A2(net31));
 sg13g2_a21oi_1 _1965_ (.A1(_0643_),
    .A2(_0644_),
    .Y(_0237_),
    .B1(_0645_));
 sg13g2_mux2_1 _1966_ (.A0(\state[110] ),
    .A1(\daisychain[110] ),
    .S(net144),
    .X(_0646_));
 sg13g2_nand2_1 _1967_ (.Y(_0647_),
    .A(net164),
    .B(_0646_));
 sg13g2_a21oi_1 _1968_ (.A1(net109),
    .A2(\daisychain[109] ),
    .Y(_0648_),
    .B1(net56));
 sg13g2_o21ai_1 _1969_ (.B1(net186),
    .Y(_0649_),
    .A1(\daisychain[110] ),
    .A2(net31));
 sg13g2_a21oi_1 _1970_ (.A1(_0647_),
    .A2(_0648_),
    .Y(_0238_),
    .B1(_0649_));
 sg13g2_mux2_1 _1971_ (.A0(\state[111] ),
    .A1(\daisychain[111] ),
    .S(net144),
    .X(_0650_));
 sg13g2_nand2_1 _1972_ (.Y(_0651_),
    .A(net164),
    .B(_0650_));
 sg13g2_a21oi_1 _1973_ (.A1(net109),
    .A2(\daisychain[110] ),
    .Y(_0652_),
    .B1(net56));
 sg13g2_o21ai_1 _1974_ (.B1(net186),
    .Y(_0653_),
    .A1(\daisychain[111] ),
    .A2(net31));
 sg13g2_a21oi_1 _1975_ (.A1(_0651_),
    .A2(_0652_),
    .Y(_0239_),
    .B1(_0653_));
 sg13g2_mux2_1 _1976_ (.A0(\state[112] ),
    .A1(\daisychain[112] ),
    .S(net141),
    .X(_0654_));
 sg13g2_nand2_1 _1977_ (.Y(_0655_),
    .A(net163),
    .B(_0654_));
 sg13g2_a21oi_1 _1978_ (.A1(net107),
    .A2(\daisychain[111] ),
    .Y(_0656_),
    .B1(net53));
 sg13g2_o21ai_1 _1979_ (.B1(net185),
    .Y(_0657_),
    .A1(\daisychain[112] ),
    .A2(net30));
 sg13g2_a21oi_1 _1980_ (.A1(_0655_),
    .A2(_0656_),
    .Y(_0240_),
    .B1(_0657_));
 sg13g2_mux2_1 _1981_ (.A0(\state[113] ),
    .A1(\daisychain[113] ),
    .S(net134),
    .X(_0658_));
 sg13g2_nand2_1 _1982_ (.Y(_0659_),
    .A(net163),
    .B(_0658_));
 sg13g2_a21oi_1 _1983_ (.A1(net95),
    .A2(\daisychain[112] ),
    .Y(_0660_),
    .B1(net53));
 sg13g2_o21ai_1 _1984_ (.B1(net185),
    .Y(_0661_),
    .A1(\daisychain[113] ),
    .A2(net30));
 sg13g2_a21oi_1 _1985_ (.A1(_0659_),
    .A2(_0660_),
    .Y(_0241_),
    .B1(_0661_));
 sg13g2_mux2_1 _1986_ (.A0(\state[114] ),
    .A1(\daisychain[114] ),
    .S(net141),
    .X(_0662_));
 sg13g2_nand2_1 _1987_ (.Y(_0663_),
    .A(net163),
    .B(_0662_));
 sg13g2_a21oi_1 _1988_ (.A1(net96),
    .A2(\daisychain[113] ),
    .Y(_0664_),
    .B1(net46));
 sg13g2_o21ai_1 _1989_ (.B1(net179),
    .Y(_0665_),
    .A1(\daisychain[114] ),
    .A2(net24));
 sg13g2_a21oi_1 _1990_ (.A1(_0663_),
    .A2(_0664_),
    .Y(_0242_),
    .B1(_0665_));
 sg13g2_mux2_1 _1991_ (.A0(\state[115] ),
    .A1(\daisychain[115] ),
    .S(net134),
    .X(_0666_));
 sg13g2_nand2_1 _1992_ (.Y(_0667_),
    .A(net157),
    .B(_0666_));
 sg13g2_a21oi_1 _1993_ (.A1(net96),
    .A2(\daisychain[114] ),
    .Y(_0668_),
    .B1(net46));
 sg13g2_o21ai_1 _1994_ (.B1(net179),
    .Y(_0669_),
    .A1(\daisychain[115] ),
    .A2(net24));
 sg13g2_a21oi_1 _1995_ (.A1(_0667_),
    .A2(_0668_),
    .Y(_0243_),
    .B1(_0669_));
 sg13g2_mux2_1 _1996_ (.A0(\state[116] ),
    .A1(\daisychain[116] ),
    .S(net134),
    .X(_0670_));
 sg13g2_nand2_1 _1997_ (.Y(_0671_),
    .A(net157),
    .B(_0670_));
 sg13g2_a21oi_1 _1998_ (.A1(net96),
    .A2(\daisychain[115] ),
    .Y(_0672_),
    .B1(net46));
 sg13g2_o21ai_1 _1999_ (.B1(net179),
    .Y(_0673_),
    .A1(\daisychain[116] ),
    .A2(net24));
 sg13g2_a21oi_1 _2000_ (.A1(_0671_),
    .A2(_0672_),
    .Y(_0244_),
    .B1(_0673_));
 sg13g2_mux2_1 _2001_ (.A0(\state[117] ),
    .A1(\daisychain[117] ),
    .S(net136),
    .X(_0674_));
 sg13g2_nand2_1 _2002_ (.Y(_0675_),
    .A(net157),
    .B(_0674_));
 sg13g2_a21oi_1 _2003_ (.A1(net95),
    .A2(\daisychain[116] ),
    .Y(_0676_),
    .B1(net46));
 sg13g2_o21ai_1 _2004_ (.B1(net179),
    .Y(_0677_),
    .A1(\daisychain[117] ),
    .A2(net24));
 sg13g2_a21oi_1 _2005_ (.A1(_0675_),
    .A2(_0676_),
    .Y(_0245_),
    .B1(_0677_));
 sg13g2_mux2_1 _2006_ (.A0(\state[118] ),
    .A1(\daisychain[118] ),
    .S(net136),
    .X(_0678_));
 sg13g2_nand2_1 _2007_ (.Y(_0679_),
    .A(net157),
    .B(_0678_));
 sg13g2_a21oi_1 _2008_ (.A1(net95),
    .A2(\daisychain[117] ),
    .Y(_0680_),
    .B1(net47));
 sg13g2_o21ai_1 _2009_ (.B1(net179),
    .Y(_0681_),
    .A1(\daisychain[118] ),
    .A2(net24));
 sg13g2_a21oi_1 _2010_ (.A1(_0679_),
    .A2(_0680_),
    .Y(_0246_),
    .B1(_0681_));
 sg13g2_mux2_1 _2011_ (.A0(\state[119] ),
    .A1(\daisychain[119] ),
    .S(net136),
    .X(_0682_));
 sg13g2_nand2_1 _2012_ (.Y(_0683_),
    .A(net157),
    .B(_0682_));
 sg13g2_a21oi_1 _2013_ (.A1(net97),
    .A2(\daisychain[118] ),
    .Y(_0684_),
    .B1(net46));
 sg13g2_o21ai_1 _2014_ (.B1(net179),
    .Y(_0685_),
    .A1(\daisychain[119] ),
    .A2(net24));
 sg13g2_a21oi_1 _2015_ (.A1(_0683_),
    .A2(_0684_),
    .Y(_0247_),
    .B1(_0685_));
 sg13g2_mux2_1 _2016_ (.A0(\state[120] ),
    .A1(\daisychain[120] ),
    .S(net135),
    .X(_0686_));
 sg13g2_nand2_1 _2017_ (.Y(_0687_),
    .A(net155),
    .B(_0686_));
 sg13g2_a21oi_1 _2018_ (.A1(net97),
    .A2(\daisychain[119] ),
    .Y(_0688_),
    .B1(net46));
 sg13g2_o21ai_1 _2019_ (.B1(net177),
    .Y(_0689_),
    .A1(\daisychain[120] ),
    .A2(net25));
 sg13g2_a21oi_1 _2020_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0248_),
    .B1(_0689_));
 sg13g2_mux2_1 _2021_ (.A0(\state[121] ),
    .A1(\daisychain[121] ),
    .S(net135),
    .X(_0690_));
 sg13g2_nand2_1 _2022_ (.Y(_0691_),
    .A(net155),
    .B(_0690_));
 sg13g2_a21oi_1 _2023_ (.A1(net90),
    .A2(\daisychain[120] ),
    .Y(_0692_),
    .B1(net48));
 sg13g2_o21ai_1 _2024_ (.B1(net177),
    .Y(_0693_),
    .A1(\daisychain[121] ),
    .A2(net25));
 sg13g2_a21oi_1 _2025_ (.A1(_0691_),
    .A2(_0692_),
    .Y(_0249_),
    .B1(_0693_));
 sg13g2_mux2_1 _2026_ (.A0(\state[122] ),
    .A1(\daisychain[122] ),
    .S(net135),
    .X(_0694_));
 sg13g2_nand2_1 _2027_ (.Y(_0695_),
    .A(net155),
    .B(_0694_));
 sg13g2_a21oi_1 _2028_ (.A1(net90),
    .A2(\daisychain[121] ),
    .Y(_0696_),
    .B1(net48));
 sg13g2_o21ai_1 _2029_ (.B1(net177),
    .Y(_0697_),
    .A1(\daisychain[122] ),
    .A2(net25));
 sg13g2_a21oi_1 _2030_ (.A1(_0695_),
    .A2(_0696_),
    .Y(_0250_),
    .B1(_0697_));
 sg13g2_mux2_1 _2031_ (.A0(\state[123] ),
    .A1(\daisychain[123] ),
    .S(net135),
    .X(_0698_));
 sg13g2_nand2_1 _2032_ (.Y(_0699_),
    .A(net155),
    .B(_0698_));
 sg13g2_a21oi_1 _2033_ (.A1(net90),
    .A2(\daisychain[122] ),
    .Y(_0700_),
    .B1(net48));
 sg13g2_o21ai_1 _2034_ (.B1(net177),
    .Y(_0701_),
    .A1(\daisychain[123] ),
    .A2(net25));
 sg13g2_a21oi_1 _2035_ (.A1(_0699_),
    .A2(_0700_),
    .Y(_0251_),
    .B1(_0701_));
 sg13g2_mux2_1 _2036_ (.A0(\state[124] ),
    .A1(\daisychain[124] ),
    .S(net135),
    .X(_0702_));
 sg13g2_nand2_1 _2037_ (.Y(_0703_),
    .A(net155),
    .B(_0702_));
 sg13g2_a21oi_1 _2038_ (.A1(net90),
    .A2(\daisychain[123] ),
    .Y(_0704_),
    .B1(net48));
 sg13g2_o21ai_1 _2039_ (.B1(net177),
    .Y(_0705_),
    .A1(\daisychain[124] ),
    .A2(net25));
 sg13g2_a21oi_1 _2040_ (.A1(_0703_),
    .A2(_0704_),
    .Y(_0252_),
    .B1(_0705_));
 sg13g2_mux2_1 _2041_ (.A0(\state[125] ),
    .A1(\daisychain[125] ),
    .S(net135),
    .X(_0706_));
 sg13g2_nand2_1 _2042_ (.Y(_0707_),
    .A(net155),
    .B(_0706_));
 sg13g2_a21oi_1 _2043_ (.A1(net90),
    .A2(\daisychain[124] ),
    .Y(_0708_),
    .B1(net48));
 sg13g2_o21ai_1 _2044_ (.B1(net177),
    .Y(_0709_),
    .A1(\daisychain[125] ),
    .A2(net25));
 sg13g2_a21oi_1 _2045_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0253_),
    .B1(_0709_));
 sg13g2_mux2_1 _2046_ (.A0(\state[126] ),
    .A1(\daisychain[126] ),
    .S(net135),
    .X(_0710_));
 sg13g2_nand2_1 _2047_ (.Y(_0711_),
    .A(net155),
    .B(_0710_));
 sg13g2_a21oi_1 _2048_ (.A1(net91),
    .A2(\daisychain[125] ),
    .Y(_0712_),
    .B1(net48));
 sg13g2_o21ai_1 _2049_ (.B1(net177),
    .Y(_0713_),
    .A1(\daisychain[126] ),
    .A2(net25));
 sg13g2_a21oi_1 _2050_ (.A1(_0711_),
    .A2(_0712_),
    .Y(_0254_),
    .B1(_0713_));
 sg13g2_mux2_1 _2051_ (.A0(\state[127] ),
    .A1(\daisychain[127] ),
    .S(net135),
    .X(_0714_));
 sg13g2_nand2_1 _2052_ (.Y(_0715_),
    .A(net155),
    .B(_0714_));
 sg13g2_a21oi_1 _2053_ (.A1(net91),
    .A2(\daisychain[126] ),
    .Y(_0716_),
    .B1(net48));
 sg13g2_o21ai_1 _2054_ (.B1(net180),
    .Y(_0717_),
    .A1(\daisychain[127] ),
    .A2(net25));
 sg13g2_a21oi_1 _2055_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0255_),
    .B1(_0717_));
 sg13g2_nand2_1 _2056_ (.Y(_0718_),
    .A(net94),
    .B(\state[0] ));
 sg13g2_a21oi_1 _2057_ (.A1(_0849_),
    .A2(_0718_),
    .Y(_0256_),
    .B1(net67));
 sg13g2_nand2_1 _2058_ (.Y(_0719_),
    .A(net94),
    .B(\state[1] ));
 sg13g2_a21oi_1 _2059_ (.A1(_0855_),
    .A2(_0719_),
    .Y(_0257_),
    .B1(net67));
 sg13g2_nand2_1 _2060_ (.Y(_0720_),
    .A(net92),
    .B(\state[2] ));
 sg13g2_a21oi_1 _2061_ (.A1(_0859_),
    .A2(_0720_),
    .Y(_0258_),
    .B1(net67));
 sg13g2_nand2_1 _2062_ (.Y(_0721_),
    .A(net92),
    .B(\state[3] ));
 sg13g2_a21oi_1 _2063_ (.A1(_0863_),
    .A2(_0721_),
    .Y(_0259_),
    .B1(net67));
 sg13g2_nand2_1 _2064_ (.Y(_0722_),
    .A(net93),
    .B(\state[4] ));
 sg13g2_a21oi_1 _2065_ (.A1(_0867_),
    .A2(_0722_),
    .Y(_0260_),
    .B1(net67));
 sg13g2_nand2_1 _2066_ (.Y(_0723_),
    .A(net93),
    .B(\state[5] ));
 sg13g2_a21oi_1 _2067_ (.A1(_0871_),
    .A2(_0723_),
    .Y(_0261_),
    .B1(net67));
 sg13g2_nand2_1 _2068_ (.Y(_0724_),
    .A(net101),
    .B(\state[6] ));
 sg13g2_a21oi_1 _2069_ (.A1(_0875_),
    .A2(_0724_),
    .Y(_0262_),
    .B1(net71));
 sg13g2_nand2_1 _2070_ (.Y(_0725_),
    .A(net101),
    .B(\state[7] ));
 sg13g2_a21oi_1 _2071_ (.A1(_0879_),
    .A2(_0725_),
    .Y(_0263_),
    .B1(net71));
 sg13g2_nand2_1 _2072_ (.Y(_0726_),
    .A(net101),
    .B(\state[8] ));
 sg13g2_a21oi_1 _2073_ (.A1(_0883_),
    .A2(_0726_),
    .Y(_0264_),
    .B1(net71));
 sg13g2_nand2_1 _2074_ (.Y(_0727_),
    .A(net101),
    .B(\state[9] ));
 sg13g2_a21oi_1 _2075_ (.A1(_0887_),
    .A2(_0727_),
    .Y(_0265_),
    .B1(net67));
 sg13g2_nand2_1 _2076_ (.Y(_0728_),
    .A(net93),
    .B(\state[10] ));
 sg13g2_a21oi_1 _2077_ (.A1(_0891_),
    .A2(_0728_),
    .Y(_0266_),
    .B1(net68));
 sg13g2_nand2_1 _2078_ (.Y(_0729_),
    .A(net92),
    .B(\state[11] ));
 sg13g2_a21oi_1 _2079_ (.A1(_0895_),
    .A2(_0729_),
    .Y(_0267_),
    .B1(net68));
 sg13g2_nand2_1 _2080_ (.Y(_0730_),
    .A(net92),
    .B(\state[12] ));
 sg13g2_a21oi_1 _2081_ (.A1(_0899_),
    .A2(_0730_),
    .Y(_0268_),
    .B1(net67));
 sg13g2_nand2_1 _2082_ (.Y(_0731_),
    .A(net93),
    .B(\state[13] ));
 sg13g2_a21oi_1 _2083_ (.A1(_0903_),
    .A2(_0731_),
    .Y(_0269_),
    .B1(net68));
 sg13g2_nand2_1 _2084_ (.Y(_0732_),
    .A(net93),
    .B(\state[14] ));
 sg13g2_a21oi_1 _2085_ (.A1(_0907_),
    .A2(_0732_),
    .Y(_0270_),
    .B1(net68));
 sg13g2_nand2_1 _2086_ (.Y(_0733_),
    .A(net101),
    .B(\state[15] ));
 sg13g2_a21oi_1 _2087_ (.A1(_0911_),
    .A2(_0733_),
    .Y(_0271_),
    .B1(net71));
 sg13g2_nand2_1 _2088_ (.Y(_0734_),
    .A(net99),
    .B(\state[16] ));
 sg13g2_a21oi_1 _2089_ (.A1(_0915_),
    .A2(_0734_),
    .Y(_0272_),
    .B1(net71));
 sg13g2_nand2_1 _2090_ (.Y(_0735_),
    .A(net99),
    .B(\state[17] ));
 sg13g2_a21oi_1 _2091_ (.A1(_0919_),
    .A2(_0735_),
    .Y(_0273_),
    .B1(net71));
 sg13g2_nand2_1 _2092_ (.Y(_0736_),
    .A(net99),
    .B(\state[18] ));
 sg13g2_a21oi_1 _2093_ (.A1(_0923_),
    .A2(_0736_),
    .Y(_0274_),
    .B1(net71));
 sg13g2_nand2_1 _2094_ (.Y(_0737_),
    .A(net102),
    .B(\state[19] ));
 sg13g2_a21oi_1 _2095_ (.A1(_0927_),
    .A2(_0737_),
    .Y(_0275_),
    .B1(net71));
 sg13g2_nand2_1 _2096_ (.Y(_0738_),
    .A(net104),
    .B(\state[20] ));
 sg13g2_a21oi_1 _2097_ (.A1(_0931_),
    .A2(_0738_),
    .Y(_0276_),
    .B1(net73));
 sg13g2_nand2_1 _2098_ (.Y(_0739_),
    .A(net103),
    .B(\state[21] ));
 sg13g2_a21oi_1 _2099_ (.A1(_0935_),
    .A2(_0739_),
    .Y(_0277_),
    .B1(net73));
 sg13g2_nand2_1 _2100_ (.Y(_0740_),
    .A(net104),
    .B(\state[22] ));
 sg13g2_a21oi_1 _2101_ (.A1(_0939_),
    .A2(_0740_),
    .Y(_0278_),
    .B1(net73));
 sg13g2_nand2_1 _2102_ (.Y(_0741_),
    .A(net104),
    .B(\state[23] ));
 sg13g2_a21oi_1 _2103_ (.A1(_0943_),
    .A2(_0741_),
    .Y(_0279_),
    .B1(net73));
 sg13g2_nand2_1 _2104_ (.Y(_0742_),
    .A(net105),
    .B(\state[24] ));
 sg13g2_a21oi_1 _2105_ (.A1(_0947_),
    .A2(_0742_),
    .Y(_0280_),
    .B1(net73));
 sg13g2_nand2_1 _2106_ (.Y(_0743_),
    .A(net100),
    .B(\state[25] ));
 sg13g2_a21oi_1 _2107_ (.A1(_0951_),
    .A2(_0743_),
    .Y(_0281_),
    .B1(net72));
 sg13g2_nand2_1 _2108_ (.Y(_0744_),
    .A(net100),
    .B(\state[26] ));
 sg13g2_a21oi_1 _2109_ (.A1(_0955_),
    .A2(_0744_),
    .Y(_0282_),
    .B1(net72));
 sg13g2_nand2_1 _2110_ (.Y(_0745_),
    .A(net100),
    .B(\state[27] ));
 sg13g2_a21oi_1 _2111_ (.A1(_0959_),
    .A2(_0745_),
    .Y(_0283_),
    .B1(net72));
 sg13g2_nand2_1 _2112_ (.Y(_0746_),
    .A(net102),
    .B(\state[28] ));
 sg13g2_a21oi_1 _2113_ (.A1(_0963_),
    .A2(_0746_),
    .Y(_0284_),
    .B1(net72));
 sg13g2_nand2_1 _2114_ (.Y(_0747_),
    .A(net105),
    .B(\state[29] ));
 sg13g2_a21oi_1 _2115_ (.A1(_0967_),
    .A2(_0747_),
    .Y(_0285_),
    .B1(net73));
 sg13g2_nand2_1 _2116_ (.Y(_0748_),
    .A(net105),
    .B(\state[30] ));
 sg13g2_a21oi_1 _2117_ (.A1(_0971_),
    .A2(_0748_),
    .Y(_0286_),
    .B1(net74));
 sg13g2_nand2_1 _2118_ (.Y(_0749_),
    .A(net105),
    .B(\state[31] ));
 sg13g2_a21oi_1 _2119_ (.A1(_0975_),
    .A2(_0749_),
    .Y(_0287_),
    .B1(net74));
 sg13g2_nand2_1 _2120_ (.Y(_0750_),
    .A(net106),
    .B(\state[32] ));
 sg13g2_a21oi_1 _2121_ (.A1(_0979_),
    .A2(_0750_),
    .Y(_0288_),
    .B1(net74));
 sg13g2_nand2_1 _2122_ (.Y(_0751_),
    .A(net117),
    .B(\state[33] ));
 sg13g2_a21oi_1 _2123_ (.A1(_0983_),
    .A2(_0751_),
    .Y(_0289_),
    .B1(net74));
 sg13g2_nand2_1 _2124_ (.Y(_0752_),
    .A(net116),
    .B(\state[34] ));
 sg13g2_a21oi_1 _2125_ (.A1(_0987_),
    .A2(_0752_),
    .Y(_0290_),
    .B1(net80));
 sg13g2_nand2_1 _2126_ (.Y(_0753_),
    .A(net116),
    .B(\state[35] ));
 sg13g2_a21oi_1 _2127_ (.A1(_0991_),
    .A2(_0753_),
    .Y(_0291_),
    .B1(net80));
 sg13g2_nand2_1 _2128_ (.Y(_0754_),
    .A(net116),
    .B(\state[36] ));
 sg13g2_a21oi_1 _2129_ (.A1(_0995_),
    .A2(_0754_),
    .Y(_0292_),
    .B1(net80));
 sg13g2_nand2_1 _2130_ (.Y(_0755_),
    .A(net103),
    .B(\state[37] ));
 sg13g2_a21oi_1 _2131_ (.A1(_0999_),
    .A2(_0755_),
    .Y(_0293_),
    .B1(net73));
 sg13g2_nand2_1 _2132_ (.Y(_0756_),
    .A(net103),
    .B(\state[38] ));
 sg13g2_a21oi_1 _2133_ (.A1(_1003_),
    .A2(_0756_),
    .Y(_0294_),
    .B1(net73));
 sg13g2_nand2_1 _2134_ (.Y(_0757_),
    .A(net116),
    .B(\state[39] ));
 sg13g2_a21oi_1 _2135_ (.A1(_1007_),
    .A2(_0757_),
    .Y(_0295_),
    .B1(net80));
 sg13g2_nand2_1 _2136_ (.Y(_0758_),
    .A(net115),
    .B(\state[40] ));
 sg13g2_a21oi_1 _2137_ (.A1(_1011_),
    .A2(_0758_),
    .Y(_0296_),
    .B1(net80));
 sg13g2_nand2_1 _2138_ (.Y(_0759_),
    .A(net115),
    .B(\state[41] ));
 sg13g2_a21oi_1 _2139_ (.A1(_1015_),
    .A2(_0759_),
    .Y(_0297_),
    .B1(net80));
 sg13g2_nand2_1 _2140_ (.Y(_0760_),
    .A(net115),
    .B(\state[42] ));
 sg13g2_a21oi_1 _2141_ (.A1(_1019_),
    .A2(_0760_),
    .Y(_0298_),
    .B1(net80));
 sg13g2_nand2_1 _2142_ (.Y(_0761_),
    .A(net115),
    .B(\state[43] ));
 sg13g2_a21oi_1 _2143_ (.A1(_1023_),
    .A2(_0761_),
    .Y(_0299_),
    .B1(net80));
 sg13g2_nand2_1 _2144_ (.Y(_0762_),
    .A(net117),
    .B(\state[44] ));
 sg13g2_a21oi_1 _2145_ (.A1(_1027_),
    .A2(_0762_),
    .Y(_0300_),
    .B1(net81));
 sg13g2_nand2_1 _2146_ (.Y(_0763_),
    .A(net117),
    .B(\state[45] ));
 sg13g2_a21oi_1 _2147_ (.A1(_0387_),
    .A2(_0763_),
    .Y(_0301_),
    .B1(net81));
 sg13g2_nand2_1 _2148_ (.Y(_0764_),
    .A(net117),
    .B(\state[46] ));
 sg13g2_a21oi_1 _2149_ (.A1(_0391_),
    .A2(_0764_),
    .Y(_0302_),
    .B1(net81));
 sg13g2_nand2_1 _2150_ (.Y(_0765_),
    .A(net123),
    .B(\state[47] ));
 sg13g2_a21oi_1 _2151_ (.A1(_0395_),
    .A2(_0765_),
    .Y(_0303_),
    .B1(net81));
 sg13g2_nand2_1 _2152_ (.Y(_0766_),
    .A(net122),
    .B(\state[48] ));
 sg13g2_a21oi_1 _2153_ (.A1(_0399_),
    .A2(_0766_),
    .Y(_0304_),
    .B1(net83));
 sg13g2_nand2_1 _2154_ (.Y(_0767_),
    .A(net122),
    .B(\state[49] ));
 sg13g2_a21oi_1 _2155_ (.A1(_0403_),
    .A2(_0767_),
    .Y(_0305_),
    .B1(net83));
 sg13g2_nand2_1 _2156_ (.Y(_0768_),
    .A(net118),
    .B(\state[50] ));
 sg13g2_a21oi_1 _2157_ (.A1(_0407_),
    .A2(_0768_),
    .Y(_0306_),
    .B1(net82));
 sg13g2_nand2_1 _2158_ (.Y(_0769_),
    .A(net121),
    .B(\state[51] ));
 sg13g2_a21oi_1 _2159_ (.A1(_0411_),
    .A2(_0769_),
    .Y(_0307_),
    .B1(net82));
 sg13g2_nand2_1 _2160_ (.Y(_0770_),
    .A(net121),
    .B(\state[52] ));
 sg13g2_a21oi_1 _2161_ (.A1(_0415_),
    .A2(_0770_),
    .Y(_0308_),
    .B1(net82));
 sg13g2_nand2_1 _2162_ (.Y(_0771_),
    .A(net118),
    .B(\state[53] ));
 sg13g2_a21oi_1 _2163_ (.A1(_0419_),
    .A2(_0771_),
    .Y(_0309_),
    .B1(net82));
 sg13g2_nand2_1 _2164_ (.Y(_0772_),
    .A(net118),
    .B(\state[54] ));
 sg13g2_a21oi_1 _2165_ (.A1(_0423_),
    .A2(_0772_),
    .Y(_0310_),
    .B1(net82));
 sg13g2_nand2_1 _2166_ (.Y(_0773_),
    .A(net119),
    .B(\state[55] ));
 sg13g2_a21oi_1 _2167_ (.A1(_0427_),
    .A2(_0773_),
    .Y(_0311_),
    .B1(net82));
 sg13g2_nand2_1 _2168_ (.Y(_0774_),
    .A(net119),
    .B(\state[56] ));
 sg13g2_a21oi_1 _2169_ (.A1(_0431_),
    .A2(_0774_),
    .Y(_0312_),
    .B1(net82));
 sg13g2_nand2_1 _2170_ (.Y(_0775_),
    .A(net119),
    .B(\state[57] ));
 sg13g2_a21oi_1 _2171_ (.A1(_0435_),
    .A2(_0775_),
    .Y(_0313_),
    .B1(net82));
 sg13g2_nand2_1 _2172_ (.Y(_0776_),
    .A(net120),
    .B(\state[58] ));
 sg13g2_a21oi_1 _2173_ (.A1(_0439_),
    .A2(_0776_),
    .Y(_0314_),
    .B1(net83));
 sg13g2_nand2_1 _2174_ (.Y(_0777_),
    .A(net120),
    .B(\state[59] ));
 sg13g2_a21oi_1 _2175_ (.A1(_0443_),
    .A2(_0777_),
    .Y(_0315_),
    .B1(net83));
 sg13g2_nand2_1 _2176_ (.Y(_0778_),
    .A(net120),
    .B(\state[60] ));
 sg13g2_a21oi_1 _2177_ (.A1(_0447_),
    .A2(_0778_),
    .Y(_0316_),
    .B1(net83));
 sg13g2_nand2_1 _2178_ (.Y(_0779_),
    .A(net122),
    .B(\state[61] ));
 sg13g2_a21oi_1 _2179_ (.A1(_0451_),
    .A2(_0779_),
    .Y(_0317_),
    .B1(net83));
 sg13g2_nand2_1 _2180_ (.Y(_0780_),
    .A(net122),
    .B(\state[62] ));
 sg13g2_a21oi_1 _2181_ (.A1(_0455_),
    .A2(_0780_),
    .Y(_0318_),
    .B1(net83));
 sg13g2_nand2_1 _2182_ (.Y(_0781_),
    .A(net123),
    .B(\state[63] ));
 sg13g2_a21oi_1 _2183_ (.A1(_0459_),
    .A2(_0781_),
    .Y(_0319_),
    .B1(net88));
 sg13g2_nand2_1 _2184_ (.Y(_0782_),
    .A(net127),
    .B(\state[64] ));
 sg13g2_a21oi_1 _2185_ (.A1(_0463_),
    .A2(_0782_),
    .Y(_0320_),
    .B1(net87));
 sg13g2_nand2_1 _2186_ (.Y(_0783_),
    .A(net131),
    .B(\state[65] ));
 sg13g2_a21oi_1 _2187_ (.A1(_0467_),
    .A2(_0783_),
    .Y(_0321_),
    .B1(net87));
 sg13g2_nand2_1 _2188_ (.Y(_0784_),
    .A(net129),
    .B(\state[66] ));
 sg13g2_a21oi_1 _2189_ (.A1(_0471_),
    .A2(_0784_),
    .Y(_0322_),
    .B1(net86));
 sg13g2_nand2_1 _2190_ (.Y(_0785_),
    .A(net129),
    .B(\state[67] ));
 sg13g2_a21oi_1 _2191_ (.A1(_0475_),
    .A2(_0785_),
    .Y(_0323_),
    .B1(net86));
 sg13g2_nand2_1 _2192_ (.Y(_0786_),
    .A(net129),
    .B(\state[68] ));
 sg13g2_a21oi_1 _2193_ (.A1(_0479_),
    .A2(_0786_),
    .Y(_0324_),
    .B1(net86));
 sg13g2_nand2_1 _2194_ (.Y(_0787_),
    .A(net130),
    .B(\state[69] ));
 sg13g2_a21oi_1 _2195_ (.A1(_0483_),
    .A2(_0787_),
    .Y(_0325_),
    .B1(net86));
 sg13g2_nand2_1 _2196_ (.Y(_0788_),
    .A(net130),
    .B(\state[70] ));
 sg13g2_a21oi_1 _2197_ (.A1(_0487_),
    .A2(_0788_),
    .Y(_0326_),
    .B1(net87));
 sg13g2_nand2_1 _2198_ (.Y(_0789_),
    .A(net130),
    .B(\state[71] ));
 sg13g2_a21oi_1 _2199_ (.A1(_0491_),
    .A2(_0789_),
    .Y(_0327_),
    .B1(net87));
 sg13g2_nand2_1 _2200_ (.Y(_0790_),
    .A(net128),
    .B(\state[72] ));
 sg13g2_a21oi_1 _2201_ (.A1(_0495_),
    .A2(_0790_),
    .Y(_0328_),
    .B1(net86));
 sg13g2_nand2_1 _2202_ (.Y(_0791_),
    .A(net130),
    .B(\state[73] ));
 sg13g2_a21oi_1 _2203_ (.A1(_0499_),
    .A2(_0791_),
    .Y(_0329_),
    .B1(net86));
 sg13g2_nand2_1 _2204_ (.Y(_0792_),
    .A(net125),
    .B(\state[74] ));
 sg13g2_a21oi_1 _2205_ (.A1(_0503_),
    .A2(_0792_),
    .Y(_0330_),
    .B1(net84));
 sg13g2_nand2_1 _2206_ (.Y(_0793_),
    .A(net125),
    .B(\state[75] ));
 sg13g2_a21oi_1 _2207_ (.A1(_0507_),
    .A2(_0793_),
    .Y(_0331_),
    .B1(net84));
 sg13g2_nand2_1 _2208_ (.Y(_0794_),
    .A(net128),
    .B(\state[76] ));
 sg13g2_a21oi_1 _2209_ (.A1(_0511_),
    .A2(_0794_),
    .Y(_0332_),
    .B1(net86));
 sg13g2_nand2_1 _2210_ (.Y(_0795_),
    .A(net128),
    .B(\state[77] ));
 sg13g2_a21oi_1 _2211_ (.A1(_0515_),
    .A2(_0795_),
    .Y(_0333_),
    .B1(net86));
 sg13g2_nand2_1 _2212_ (.Y(_0796_),
    .A(net127),
    .B(\state[78] ));
 sg13g2_a21oi_1 _2213_ (.A1(_0519_),
    .A2(_0796_),
    .Y(_0334_),
    .B1(net87));
 sg13g2_nand2_1 _2214_ (.Y(_0797_),
    .A(net127),
    .B(\state[79] ));
 sg13g2_a21oi_1 _2215_ (.A1(_0523_),
    .A2(_0797_),
    .Y(_0335_),
    .B1(net87));
 sg13g2_nand2_1 _2216_ (.Y(_0798_),
    .A(net126),
    .B(\state[80] ));
 sg13g2_a21oi_1 _2217_ (.A1(_0527_),
    .A2(_0798_),
    .Y(_0336_),
    .B1(net84));
 sg13g2_nand2_1 _2218_ (.Y(_0799_),
    .A(net126),
    .B(\state[81] ));
 sg13g2_a21oi_1 _2219_ (.A1(_0531_),
    .A2(_0799_),
    .Y(_0337_),
    .B1(net84));
 sg13g2_nand2_1 _2220_ (.Y(_0800_),
    .A(net126),
    .B(\state[82] ));
 sg13g2_a21oi_1 _2221_ (.A1(_0535_),
    .A2(_0800_),
    .Y(_0338_),
    .B1(net84));
 sg13g2_nand2_1 _2222_ (.Y(_0801_),
    .A(net131),
    .B(\state[83] ));
 sg13g2_a21oi_1 _2223_ (.A1(_0539_),
    .A2(_0801_),
    .Y(_0339_),
    .B1(net84));
 sg13g2_nand2_1 _2224_ (.Y(_0802_),
    .A(net124),
    .B(\state[84] ));
 sg13g2_a21oi_1 _2225_ (.A1(_0543_),
    .A2(_0802_),
    .Y(_0340_),
    .B1(net85));
 sg13g2_nand2_1 _2226_ (.Y(_0803_),
    .A(net125),
    .B(\state[85] ));
 sg13g2_a21oi_1 _2227_ (.A1(_0547_),
    .A2(_0803_),
    .Y(_0341_),
    .B1(net85));
 sg13g2_nand2_1 _2228_ (.Y(_0804_),
    .A(net131),
    .B(\state[86] ));
 sg13g2_a21oi_1 _2229_ (.A1(_0551_),
    .A2(_0804_),
    .Y(_0342_),
    .B1(net85));
 sg13g2_nand2_1 _2230_ (.Y(_0805_),
    .A(net125),
    .B(\state[87] ));
 sg13g2_a21oi_1 _2231_ (.A1(_0555_),
    .A2(_0805_),
    .Y(_0343_),
    .B1(net77));
 sg13g2_nand2_1 _2232_ (.Y(_0806_),
    .A(net111),
    .B(\state[88] ));
 sg13g2_a21oi_1 _2233_ (.A1(_0559_),
    .A2(_0806_),
    .Y(_0344_),
    .B1(net77));
 sg13g2_nand2_1 _2234_ (.Y(_0807_),
    .A(net111),
    .B(\state[89] ));
 sg13g2_a21oi_1 _2235_ (.A1(_0563_),
    .A2(_0807_),
    .Y(_0345_),
    .B1(net77));
 sg13g2_nand2_1 _2236_ (.Y(_0808_),
    .A(net124),
    .B(\state[90] ));
 sg13g2_a21oi_1 _2237_ (.A1(_0567_),
    .A2(_0808_),
    .Y(_0346_),
    .B1(net85));
 sg13g2_nand2_1 _2238_ (.Y(_0809_),
    .A(net126),
    .B(\state[91] ));
 sg13g2_a21oi_1 _2239_ (.A1(_0571_),
    .A2(_0809_),
    .Y(_0347_),
    .B1(net84));
 sg13g2_nand2_1 _2240_ (.Y(_0810_),
    .A(net126),
    .B(\state[92] ));
 sg13g2_a21oi_1 _2241_ (.A1(_0575_),
    .A2(_0810_),
    .Y(_0348_),
    .B1(net84));
 sg13g2_nand2_1 _2242_ (.Y(_0811_),
    .A(net113),
    .B(\state[93] ));
 sg13g2_a21oi_1 _2243_ (.A1(_0579_),
    .A2(_0811_),
    .Y(_0349_),
    .B1(net78));
 sg13g2_nand2_1 _2244_ (.Y(_0812_),
    .A(net111),
    .B(\state[94] ));
 sg13g2_a21oi_1 _2245_ (.A1(_0583_),
    .A2(_0812_),
    .Y(_0350_),
    .B1(net77));
 sg13g2_nand2_1 _2246_ (.Y(_0813_),
    .A(net111),
    .B(\state[95] ));
 sg13g2_a21oi_1 _2247_ (.A1(_0587_),
    .A2(_0813_),
    .Y(_0351_),
    .B1(net77));
 sg13g2_nand2_1 _2248_ (.Y(_0814_),
    .A(net112),
    .B(\state[96] ));
 sg13g2_a21oi_1 _2249_ (.A1(_0591_),
    .A2(_0814_),
    .Y(_0352_),
    .B1(net78));
 sg13g2_nand2_1 _2250_ (.Y(_0815_),
    .A(net112),
    .B(\state[97] ));
 sg13g2_a21oi_1 _2251_ (.A1(_0595_),
    .A2(_0815_),
    .Y(_0353_),
    .B1(net77));
 sg13g2_nand2_1 _2252_ (.Y(_0816_),
    .A(net109),
    .B(\state[98] ));
 sg13g2_a21oi_1 _2253_ (.A1(_0599_),
    .A2(_0816_),
    .Y(_0354_),
    .B1(net76));
 sg13g2_nand2_1 _2254_ (.Y(_0817_),
    .A(net112),
    .B(\state[99] ));
 sg13g2_a21oi_1 _2255_ (.A1(_0603_),
    .A2(_0817_),
    .Y(_0355_),
    .B1(net77));
 sg13g2_nand2_1 _2256_ (.Y(_0818_),
    .A(net112),
    .B(\state[100] ));
 sg13g2_a21oi_1 _2257_ (.A1(_0607_),
    .A2(_0818_),
    .Y(_0356_),
    .B1(net77));
 sg13g2_nand2_1 _2258_ (.Y(_0819_),
    .A(net110),
    .B(\state[101] ));
 sg13g2_a21oi_1 _2259_ (.A1(_0611_),
    .A2(_0819_),
    .Y(_0357_),
    .B1(net78));
 sg13g2_nand2_1 _2260_ (.Y(_0820_),
    .A(net110),
    .B(\state[102] ));
 sg13g2_a21oi_1 _2261_ (.A1(_0615_),
    .A2(_0820_),
    .Y(_0358_),
    .B1(net78));
 sg13g2_nand2_1 _2262_ (.Y(_0821_),
    .A(net110),
    .B(\state[103] ));
 sg13g2_a21oi_1 _2263_ (.A1(_0619_),
    .A2(_0821_),
    .Y(_0359_),
    .B1(net78));
 sg13g2_nand2_1 _2264_ (.Y(_0822_),
    .A(net110),
    .B(\state[104] ));
 sg13g2_a21oi_1 _2265_ (.A1(_0623_),
    .A2(_0822_),
    .Y(_0360_),
    .B1(net78));
 sg13g2_nand2_1 _2266_ (.Y(_0823_),
    .A(net108),
    .B(\state[105] ));
 sg13g2_a21oi_1 _2267_ (.A1(_0627_),
    .A2(_0823_),
    .Y(_0361_),
    .B1(net76));
 sg13g2_nand2_1 _2268_ (.Y(_0824_),
    .A(net108),
    .B(\state[106] ));
 sg13g2_a21oi_1 _2269_ (.A1(_0631_),
    .A2(_0824_),
    .Y(_0362_),
    .B1(net76));
 sg13g2_nand2_1 _2270_ (.Y(_0825_),
    .A(net108),
    .B(\state[107] ));
 sg13g2_a21oi_1 _2271_ (.A1(_0635_),
    .A2(_0825_),
    .Y(_0363_),
    .B1(net76));
 sg13g2_nand2_1 _2272_ (.Y(_0826_),
    .A(net108),
    .B(\state[108] ));
 sg13g2_a21oi_1 _2273_ (.A1(_0639_),
    .A2(_0826_),
    .Y(_0364_),
    .B1(net76));
 sg13g2_nand2_1 _2274_ (.Y(_0827_),
    .A(net109),
    .B(\state[109] ));
 sg13g2_a21oi_1 _2275_ (.A1(_0643_),
    .A2(_0827_),
    .Y(_0365_),
    .B1(net76));
 sg13g2_nand2_1 _2276_ (.Y(_0828_),
    .A(net114),
    .B(\state[110] ));
 sg13g2_a21oi_1 _2277_ (.A1(_0647_),
    .A2(_0828_),
    .Y(_0366_),
    .B1(net79));
 sg13g2_nand2_1 _2278_ (.Y(_0829_),
    .A(net114),
    .B(\state[111] ));
 sg13g2_a21oi_1 _2279_ (.A1(_0651_),
    .A2(_0829_),
    .Y(_0367_),
    .B1(net79));
 sg13g2_nand2_1 _2280_ (.Y(_0830_),
    .A(net107),
    .B(\state[112] ));
 sg13g2_a21oi_1 _2281_ (.A1(_0655_),
    .A2(_0830_),
    .Y(_0368_),
    .B1(net76));
 sg13g2_nand2_1 _2282_ (.Y(_0831_),
    .A(net107),
    .B(\state[113] ));
 sg13g2_a21oi_1 _2283_ (.A1(_0659_),
    .A2(_0831_),
    .Y(_0369_),
    .B1(net69));
 sg13g2_nand2_1 _2284_ (.Y(_0832_),
    .A(net107),
    .B(\state[114] ));
 sg13g2_a21oi_1 _2285_ (.A1(_0663_),
    .A2(_0832_),
    .Y(_0370_),
    .B1(net76));
 sg13g2_nand2_1 _2286_ (.Y(_0833_),
    .A(net96),
    .B(\state[115] ));
 sg13g2_a21oi_1 _2287_ (.A1(_0667_),
    .A2(_0833_),
    .Y(_0371_),
    .B1(net69));
 sg13g2_nand2_1 _2288_ (.Y(_0834_),
    .A(net96),
    .B(\state[116] ));
 sg13g2_a21oi_1 _2289_ (.A1(_0671_),
    .A2(_0834_),
    .Y(_0372_),
    .B1(net69));
 sg13g2_nand2_1 _2290_ (.Y(_0835_),
    .A(net95),
    .B(\state[117] ));
 sg13g2_a21oi_1 _2291_ (.A1(_0675_),
    .A2(_0835_),
    .Y(_0373_),
    .B1(net69));
 sg13g2_nand2_1 _2292_ (.Y(_0836_),
    .A(net95),
    .B(\state[118] ));
 sg13g2_a21oi_1 _2293_ (.A1(_0679_),
    .A2(_0836_),
    .Y(_0374_),
    .B1(net69));
 sg13g2_nand2_1 _2294_ (.Y(_0837_),
    .A(net97),
    .B(\state[119] ));
 sg13g2_a21oi_1 _2295_ (.A1(_0683_),
    .A2(_0837_),
    .Y(_0375_),
    .B1(net69));
 sg13g2_nand2_1 _2296_ (.Y(_0838_),
    .A(net91),
    .B(\state[120] ));
 sg13g2_a21oi_1 _2297_ (.A1(_0687_),
    .A2(_0838_),
    .Y(_0376_),
    .B1(net70));
 sg13g2_nand2_1 _2298_ (.Y(_0839_),
    .A(net90),
    .B(\state[121] ));
 sg13g2_a21oi_1 _2299_ (.A1(_0691_),
    .A2(_0839_),
    .Y(_0377_),
    .B1(net70));
 sg13g2_nand2_1 _2300_ (.Y(_0840_),
    .A(net90),
    .B(\state[122] ));
 sg13g2_a21oi_1 _2301_ (.A1(_0695_),
    .A2(_0840_),
    .Y(_0378_),
    .B1(net70));
 sg13g2_nand2_1 _2302_ (.Y(_0841_),
    .A(net90),
    .B(\state[123] ));
 sg13g2_a21oi_1 _2303_ (.A1(_0699_),
    .A2(_0841_),
    .Y(_0379_),
    .B1(net70));
 sg13g2_nand2_1 _2304_ (.Y(_0842_),
    .A(net91),
    .B(\state[124] ));
 sg13g2_a21oi_1 _2305_ (.A1(_0703_),
    .A2(_0842_),
    .Y(_0380_),
    .B1(net70));
 sg13g2_nand2_1 _2306_ (.Y(_0843_),
    .A(net91),
    .B(\state[125] ));
 sg13g2_a21oi_1 _2307_ (.A1(_0707_),
    .A2(_0843_),
    .Y(_0381_),
    .B1(net70));
 sg13g2_nand2_1 _2308_ (.Y(_0844_),
    .A(net91),
    .B(\state[126] ));
 sg13g2_a21oi_1 _2309_ (.A1(_0711_),
    .A2(_0844_),
    .Y(_0382_),
    .B1(net70));
 sg13g2_nand2_1 _2310_ (.Y(_0845_),
    .A(\state[127] ),
    .B(net91));
 sg13g2_a21oi_1 _2311_ (.A1(_0715_),
    .A2(_0845_),
    .Y(_0383_),
    .B1(net70));
 sg13g2_dfrbpq_1 _2312_ (.RESET_B(net325),
    .D(_0128_),
    .Q(\daisychain[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2313_ (.RESET_B(net324),
    .D(_0129_),
    .Q(\daisychain[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2314_ (.RESET_B(net322),
    .D(_0130_),
    .Q(\daisychain[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net320),
    .D(_0131_),
    .Q(\daisychain[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net318),
    .D(_0132_),
    .Q(\daisychain[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net316),
    .D(_0133_),
    .Q(\daisychain[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net314),
    .D(_0134_),
    .Q(\daisychain[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2319_ (.RESET_B(net312),
    .D(_0135_),
    .Q(\daisychain[7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net310),
    .D(_0136_),
    .Q(\daisychain[8] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net308),
    .D(_0137_),
    .Q(\daisychain[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net306),
    .D(_0138_),
    .Q(\daisychain[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2323_ (.RESET_B(net304),
    .D(_0139_),
    .Q(\daisychain[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2324_ (.RESET_B(net302),
    .D(_0140_),
    .Q(\daisychain[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2325_ (.RESET_B(net300),
    .D(_0141_),
    .Q(\daisychain[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2326_ (.RESET_B(net298),
    .D(_0142_),
    .Q(\daisychain[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2327_ (.RESET_B(net296),
    .D(_0143_),
    .Q(\daisychain[15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net294),
    .D(_0144_),
    .Q(\daisychain[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2329_ (.RESET_B(net292),
    .D(_0145_),
    .Q(\daisychain[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2330_ (.RESET_B(net290),
    .D(_0146_),
    .Q(\daisychain[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2331_ (.RESET_B(net288),
    .D(_0147_),
    .Q(\daisychain[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2332_ (.RESET_B(net286),
    .D(_0148_),
    .Q(\daisychain[20] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net284),
    .D(_0149_),
    .Q(\daisychain[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net282),
    .D(_0150_),
    .Q(\daisychain[22] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net280),
    .D(_0151_),
    .Q(\daisychain[23] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2336_ (.RESET_B(net278),
    .D(_0152_),
    .Q(\daisychain[24] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2337_ (.RESET_B(net276),
    .D(_0153_),
    .Q(\daisychain[25] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2338_ (.RESET_B(net274),
    .D(_0154_),
    .Q(\daisychain[26] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2339_ (.RESET_B(net272),
    .D(_0155_),
    .Q(\daisychain[27] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2340_ (.RESET_B(net270),
    .D(_0156_),
    .Q(\daisychain[28] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2341_ (.RESET_B(net268),
    .D(_0157_),
    .Q(\daisychain[29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2342_ (.RESET_B(net266),
    .D(_0158_),
    .Q(\daisychain[30] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2343_ (.RESET_B(net264),
    .D(_0159_),
    .Q(\daisychain[31] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net262),
    .D(_0160_),
    .Q(\daisychain[32] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net260),
    .D(_0161_),
    .Q(\daisychain[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2346_ (.RESET_B(net258),
    .D(_0162_),
    .Q(\daisychain[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2347_ (.RESET_B(net256),
    .D(_0163_),
    .Q(\daisychain[35] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net254),
    .D(_0164_),
    .Q(\daisychain[36] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net252),
    .D(_0165_),
    .Q(\daisychain[37] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net250),
    .D(_0166_),
    .Q(\daisychain[38] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2351_ (.RESET_B(net248),
    .D(_0167_),
    .Q(\daisychain[39] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2352_ (.RESET_B(net246),
    .D(_0168_),
    .Q(\daisychain[40] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2353_ (.RESET_B(net244),
    .D(_0169_),
    .Q(\daisychain[41] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2354_ (.RESET_B(net242),
    .D(_0170_),
    .Q(\daisychain[42] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2355_ (.RESET_B(net240),
    .D(_0171_),
    .Q(\daisychain[43] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2356_ (.RESET_B(net238),
    .D(_0172_),
    .Q(\daisychain[44] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2357_ (.RESET_B(net236),
    .D(_0173_),
    .Q(\daisychain[45] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2358_ (.RESET_B(net234),
    .D(_0174_),
    .Q(\daisychain[46] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2359_ (.RESET_B(net232),
    .D(_0175_),
    .Q(\daisychain[47] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2360_ (.RESET_B(net230),
    .D(_0176_),
    .Q(\daisychain[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2361_ (.RESET_B(net228),
    .D(_0177_),
    .Q(\daisychain[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2362_ (.RESET_B(net226),
    .D(_0178_),
    .Q(\daisychain[50] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2363_ (.RESET_B(net224),
    .D(_0179_),
    .Q(\daisychain[51] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2364_ (.RESET_B(net222),
    .D(_0180_),
    .Q(\daisychain[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2365_ (.RESET_B(net220),
    .D(_0181_),
    .Q(\daisychain[53] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2366_ (.RESET_B(net218),
    .D(_0182_),
    .Q(\daisychain[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2367_ (.RESET_B(net216),
    .D(_0183_),
    .Q(\daisychain[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2368_ (.RESET_B(net214),
    .D(_0184_),
    .Q(\daisychain[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2369_ (.RESET_B(net212),
    .D(_0185_),
    .Q(\daisychain[57] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2370_ (.RESET_B(net210),
    .D(_0186_),
    .Q(\daisychain[58] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2371_ (.RESET_B(net208),
    .D(_0187_),
    .Q(\daisychain[59] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2372_ (.RESET_B(net206),
    .D(_0188_),
    .Q(\daisychain[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2373_ (.RESET_B(net204),
    .D(_0189_),
    .Q(\daisychain[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2374_ (.RESET_B(net202),
    .D(_0190_),
    .Q(\daisychain[62] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2375_ (.RESET_B(net200),
    .D(_0191_),
    .Q(\daisychain[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2376_ (.RESET_B(net454),
    .D(_0192_),
    .Q(\daisychain[64] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2377_ (.RESET_B(net452),
    .D(_0193_),
    .Q(\daisychain[65] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2378_ (.RESET_B(net450),
    .D(_0194_),
    .Q(\daisychain[66] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2379_ (.RESET_B(net448),
    .D(_0195_),
    .Q(\daisychain[67] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2380_ (.RESET_B(net446),
    .D(_0196_),
    .Q(\daisychain[68] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2381_ (.RESET_B(net444),
    .D(_0197_),
    .Q(\daisychain[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2382_ (.RESET_B(net442),
    .D(_0198_),
    .Q(\daisychain[70] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2383_ (.RESET_B(net440),
    .D(_0199_),
    .Q(\daisychain[71] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2384_ (.RESET_B(net438),
    .D(_0200_),
    .Q(\daisychain[72] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2385_ (.RESET_B(net436),
    .D(_0201_),
    .Q(\daisychain[73] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2386_ (.RESET_B(net434),
    .D(_0202_),
    .Q(\daisychain[74] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2387_ (.RESET_B(net432),
    .D(_0203_),
    .Q(\daisychain[75] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2388_ (.RESET_B(net430),
    .D(_0204_),
    .Q(\daisychain[76] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2389_ (.RESET_B(net428),
    .D(_0205_),
    .Q(\daisychain[77] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2390_ (.RESET_B(net426),
    .D(_0206_),
    .Q(\daisychain[78] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2391_ (.RESET_B(net424),
    .D(_0207_),
    .Q(\daisychain[79] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2392_ (.RESET_B(net422),
    .D(_0208_),
    .Q(\daisychain[80] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2393_ (.RESET_B(net420),
    .D(_0209_),
    .Q(\daisychain[81] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2394_ (.RESET_B(net418),
    .D(_0210_),
    .Q(\daisychain[82] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2395_ (.RESET_B(net416),
    .D(_0211_),
    .Q(\daisychain[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2396_ (.RESET_B(net414),
    .D(_0212_),
    .Q(\daisychain[84] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2397_ (.RESET_B(net412),
    .D(_0213_),
    .Q(\daisychain[85] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2398_ (.RESET_B(net410),
    .D(_0214_),
    .Q(\daisychain[86] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2399_ (.RESET_B(net408),
    .D(_0215_),
    .Q(\daisychain[87] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2400_ (.RESET_B(net406),
    .D(_0216_),
    .Q(\daisychain[88] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2401_ (.RESET_B(net404),
    .D(_0217_),
    .Q(\daisychain[89] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2402_ (.RESET_B(net402),
    .D(_0218_),
    .Q(\daisychain[90] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2403_ (.RESET_B(net400),
    .D(_0219_),
    .Q(\daisychain[91] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2404_ (.RESET_B(net398),
    .D(_0220_),
    .Q(\daisychain[92] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2405_ (.RESET_B(net396),
    .D(_0221_),
    .Q(\daisychain[93] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2406_ (.RESET_B(net394),
    .D(_0222_),
    .Q(\daisychain[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2407_ (.RESET_B(net392),
    .D(_0223_),
    .Q(\daisychain[95] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2408_ (.RESET_B(net390),
    .D(_0224_),
    .Q(\daisychain[96] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2409_ (.RESET_B(net388),
    .D(_0225_),
    .Q(\daisychain[97] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2410_ (.RESET_B(net386),
    .D(_0226_),
    .Q(\daisychain[98] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2411_ (.RESET_B(net384),
    .D(_0227_),
    .Q(\daisychain[99] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2412_ (.RESET_B(net382),
    .D(_0228_),
    .Q(\daisychain[100] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2413_ (.RESET_B(net380),
    .D(_0229_),
    .Q(\daisychain[101] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2414_ (.RESET_B(net378),
    .D(_0230_),
    .Q(\daisychain[102] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2415_ (.RESET_B(net376),
    .D(_0231_),
    .Q(\daisychain[103] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2416_ (.RESET_B(net374),
    .D(_0232_),
    .Q(\daisychain[104] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2417_ (.RESET_B(net372),
    .D(_0233_),
    .Q(\daisychain[105] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2418_ (.RESET_B(net370),
    .D(_0234_),
    .Q(\daisychain[106] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2419_ (.RESET_B(net368),
    .D(_0235_),
    .Q(\daisychain[107] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2420_ (.RESET_B(net366),
    .D(_0236_),
    .Q(\daisychain[108] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2421_ (.RESET_B(net364),
    .D(_0237_),
    .Q(\daisychain[109] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2422_ (.RESET_B(net362),
    .D(_0238_),
    .Q(\daisychain[110] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2423_ (.RESET_B(net360),
    .D(_0239_),
    .Q(\daisychain[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2424_ (.RESET_B(net358),
    .D(_0240_),
    .Q(\daisychain[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2425_ (.RESET_B(net356),
    .D(_0241_),
    .Q(\daisychain[113] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2426_ (.RESET_B(net354),
    .D(_0242_),
    .Q(\daisychain[114] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2427_ (.RESET_B(net352),
    .D(_0243_),
    .Q(\daisychain[115] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2428_ (.RESET_B(net350),
    .D(_0244_),
    .Q(\daisychain[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2429_ (.RESET_B(net348),
    .D(_0245_),
    .Q(\daisychain[117] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2430_ (.RESET_B(net346),
    .D(_0246_),
    .Q(\daisychain[118] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2431_ (.RESET_B(net344),
    .D(_0247_),
    .Q(\daisychain[119] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2432_ (.RESET_B(net342),
    .D(_0248_),
    .Q(\daisychain[120] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2433_ (.RESET_B(net340),
    .D(_0249_),
    .Q(\daisychain[121] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2434_ (.RESET_B(net338),
    .D(_0250_),
    .Q(\daisychain[122] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2435_ (.RESET_B(net336),
    .D(_0251_),
    .Q(\daisychain[123] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2436_ (.RESET_B(net334),
    .D(_0252_),
    .Q(\daisychain[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2437_ (.RESET_B(net332),
    .D(_0253_),
    .Q(\daisychain[125] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2438_ (.RESET_B(net330),
    .D(_0254_),
    .Q(\daisychain[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2439_ (.RESET_B(net328),
    .D(_0255_),
    .Q(\daisychain[127] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2440_ (.RESET_B(net326),
    .D(_0256_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2441_ (.RESET_B(net323),
    .D(_0257_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2442_ (.RESET_B(net319),
    .D(_0258_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2443_ (.RESET_B(net315),
    .D(_0259_),
    .Q(\state[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2444_ (.RESET_B(net311),
    .D(_0260_),
    .Q(\state[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2445_ (.RESET_B(net307),
    .D(_0261_),
    .Q(\state[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2446_ (.RESET_B(net303),
    .D(_0262_),
    .Q(\state[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2447_ (.RESET_B(net299),
    .D(_0263_),
    .Q(\state[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2448_ (.RESET_B(net295),
    .D(_0264_),
    .Q(\state[8] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2449_ (.RESET_B(net291),
    .D(_0265_),
    .Q(\state[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2450_ (.RESET_B(net287),
    .D(_0266_),
    .Q(\state[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2451_ (.RESET_B(net283),
    .D(_0267_),
    .Q(\state[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2452_ (.RESET_B(net279),
    .D(_0268_),
    .Q(\state[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2453_ (.RESET_B(net275),
    .D(_0269_),
    .Q(\state[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2454_ (.RESET_B(net271),
    .D(_0270_),
    .Q(\state[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2455_ (.RESET_B(net267),
    .D(_0271_),
    .Q(\state[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2456_ (.RESET_B(net263),
    .D(_0272_),
    .Q(\state[16] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2457_ (.RESET_B(net259),
    .D(_0273_),
    .Q(\state[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2458_ (.RESET_B(net255),
    .D(_0274_),
    .Q(\state[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2459_ (.RESET_B(net251),
    .D(_0275_),
    .Q(\state[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2460_ (.RESET_B(net247),
    .D(_0276_),
    .Q(\state[20] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2461_ (.RESET_B(net243),
    .D(_0277_),
    .Q(\state[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2462_ (.RESET_B(net239),
    .D(_0278_),
    .Q(\state[22] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2463_ (.RESET_B(net235),
    .D(_0279_),
    .Q(\state[23] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2464_ (.RESET_B(net231),
    .D(_0280_),
    .Q(\state[24] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2465_ (.RESET_B(net227),
    .D(_0281_),
    .Q(\state[25] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2466_ (.RESET_B(net223),
    .D(_0282_),
    .Q(\state[26] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2467_ (.RESET_B(net219),
    .D(_0283_),
    .Q(\state[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2468_ (.RESET_B(net215),
    .D(_0284_),
    .Q(\state[28] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2469_ (.RESET_B(net211),
    .D(_0285_),
    .Q(\state[29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2470_ (.RESET_B(net207),
    .D(_0286_),
    .Q(\state[30] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2471_ (.RESET_B(net203),
    .D(_0287_),
    .Q(\state[31] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2472_ (.RESET_B(net),
    .D(_0288_),
    .Q(\state[32] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2473_ (.RESET_B(net451),
    .D(_0289_),
    .Q(\state[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2474_ (.RESET_B(net447),
    .D(_0290_),
    .Q(\state[34] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2475_ (.RESET_B(net443),
    .D(_0291_),
    .Q(\state[35] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2476_ (.RESET_B(net439),
    .D(_0292_),
    .Q(\state[36] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2477_ (.RESET_B(net435),
    .D(_0293_),
    .Q(\state[37] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2478_ (.RESET_B(net431),
    .D(_0294_),
    .Q(\state[38] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2479_ (.RESET_B(net427),
    .D(_0295_),
    .Q(\state[39] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2480_ (.RESET_B(net423),
    .D(_0296_),
    .Q(\state[40] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2481_ (.RESET_B(net419),
    .D(_0297_),
    .Q(\state[41] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2482_ (.RESET_B(net415),
    .D(_0298_),
    .Q(\state[42] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2483_ (.RESET_B(net411),
    .D(_0299_),
    .Q(\state[43] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2484_ (.RESET_B(net407),
    .D(_0300_),
    .Q(\state[44] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2485_ (.RESET_B(net403),
    .D(_0301_),
    .Q(\state[45] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2486_ (.RESET_B(net399),
    .D(_0302_),
    .Q(\state[46] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2487_ (.RESET_B(net395),
    .D(_0303_),
    .Q(\state[47] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2488_ (.RESET_B(net391),
    .D(_0304_),
    .Q(\state[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2489_ (.RESET_B(net387),
    .D(_0305_),
    .Q(\state[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2490_ (.RESET_B(net383),
    .D(_0306_),
    .Q(\state[50] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2491_ (.RESET_B(net379),
    .D(_0307_),
    .Q(\state[51] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2492_ (.RESET_B(net375),
    .D(_0308_),
    .Q(\state[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2493_ (.RESET_B(net371),
    .D(_0309_),
    .Q(\state[53] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2494_ (.RESET_B(net367),
    .D(_0310_),
    .Q(\state[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2495_ (.RESET_B(net363),
    .D(_0311_),
    .Q(\state[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2496_ (.RESET_B(net359),
    .D(_0312_),
    .Q(\state[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2497_ (.RESET_B(net355),
    .D(_0313_),
    .Q(\state[57] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2498_ (.RESET_B(net351),
    .D(_0314_),
    .Q(\state[58] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2499_ (.RESET_B(net347),
    .D(_0315_),
    .Q(\state[59] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2500_ (.RESET_B(net343),
    .D(_0316_),
    .Q(\state[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2501_ (.RESET_B(net339),
    .D(_0317_),
    .Q(\state[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2502_ (.RESET_B(net335),
    .D(_0318_),
    .Q(\state[62] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2503_ (.RESET_B(net331),
    .D(_0319_),
    .Q(\state[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2504_ (.RESET_B(net327),
    .D(_0320_),
    .Q(\state[64] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2505_ (.RESET_B(net321),
    .D(_0321_),
    .Q(\state[65] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2506_ (.RESET_B(net313),
    .D(_0322_),
    .Q(\state[66] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2507_ (.RESET_B(net305),
    .D(_0323_),
    .Q(\state[67] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2508_ (.RESET_B(net297),
    .D(_0324_),
    .Q(\state[68] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2509_ (.RESET_B(net289),
    .D(_0325_),
    .Q(\state[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2510_ (.RESET_B(net281),
    .D(_0326_),
    .Q(\state[70] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2511_ (.RESET_B(net273),
    .D(_0327_),
    .Q(\state[71] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2512_ (.RESET_B(net265),
    .D(_0328_),
    .Q(\state[72] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2513_ (.RESET_B(net257),
    .D(_0329_),
    .Q(\state[73] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2514_ (.RESET_B(net249),
    .D(_0330_),
    .Q(\state[74] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2515_ (.RESET_B(net241),
    .D(_0331_),
    .Q(\state[75] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2516_ (.RESET_B(net233),
    .D(_0332_),
    .Q(\state[76] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2517_ (.RESET_B(net225),
    .D(_0333_),
    .Q(\state[77] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2518_ (.RESET_B(net217),
    .D(_0334_),
    .Q(\state[78] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2519_ (.RESET_B(net209),
    .D(_0335_),
    .Q(\state[79] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2520_ (.RESET_B(net201),
    .D(_0336_),
    .Q(\state[80] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2521_ (.RESET_B(net449),
    .D(_0337_),
    .Q(\state[81] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2522_ (.RESET_B(net441),
    .D(_0338_),
    .Q(\state[82] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2523_ (.RESET_B(net433),
    .D(_0339_),
    .Q(\state[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2524_ (.RESET_B(net425),
    .D(_0340_),
    .Q(\state[84] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2525_ (.RESET_B(net417),
    .D(_0341_),
    .Q(\state[85] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2526_ (.RESET_B(net409),
    .D(_0342_),
    .Q(\state[86] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2527_ (.RESET_B(net401),
    .D(_0343_),
    .Q(\state[87] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2528_ (.RESET_B(net393),
    .D(_0344_),
    .Q(\state[88] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2529_ (.RESET_B(net385),
    .D(_0345_),
    .Q(\state[89] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2530_ (.RESET_B(net377),
    .D(_0346_),
    .Q(\state[90] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2531_ (.RESET_B(net369),
    .D(_0347_),
    .Q(\state[91] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2532_ (.RESET_B(net361),
    .D(_0348_),
    .Q(\state[92] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2533_ (.RESET_B(net353),
    .D(_0349_),
    .Q(\state[93] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2534_ (.RESET_B(net345),
    .D(_0350_),
    .Q(\state[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2535_ (.RESET_B(net337),
    .D(_0351_),
    .Q(\state[95] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2536_ (.RESET_B(net329),
    .D(_0352_),
    .Q(\state[96] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2537_ (.RESET_B(net317),
    .D(_0353_),
    .Q(\state[97] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2538_ (.RESET_B(net301),
    .D(_0354_),
    .Q(\state[98] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2539_ (.RESET_B(net285),
    .D(_0355_),
    .Q(\state[99] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2540_ (.RESET_B(net269),
    .D(_0356_),
    .Q(\state[100] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2541_ (.RESET_B(net253),
    .D(_0357_),
    .Q(\state[101] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2542_ (.RESET_B(net237),
    .D(_0358_),
    .Q(\state[102] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2543_ (.RESET_B(net221),
    .D(_0359_),
    .Q(\state[103] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2544_ (.RESET_B(net205),
    .D(_0360_),
    .Q(\state[104] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2545_ (.RESET_B(net445),
    .D(_0361_),
    .Q(\state[105] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2546_ (.RESET_B(net429),
    .D(_0362_),
    .Q(\state[106] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2547_ (.RESET_B(net413),
    .D(_0363_),
    .Q(\state[107] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2548_ (.RESET_B(net397),
    .D(_0364_),
    .Q(\state[108] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2549_ (.RESET_B(net381),
    .D(_0365_),
    .Q(\state[109] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2550_ (.RESET_B(net365),
    .D(_0366_),
    .Q(\state[110] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2551_ (.RESET_B(net349),
    .D(_0367_),
    .Q(\state[111] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2552_ (.RESET_B(net333),
    .D(_0368_),
    .Q(\state[112] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2553_ (.RESET_B(net309),
    .D(_0369_),
    .Q(\state[113] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2554_ (.RESET_B(net277),
    .D(_0370_),
    .Q(\state[114] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2555_ (.RESET_B(net245),
    .D(_0371_),
    .Q(\state[115] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2556_ (.RESET_B(net213),
    .D(_0372_),
    .Q(\state[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2557_ (.RESET_B(net437),
    .D(_0373_),
    .Q(\state[117] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2558_ (.RESET_B(net405),
    .D(_0374_),
    .Q(\state[118] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2559_ (.RESET_B(net373),
    .D(_0375_),
    .Q(\state[119] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2560_ (.RESET_B(net341),
    .D(_0376_),
    .Q(\state[120] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2561_ (.RESET_B(net293),
    .D(_0377_),
    .Q(\state[121] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2562_ (.RESET_B(net229),
    .D(_0378_),
    .Q(\state[122] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2563_ (.RESET_B(net421),
    .D(_0379_),
    .Q(\state[123] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2564_ (.RESET_B(net357),
    .D(_0380_),
    .Q(\state[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2565_ (.RESET_B(net261),
    .D(_0381_),
    .Q(\state[125] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2566_ (.RESET_B(net389),
    .D(_0382_),
    .Q(\state[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2567_ (.RESET_B(net453),
    .D(_0383_),
    .Q(\state[127] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_tiehi _2375__201 (.L_HI(net200));
 sg13g2_tiehi _2520__202 (.L_HI(net201));
 sg13g2_tiehi _2374__203 (.L_HI(net202));
 sg13g2_tiehi _2471__204 (.L_HI(net203));
 sg13g2_tiehi _2373__205 (.L_HI(net204));
 sg13g2_tiehi _2544__206 (.L_HI(net205));
 sg13g2_tiehi _2372__207 (.L_HI(net206));
 sg13g2_tiehi _2470__208 (.L_HI(net207));
 sg13g2_tiehi _2371__209 (.L_HI(net208));
 sg13g2_tiehi _2519__210 (.L_HI(net209));
 sg13g2_tiehi _2370__211 (.L_HI(net210));
 sg13g2_tiehi _2469__212 (.L_HI(net211));
 sg13g2_tiehi _2369__213 (.L_HI(net212));
 sg13g2_tiehi _2556__214 (.L_HI(net213));
 sg13g2_tiehi _2368__215 (.L_HI(net214));
 sg13g2_tiehi _2468__216 (.L_HI(net215));
 sg13g2_tiehi _2367__217 (.L_HI(net216));
 sg13g2_tiehi _2518__218 (.L_HI(net217));
 sg13g2_tiehi _2366__219 (.L_HI(net218));
 sg13g2_tiehi _2467__220 (.L_HI(net219));
 sg13g2_tiehi _2365__221 (.L_HI(net220));
 sg13g2_tiehi _2543__222 (.L_HI(net221));
 sg13g2_tiehi _2364__223 (.L_HI(net222));
 sg13g2_tiehi _2466__224 (.L_HI(net223));
 sg13g2_tiehi _2363__225 (.L_HI(net224));
 sg13g2_tiehi _2517__226 (.L_HI(net225));
 sg13g2_tiehi _2362__227 (.L_HI(net226));
 sg13g2_tiehi _2465__228 (.L_HI(net227));
 sg13g2_tiehi _2361__229 (.L_HI(net228));
 sg13g2_tiehi _2562__230 (.L_HI(net229));
 sg13g2_tiehi _2360__231 (.L_HI(net230));
 sg13g2_tiehi _2464__232 (.L_HI(net231));
 sg13g2_tiehi _2359__233 (.L_HI(net232));
 sg13g2_tiehi _2516__234 (.L_HI(net233));
 sg13g2_tiehi _2358__235 (.L_HI(net234));
 sg13g2_tiehi _2463__236 (.L_HI(net235));
 sg13g2_tiehi _2357__237 (.L_HI(net236));
 sg13g2_tiehi _2542__238 (.L_HI(net237));
 sg13g2_tiehi _2356__239 (.L_HI(net238));
 sg13g2_tiehi _2462__240 (.L_HI(net239));
 sg13g2_tiehi _2355__241 (.L_HI(net240));
 sg13g2_tiehi _2515__242 (.L_HI(net241));
 sg13g2_tiehi _2354__243 (.L_HI(net242));
 sg13g2_tiehi _2461__244 (.L_HI(net243));
 sg13g2_tiehi _2353__245 (.L_HI(net244));
 sg13g2_tiehi _2555__246 (.L_HI(net245));
 sg13g2_tiehi _2352__247 (.L_HI(net246));
 sg13g2_tiehi _2460__248 (.L_HI(net247));
 sg13g2_tiehi _2351__249 (.L_HI(net248));
 sg13g2_tiehi _2514__250 (.L_HI(net249));
 sg13g2_tiehi _2350__251 (.L_HI(net250));
 sg13g2_tiehi _2459__252 (.L_HI(net251));
 sg13g2_tiehi _2349__253 (.L_HI(net252));
 sg13g2_tiehi _2541__254 (.L_HI(net253));
 sg13g2_tiehi _2348__255 (.L_HI(net254));
 sg13g2_tiehi _2458__256 (.L_HI(net255));
 sg13g2_tiehi _2347__257 (.L_HI(net256));
 sg13g2_tiehi _2513__258 (.L_HI(net257));
 sg13g2_tiehi _2346__259 (.L_HI(net258));
 sg13g2_tiehi _2457__260 (.L_HI(net259));
 sg13g2_tiehi _2345__261 (.L_HI(net260));
 sg13g2_tiehi _2565__262 (.L_HI(net261));
 sg13g2_tiehi _2344__263 (.L_HI(net262));
 sg13g2_tiehi _2456__264 (.L_HI(net263));
 sg13g2_tiehi _2343__265 (.L_HI(net264));
 sg13g2_tiehi _2512__266 (.L_HI(net265));
 sg13g2_tiehi _2342__267 (.L_HI(net266));
 sg13g2_tiehi _2455__268 (.L_HI(net267));
 sg13g2_tiehi _2341__269 (.L_HI(net268));
 sg13g2_tiehi _2540__270 (.L_HI(net269));
 sg13g2_tiehi _2340__271 (.L_HI(net270));
 sg13g2_tiehi _2454__272 (.L_HI(net271));
 sg13g2_tiehi _2339__273 (.L_HI(net272));
 sg13g2_tiehi _2511__274 (.L_HI(net273));
 sg13g2_tiehi _2338__275 (.L_HI(net274));
 sg13g2_tiehi _2453__276 (.L_HI(net275));
 sg13g2_tiehi _2337__277 (.L_HI(net276));
 sg13g2_tiehi _2554__278 (.L_HI(net277));
 sg13g2_tiehi _2336__279 (.L_HI(net278));
 sg13g2_tiehi _2452__280 (.L_HI(net279));
 sg13g2_tiehi _2335__281 (.L_HI(net280));
 sg13g2_tiehi _2510__282 (.L_HI(net281));
 sg13g2_tiehi _2334__283 (.L_HI(net282));
 sg13g2_tiehi _2451__284 (.L_HI(net283));
 sg13g2_tiehi _2333__285 (.L_HI(net284));
 sg13g2_tiehi _2539__286 (.L_HI(net285));
 sg13g2_tiehi _2332__287 (.L_HI(net286));
 sg13g2_tiehi _2450__288 (.L_HI(net287));
 sg13g2_tiehi _2331__289 (.L_HI(net288));
 sg13g2_tiehi _2509__290 (.L_HI(net289));
 sg13g2_tiehi _2330__291 (.L_HI(net290));
 sg13g2_tiehi _2449__292 (.L_HI(net291));
 sg13g2_tiehi _2329__293 (.L_HI(net292));
 sg13g2_tiehi _2561__294 (.L_HI(net293));
 sg13g2_tiehi _2328__295 (.L_HI(net294));
 sg13g2_tiehi _2448__296 (.L_HI(net295));
 sg13g2_tiehi _2327__297 (.L_HI(net296));
 sg13g2_tiehi _2508__298 (.L_HI(net297));
 sg13g2_tiehi _2326__299 (.L_HI(net298));
 sg13g2_tiehi _2447__300 (.L_HI(net299));
 sg13g2_tiehi _2325__301 (.L_HI(net300));
 sg13g2_tiehi _2538__302 (.L_HI(net301));
 sg13g2_tiehi _2324__303 (.L_HI(net302));
 sg13g2_tiehi _2446__304 (.L_HI(net303));
 sg13g2_tiehi _2323__305 (.L_HI(net304));
 sg13g2_tiehi _2507__306 (.L_HI(net305));
 sg13g2_tiehi _2322__307 (.L_HI(net306));
 sg13g2_tiehi _2445__308 (.L_HI(net307));
 sg13g2_tiehi _2321__309 (.L_HI(net308));
 sg13g2_tiehi _2553__310 (.L_HI(net309));
 sg13g2_tiehi _2320__311 (.L_HI(net310));
 sg13g2_tiehi _2444__312 (.L_HI(net311));
 sg13g2_tiehi _2319__313 (.L_HI(net312));
 sg13g2_tiehi _2506__314 (.L_HI(net313));
 sg13g2_tiehi _2318__315 (.L_HI(net314));
 sg13g2_tiehi _2443__316 (.L_HI(net315));
 sg13g2_tiehi _2317__317 (.L_HI(net316));
 sg13g2_tiehi _2537__318 (.L_HI(net317));
 sg13g2_tiehi _2316__319 (.L_HI(net318));
 sg13g2_tiehi _2442__320 (.L_HI(net319));
 sg13g2_tiehi _2315__321 (.L_HI(net320));
 sg13g2_tiehi _2505__322 (.L_HI(net321));
 sg13g2_tiehi _2314__323 (.L_HI(net322));
 sg13g2_tiehi _2441__324 (.L_HI(net323));
 sg13g2_tiehi _2313__325 (.L_HI(net324));
 sg13g2_tiehi _2312__326 (.L_HI(net325));
 sg13g2_tiehi _2440__327 (.L_HI(net326));
 sg13g2_tiehi _2504__328 (.L_HI(net327));
 sg13g2_tiehi _2439__329 (.L_HI(net328));
 sg13g2_tiehi _2536__330 (.L_HI(net329));
 sg13g2_tiehi _2438__331 (.L_HI(net330));
 sg13g2_tiehi _2503__332 (.L_HI(net331));
 sg13g2_tiehi _2437__333 (.L_HI(net332));
 sg13g2_tiehi _2552__334 (.L_HI(net333));
 sg13g2_tiehi _2436__335 (.L_HI(net334));
 sg13g2_tiehi _2502__336 (.L_HI(net335));
 sg13g2_tiehi _2435__337 (.L_HI(net336));
 sg13g2_tiehi _2535__338 (.L_HI(net337));
 sg13g2_tiehi _2434__339 (.L_HI(net338));
 sg13g2_tiehi _2501__340 (.L_HI(net339));
 sg13g2_tiehi _2433__341 (.L_HI(net340));
 sg13g2_tiehi _2560__342 (.L_HI(net341));
 sg13g2_tiehi _2432__343 (.L_HI(net342));
 sg13g2_tiehi _2500__344 (.L_HI(net343));
 sg13g2_tiehi _2431__345 (.L_HI(net344));
 sg13g2_tiehi _2534__346 (.L_HI(net345));
 sg13g2_tiehi _2430__347 (.L_HI(net346));
 sg13g2_tiehi _2499__348 (.L_HI(net347));
 sg13g2_tiehi _2429__349 (.L_HI(net348));
 sg13g2_tiehi _2551__350 (.L_HI(net349));
 sg13g2_tiehi _2428__351 (.L_HI(net350));
 sg13g2_tiehi _2498__352 (.L_HI(net351));
 sg13g2_tiehi _2427__353 (.L_HI(net352));
 sg13g2_tiehi _2533__354 (.L_HI(net353));
 sg13g2_tiehi _2426__355 (.L_HI(net354));
 sg13g2_tiehi _2497__356 (.L_HI(net355));
 sg13g2_tiehi _2425__357 (.L_HI(net356));
 sg13g2_tiehi _2564__358 (.L_HI(net357));
 sg13g2_tiehi _2424__359 (.L_HI(net358));
 sg13g2_tiehi _2496__360 (.L_HI(net359));
 sg13g2_tiehi _2423__361 (.L_HI(net360));
 sg13g2_tiehi _2532__362 (.L_HI(net361));
 sg13g2_tiehi _2422__363 (.L_HI(net362));
 sg13g2_tiehi _2495__364 (.L_HI(net363));
 sg13g2_tiehi _2421__365 (.L_HI(net364));
 sg13g2_tiehi _2550__366 (.L_HI(net365));
 sg13g2_tiehi _2420__367 (.L_HI(net366));
 sg13g2_tiehi _2494__368 (.L_HI(net367));
 sg13g2_tiehi _2419__369 (.L_HI(net368));
 sg13g2_tiehi _2531__370 (.L_HI(net369));
 sg13g2_tiehi _2418__371 (.L_HI(net370));
 sg13g2_tiehi _2493__372 (.L_HI(net371));
 sg13g2_tiehi _2417__373 (.L_HI(net372));
 sg13g2_tiehi _2559__374 (.L_HI(net373));
 sg13g2_tiehi _2416__375 (.L_HI(net374));
 sg13g2_tiehi _2492__376 (.L_HI(net375));
 sg13g2_tiehi _2415__377 (.L_HI(net376));
 sg13g2_tiehi _2530__378 (.L_HI(net377));
 sg13g2_tiehi _2414__379 (.L_HI(net378));
 sg13g2_tiehi _2491__380 (.L_HI(net379));
 sg13g2_tiehi _2413__381 (.L_HI(net380));
 sg13g2_tiehi _2549__382 (.L_HI(net381));
 sg13g2_tiehi _2412__383 (.L_HI(net382));
 sg13g2_tiehi _2490__384 (.L_HI(net383));
 sg13g2_tiehi _2411__385 (.L_HI(net384));
 sg13g2_tiehi _2529__386 (.L_HI(net385));
 sg13g2_tiehi _2410__387 (.L_HI(net386));
 sg13g2_tiehi _2489__388 (.L_HI(net387));
 sg13g2_tiehi _2409__389 (.L_HI(net388));
 sg13g2_tiehi _2566__390 (.L_HI(net389));
 sg13g2_tiehi _2408__391 (.L_HI(net390));
 sg13g2_tiehi _2488__392 (.L_HI(net391));
 sg13g2_tiehi _2407__393 (.L_HI(net392));
 sg13g2_tiehi _2528__394 (.L_HI(net393));
 sg13g2_tiehi _2406__395 (.L_HI(net394));
 sg13g2_tiehi _2487__396 (.L_HI(net395));
 sg13g2_tiehi _2405__397 (.L_HI(net396));
 sg13g2_tiehi _2548__398 (.L_HI(net397));
 sg13g2_tiehi _2404__399 (.L_HI(net398));
 sg13g2_tiehi _2486__400 (.L_HI(net399));
 sg13g2_tiehi _2403__401 (.L_HI(net400));
 sg13g2_tiehi _2527__402 (.L_HI(net401));
 sg13g2_tiehi _2402__403 (.L_HI(net402));
 sg13g2_tiehi _2485__404 (.L_HI(net403));
 sg13g2_tiehi _2401__405 (.L_HI(net404));
 sg13g2_tiehi _2558__406 (.L_HI(net405));
 sg13g2_tiehi _2400__407 (.L_HI(net406));
 sg13g2_tiehi _2484__408 (.L_HI(net407));
 sg13g2_tiehi _2399__409 (.L_HI(net408));
 sg13g2_tiehi _2526__410 (.L_HI(net409));
 sg13g2_tiehi _2398__411 (.L_HI(net410));
 sg13g2_tiehi _2483__412 (.L_HI(net411));
 sg13g2_tiehi _2397__413 (.L_HI(net412));
 sg13g2_tiehi _2547__414 (.L_HI(net413));
 sg13g2_tiehi _2396__415 (.L_HI(net414));
 sg13g2_tiehi _2482__416 (.L_HI(net415));
 sg13g2_tiehi _2395__417 (.L_HI(net416));
 sg13g2_tiehi _2525__418 (.L_HI(net417));
 sg13g2_tiehi _2394__419 (.L_HI(net418));
 sg13g2_tiehi _2481__420 (.L_HI(net419));
 sg13g2_tiehi _2393__421 (.L_HI(net420));
 sg13g2_tiehi _2563__422 (.L_HI(net421));
 sg13g2_tiehi _2392__423 (.L_HI(net422));
 sg13g2_tiehi _2480__424 (.L_HI(net423));
 sg13g2_tiehi _2391__425 (.L_HI(net424));
 sg13g2_tiehi _2524__426 (.L_HI(net425));
 sg13g2_tiehi _2390__427 (.L_HI(net426));
 sg13g2_tiehi _2479__428 (.L_HI(net427));
 sg13g2_tiehi _2389__429 (.L_HI(net428));
 sg13g2_tiehi _2546__430 (.L_HI(net429));
 sg13g2_tiehi _2388__431 (.L_HI(net430));
 sg13g2_tiehi _2478__432 (.L_HI(net431));
 sg13g2_tiehi _2387__433 (.L_HI(net432));
 sg13g2_tiehi _2523__434 (.L_HI(net433));
 sg13g2_tiehi _2386__435 (.L_HI(net434));
 sg13g2_tiehi _2477__436 (.L_HI(net435));
 sg13g2_tiehi _2385__437 (.L_HI(net436));
 sg13g2_tiehi _2557__438 (.L_HI(net437));
 sg13g2_tiehi _2384__439 (.L_HI(net438));
 sg13g2_tiehi _2476__440 (.L_HI(net439));
 sg13g2_tiehi _2383__441 (.L_HI(net440));
 sg13g2_tiehi _2522__442 (.L_HI(net441));
 sg13g2_tiehi _2382__443 (.L_HI(net442));
 sg13g2_tiehi _2475__444 (.L_HI(net443));
 sg13g2_tiehi _2381__445 (.L_HI(net444));
 sg13g2_tiehi _2545__446 (.L_HI(net445));
 sg13g2_tiehi _2380__447 (.L_HI(net446));
 sg13g2_tiehi _2474__448 (.L_HI(net447));
 sg13g2_tiehi _2379__449 (.L_HI(net448));
 sg13g2_tiehi _2521__450 (.L_HI(net449));
 sg13g2_tiehi _2378__451 (.L_HI(net450));
 sg13g2_tiehi _2473__452 (.L_HI(net451));
 sg13g2_tiehi _2377__453 (.L_HI(net452));
 sg13g2_tiehi _2567__454 (.L_HI(net453));
 sg13g2_tiehi _2376__455 (.L_HI(net454));
 sg13g2_tiehi heichips25_pudding (.L_HI(net455));
 sg13g2_tiehi heichips25_pudding_456 (.L_HI(net456));
 sg13g2_tiehi heichips25_pudding_457 (.L_HI(net457));
 sg13g2_tiehi heichips25_pudding_458 (.L_HI(net458));
 sg13g2_tiehi heichips25_pudding_459 (.L_HI(net459));
 sg13g2_tiehi heichips25_pudding_460 (.L_HI(net460));
 sg13g2_tiehi heichips25_pudding_461 (.L_HI(net461));
 sg13g2_tiehi heichips25_pudding_462 (.L_HI(net462));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _2832_ (.A(\state[120] ),
    .X(net7));
 sg13g2_buf_1 _2833_ (.A(\state[121] ),
    .X(net8));
 sg13g2_buf_1 _2834_ (.A(\state[122] ),
    .X(net9));
 sg13g2_buf_1 _2835_ (.A(\state[123] ),
    .X(net10));
 sg13g2_buf_1 _2836_ (.A(\state[124] ),
    .X(net11));
 sg13g2_buf_1 _2837_ (.A(\state[125] ),
    .X(net12));
 sg13g2_buf_1 _2838_ (.A(\state[126] ),
    .X(net13));
 sg13g2_buf_1 _2839_ (.A(\state[127] ),
    .X(net14));
 sg13g2_buf_1 _2840_ (.A(\daisychain[120] ),
    .X(net15));
 sg13g2_buf_1 _2841_ (.A(\daisychain[121] ),
    .X(net16));
 sg13g2_buf_1 _2842_ (.A(\daisychain[122] ),
    .X(net17));
 sg13g2_buf_1 _2843_ (.A(\daisychain[123] ),
    .X(net18));
 sg13g2_buf_1 _2844_ (.A(\daisychain[124] ),
    .X(net19));
 sg13g2_buf_1 _2845_ (.A(\daisychain[125] ),
    .X(net20));
 sg13g2_buf_1 _2846_ (.A(\daisychain[126] ),
    .X(net21));
 sg13g2_buf_1 _2847_ (.A(\daisychain[127] ),
    .X(net22));
 dac128module dac (.IOUT(dacout),
    .EN({\digitalen.g[3].u.OUTP ,
    \digitalen.g[2].u.OUTP ,
    \digitalen.g[1].u.OUTP ,
    \digitalen.g[0].u.OUTP }),
    .ENB({\digitalen.g[3].u.OUTN ,
    \digitalen.g[2].u.OUTN ,
    \digitalen.g[1].u.OUTN ,
    \digitalen.g[0].u.OUTN }),
    .ON({\state[127] ,
    \state[126] ,
    \state[125] ,
    \state[124] ,
    \state[123] ,
    \state[122] ,
    \state[121] ,
    \state[120] ,
    \state[119] ,
    \state[118] ,
    \state[117] ,
    \state[116] ,
    \state[115] ,
    \state[114] ,
    \state[113] ,
    \state[112] ,
    \state[111] ,
    \state[110] ,
    \state[109] ,
    \state[108] ,
    \state[107] ,
    \state[106] ,
    \state[105] ,
    \state[104] ,
    \state[103] ,
    \state[102] ,
    \state[101] ,
    \state[100] ,
    \state[99] ,
    \state[98] ,
    \state[97] ,
    \state[96] ,
    \state[95] ,
    \state[94] ,
    \state[93] ,
    \state[92] ,
    \state[91] ,
    \state[90] ,
    \state[89] ,
    \state[88] ,
    \state[87] ,
    \state[86] ,
    \state[85] ,
    \state[84] ,
    \state[83] ,
    \state[82] ,
    \state[81] ,
    \state[80] ,
    \state[79] ,
    \state[78] ,
    \state[77] ,
    \state[76] ,
    \state[75] ,
    \state[74] ,
    \state[73] ,
    \state[72] ,
    \state[71] ,
    \state[70] ,
    \state[69] ,
    \state[68] ,
    \state[67] ,
    \state[66] ,
    \state[65] ,
    \state[64] ,
    \state[63] ,
    \state[62] ,
    \state[61] ,
    \state[60] ,
    \state[59] ,
    \state[58] ,
    \state[57] ,
    \state[56] ,
    \state[55] ,
    \state[54] ,
    \state[53] ,
    \state[52] ,
    \state[51] ,
    \state[50] ,
    \state[49] ,
    \state[48] ,
    \state[47] ,
    \state[46] ,
    \state[45] ,
    \state[44] ,
    \state[43] ,
    \state[42] ,
    \state[41] ,
    \state[40] ,
    \state[39] ,
    \state[38] ,
    \state[37] ,
    \state[36] ,
    \state[35] ,
    \state[34] ,
    \state[33] ,
    \state[32] ,
    \state[31] ,
    \state[30] ,
    \state[29] ,
    \state[28] ,
    \state[27] ,
    \state[26] ,
    \state[25] ,
    \state[24] ,
    \state[23] ,
    \state[22] ,
    \state[21] ,
    \state[20] ,
    \state[19] ,
    \state[18] ,
    \state[17] ,
    \state[16] ,
    \state[15] ,
    \state[14] ,
    \state[13] ,
    \state[12] ,
    \state[11] ,
    \state[10] ,
    \state[9] ,
    \state[8] ,
    \state[7] ,
    \state[6] ,
    \state[5] ,
    \state[4] ,
    \state[3] ,
    \state[2] ,
    \state[1] ,
    \state[0] }),
    .ONB({_0030_,
    _0029_,
    _0028_,
    _0027_,
    _0026_,
    _0025_,
    _0024_,
    _0023_,
    _0021_,
    _0020_,
    _0019_,
    _0018_,
    _0017_,
    _0016_,
    _0015_,
    _0014_,
    _0013_,
    _0012_,
    _0010_,
    _0009_,
    _0008_,
    _0007_,
    _0006_,
    _0005_,
    _0004_,
    _0003_,
    _0002_,
    _0001_,
    _0126_,
    _0125_,
    _0124_,
    _0123_,
    _0122_,
    _0121_,
    _0120_,
    _0119_,
    _0118_,
    _0117_,
    _0115_,
    _0114_,
    _0113_,
    _0112_,
    _0111_,
    _0110_,
    _0109_,
    _0108_,
    _0107_,
    _0106_,
    _0104_,
    _0103_,
    _0102_,
    _0101_,
    _0100_,
    _0099_,
    _0098_,
    _0097_,
    _0096_,
    _0095_,
    _0093_,
    _0092_,
    _0091_,
    _0090_,
    _0089_,
    _0088_,
    _0087_,
    _0086_,
    _0085_,
    _0084_,
    _0082_,
    _0081_,
    _0080_,
    _0079_,
    _0078_,
    _0077_,
    _0076_,
    _0075_,
    _0074_,
    _0073_,
    _0071_,
    _0070_,
    _0069_,
    _0068_,
    _0067_,
    _0066_,
    _0065_,
    _0064_,
    _0063_,
    _0062_,
    _0060_,
    _0059_,
    _0058_,
    _0057_,
    _0056_,
    _0055_,
    _0054_,
    _0053_,
    _0052_,
    _0051_,
    _0049_,
    _0048_,
    _0047_,
    _0046_,
    _0045_,
    _0044_,
    _0043_,
    _0042_,
    _0041_,
    _0040_,
    _0038_,
    _0037_,
    _0036_,
    _0035_,
    _0034_,
    _0033_,
    _0032_,
    _0031_,
    _0022_,
    _0011_,
    _0127_,
    _0116_,
    _0105_,
    _0094_,
    _0083_,
    _0072_,
    _0061_,
    _0050_,
    _0039_,
    _0000_}),
    .VbiasP({\bias[1] ,
    \bias[0] }),
    .VcascP({\iref[1] ,
    \iref[0] }));
 sg13g2_inv_1 \digitalen.g[0].u.inv1  (.Y(\digitalen.g[0].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[0].u.inv2  (.Y(\digitalen.g[0].u.OUTP ),
    .A(\digitalen.g[0].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[1].u.inv1  (.Y(\digitalen.g[1].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[1].u.inv2  (.Y(\digitalen.g[1].u.OUTP ),
    .A(\digitalen.g[1].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[2].u.inv1  (.Y(\digitalen.g[2].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[2].u.inv2  (.Y(\digitalen.g[2].u.OUTP ),
    .A(\digitalen.g[2].u.OUTN ));
 sg13g2_inv_1 \digitalen.g[3].u.inv1  (.Y(\digitalen.g[3].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalen.g[3].u.inv2  (.Y(\digitalen.g[3].u.OUTP ),
    .A(\digitalen.g[3].u.OUTN ));
 analog_wires wires (.Iout(dacout),
    .i_in(i_in),
    .i_out(i_out),
    .VcascP({\iref[1] ,
    \iref[0] }));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]));
 sg13g2_buf_1 fanout23 (.A(net44),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net44),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(net44),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net29),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(net29),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(net29),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(net44),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net34),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net34),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net34),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net34),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net44),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net36),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net43),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net38),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net43),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net40),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net43),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net42),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(_0851_),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net47),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(net66),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(net66),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net52),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net52),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net52),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net66),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(net56),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net56),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(net66),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net58),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(net65),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net65),
    .X(net60));
 sg13g2_buf_1 fanout61 (.A(net64),
    .X(net61));
 sg13g2_buf_1 fanout62 (.A(net63),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(net64),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(net65),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(_0850_),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(net69),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(net69),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(net89),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net89),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(net75),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net75),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net75),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(net89),
    .X(net75));
 sg13g2_buf_1 fanout76 (.A(net79),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net78),
    .X(net77));
 sg13g2_buf_1 fanout78 (.A(net79),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net89),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net88),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_1 fanout83 (.A(net88),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(net88),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net88),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(_0847_),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(net98),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net94),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(net98),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(_0846_),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net102),
    .X(net99));
 sg13g2_buf_1 fanout100 (.A(net102),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(net106),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net106),
    .X(net104));
 sg13g2_buf_1 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net132),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net109),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_1 fanout109 (.A(net114),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net113),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(net132),
    .X(net114));
 sg13g2_buf_1 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net123),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(net121),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(net123),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(net132),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(net131),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net131),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net130),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(_0846_),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net154),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net154),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net140),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net140),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(net154),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net144),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net154),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(net153),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(net153),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(net153),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net153),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net5),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net158),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(net4),
    .X(net158));
 sg13g2_buf_1 fanout159 (.A(net162),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(net162),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_1 fanout162 (.A(net167),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net4),
    .X(net167));
 sg13g2_buf_1 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net176),
    .X(net169));
 sg13g2_buf_1 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_1 fanout171 (.A(net176),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net176),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net4),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net180),
    .X(net177));
 sg13g2_buf_1 fanout178 (.A(net180),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net199),
    .X(net180));
 sg13g2_buf_1 fanout181 (.A(net184),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net199),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net189),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(net189),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net189),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_1 fanout189 (.A(net199),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net198),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_1 fanout193 (.A(net198),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_1 fanout195 (.A(net198),
    .X(net195));
 sg13g2_buf_1 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_1 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net1),
    .X(net199));
 sg13g2_tiehi _2472__200 (.L_HI(net));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_16 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_15_clk));
 sg13g2_inv_8 clkload4 (.A(clknet_leaf_0_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_16_clk));
 sg13g2_inv_8 clkload6 (.A(clknet_leaf_17_clk));
 sg13g2_inv_16 clkload7 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_11_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_9_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_4 FILLER_0_567 ();
 sg13g2_fill_1 FILLER_0_576 ();
 sg13g2_fill_1 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_4 FILLER_0_631 ();
 sg13g2_fill_1 FILLER_0_635 ();
 sg13g2_decap_4 FILLER_0_651 ();
 sg13g2_fill_2 FILLER_0_655 ();
 sg13g2_decap_4 FILLER_0_675 ();
 sg13g2_fill_2 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_4 FILLER_0_724 ();
 sg13g2_fill_1 FILLER_0_728 ();
 sg13g2_fill_2 FILLER_0_784 ();
 sg13g2_fill_1 FILLER_0_786 ();
 sg13g2_fill_1 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_4 FILLER_1_546 ();
 sg13g2_fill_1 FILLER_1_550 ();
 sg13g2_fill_1 FILLER_1_664 ();
 sg13g2_decap_4 FILLER_1_692 ();
 sg13g2_fill_2 FILLER_1_775 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_fill_2 FILLER_1_821 ();
 sg13g2_fill_1 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_13 ();
 sg13g2_decap_4 FILLER_2_20 ();
 sg13g2_fill_1 FILLER_2_24 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_fill_2 FILLER_2_553 ();
 sg13g2_fill_1 FILLER_2_555 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_fill_1 FILLER_2_579 ();
 sg13g2_decap_8 FILLER_2_593 ();
 sg13g2_decap_4 FILLER_2_600 ();
 sg13g2_fill_2 FILLER_2_604 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_decap_8 FILLER_2_632 ();
 sg13g2_fill_2 FILLER_2_639 ();
 sg13g2_decap_8 FILLER_2_645 ();
 sg13g2_decap_4 FILLER_2_652 ();
 sg13g2_fill_1 FILLER_2_656 ();
 sg13g2_decap_8 FILLER_2_671 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_fill_1 FILLER_2_685 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_fill_2 FILLER_2_713 ();
 sg13g2_fill_1 FILLER_2_715 ();
 sg13g2_decap_8 FILLER_2_720 ();
 sg13g2_decap_8 FILLER_2_727 ();
 sg13g2_fill_1 FILLER_2_734 ();
 sg13g2_decap_8 FILLER_2_775 ();
 sg13g2_decap_8 FILLER_2_810 ();
 sg13g2_decap_4 FILLER_2_817 ();
 sg13g2_fill_2 FILLER_2_821 ();
 sg13g2_fill_2 FILLER_3_31 ();
 sg13g2_fill_1 FILLER_3_33 ();
 sg13g2_decap_4 FILLER_3_39 ();
 sg13g2_fill_2 FILLER_3_43 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_4 FILLER_3_511 ();
 sg13g2_fill_1 FILLER_3_515 ();
 sg13g2_fill_2 FILLER_3_526 ();
 sg13g2_fill_1 FILLER_3_528 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_4 FILLER_3_550 ();
 sg13g2_fill_2 FILLER_3_581 ();
 sg13g2_fill_1 FILLER_3_583 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_fill_2 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_642 ();
 sg13g2_decap_4 FILLER_3_649 ();
 sg13g2_fill_1 FILLER_3_657 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_687 ();
 sg13g2_decap_8 FILLER_3_694 ();
 sg13g2_decap_8 FILLER_3_701 ();
 sg13g2_fill_1 FILLER_3_713 ();
 sg13g2_fill_1 FILLER_3_719 ();
 sg13g2_decap_4 FILLER_3_725 ();
 sg13g2_fill_1 FILLER_3_744 ();
 sg13g2_fill_2 FILLER_3_762 ();
 sg13g2_fill_1 FILLER_3_764 ();
 sg13g2_decap_8 FILLER_3_769 ();
 sg13g2_decap_8 FILLER_3_776 ();
 sg13g2_decap_8 FILLER_3_806 ();
 sg13g2_decap_8 FILLER_3_813 ();
 sg13g2_fill_2 FILLER_3_820 ();
 sg13g2_fill_1 FILLER_3_822 ();
 sg13g2_fill_1 FILLER_4_8 ();
 sg13g2_decap_4 FILLER_4_13 ();
 sg13g2_fill_2 FILLER_4_17 ();
 sg13g2_fill_1 FILLER_4_24 ();
 sg13g2_fill_2 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_73 ();
 sg13g2_decap_8 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_87 ();
 sg13g2_decap_8 FILLER_4_94 ();
 sg13g2_decap_8 FILLER_4_101 ();
 sg13g2_decap_8 FILLER_4_108 ();
 sg13g2_decap_8 FILLER_4_115 ();
 sg13g2_decap_8 FILLER_4_122 ();
 sg13g2_decap_8 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_136 ();
 sg13g2_decap_8 FILLER_4_143 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_206 ();
 sg13g2_decap_8 FILLER_4_213 ();
 sg13g2_decap_8 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_227 ();
 sg13g2_decap_8 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_241 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_8 FILLER_4_255 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_4_430 ();
 sg13g2_decap_8 FILLER_4_437 ();
 sg13g2_decap_8 FILLER_4_444 ();
 sg13g2_decap_8 FILLER_4_451 ();
 sg13g2_decap_8 FILLER_4_458 ();
 sg13g2_decap_8 FILLER_4_465 ();
 sg13g2_decap_8 FILLER_4_472 ();
 sg13g2_decap_8 FILLER_4_479 ();
 sg13g2_fill_2 FILLER_4_486 ();
 sg13g2_decap_8 FILLER_4_493 ();
 sg13g2_decap_4 FILLER_4_505 ();
 sg13g2_fill_2 FILLER_4_509 ();
 sg13g2_decap_8 FILLER_4_565 ();
 sg13g2_decap_4 FILLER_4_592 ();
 sg13g2_fill_1 FILLER_4_596 ();
 sg13g2_decap_4 FILLER_4_602 ();
 sg13g2_fill_2 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_624 ();
 sg13g2_decap_8 FILLER_4_631 ();
 sg13g2_decap_8 FILLER_4_638 ();
 sg13g2_fill_2 FILLER_4_645 ();
 sg13g2_fill_1 FILLER_4_647 ();
 sg13g2_fill_2 FILLER_4_739 ();
 sg13g2_fill_1 FILLER_4_741 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_decap_4 FILLER_5_20 ();
 sg13g2_fill_1 FILLER_5_34 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_fill_1 FILLER_5_469 ();
 sg13g2_decap_4 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_505 ();
 sg13g2_decap_4 FILLER_5_512 ();
 sg13g2_decap_8 FILLER_5_520 ();
 sg13g2_fill_2 FILLER_5_527 ();
 sg13g2_fill_1 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_548 ();
 sg13g2_decap_4 FILLER_5_555 ();
 sg13g2_decap_8 FILLER_5_563 ();
 sg13g2_fill_2 FILLER_5_570 ();
 sg13g2_fill_1 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_605 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_fill_1 FILLER_5_648 ();
 sg13g2_fill_1 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_fill_2 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_719 ();
 sg13g2_decap_8 FILLER_5_726 ();
 sg13g2_fill_2 FILLER_5_733 ();
 sg13g2_fill_2 FILLER_5_744 ();
 sg13g2_fill_1 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_fill_2 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_decap_4 FILLER_5_778 ();
 sg13g2_fill_2 FILLER_5_782 ();
 sg13g2_fill_2 FILLER_5_794 ();
 sg13g2_fill_1 FILLER_5_796 ();
 sg13g2_fill_2 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_808 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_fill_1 FILLER_5_822 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_32 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_decap_8 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_65 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_decap_8 FILLER_6_93 ();
 sg13g2_decap_8 FILLER_6_100 ();
 sg13g2_decap_8 FILLER_6_107 ();
 sg13g2_decap_8 FILLER_6_114 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_decap_8 FILLER_6_198 ();
 sg13g2_decap_8 FILLER_6_205 ();
 sg13g2_decap_8 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_219 ();
 sg13g2_decap_8 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_233 ();
 sg13g2_decap_8 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_decap_8 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_6_436 ();
 sg13g2_decap_8 FILLER_6_443 ();
 sg13g2_decap_8 FILLER_6_450 ();
 sg13g2_decap_8 FILLER_6_457 ();
 sg13g2_decap_8 FILLER_6_464 ();
 sg13g2_decap_4 FILLER_6_471 ();
 sg13g2_decap_4 FILLER_6_479 ();
 sg13g2_fill_2 FILLER_6_483 ();
 sg13g2_fill_2 FILLER_6_490 ();
 sg13g2_fill_1 FILLER_6_492 ();
 sg13g2_decap_8 FILLER_6_512 ();
 sg13g2_decap_8 FILLER_6_519 ();
 sg13g2_decap_8 FILLER_6_526 ();
 sg13g2_decap_4 FILLER_6_533 ();
 sg13g2_decap_4 FILLER_6_547 ();
 sg13g2_fill_2 FILLER_6_551 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_4 FILLER_6_574 ();
 sg13g2_fill_1 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_587 ();
 sg13g2_decap_8 FILLER_6_594 ();
 sg13g2_decap_8 FILLER_6_601 ();
 sg13g2_fill_2 FILLER_6_608 ();
 sg13g2_fill_2 FILLER_6_619 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_fill_1 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_fill_1 FILLER_6_683 ();
 sg13g2_fill_2 FILLER_6_689 ();
 sg13g2_fill_1 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_696 ();
 sg13g2_decap_8 FILLER_6_703 ();
 sg13g2_decap_4 FILLER_6_710 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_4 FILLER_6_756 ();
 sg13g2_fill_1 FILLER_6_760 ();
 sg13g2_decap_4 FILLER_6_793 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_13 ();
 sg13g2_decap_8 FILLER_7_24 ();
 sg13g2_fill_2 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_37 ();
 sg13g2_decap_8 FILLER_7_71 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_decap_8 FILLER_7_85 ();
 sg13g2_decap_8 FILLER_7_92 ();
 sg13g2_decap_8 FILLER_7_99 ();
 sg13g2_decap_8 FILLER_7_106 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_decap_8 FILLER_7_120 ();
 sg13g2_decap_8 FILLER_7_127 ();
 sg13g2_decap_8 FILLER_7_134 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_decap_8 FILLER_7_148 ();
 sg13g2_decap_8 FILLER_7_155 ();
 sg13g2_decap_8 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_169 ();
 sg13g2_decap_8 FILLER_7_176 ();
 sg13g2_decap_8 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_190 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_225 ();
 sg13g2_decap_8 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_239 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_8 FILLER_7_253 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_decap_8 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_7_435 ();
 sg13g2_decap_8 FILLER_7_442 ();
 sg13g2_decap_8 FILLER_7_449 ();
 sg13g2_decap_8 FILLER_7_456 ();
 sg13g2_decap_8 FILLER_7_463 ();
 sg13g2_decap_8 FILLER_7_470 ();
 sg13g2_decap_8 FILLER_7_477 ();
 sg13g2_decap_4 FILLER_7_494 ();
 sg13g2_fill_1 FILLER_7_556 ();
 sg13g2_fill_1 FILLER_7_589 ();
 sg13g2_decap_4 FILLER_7_594 ();
 sg13g2_fill_2 FILLER_7_608 ();
 sg13g2_decap_4 FILLER_7_615 ();
 sg13g2_decap_4 FILLER_7_623 ();
 sg13g2_fill_2 FILLER_7_627 ();
 sg13g2_fill_2 FILLER_7_634 ();
 sg13g2_decap_8 FILLER_7_640 ();
 sg13g2_decap_8 FILLER_7_647 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_4 FILLER_7_672 ();
 sg13g2_fill_1 FILLER_7_686 ();
 sg13g2_fill_2 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_774 ();
 sg13g2_decap_4 FILLER_8_4 ();
 sg13g2_fill_2 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_37 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_48 ();
 sg13g2_decap_8 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_decap_8 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_76 ();
 sg13g2_decap_8 FILLER_8_83 ();
 sg13g2_decap_8 FILLER_8_90 ();
 sg13g2_decap_8 FILLER_8_97 ();
 sg13g2_decap_8 FILLER_8_104 ();
 sg13g2_decap_8 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_118 ();
 sg13g2_decap_8 FILLER_8_125 ();
 sg13g2_decap_8 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_139 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_174 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_412 ();
 sg13g2_decap_8 FILLER_8_419 ();
 sg13g2_decap_8 FILLER_8_426 ();
 sg13g2_decap_8 FILLER_8_433 ();
 sg13g2_decap_8 FILLER_8_440 ();
 sg13g2_decap_8 FILLER_8_447 ();
 sg13g2_decap_8 FILLER_8_454 ();
 sg13g2_decap_4 FILLER_8_461 ();
 sg13g2_fill_1 FILLER_8_465 ();
 sg13g2_decap_4 FILLER_8_493 ();
 sg13g2_decap_4 FILLER_8_528 ();
 sg13g2_fill_2 FILLER_8_532 ();
 sg13g2_decap_4 FILLER_8_538 ();
 sg13g2_fill_1 FILLER_8_542 ();
 sg13g2_decap_4 FILLER_8_553 ();
 sg13g2_fill_2 FILLER_8_557 ();
 sg13g2_fill_2 FILLER_8_563 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_decap_4 FILLER_8_580 ();
 sg13g2_fill_1 FILLER_8_584 ();
 sg13g2_fill_1 FILLER_8_612 ();
 sg13g2_decap_8 FILLER_8_632 ();
 sg13g2_fill_2 FILLER_8_639 ();
 sg13g2_fill_2 FILLER_8_677 ();
 sg13g2_decap_8 FILLER_8_691 ();
 sg13g2_decap_8 FILLER_8_698 ();
 sg13g2_decap_8 FILLER_8_705 ();
 sg13g2_decap_4 FILLER_8_712 ();
 sg13g2_fill_1 FILLER_8_716 ();
 sg13g2_decap_8 FILLER_8_727 ();
 sg13g2_fill_2 FILLER_8_734 ();
 sg13g2_fill_2 FILLER_8_745 ();
 sg13g2_fill_1 FILLER_8_747 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_759 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_decap_4 FILLER_8_773 ();
 sg13g2_fill_2 FILLER_8_777 ();
 sg13g2_decap_4 FILLER_8_789 ();
 sg13g2_fill_2 FILLER_8_793 ();
 sg13g2_fill_1 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_808 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_822 ();
 sg13g2_fill_2 FILLER_9_17 ();
 sg13g2_fill_1 FILLER_9_19 ();
 sg13g2_decap_4 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_decap_8 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_120 ();
 sg13g2_decap_8 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_134 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_155 ();
 sg13g2_decap_8 FILLER_9_162 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_decap_8 FILLER_9_183 ();
 sg13g2_decap_8 FILLER_9_190 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_decap_8 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_9_414 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_decap_8 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_9_435 ();
 sg13g2_decap_8 FILLER_9_442 ();
 sg13g2_fill_2 FILLER_9_449 ();
 sg13g2_fill_1 FILLER_9_451 ();
 sg13g2_fill_1 FILLER_9_457 ();
 sg13g2_fill_2 FILLER_9_463 ();
 sg13g2_fill_1 FILLER_9_470 ();
 sg13g2_decap_4 FILLER_9_475 ();
 sg13g2_fill_2 FILLER_9_489 ();
 sg13g2_decap_4 FILLER_9_551 ();
 sg13g2_fill_1 FILLER_9_555 ();
 sg13g2_decap_8 FILLER_9_561 ();
 sg13g2_decap_8 FILLER_9_568 ();
 sg13g2_fill_1 FILLER_9_575 ();
 sg13g2_decap_8 FILLER_9_608 ();
 sg13g2_decap_4 FILLER_9_615 ();
 sg13g2_fill_2 FILLER_9_654 ();
 sg13g2_fill_2 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_fill_2 FILLER_9_756 ();
 sg13g2_fill_1 FILLER_9_758 ();
 sg13g2_fill_2 FILLER_9_800 ();
 sg13g2_fill_1 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_fill_2 FILLER_9_821 ();
 sg13g2_fill_2 FILLER_10_8 ();
 sg13g2_fill_1 FILLER_10_10 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_41 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_fill_1 FILLER_10_424 ();
 sg13g2_fill_1 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_514 ();
 sg13g2_fill_2 FILLER_10_521 ();
 sg13g2_fill_1 FILLER_10_523 ();
 sg13g2_decap_8 FILLER_10_533 ();
 sg13g2_decap_8 FILLER_10_540 ();
 sg13g2_fill_2 FILLER_10_557 ();
 sg13g2_fill_1 FILLER_10_559 ();
 sg13g2_decap_8 FILLER_10_587 ();
 sg13g2_fill_2 FILLER_10_594 ();
 sg13g2_fill_1 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_fill_1 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_fill_1 FILLER_10_704 ();
 sg13g2_fill_1 FILLER_10_723 ();
 sg13g2_fill_2 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_771 ();
 sg13g2_fill_2 FILLER_10_778 ();
 sg13g2_fill_1 FILLER_10_780 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_37 ();
 sg13g2_fill_1 FILLER_11_39 ();
 sg13g2_decap_4 FILLER_11_45 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_89 ();
 sg13g2_decap_8 FILLER_11_96 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_194 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_decap_8 FILLER_11_208 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_229 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_413 ();
 sg13g2_fill_2 FILLER_11_419 ();
 sg13g2_fill_1 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_fill_2 FILLER_11_455 ();
 sg13g2_fill_1 FILLER_11_457 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_fill_2 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_489 ();
 sg13g2_decap_8 FILLER_11_496 ();
 sg13g2_decap_8 FILLER_11_503 ();
 sg13g2_decap_4 FILLER_11_510 ();
 sg13g2_fill_1 FILLER_11_514 ();
 sg13g2_fill_2 FILLER_11_562 ();
 sg13g2_fill_1 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_569 ();
 sg13g2_decap_4 FILLER_11_576 ();
 sg13g2_fill_1 FILLER_11_580 ();
 sg13g2_decap_4 FILLER_11_585 ();
 sg13g2_fill_2 FILLER_11_589 ();
 sg13g2_decap_8 FILLER_11_678 ();
 sg13g2_decap_4 FILLER_11_685 ();
 sg13g2_fill_1 FILLER_11_689 ();
 sg13g2_fill_2 FILLER_11_734 ();
 sg13g2_fill_1 FILLER_11_744 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_4 FILLER_11_774 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_fill_2 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_fill_1 FILLER_12_8 ();
 sg13g2_fill_2 FILLER_12_17 ();
 sg13g2_decap_8 FILLER_12_29 ();
 sg13g2_decap_4 FILLER_12_36 ();
 sg13g2_fill_1 FILLER_12_40 ();
 sg13g2_decap_8 FILLER_12_72 ();
 sg13g2_decap_8 FILLER_12_79 ();
 sg13g2_decap_8 FILLER_12_86 ();
 sg13g2_decap_8 FILLER_12_93 ();
 sg13g2_decap_8 FILLER_12_100 ();
 sg13g2_decap_8 FILLER_12_107 ();
 sg13g2_decap_8 FILLER_12_114 ();
 sg13g2_decap_8 FILLER_12_121 ();
 sg13g2_decap_8 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_decap_8 FILLER_12_142 ();
 sg13g2_decap_8 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_8 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_375 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_4 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_4 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_fill_2 FILLER_12_473 ();
 sg13g2_decap_4 FILLER_12_507 ();
 sg13g2_fill_1 FILLER_12_511 ();
 sg13g2_fill_2 FILLER_12_539 ();
 sg13g2_decap_4 FILLER_12_555 ();
 sg13g2_decap_8 FILLER_12_563 ();
 sg13g2_decap_8 FILLER_12_570 ();
 sg13g2_decap_8 FILLER_12_577 ();
 sg13g2_decap_8 FILLER_12_584 ();
 sg13g2_decap_8 FILLER_12_625 ();
 sg13g2_decap_8 FILLER_12_632 ();
 sg13g2_fill_2 FILLER_12_639 ();
 sg13g2_decap_8 FILLER_12_645 ();
 sg13g2_fill_2 FILLER_12_652 ();
 sg13g2_fill_2 FILLER_12_659 ();
 sg13g2_fill_1 FILLER_12_661 ();
 sg13g2_fill_2 FILLER_12_672 ();
 sg13g2_fill_2 FILLER_12_701 ();
 sg13g2_fill_1 FILLER_12_703 ();
 sg13g2_fill_2 FILLER_12_724 ();
 sg13g2_fill_1 FILLER_12_726 ();
 sg13g2_decap_4 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_785 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_34 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_fill_2 FILLER_13_364 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_4 FILLER_13_419 ();
 sg13g2_fill_1 FILLER_13_423 ();
 sg13g2_decap_4 FILLER_13_438 ();
 sg13g2_fill_1 FILLER_13_442 ();
 sg13g2_fill_2 FILLER_13_479 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_fill_1 FILLER_13_492 ();
 sg13g2_fill_1 FILLER_13_520 ();
 sg13g2_decap_4 FILLER_13_535 ();
 sg13g2_fill_1 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_618 ();
 sg13g2_fill_2 FILLER_13_625 ();
 sg13g2_fill_1 FILLER_13_627 ();
 sg13g2_decap_4 FILLER_13_655 ();
 sg13g2_fill_2 FILLER_13_663 ();
 sg13g2_fill_1 FILLER_13_665 ();
 sg13g2_decap_4 FILLER_13_675 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_4 FILLER_13_690 ();
 sg13g2_fill_1 FILLER_13_694 ();
 sg13g2_decap_8 FILLER_13_699 ();
 sg13g2_fill_2 FILLER_13_706 ();
 sg13g2_fill_1 FILLER_13_721 ();
 sg13g2_fill_2 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_4 FILLER_13_747 ();
 sg13g2_fill_2 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_757 ();
 sg13g2_decap_8 FILLER_13_764 ();
 sg13g2_fill_2 FILLER_13_794 ();
 sg13g2_fill_2 FILLER_13_800 ();
 sg13g2_decap_8 FILLER_13_806 ();
 sg13g2_decap_8 FILLER_13_813 ();
 sg13g2_fill_2 FILLER_13_820 ();
 sg13g2_fill_1 FILLER_13_822 ();
 sg13g2_decap_4 FILLER_14_4 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_58 ();
 sg13g2_decap_8 FILLER_14_65 ();
 sg13g2_decap_8 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_79 ();
 sg13g2_decap_8 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_decap_8 FILLER_14_107 ();
 sg13g2_decap_8 FILLER_14_114 ();
 sg13g2_decap_8 FILLER_14_121 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_4 FILLER_14_345 ();
 sg13g2_fill_2 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_366 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_fill_2 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_464 ();
 sg13g2_fill_1 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_4 FILLER_14_490 ();
 sg13g2_fill_2 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_510 ();
 sg13g2_fill_2 FILLER_14_517 ();
 sg13g2_fill_1 FILLER_14_519 ();
 sg13g2_decap_8 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_550 ();
 sg13g2_decap_8 FILLER_14_557 ();
 sg13g2_decap_4 FILLER_14_564 ();
 sg13g2_fill_1 FILLER_14_568 ();
 sg13g2_decap_4 FILLER_14_573 ();
 sg13g2_fill_1 FILLER_14_577 ();
 sg13g2_fill_2 FILLER_14_587 ();
 sg13g2_fill_1 FILLER_14_589 ();
 sg13g2_fill_2 FILLER_14_604 ();
 sg13g2_decap_4 FILLER_14_642 ();
 sg13g2_fill_1 FILLER_14_646 ();
 sg13g2_fill_1 FILLER_14_652 ();
 sg13g2_decap_4 FILLER_14_668 ();
 sg13g2_fill_2 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_fill_2 FILLER_14_692 ();
 sg13g2_fill_1 FILLER_14_694 ();
 sg13g2_decap_8 FILLER_14_699 ();
 sg13g2_decap_4 FILLER_14_706 ();
 sg13g2_fill_2 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_738 ();
 sg13g2_fill_2 FILLER_14_745 ();
 sg13g2_fill_1 FILLER_14_747 ();
 sg13g2_fill_2 FILLER_14_775 ();
 sg13g2_fill_2 FILLER_14_787 ();
 sg13g2_fill_1 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_4 FILLER_14_817 ();
 sg13g2_fill_2 FILLER_14_821 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_13 ();
 sg13g2_fill_1 FILLER_15_15 ();
 sg13g2_decap_8 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_381 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_fill_1 FILLER_15_389 ();
 sg13g2_decap_4 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_431 ();
 sg13g2_fill_2 FILLER_15_436 ();
 sg13g2_decap_8 FILLER_15_442 ();
 sg13g2_decap_8 FILLER_15_449 ();
 sg13g2_decap_8 FILLER_15_456 ();
 sg13g2_decap_4 FILLER_15_463 ();
 sg13g2_decap_8 FILLER_15_517 ();
 sg13g2_decap_4 FILLER_15_524 ();
 sg13g2_fill_2 FILLER_15_528 ();
 sg13g2_fill_2 FILLER_15_561 ();
 sg13g2_fill_1 FILLER_15_563 ();
 sg13g2_decap_4 FILLER_15_591 ();
 sg13g2_fill_1 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_604 ();
 sg13g2_fill_1 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_4 FILLER_15_627 ();
 sg13g2_fill_1 FILLER_15_631 ();
 sg13g2_fill_2 FILLER_15_637 ();
 sg13g2_decap_4 FILLER_15_644 ();
 sg13g2_fill_2 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_fill_2 FILLER_15_662 ();
 sg13g2_fill_1 FILLER_15_664 ();
 sg13g2_decap_8 FILLER_15_755 ();
 sg13g2_decap_4 FILLER_15_762 ();
 sg13g2_fill_1 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_fill_1 FILLER_15_784 ();
 sg13g2_decap_4 FILLER_15_789 ();
 sg13g2_fill_1 FILLER_15_793 ();
 sg13g2_fill_2 FILLER_15_821 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_decap_4 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_48 ();
 sg13g2_decap_8 FILLER_16_54 ();
 sg13g2_decap_8 FILLER_16_61 ();
 sg13g2_decap_8 FILLER_16_68 ();
 sg13g2_decap_8 FILLER_16_75 ();
 sg13g2_decap_8 FILLER_16_82 ();
 sg13g2_decap_8 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_96 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_decap_8 FILLER_16_117 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_decap_8 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_8 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_159 ();
 sg13g2_decap_8 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_decap_8 FILLER_16_236 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_278 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_decap_8 FILLER_16_313 ();
 sg13g2_decap_4 FILLER_16_320 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_416 ();
 sg13g2_decap_4 FILLER_16_422 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_473 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_491 ();
 sg13g2_fill_2 FILLER_16_497 ();
 sg13g2_fill_1 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_535 ();
 sg13g2_decap_8 FILLER_16_542 ();
 sg13g2_decap_8 FILLER_16_549 ();
 sg13g2_decap_4 FILLER_16_556 ();
 sg13g2_fill_2 FILLER_16_565 ();
 sg13g2_decap_4 FILLER_16_572 ();
 sg13g2_fill_1 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_587 ();
 sg13g2_fill_1 FILLER_16_594 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_decap_8 FILLER_16_617 ();
 sg13g2_decap_4 FILLER_16_624 ();
 sg13g2_fill_1 FILLER_16_628 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_fill_2 FILLER_16_655 ();
 sg13g2_fill_1 FILLER_16_657 ();
 sg13g2_decap_4 FILLER_16_668 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_4 FILLER_16_704 ();
 sg13g2_fill_1 FILLER_16_718 ();
 sg13g2_decap_4 FILLER_16_727 ();
 sg13g2_fill_2 FILLER_16_731 ();
 sg13g2_decap_4 FILLER_16_737 ();
 sg13g2_fill_1 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_788 ();
 sg13g2_fill_1 FILLER_16_799 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_4 FILLER_16_818 ();
 sg13g2_fill_1 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_22 ();
 sg13g2_fill_2 FILLER_17_38 ();
 sg13g2_decap_8 FILLER_17_72 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_93 ();
 sg13g2_decap_8 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_107 ();
 sg13g2_decap_8 FILLER_17_114 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_decap_8 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_4 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_4 FILLER_17_371 ();
 sg13g2_decap_4 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_17_454 ();
 sg13g2_fill_1 FILLER_17_456 ();
 sg13g2_decap_4 FILLER_17_484 ();
 sg13g2_decap_8 FILLER_17_493 ();
 sg13g2_decap_8 FILLER_17_500 ();
 sg13g2_decap_8 FILLER_17_507 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_521 ();
 sg13g2_fill_1 FILLER_17_580 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_fill_2 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_594 ();
 sg13g2_fill_1 FILLER_17_626 ();
 sg13g2_decap_4 FILLER_17_663 ();
 sg13g2_fill_2 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_701 ();
 sg13g2_fill_2 FILLER_17_716 ();
 sg13g2_decap_8 FILLER_17_736 ();
 sg13g2_fill_2 FILLER_17_743 ();
 sg13g2_decap_4 FILLER_17_777 ();
 sg13g2_fill_2 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_fill_1 FILLER_17_794 ();
 sg13g2_fill_1 FILLER_17_822 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_decap_4 FILLER_18_13 ();
 sg13g2_decap_8 FILLER_18_31 ();
 sg13g2_decap_8 FILLER_18_38 ();
 sg13g2_decap_8 FILLER_18_45 ();
 sg13g2_decap_8 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_73 ();
 sg13g2_decap_8 FILLER_18_80 ();
 sg13g2_decap_8 FILLER_18_87 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_decap_8 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_decap_4 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_4 FILLER_18_419 ();
 sg13g2_decap_8 FILLER_18_428 ();
 sg13g2_decap_4 FILLER_18_435 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_4 FILLER_18_455 ();
 sg13g2_fill_1 FILLER_18_491 ();
 sg13g2_fill_2 FILLER_18_519 ();
 sg13g2_decap_4 FILLER_18_552 ();
 sg13g2_fill_2 FILLER_18_556 ();
 sg13g2_decap_8 FILLER_18_562 ();
 sg13g2_decap_8 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_fill_2 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_608 ();
 sg13g2_decap_8 FILLER_18_615 ();
 sg13g2_fill_2 FILLER_18_622 ();
 sg13g2_decap_8 FILLER_18_649 ();
 sg13g2_fill_1 FILLER_18_656 ();
 sg13g2_decap_4 FILLER_18_676 ();
 sg13g2_decap_8 FILLER_18_684 ();
 sg13g2_fill_2 FILLER_18_691 ();
 sg13g2_fill_2 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_fill_2 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_fill_2 FILLER_18_821 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_36 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_50 ();
 sg13g2_decap_8 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_71 ();
 sg13g2_decap_8 FILLER_19_78 ();
 sg13g2_decap_8 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_99 ();
 sg13g2_decap_8 FILLER_19_106 ();
 sg13g2_decap_8 FILLER_19_113 ();
 sg13g2_decap_8 FILLER_19_120 ();
 sg13g2_decap_8 FILLER_19_127 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_decap_8 FILLER_19_148 ();
 sg13g2_decap_8 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_162 ();
 sg13g2_decap_8 FILLER_19_169 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_8 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_4 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_fill_2 FILLER_19_399 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_19_435 ();
 sg13g2_decap_8 FILLER_19_442 ();
 sg13g2_decap_8 FILLER_19_453 ();
 sg13g2_decap_4 FILLER_19_460 ();
 sg13g2_fill_2 FILLER_19_464 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_fill_2 FILLER_19_495 ();
 sg13g2_fill_1 FILLER_19_497 ();
 sg13g2_fill_2 FILLER_19_502 ();
 sg13g2_decap_4 FILLER_19_508 ();
 sg13g2_fill_1 FILLER_19_512 ();
 sg13g2_decap_4 FILLER_19_517 ();
 sg13g2_fill_1 FILLER_19_521 ();
 sg13g2_fill_2 FILLER_19_527 ();
 sg13g2_fill_2 FILLER_19_534 ();
 sg13g2_fill_1 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_fill_2 FILLER_19_622 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_fill_2 FILLER_19_665 ();
 sg13g2_fill_1 FILLER_19_667 ();
 sg13g2_fill_2 FILLER_19_672 ();
 sg13g2_fill_1 FILLER_19_674 ();
 sg13g2_fill_2 FILLER_19_706 ();
 sg13g2_fill_1 FILLER_19_708 ();
 sg13g2_decap_4 FILLER_19_713 ();
 sg13g2_fill_2 FILLER_19_717 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_fill_2 FILLER_19_747 ();
 sg13g2_fill_1 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_fill_1 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_decap_4 FILLER_19_787 ();
 sg13g2_fill_1 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_fill_2 FILLER_19_817 ();
 sg13g2_fill_1 FILLER_19_819 ();
 sg13g2_decap_4 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_8 ();
 sg13g2_fill_2 FILLER_20_27 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_4 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_2 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_20_441 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_1 FILLER_20_471 ();
 sg13g2_fill_2 FILLER_20_477 ();
 sg13g2_fill_1 FILLER_20_479 ();
 sg13g2_decap_8 FILLER_20_484 ();
 sg13g2_decap_8 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_498 ();
 sg13g2_fill_1 FILLER_20_530 ();
 sg13g2_decap_4 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_539 ();
 sg13g2_fill_2 FILLER_20_550 ();
 sg13g2_decap_4 FILLER_20_556 ();
 sg13g2_fill_1 FILLER_20_563 ();
 sg13g2_fill_2 FILLER_20_567 ();
 sg13g2_fill_1 FILLER_20_572 ();
 sg13g2_fill_2 FILLER_20_576 ();
 sg13g2_fill_1 FILLER_20_581 ();
 sg13g2_fill_1 FILLER_20_585 ();
 sg13g2_fill_1 FILLER_20_589 ();
 sg13g2_fill_1 FILLER_20_606 ();
 sg13g2_fill_1 FILLER_20_610 ();
 sg13g2_fill_1 FILLER_20_614 ();
 sg13g2_fill_1 FILLER_20_618 ();
 sg13g2_fill_2 FILLER_20_622 ();
 sg13g2_fill_2 FILLER_20_627 ();
 sg13g2_fill_1 FILLER_20_664 ();
 sg13g2_fill_2 FILLER_20_668 ();
 sg13g2_fill_1 FILLER_20_673 ();
 sg13g2_fill_1 FILLER_20_677 ();
 sg13g2_fill_1 FILLER_20_681 ();
 sg13g2_fill_1 FILLER_20_685 ();
 sg13g2_fill_2 FILLER_20_689 ();
 sg13g2_fill_1 FILLER_20_694 ();
 sg13g2_fill_1 FILLER_20_698 ();
 sg13g2_fill_1 FILLER_20_702 ();
 sg13g2_fill_1 FILLER_20_706 ();
 sg13g2_fill_1 FILLER_20_710 ();
 sg13g2_fill_2 FILLER_20_714 ();
 sg13g2_fill_1 FILLER_20_719 ();
 sg13g2_fill_1 FILLER_20_723 ();
 sg13g2_fill_1 FILLER_20_727 ();
 sg13g2_fill_1 FILLER_20_731 ();
 sg13g2_fill_1 FILLER_20_735 ();
 sg13g2_fill_2 FILLER_20_739 ();
 sg13g2_fill_1 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_748 ();
 sg13g2_fill_1 FILLER_20_752 ();
 sg13g2_fill_1 FILLER_20_756 ();
 sg13g2_fill_1 FILLER_20_760 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_769 ();
 sg13g2_fill_1 FILLER_20_773 ();
 sg13g2_fill_1 FILLER_20_777 ();
 sg13g2_fill_1 FILLER_20_781 ();
 sg13g2_decap_4 FILLER_20_785 ();
 sg13g2_fill_1 FILLER_20_789 ();
 sg13g2_fill_1 FILLER_20_793 ();
 sg13g2_fill_1 FILLER_20_803 ();
 sg13g2_fill_1 FILLER_20_807 ();
 sg13g2_fill_1 FILLER_20_811 ();
 sg13g2_fill_2 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_45 ();
 sg13g2_decap_8 FILLER_21_52 ();
 sg13g2_decap_8 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_66 ();
 sg13g2_decap_8 FILLER_21_73 ();
 sg13g2_decap_8 FILLER_21_80 ();
 sg13g2_decap_8 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_185 ();
 sg13g2_decap_8 FILLER_21_192 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_4 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_4 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_377 ();
 sg13g2_decap_4 FILLER_21_410 ();
 sg13g2_fill_1 FILLER_21_418 ();
 sg13g2_fill_2 FILLER_21_446 ();
 sg13g2_fill_1 FILLER_21_448 ();
 sg13g2_fill_2 FILLER_21_502 ();
 sg13g2_fill_1 FILLER_21_504 ();
 sg13g2_fill_2 FILLER_21_515 ();
 sg13g2_fill_2 FILLER_21_539 ();
 sg13g2_decap_4 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_8 ();
 sg13g2_decap_8 FILLER_22_13 ();
 sg13g2_decap_8 FILLER_22_20 ();
 sg13g2_decap_8 FILLER_22_27 ();
 sg13g2_decap_8 FILLER_22_34 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_decap_8 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_decap_8 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_83 ();
 sg13g2_decap_8 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_decap_8 FILLER_22_124 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_decap_8 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_4 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_decap_4 FILLER_22_337 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_4 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_22_436 ();
 sg13g2_fill_2 FILLER_22_470 ();
 sg13g2_fill_1 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_486 ();
 sg13g2_fill_2 FILLER_22_493 ();
 sg13g2_fill_1 FILLER_22_495 ();
 sg13g2_fill_2 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_507 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_194 ();
 sg13g2_decap_8 FILLER_23_201 ();
 sg13g2_decap_8 FILLER_23_208 ();
 sg13g2_decap_4 FILLER_23_215 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_decap_4 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_fill_2 FILLER_23_423 ();
 sg13g2_fill_1 FILLER_23_425 ();
 sg13g2_decap_8 FILLER_23_461 ();
 sg13g2_decap_8 FILLER_23_468 ();
 sg13g2_fill_1 FILLER_23_475 ();
 sg13g2_fill_2 FILLER_23_485 ();
 sg13g2_decap_4 FILLER_23_492 ();
 sg13g2_fill_1 FILLER_23_496 ();
 sg13g2_fill_2 FILLER_23_519 ();
 sg13g2_fill_1 FILLER_23_521 ();
 sg13g2_decap_4 FILLER_23_530 ();
 sg13g2_fill_1 FILLER_23_534 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_fill_1 FILLER_24_420 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_1 FILLER_24_503 ();
 sg13g2_fill_1 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_537 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_4 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_decap_8 FILLER_25_52 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_8 FILLER_25_73 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_87 ();
 sg13g2_decap_8 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_108 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_decap_8 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_4 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_346 ();
 sg13g2_decap_4 FILLER_25_353 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_418 ();
 sg13g2_fill_2 FILLER_25_452 ();
 sg13g2_fill_2 FILLER_25_458 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_decap_8 FILLER_25_471 ();
 sg13g2_fill_2 FILLER_25_478 ();
 sg13g2_fill_1 FILLER_25_480 ();
 sg13g2_fill_1 FILLER_25_485 ();
 sg13g2_decap_8 FILLER_25_494 ();
 sg13g2_decap_4 FILLER_25_501 ();
 sg13g2_fill_1 FILLER_25_505 ();
 sg13g2_decap_4 FILLER_25_510 ();
 sg13g2_fill_2 FILLER_25_514 ();
 sg13g2_decap_8 FILLER_25_521 ();
 sg13g2_decap_8 FILLER_25_528 ();
 sg13g2_decap_8 FILLER_25_535 ();
 sg13g2_fill_2 FILLER_25_542 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_4 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_34 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_4 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_decap_4 FILLER_26_358 ();
 sg13g2_decap_4 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_425 ();
 sg13g2_decap_4 FILLER_26_435 ();
 sg13g2_fill_1 FILLER_26_439 ();
 sg13g2_fill_1 FILLER_26_444 ();
 sg13g2_decap_4 FILLER_26_457 ();
 sg13g2_fill_1 FILLER_26_461 ();
 sg13g2_decap_4 FILLER_26_471 ();
 sg13g2_fill_1 FILLER_26_475 ();
 sg13g2_decap_8 FILLER_26_481 ();
 sg13g2_fill_2 FILLER_26_488 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_40 ();
 sg13g2_decap_8 FILLER_27_47 ();
 sg13g2_decap_8 FILLER_27_54 ();
 sg13g2_decap_8 FILLER_27_61 ();
 sg13g2_decap_8 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_75 ();
 sg13g2_decap_8 FILLER_27_82 ();
 sg13g2_decap_8 FILLER_27_89 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_8 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_117 ();
 sg13g2_decap_8 FILLER_27_124 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_decap_8 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_decap_4 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_decap_4 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_355 ();
 sg13g2_decap_4 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_27_414 ();
 sg13g2_fill_1 FILLER_27_418 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_decap_8 FILLER_27_430 ();
 sg13g2_fill_2 FILLER_27_437 ();
 sg13g2_decap_8 FILLER_27_443 ();
 sg13g2_decap_4 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_fill_1 FILLER_27_508 ();
 sg13g2_decap_8 FILLER_27_531 ();
 sg13g2_fill_2 FILLER_27_538 ();
 sg13g2_fill_1 FILLER_27_540 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_4 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_4 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_decap_4 FILLER_28_360 ();
 sg13g2_decap_4 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_fill_2 FILLER_28_412 ();
 sg13g2_decap_4 FILLER_28_428 ();
 sg13g2_fill_2 FILLER_28_432 ();
 sg13g2_fill_2 FILLER_28_461 ();
 sg13g2_decap_4 FILLER_28_472 ();
 sg13g2_fill_1 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_488 ();
 sg13g2_decap_4 FILLER_28_495 ();
 sg13g2_decap_4 FILLER_28_504 ();
 sg13g2_fill_2 FILLER_28_513 ();
 sg13g2_decap_4 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_17 ();
 sg13g2_decap_8 FILLER_29_24 ();
 sg13g2_decap_8 FILLER_29_31 ();
 sg13g2_decap_8 FILLER_29_38 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_59 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_decap_8 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_129 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_192 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_4 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_decap_4 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_fill_2 FILLER_29_455 ();
 sg13g2_decap_4 FILLER_29_462 ();
 sg13g2_fill_1 FILLER_29_466 ();
 sg13g2_fill_1 FILLER_29_476 ();
 sg13g2_decap_4 FILLER_29_504 ();
 sg13g2_decap_4 FILLER_29_535 ();
 sg13g2_fill_2 FILLER_29_539 ();
 sg13g2_decap_4 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_8 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_4 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_30_412 ();
 sg13g2_fill_2 FILLER_30_423 ();
 sg13g2_fill_1 FILLER_30_425 ();
 sg13g2_decap_8 FILLER_30_430 ();
 sg13g2_fill_2 FILLER_30_437 ();
 sg13g2_decap_8 FILLER_30_443 ();
 sg13g2_fill_1 FILLER_30_450 ();
 sg13g2_decap_8 FILLER_30_475 ();
 sg13g2_decap_8 FILLER_30_486 ();
 sg13g2_fill_1 FILLER_30_525 ();
 sg13g2_fill_1 FILLER_30_531 ();
 sg13g2_decap_4 FILLER_30_559 ();
 sg13g2_fill_1 FILLER_30_563 ();
 sg13g2_fill_1 FILLER_30_567 ();
 sg13g2_fill_2 FILLER_30_571 ();
 sg13g2_fill_1 FILLER_30_589 ();
 sg13g2_fill_1 FILLER_30_593 ();
 sg13g2_fill_1 FILLER_30_597 ();
 sg13g2_fill_1 FILLER_30_601 ();
 sg13g2_fill_2 FILLER_30_605 ();
 sg13g2_fill_1 FILLER_30_610 ();
 sg13g2_fill_1 FILLER_30_614 ();
 sg13g2_fill_1 FILLER_30_618 ();
 sg13g2_fill_1 FILLER_30_622 ();
 sg13g2_fill_1 FILLER_30_626 ();
 sg13g2_fill_2 FILLER_30_630 ();
 sg13g2_fill_1 FILLER_30_635 ();
 sg13g2_fill_1 FILLER_30_639 ();
 sg13g2_fill_1 FILLER_30_643 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_fill_1 FILLER_30_651 ();
 sg13g2_fill_2 FILLER_30_655 ();
 sg13g2_fill_1 FILLER_30_660 ();
 sg13g2_fill_1 FILLER_30_664 ();
 sg13g2_fill_1 FILLER_30_668 ();
 sg13g2_fill_1 FILLER_30_672 ();
 sg13g2_fill_2 FILLER_30_676 ();
 sg13g2_fill_1 FILLER_30_681 ();
 sg13g2_fill_1 FILLER_30_685 ();
 sg13g2_fill_1 FILLER_30_689 ();
 sg13g2_fill_1 FILLER_30_693 ();
 sg13g2_fill_2 FILLER_30_697 ();
 sg13g2_fill_1 FILLER_30_702 ();
 sg13g2_fill_1 FILLER_30_706 ();
 sg13g2_fill_1 FILLER_30_710 ();
 sg13g2_fill_1 FILLER_30_714 ();
 sg13g2_fill_2 FILLER_30_718 ();
 sg13g2_fill_1 FILLER_30_723 ();
 sg13g2_fill_1 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_731 ();
 sg13g2_fill_1 FILLER_30_735 ();
 sg13g2_fill_1 FILLER_30_739 ();
 sg13g2_fill_1 FILLER_30_743 ();
 sg13g2_fill_1 FILLER_30_747 ();
 sg13g2_fill_1 FILLER_30_751 ();
 sg13g2_fill_2 FILLER_30_755 ();
 sg13g2_fill_1 FILLER_30_760 ();
 sg13g2_fill_1 FILLER_30_764 ();
 sg13g2_fill_1 FILLER_30_768 ();
 sg13g2_fill_1 FILLER_30_772 ();
 sg13g2_fill_1 FILLER_30_776 ();
 sg13g2_fill_1 FILLER_30_780 ();
 sg13g2_fill_2 FILLER_30_784 ();
 sg13g2_decap_4 FILLER_30_789 ();
 sg13g2_fill_1 FILLER_30_793 ();
 sg13g2_fill_1 FILLER_30_806 ();
 sg13g2_fill_1 FILLER_30_810 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_decap_4 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_fill_1 FILLER_31_414 ();
 sg13g2_fill_1 FILLER_31_419 ();
 sg13g2_decap_4 FILLER_31_428 ();
 sg13g2_fill_2 FILLER_31_432 ();
 sg13g2_decap_4 FILLER_31_475 ();
 sg13g2_fill_2 FILLER_31_479 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_fill_2 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_503 ();
 sg13g2_decap_4 FILLER_31_510 ();
 sg13g2_fill_2 FILLER_31_523 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_decap_4 FILLER_31_530 ();
 sg13g2_fill_2 FILLER_31_534 ();
 sg13g2_decap_8 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_decap_8 FILLER_31_559 ();
 sg13g2_decap_4 FILLER_31_593 ();
 sg13g2_fill_1 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_675 ();
 sg13g2_decap_8 FILLER_31_682 ();
 sg13g2_decap_8 FILLER_31_689 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_decap_8 FILLER_31_711 ();
 sg13g2_decap_8 FILLER_31_718 ();
 sg13g2_decap_4 FILLER_31_725 ();
 sg13g2_fill_1 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_fill_2 FILLER_31_764 ();
 sg13g2_fill_1 FILLER_31_766 ();
 sg13g2_decap_4 FILLER_31_772 ();
 sg13g2_fill_2 FILLER_31_776 ();
 sg13g2_fill_1 FILLER_31_788 ();
 sg13g2_decap_4 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_fill_1 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_446 ();
 sg13g2_fill_1 FILLER_32_450 ();
 sg13g2_fill_1 FILLER_32_473 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_decap_4 FILLER_32_525 ();
 sg13g2_fill_2 FILLER_32_566 ();
 sg13g2_fill_1 FILLER_32_568 ();
 sg13g2_decap_8 FILLER_32_582 ();
 sg13g2_fill_2 FILLER_32_589 ();
 sg13g2_fill_2 FILLER_32_618 ();
 sg13g2_fill_2 FILLER_32_647 ();
 sg13g2_fill_1 FILLER_32_649 ();
 sg13g2_fill_1 FILLER_32_687 ();
 sg13g2_decap_4 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_81 ();
 sg13g2_decap_8 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_436 ();
 sg13g2_decap_4 FILLER_33_443 ();
 sg13g2_fill_2 FILLER_33_447 ();
 sg13g2_fill_1 FILLER_33_481 ();
 sg13g2_fill_2 FILLER_33_499 ();
 sg13g2_fill_1 FILLER_33_501 ();
 sg13g2_fill_2 FILLER_33_529 ();
 sg13g2_fill_1 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_decap_8 FILLER_33_555 ();
 sg13g2_fill_1 FILLER_33_562 ();
 sg13g2_fill_2 FILLER_33_567 ();
 sg13g2_fill_1 FILLER_33_569 ();
 sg13g2_fill_2 FILLER_33_590 ();
 sg13g2_fill_1 FILLER_33_600 ();
 sg13g2_fill_2 FILLER_33_631 ();
 sg13g2_fill_1 FILLER_33_633 ();
 sg13g2_fill_2 FILLER_33_671 ();
 sg13g2_fill_1 FILLER_33_673 ();
 sg13g2_fill_2 FILLER_33_679 ();
 sg13g2_fill_1 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_fill_2 FILLER_33_703 ();
 sg13g2_decap_8 FILLER_33_710 ();
 sg13g2_fill_1 FILLER_33_717 ();
 sg13g2_decap_4 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_745 ();
 sg13g2_decap_4 FILLER_33_752 ();
 sg13g2_decap_4 FILLER_33_760 ();
 sg13g2_fill_2 FILLER_33_764 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_4 FILLER_33_788 ();
 sg13g2_fill_2 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_8 FILLER_33_813 ();
 sg13g2_fill_2 FILLER_33_820 ();
 sg13g2_fill_1 FILLER_33_822 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_4 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_34_390 ();
 sg13g2_fill_1 FILLER_34_426 ();
 sg13g2_decap_4 FILLER_34_454 ();
 sg13g2_decap_4 FILLER_34_510 ();
 sg13g2_fill_1 FILLER_34_514 ();
 sg13g2_fill_1 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_540 ();
 sg13g2_fill_2 FILLER_34_547 ();
 sg13g2_decap_4 FILLER_34_553 ();
 sg13g2_fill_1 FILLER_34_557 ();
 sg13g2_decap_8 FILLER_34_585 ();
 sg13g2_decap_8 FILLER_34_592 ();
 sg13g2_fill_2 FILLER_34_599 ();
 sg13g2_fill_2 FILLER_34_610 ();
 sg13g2_decap_4 FILLER_34_634 ();
 sg13g2_fill_1 FILLER_34_638 ();
 sg13g2_decap_8 FILLER_34_643 ();
 sg13g2_decap_8 FILLER_34_650 ();
 sg13g2_decap_8 FILLER_34_662 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_fill_1 FILLER_34_676 ();
 sg13g2_fill_1 FILLER_34_704 ();
 sg13g2_decap_4 FILLER_34_749 ();
 sg13g2_fill_1 FILLER_34_753 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_4 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_35_433 ();
 sg13g2_decap_8 FILLER_35_440 ();
 sg13g2_decap_4 FILLER_35_493 ();
 sg13g2_fill_1 FILLER_35_497 ();
 sg13g2_fill_2 FILLER_35_529 ();
 sg13g2_decap_4 FILLER_35_563 ();
 sg13g2_decap_8 FILLER_35_577 ();
 sg13g2_decap_4 FILLER_35_584 ();
 sg13g2_fill_1 FILLER_35_588 ();
 sg13g2_fill_2 FILLER_35_621 ();
 sg13g2_decap_8 FILLER_35_650 ();
 sg13g2_decap_4 FILLER_35_662 ();
 sg13g2_fill_2 FILLER_35_666 ();
 sg13g2_fill_1 FILLER_35_681 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_fill_2 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_699 ();
 sg13g2_fill_2 FILLER_35_706 ();
 sg13g2_fill_2 FILLER_35_712 ();
 sg13g2_fill_1 FILLER_35_714 ();
 sg13g2_decap_4 FILLER_35_724 ();
 sg13g2_fill_1 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_4 FILLER_35_753 ();
 sg13g2_fill_2 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_fill_2 FILLER_35_770 ();
 sg13g2_fill_1 FILLER_35_772 ();
 sg13g2_decap_8 FILLER_35_783 ();
 sg13g2_fill_2 FILLER_35_790 ();
 sg13g2_fill_1 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_4 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_38 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_decap_8 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_59 ();
 sg13g2_decap_8 FILLER_36_66 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_decap_8 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_87 ();
 sg13g2_decap_8 FILLER_36_94 ();
 sg13g2_decap_8 FILLER_36_101 ();
 sg13g2_decap_8 FILLER_36_108 ();
 sg13g2_decap_8 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_122 ();
 sg13g2_decap_8 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_decap_8 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_4 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_476 ();
 sg13g2_decap_4 FILLER_36_482 ();
 sg13g2_fill_2 FILLER_36_486 ();
 sg13g2_decap_8 FILLER_36_492 ();
 sg13g2_decap_4 FILLER_36_499 ();
 sg13g2_fill_1 FILLER_36_503 ();
 sg13g2_decap_8 FILLER_36_523 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_583 ();
 sg13g2_decap_4 FILLER_36_588 ();
 sg13g2_fill_2 FILLER_36_592 ();
 sg13g2_decap_4 FILLER_36_598 ();
 sg13g2_decap_4 FILLER_36_632 ();
 sg13g2_fill_2 FILLER_36_636 ();
 sg13g2_fill_2 FILLER_36_675 ();
 sg13g2_decap_8 FILLER_36_708 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_fill_2 FILLER_36_722 ();
 sg13g2_fill_2 FILLER_36_734 ();
 sg13g2_fill_1 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_decap_4 FILLER_36_771 ();
 sg13g2_fill_2 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_4 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_fill_2 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_440 ();
 sg13g2_decap_4 FILLER_37_447 ();
 sg13g2_fill_1 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_460 ();
 sg13g2_fill_2 FILLER_37_466 ();
 sg13g2_decap_8 FILLER_37_478 ();
 sg13g2_decap_8 FILLER_37_485 ();
 sg13g2_decap_8 FILLER_37_492 ();
 sg13g2_decap_8 FILLER_37_499 ();
 sg13g2_decap_8 FILLER_37_506 ();
 sg13g2_fill_1 FILLER_37_513 ();
 sg13g2_decap_8 FILLER_37_531 ();
 sg13g2_decap_4 FILLER_37_538 ();
 sg13g2_fill_2 FILLER_37_542 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_fill_1 FILLER_37_578 ();
 sg13g2_decap_8 FILLER_37_606 ();
 sg13g2_decap_8 FILLER_37_631 ();
 sg13g2_decap_4 FILLER_37_638 ();
 sg13g2_fill_2 FILLER_37_642 ();
 sg13g2_decap_8 FILLER_37_648 ();
 sg13g2_fill_2 FILLER_37_655 ();
 sg13g2_fill_1 FILLER_37_657 ();
 sg13g2_decap_8 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_675 ();
 sg13g2_decap_8 FILLER_37_682 ();
 sg13g2_decap_8 FILLER_37_689 ();
 sg13g2_fill_2 FILLER_37_696 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_fill_2 FILLER_37_756 ();
 sg13g2_fill_1 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_2 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_424 ();
 sg13g2_decap_8 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_38_436 ();
 sg13g2_fill_2 FILLER_38_443 ();
 sg13g2_fill_1 FILLER_38_445 ();
 sg13g2_fill_2 FILLER_38_504 ();
 sg13g2_fill_2 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_554 ();
 sg13g2_fill_1 FILLER_38_561 ();
 sg13g2_fill_2 FILLER_38_572 ();
 sg13g2_decap_8 FILLER_38_587 ();
 sg13g2_decap_8 FILLER_38_594 ();
 sg13g2_fill_1 FILLER_38_601 ();
 sg13g2_decap_4 FILLER_38_662 ();
 sg13g2_fill_1 FILLER_38_666 ();
 sg13g2_decap_4 FILLER_38_708 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_fill_1 FILLER_38_745 ();
 sg13g2_decap_8 FILLER_38_750 ();
 sg13g2_decap_4 FILLER_38_757 ();
 sg13g2_fill_2 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_fill_2 FILLER_38_774 ();
 sg13g2_fill_1 FILLER_38_776 ();
 sg13g2_fill_1 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_4 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_fill_2 FILLER_39_413 ();
 sg13g2_decap_4 FILLER_39_423 ();
 sg13g2_decap_4 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_450 ();
 sg13g2_decap_8 FILLER_39_457 ();
 sg13g2_fill_1 FILLER_39_469 ();
 sg13g2_fill_2 FILLER_39_479 ();
 sg13g2_fill_1 FILLER_39_481 ();
 sg13g2_decap_4 FILLER_39_486 ();
 sg13g2_fill_2 FILLER_39_490 ();
 sg13g2_fill_1 FILLER_39_519 ();
 sg13g2_fill_1 FILLER_39_524 ();
 sg13g2_decap_8 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_548 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_fill_2 FILLER_39_560 ();
 sg13g2_fill_2 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_583 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_fill_2 FILLER_39_595 ();
 sg13g2_decap_4 FILLER_39_640 ();
 sg13g2_fill_2 FILLER_39_644 ();
 sg13g2_fill_2 FILLER_39_678 ();
 sg13g2_fill_2 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_690 ();
 sg13g2_decap_8 FILLER_39_697 ();
 sg13g2_fill_1 FILLER_39_704 ();
 sg13g2_decap_4 FILLER_39_768 ();
 sg13g2_fill_1 FILLER_39_772 ();
 sg13g2_fill_2 FILLER_39_783 ();
 sg13g2_fill_1 FILLER_39_785 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_fill_1 FILLER_40_501 ();
 sg13g2_decap_8 FILLER_40_535 ();
 sg13g2_fill_2 FILLER_40_542 ();
 sg13g2_fill_2 FILLER_40_571 ();
 sg13g2_fill_1 FILLER_40_573 ();
 sg13g2_decap_8 FILLER_40_606 ();
 sg13g2_fill_1 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_627 ();
 sg13g2_decap_4 FILLER_40_634 ();
 sg13g2_fill_1 FILLER_40_638 ();
 sg13g2_fill_2 FILLER_40_654 ();
 sg13g2_decap_8 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_667 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_decap_4 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_decap_4 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_fill_1 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_747 ();
 sg13g2_decap_4 FILLER_40_754 ();
 sg13g2_fill_2 FILLER_40_758 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_fill_1 FILLER_40_794 ();
 sg13g2_fill_1 FILLER_40_799 ();
 sg13g2_decap_8 FILLER_40_808 ();
 sg13g2_decap_8 FILLER_40_815 ();
 sg13g2_fill_1 FILLER_40_822 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_4 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_417 ();
 sg13g2_decap_8 FILLER_41_422 ();
 sg13g2_decap_4 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_41_433 ();
 sg13g2_fill_1 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_485 ();
 sg13g2_decap_4 FILLER_41_492 ();
 sg13g2_fill_1 FILLER_41_496 ();
 sg13g2_fill_2 FILLER_41_524 ();
 sg13g2_decap_4 FILLER_41_553 ();
 sg13g2_decap_4 FILLER_41_567 ();
 sg13g2_fill_2 FILLER_41_571 ();
 sg13g2_decap_8 FILLER_41_577 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_fill_1 FILLER_41_598 ();
 sg13g2_fill_2 FILLER_41_613 ();
 sg13g2_fill_1 FILLER_41_620 ();
 sg13g2_decap_4 FILLER_41_716 ();
 sg13g2_fill_1 FILLER_41_730 ();
 sg13g2_fill_2 FILLER_41_736 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_fill_2 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_769 ();
 sg13g2_decap_8 FILLER_41_776 ();
 sg13g2_decap_4 FILLER_41_788 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_4 FILLER_42_448 ();
 sg13g2_fill_1 FILLER_42_452 ();
 sg13g2_decap_8 FILLER_42_457 ();
 sg13g2_fill_2 FILLER_42_464 ();
 sg13g2_fill_1 FILLER_42_466 ();
 sg13g2_fill_2 FILLER_42_529 ();
 sg13g2_decap_8 FILLER_42_535 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_fill_2 FILLER_42_549 ();
 sg13g2_decap_4 FILLER_42_556 ();
 sg13g2_fill_2 FILLER_42_560 ();
 sg13g2_fill_1 FILLER_42_598 ();
 sg13g2_decap_8 FILLER_42_635 ();
 sg13g2_fill_2 FILLER_42_642 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_fill_1 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_decap_4 FILLER_42_705 ();
 sg13g2_fill_1 FILLER_42_709 ();
 sg13g2_fill_2 FILLER_42_742 ();
 sg13g2_fill_1 FILLER_42_744 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_fill_2 FILLER_42_820 ();
 sg13g2_fill_1 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_fill_2 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_489 ();
 sg13g2_decap_4 FILLER_43_496 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_fill_2 FILLER_43_530 ();
 sg13g2_fill_2 FILLER_43_573 ();
 sg13g2_fill_1 FILLER_43_575 ();
 sg13g2_decap_8 FILLER_43_580 ();
 sg13g2_decap_8 FILLER_43_587 ();
 sg13g2_fill_2 FILLER_43_594 ();
 sg13g2_fill_1 FILLER_43_596 ();
 sg13g2_decap_8 FILLER_43_610 ();
 sg13g2_decap_8 FILLER_43_617 ();
 sg13g2_decap_8 FILLER_43_624 ();
 sg13g2_decap_8 FILLER_43_631 ();
 sg13g2_fill_2 FILLER_43_638 ();
 sg13g2_decap_8 FILLER_43_653 ();
 sg13g2_decap_8 FILLER_43_660 ();
 sg13g2_decap_8 FILLER_43_667 ();
 sg13g2_decap_4 FILLER_43_674 ();
 sg13g2_decap_8 FILLER_43_710 ();
 sg13g2_fill_2 FILLER_43_717 ();
 sg13g2_fill_1 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_724 ();
 sg13g2_decap_8 FILLER_43_731 ();
 sg13g2_decap_4 FILLER_43_738 ();
 sg13g2_fill_1 FILLER_43_742 ();
 sg13g2_fill_2 FILLER_43_748 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_4 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_772 ();
 sg13g2_decap_4 FILLER_43_777 ();
 sg13g2_fill_1 FILLER_43_781 ();
 sg13g2_fill_1 FILLER_43_797 ();
 sg13g2_fill_1 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_808 ();
 sg13g2_decap_8 FILLER_43_815 ();
 sg13g2_fill_1 FILLER_43_822 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_fill_1 FILLER_44_517 ();
 sg13g2_decap_4 FILLER_44_528 ();
 sg13g2_fill_1 FILLER_44_532 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_decap_4 FILLER_44_549 ();
 sg13g2_fill_2 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_4 FILLER_44_567 ();
 sg13g2_fill_1 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_582 ();
 sg13g2_fill_2 FILLER_44_589 ();
 sg13g2_fill_1 FILLER_44_591 ();
 sg13g2_decap_8 FILLER_44_624 ();
 sg13g2_decap_4 FILLER_44_631 ();
 sg13g2_fill_2 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_642 ();
 sg13g2_fill_1 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_677 ();
 sg13g2_decap_4 FILLER_44_684 ();
 sg13g2_decap_8 FILLER_44_723 ();
 sg13g2_fill_1 FILLER_44_730 ();
 sg13g2_decap_8 FILLER_44_776 ();
 sg13g2_fill_2 FILLER_44_783 ();
 sg13g2_decap_8 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_fill_1 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_fill_2 FILLER_45_476 ();
 sg13g2_fill_1 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_488 ();
 sg13g2_fill_2 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_544 ();
 sg13g2_decap_8 FILLER_45_551 ();
 sg13g2_decap_8 FILLER_45_558 ();
 sg13g2_decap_8 FILLER_45_606 ();
 sg13g2_fill_2 FILLER_45_613 ();
 sg13g2_fill_1 FILLER_45_615 ();
 sg13g2_fill_2 FILLER_45_653 ();
 sg13g2_decap_8 FILLER_45_659 ();
 sg13g2_fill_1 FILLER_45_666 ();
 sg13g2_decap_8 FILLER_45_671 ();
 sg13g2_fill_1 FILLER_45_678 ();
 sg13g2_decap_4 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_fill_2 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_508 ();
 sg13g2_decap_4 FILLER_46_515 ();
 sg13g2_fill_2 FILLER_46_519 ();
 sg13g2_fill_1 FILLER_46_525 ();
 sg13g2_fill_1 FILLER_46_530 ();
 sg13g2_decap_8 FILLER_46_562 ();
 sg13g2_fill_2 FILLER_46_569 ();
 sg13g2_fill_1 FILLER_46_571 ();
 sg13g2_fill_2 FILLER_46_584 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_decap_8 FILLER_46_598 ();
 sg13g2_fill_2 FILLER_46_605 ();
 sg13g2_fill_1 FILLER_46_607 ();
 sg13g2_decap_8 FILLER_46_613 ();
 sg13g2_fill_1 FILLER_46_620 ();
 sg13g2_decap_8 FILLER_46_625 ();
 sg13g2_decap_4 FILLER_46_632 ();
 sg13g2_fill_1 FILLER_46_636 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_fill_1 FILLER_46_661 ();
 sg13g2_decap_8 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_701 ();
 sg13g2_decap_8 FILLER_46_708 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_4 FILLER_46_731 ();
 sg13g2_fill_2 FILLER_46_740 ();
 sg13g2_fill_2 FILLER_46_747 ();
 sg13g2_fill_1 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_768 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_fill_2 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_784 ();
 sg13g2_fill_2 FILLER_46_795 ();
 sg13g2_fill_2 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_4 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_4 FILLER_47_560 ();
 sg13g2_fill_1 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_579 ();
 sg13g2_decap_8 FILLER_47_626 ();
 sg13g2_fill_2 FILLER_47_633 ();
 sg13g2_decap_4 FILLER_47_645 ();
 sg13g2_fill_2 FILLER_47_649 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_4 FILLER_47_672 ();
 sg13g2_fill_2 FILLER_47_676 ();
 sg13g2_fill_1 FILLER_47_705 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_fill_2 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_fill_1 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_fill_2 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_691 ();
 sg13g2_fill_2 FILLER_48_711 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_4 FILLER_48_747 ();
 sg13g2_fill_1 FILLER_48_766 ();
 sg13g2_fill_2 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_fill_2 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_fill_2 FILLER_49_564 ();
 sg13g2_decap_8 FILLER_49_570 ();
 sg13g2_decap_8 FILLER_49_577 ();
 sg13g2_fill_1 FILLER_49_584 ();
 sg13g2_decap_4 FILLER_49_589 ();
 sg13g2_fill_1 FILLER_49_593 ();
 sg13g2_decap_8 FILLER_49_624 ();
 sg13g2_decap_4 FILLER_49_631 ();
 sg13g2_fill_2 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_fill_1 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_687 ();
 sg13g2_fill_1 FILLER_49_694 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_fill_1 FILLER_49_714 ();
 sg13g2_fill_2 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_4 FILLER_49_788 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_4 FILLER_49_817 ();
 sg13g2_fill_2 FILLER_49_821 ();
 assign uio_oe[0] = net455;
 assign uio_oe[1] = net456;
 assign uio_oe[2] = net457;
 assign uio_oe[3] = net458;
 assign uio_oe[4] = net459;
 assign uio_oe[5] = net460;
 assign uio_oe[6] = net461;
 assign uio_oe[7] = net462;
endmodule
