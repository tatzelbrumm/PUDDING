* Extracted by KLayout with SG13G2 LVS runset on : 27/08/2025 22:00

.SUBCKT CASCODEDRIVE
M$1 \$3 \$4 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$2 \$1 \$3 \$4 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$3 \$3 \$5 \$2 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p PS=1.75u
+ PD=0.68u
M$4 \$2 \$6 \$4 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p PS=0.68u
+ PD=1.75u
M$5 \$7 \$3 \$8 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u
+ PD=0.68u
M$6 \$8 \$4 \$2 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u
+ PD=1.28u
.ENDS CASCODEDRIVE
