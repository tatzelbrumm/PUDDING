magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771280484
<< metal1 >>
rect 576 38576 79584 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79584 38576
rect 576 38512 79584 38536
rect 63435 38324 63477 38333
rect 63435 38284 63436 38324
rect 63476 38284 63477 38324
rect 63435 38275 63477 38284
rect 63531 38240 63573 38249
rect 63339 38229 63381 38238
rect 63339 38189 63340 38229
rect 63380 38189 63381 38229
rect 63531 38200 63532 38240
rect 63572 38200 63573 38240
rect 63531 38191 63573 38200
rect 63619 38240 63677 38241
rect 63619 38200 63628 38240
rect 63668 38200 63677 38240
rect 63619 38199 63677 38200
rect 67467 38240 67509 38249
rect 67467 38200 67468 38240
rect 67508 38200 67509 38240
rect 67467 38191 67509 38200
rect 67659 38240 67701 38249
rect 67659 38200 67660 38240
rect 67700 38200 67701 38240
rect 67659 38191 67701 38200
rect 67747 38240 67805 38241
rect 67747 38200 67756 38240
rect 67796 38200 67805 38240
rect 67747 38199 67805 38200
rect 67947 38240 67989 38249
rect 67947 38200 67948 38240
rect 67988 38200 67989 38240
rect 67947 38191 67989 38200
rect 68043 38240 68085 38249
rect 68043 38200 68044 38240
rect 68084 38200 68085 38240
rect 68043 38191 68085 38200
rect 68139 38240 68181 38249
rect 68139 38200 68140 38240
rect 68180 38200 68181 38240
rect 68139 38191 68181 38200
rect 68235 38240 68277 38249
rect 68235 38200 68236 38240
rect 68276 38200 68277 38240
rect 68235 38191 68277 38200
rect 69291 38240 69333 38249
rect 69291 38200 69292 38240
rect 69332 38200 69333 38240
rect 69291 38191 69333 38200
rect 70635 38240 70677 38249
rect 70635 38200 70636 38240
rect 70676 38200 70677 38240
rect 70635 38191 70677 38200
rect 71019 38240 71061 38249
rect 71019 38200 71020 38240
rect 71060 38200 71061 38240
rect 71019 38191 71061 38200
rect 71203 38240 71261 38241
rect 71203 38200 71212 38240
rect 71252 38200 71261 38240
rect 71203 38199 71261 38200
rect 74275 38240 74333 38241
rect 74275 38200 74284 38240
rect 74324 38200 74333 38240
rect 74275 38199 74333 38200
rect 75235 38240 75293 38241
rect 75235 38200 75244 38240
rect 75284 38200 75293 38240
rect 75235 38199 75293 38200
rect 76963 38240 77021 38241
rect 76963 38200 76972 38240
rect 77012 38200 77021 38240
rect 76963 38199 77021 38200
rect 77259 38240 77301 38249
rect 77259 38200 77260 38240
rect 77300 38200 77301 38240
rect 77259 38191 77301 38200
rect 77355 38240 77397 38249
rect 77355 38200 77356 38240
rect 77396 38200 77397 38240
rect 77355 38191 77397 38200
rect 63339 38180 63381 38189
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 58339 38156 58397 38157
rect 58339 38116 58348 38156
rect 58388 38116 58397 38156
rect 58339 38115 58397 38116
rect 58915 38156 58973 38157
rect 58915 38116 58924 38156
rect 58964 38116 58973 38156
rect 58915 38115 58973 38116
rect 59299 38156 59357 38157
rect 59299 38116 59308 38156
rect 59348 38116 59357 38156
rect 59299 38115 59357 38116
rect 67075 38156 67133 38157
rect 67075 38116 67084 38156
rect 67124 38116 67133 38156
rect 67075 38115 67133 38116
rect 56907 38072 56949 38081
rect 56907 38032 56908 38072
rect 56948 38032 56949 38072
rect 56907 38023 56949 38032
rect 58539 38072 58581 38081
rect 58539 38032 58540 38072
rect 58580 38032 58581 38072
rect 58539 38023 58581 38032
rect 61611 38072 61653 38081
rect 61611 38032 61612 38072
rect 61652 38032 61653 38072
rect 61611 38023 61653 38032
rect 64203 38072 64245 38081
rect 64203 38032 64204 38072
rect 64244 38032 64245 38072
rect 64203 38023 64245 38032
rect 66507 38072 66549 38081
rect 66507 38032 66508 38072
rect 66548 38032 66549 38072
rect 66507 38023 66549 38032
rect 71403 38072 71445 38081
rect 71403 38032 71404 38072
rect 71444 38032 71445 38072
rect 71403 38023 71445 38032
rect 71979 38072 72021 38081
rect 71979 38032 71980 38072
rect 72020 38032 72021 38072
rect 71979 38023 72021 38032
rect 75915 38072 75957 38081
rect 75915 38032 75916 38072
rect 75956 38032 75957 38072
rect 75915 38023 75957 38032
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 58731 37988 58773 37997
rect 58731 37948 58732 37988
rect 58772 37948 58773 37988
rect 58731 37939 58773 37948
rect 59115 37988 59157 37997
rect 59115 37948 59116 37988
rect 59156 37948 59157 37988
rect 59115 37939 59157 37948
rect 67275 37988 67317 37997
rect 67275 37948 67276 37988
rect 67316 37948 67317 37988
rect 67275 37939 67317 37948
rect 67467 37988 67509 37997
rect 67467 37948 67468 37988
rect 67508 37948 67509 37988
rect 67467 37939 67509 37948
rect 69099 37988 69141 37997
rect 69099 37948 69100 37988
rect 69140 37948 69141 37988
rect 69099 37939 69141 37948
rect 70059 37988 70101 37997
rect 70059 37948 70060 37988
rect 70100 37948 70101 37988
rect 70059 37939 70101 37948
rect 71115 37988 71157 37997
rect 71115 37948 71116 37988
rect 71156 37948 71157 37988
rect 71115 37939 71157 37948
rect 77635 37988 77693 37989
rect 77635 37948 77644 37988
rect 77684 37948 77693 37988
rect 77635 37947 77693 37948
rect 576 37820 79584 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79584 37820
rect 576 37756 79584 37780
rect 55179 37568 55221 37577
rect 55179 37528 55180 37568
rect 55220 37528 55221 37568
rect 55179 37519 55221 37528
rect 59787 37568 59829 37577
rect 59787 37528 59788 37568
rect 59828 37528 59829 37568
rect 59787 37519 59829 37528
rect 74283 37568 74325 37577
rect 74283 37528 74284 37568
rect 74324 37528 74325 37568
rect 74283 37519 74325 37528
rect 78411 37568 78453 37577
rect 78411 37528 78412 37568
rect 78452 37528 78453 37568
rect 78411 37519 78453 37528
rect 55755 37400 55797 37409
rect 55755 37360 55756 37400
rect 55796 37360 55797 37400
rect 55755 37351 55797 37360
rect 55947 37400 55989 37409
rect 55947 37360 55948 37400
rect 55988 37360 55989 37400
rect 55947 37351 55989 37360
rect 56035 37400 56093 37401
rect 56035 37360 56044 37400
rect 56084 37360 56093 37400
rect 56035 37359 56093 37360
rect 57379 37400 57437 37401
rect 57379 37360 57388 37400
rect 57428 37360 57437 37400
rect 57379 37359 57437 37360
rect 58243 37400 58301 37401
rect 58243 37360 58252 37400
rect 58292 37360 58301 37400
rect 58243 37359 58301 37360
rect 58827 37400 58869 37409
rect 58827 37360 58828 37400
rect 58868 37360 58869 37400
rect 58827 37351 58869 37360
rect 58923 37400 58965 37409
rect 58923 37360 58924 37400
rect 58964 37360 58965 37400
rect 58923 37351 58965 37360
rect 59019 37400 59061 37409
rect 59019 37360 59020 37400
rect 59060 37360 59061 37400
rect 59019 37351 59061 37360
rect 59115 37400 59157 37409
rect 59115 37360 59116 37400
rect 59156 37360 59157 37400
rect 59115 37351 59157 37360
rect 59307 37400 59349 37409
rect 59307 37360 59308 37400
rect 59348 37360 59349 37400
rect 59307 37351 59349 37360
rect 59499 37400 59541 37409
rect 59499 37360 59500 37400
rect 59540 37360 59541 37400
rect 59499 37351 59541 37360
rect 59587 37400 59645 37401
rect 59587 37360 59596 37400
rect 59636 37360 59645 37400
rect 59587 37359 59645 37360
rect 60171 37400 60213 37409
rect 60171 37360 60172 37400
rect 60212 37360 60213 37400
rect 60171 37351 60213 37360
rect 60363 37400 60405 37409
rect 60363 37360 60364 37400
rect 60404 37360 60405 37400
rect 60451 37402 60509 37403
rect 60451 37362 60460 37402
rect 60500 37362 60509 37402
rect 60451 37361 60509 37362
rect 61507 37400 61565 37401
rect 60363 37351 60405 37360
rect 61507 37360 61516 37400
rect 61556 37360 61565 37400
rect 61507 37359 61565 37360
rect 62371 37400 62429 37401
rect 62371 37360 62380 37400
rect 62420 37360 62429 37400
rect 62371 37359 62429 37360
rect 63723 37400 63765 37409
rect 63723 37360 63724 37400
rect 63764 37360 63765 37400
rect 63723 37351 63765 37360
rect 64099 37400 64157 37401
rect 64099 37360 64108 37400
rect 64148 37360 64157 37400
rect 64099 37359 64157 37360
rect 64963 37400 65021 37401
rect 64963 37360 64972 37400
rect 65012 37360 65021 37400
rect 64963 37359 65021 37360
rect 66315 37400 66357 37409
rect 66315 37360 66316 37400
rect 66356 37360 66357 37400
rect 66315 37351 66357 37360
rect 66691 37400 66749 37401
rect 66691 37360 66700 37400
rect 66740 37360 66749 37400
rect 66691 37359 66749 37360
rect 67555 37400 67613 37401
rect 67555 37360 67564 37400
rect 67604 37360 67613 37400
rect 67555 37359 67613 37360
rect 69571 37400 69629 37401
rect 69571 37360 69580 37400
rect 69620 37360 69629 37400
rect 69571 37359 69629 37360
rect 70435 37400 70493 37401
rect 70435 37360 70444 37400
rect 70484 37360 70493 37400
rect 70435 37359 70493 37360
rect 72843 37400 72885 37409
rect 72843 37360 72844 37400
rect 72884 37360 72885 37400
rect 72843 37351 72885 37360
rect 72939 37400 72981 37409
rect 72939 37360 72940 37400
rect 72980 37360 72981 37400
rect 72939 37351 72981 37360
rect 73035 37400 73077 37409
rect 73035 37360 73036 37400
rect 73076 37360 73077 37400
rect 73035 37351 73077 37360
rect 73131 37400 73173 37409
rect 73131 37360 73132 37400
rect 73172 37360 73173 37400
rect 73131 37351 73173 37360
rect 73323 37400 73365 37409
rect 73323 37360 73324 37400
rect 73364 37360 73365 37400
rect 73323 37351 73365 37360
rect 73515 37400 73557 37409
rect 73515 37360 73516 37400
rect 73556 37360 73557 37400
rect 73515 37351 73557 37360
rect 73603 37400 73661 37401
rect 73603 37360 73612 37400
rect 73652 37360 73661 37400
rect 73603 37359 73661 37360
rect 73803 37400 73845 37409
rect 73803 37360 73804 37400
rect 73844 37360 73845 37400
rect 73803 37351 73845 37360
rect 73995 37400 74037 37409
rect 73995 37360 73996 37400
rect 74036 37360 74037 37400
rect 73995 37351 74037 37360
rect 74083 37400 74141 37401
rect 74083 37360 74092 37400
rect 74132 37360 74141 37400
rect 74083 37359 74141 37360
rect 74283 37400 74325 37409
rect 74283 37360 74284 37400
rect 74324 37360 74325 37400
rect 74283 37351 74325 37360
rect 74475 37400 74517 37409
rect 74475 37360 74476 37400
rect 74516 37360 74517 37400
rect 74475 37351 74517 37360
rect 74563 37400 74621 37401
rect 74563 37360 74572 37400
rect 74612 37360 74621 37400
rect 74563 37359 74621 37360
rect 74955 37400 74997 37409
rect 74955 37360 74956 37400
rect 74996 37360 74997 37400
rect 74955 37351 74997 37360
rect 75051 37400 75093 37409
rect 75051 37360 75052 37400
rect 75092 37360 75093 37400
rect 75051 37351 75093 37360
rect 75147 37400 75189 37409
rect 75147 37360 75148 37400
rect 75188 37360 75189 37400
rect 75147 37351 75189 37360
rect 75811 37400 75869 37401
rect 75811 37360 75820 37400
rect 75860 37360 75869 37400
rect 75811 37359 75869 37360
rect 76675 37400 76733 37401
rect 76675 37360 76684 37400
rect 76724 37360 76733 37400
rect 76675 37359 76733 37360
rect 78019 37400 78077 37401
rect 78019 37360 78028 37400
rect 78068 37360 78077 37400
rect 78019 37359 78077 37360
rect 78219 37400 78261 37409
rect 78219 37360 78220 37400
rect 78260 37360 78261 37400
rect 78219 37351 78261 37360
rect 58635 37316 58677 37325
rect 58635 37276 58636 37316
rect 58676 37276 58677 37316
rect 58635 37267 58677 37276
rect 59403 37316 59445 37325
rect 59403 37276 59404 37316
rect 59444 37276 59445 37316
rect 59403 37267 59445 37276
rect 60267 37316 60309 37325
rect 60267 37276 60268 37316
rect 60308 37276 60309 37316
rect 60267 37267 60309 37276
rect 61131 37316 61173 37325
rect 61131 37276 61132 37316
rect 61172 37276 61173 37316
rect 61131 37267 61173 37276
rect 69195 37316 69237 37325
rect 69195 37276 69196 37316
rect 69236 37276 69237 37316
rect 69195 37267 69237 37276
rect 75435 37316 75477 37325
rect 75435 37276 75436 37316
rect 75476 37276 75477 37316
rect 75435 37267 75477 37276
rect 78123 37316 78165 37325
rect 78123 37276 78124 37316
rect 78164 37276 78165 37316
rect 78123 37267 78165 37276
rect 55843 37232 55901 37233
rect 55843 37192 55852 37232
rect 55892 37192 55901 37232
rect 55843 37191 55901 37192
rect 56227 37232 56285 37233
rect 56227 37192 56236 37232
rect 56276 37192 56285 37232
rect 56227 37191 56285 37192
rect 63523 37232 63581 37233
rect 63523 37192 63532 37232
rect 63572 37192 63581 37232
rect 63523 37191 63581 37192
rect 66115 37232 66173 37233
rect 66115 37192 66124 37232
rect 66164 37192 66173 37232
rect 66115 37191 66173 37192
rect 68707 37232 68765 37233
rect 68707 37192 68716 37232
rect 68756 37192 68765 37232
rect 68707 37191 68765 37192
rect 71587 37232 71645 37233
rect 71587 37192 71596 37232
rect 71636 37192 71645 37232
rect 71587 37191 71645 37192
rect 73411 37232 73469 37233
rect 73411 37192 73420 37232
rect 73460 37192 73469 37232
rect 73411 37191 73469 37192
rect 73891 37232 73949 37233
rect 73891 37192 73900 37232
rect 73940 37192 73949 37232
rect 73891 37191 73949 37192
rect 75235 37232 75293 37233
rect 75235 37192 75244 37232
rect 75284 37192 75293 37232
rect 75235 37191 75293 37192
rect 77827 37232 77885 37233
rect 77827 37192 77836 37232
rect 77876 37192 77885 37232
rect 77827 37191 77885 37192
rect 576 37064 79584 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79584 37064
rect 576 37000 79584 37024
rect 62275 36896 62333 36897
rect 62275 36856 62284 36896
rect 62324 36856 62333 36896
rect 62275 36855 62333 36856
rect 67947 36896 67989 36905
rect 67947 36856 67948 36896
rect 67988 36856 67989 36896
rect 67947 36847 67989 36856
rect 79459 36896 79517 36897
rect 79459 36856 79468 36896
rect 79508 36856 79517 36896
rect 79459 36855 79517 36856
rect 54699 36812 54741 36821
rect 54699 36772 54700 36812
rect 54740 36772 54741 36812
rect 54699 36763 54741 36772
rect 58443 36812 58485 36821
rect 58443 36772 58444 36812
rect 58484 36772 58485 36812
rect 58443 36763 58485 36772
rect 63339 36812 63381 36821
rect 63339 36772 63340 36812
rect 63380 36772 63381 36812
rect 63339 36763 63381 36772
rect 63915 36812 63957 36821
rect 63915 36772 63916 36812
rect 63956 36772 63957 36812
rect 63915 36763 63957 36772
rect 64299 36812 64341 36821
rect 64299 36772 64300 36812
rect 64340 36772 64341 36812
rect 64299 36763 64341 36772
rect 73323 36812 73365 36821
rect 73323 36772 73324 36812
rect 73364 36772 73365 36812
rect 73323 36763 73365 36772
rect 73515 36812 73557 36821
rect 73515 36772 73516 36812
rect 73556 36772 73557 36812
rect 73515 36763 73557 36772
rect 55075 36728 55133 36729
rect 55075 36688 55084 36728
rect 55124 36688 55133 36728
rect 55075 36687 55133 36688
rect 55939 36728 55997 36729
rect 55939 36688 55948 36728
rect 55988 36688 55997 36728
rect 55939 36687 55997 36688
rect 57291 36728 57333 36737
rect 57291 36688 57292 36728
rect 57332 36688 57333 36728
rect 57291 36679 57333 36688
rect 57483 36728 57525 36737
rect 57483 36688 57484 36728
rect 57524 36688 57525 36728
rect 57483 36679 57525 36688
rect 57571 36728 57629 36729
rect 57571 36688 57580 36728
rect 57620 36688 57629 36728
rect 57571 36687 57629 36688
rect 58539 36728 58581 36737
rect 58539 36688 58540 36728
rect 58580 36688 58581 36728
rect 58539 36679 58581 36688
rect 58819 36728 58877 36729
rect 58819 36688 58828 36728
rect 58868 36688 58877 36728
rect 58819 36687 58877 36688
rect 59115 36728 59157 36737
rect 59115 36688 59116 36728
rect 59156 36688 59157 36728
rect 59115 36679 59157 36688
rect 59491 36728 59549 36729
rect 59491 36688 59500 36728
rect 59540 36688 59549 36728
rect 59491 36687 59549 36688
rect 60355 36728 60413 36729
rect 60355 36688 60364 36728
rect 60404 36688 60413 36728
rect 60355 36687 60413 36688
rect 61707 36728 61749 36737
rect 61707 36688 61708 36728
rect 61748 36688 61749 36728
rect 61707 36679 61749 36688
rect 61803 36728 61845 36737
rect 61803 36688 61804 36728
rect 61844 36688 61845 36728
rect 61803 36679 61845 36688
rect 61899 36728 61941 36737
rect 61899 36688 61900 36728
rect 61940 36688 61941 36728
rect 61899 36679 61941 36688
rect 61995 36728 62037 36737
rect 61995 36688 61996 36728
rect 62036 36688 62037 36728
rect 61995 36679 62037 36688
rect 62187 36728 62229 36737
rect 62187 36688 62188 36728
rect 62228 36688 62229 36728
rect 62187 36679 62229 36688
rect 62379 36728 62421 36737
rect 62379 36688 62380 36728
rect 62420 36688 62421 36728
rect 62379 36679 62421 36688
rect 62467 36728 62525 36729
rect 62467 36688 62476 36728
rect 62516 36688 62525 36728
rect 62467 36687 62525 36688
rect 62947 36728 63005 36729
rect 62947 36688 62956 36728
rect 62996 36688 63005 36728
rect 62947 36687 63005 36688
rect 63243 36728 63285 36737
rect 63243 36688 63244 36728
rect 63284 36688 63285 36728
rect 63243 36679 63285 36688
rect 63819 36728 63861 36737
rect 63819 36688 63820 36728
rect 63860 36688 63861 36728
rect 63819 36679 63861 36688
rect 64003 36728 64061 36729
rect 64003 36688 64012 36728
rect 64052 36688 64061 36728
rect 64003 36687 64061 36688
rect 64195 36728 64253 36729
rect 64195 36688 64204 36728
rect 64244 36688 64253 36728
rect 64195 36687 64253 36688
rect 64395 36728 64437 36737
rect 64395 36688 64396 36728
rect 64436 36688 64437 36728
rect 64395 36679 64437 36688
rect 66507 36728 66549 36737
rect 66507 36688 66508 36728
rect 66548 36688 66549 36728
rect 66507 36679 66549 36688
rect 66699 36728 66741 36737
rect 66699 36688 66700 36728
rect 66740 36688 66741 36728
rect 66699 36679 66741 36688
rect 66787 36728 66845 36729
rect 66787 36688 66796 36728
rect 66836 36688 66845 36728
rect 66787 36687 66845 36688
rect 67179 36728 67221 36737
rect 67179 36688 67180 36728
rect 67220 36688 67221 36728
rect 67179 36679 67221 36688
rect 67371 36728 67413 36737
rect 67371 36688 67372 36728
rect 67412 36688 67413 36728
rect 67371 36679 67413 36688
rect 67459 36728 67517 36729
rect 67459 36688 67468 36728
rect 67508 36688 67517 36728
rect 67459 36687 67517 36688
rect 68227 36728 68285 36729
rect 68227 36688 68236 36728
rect 68276 36688 68285 36728
rect 68227 36687 68285 36688
rect 68523 36728 68565 36737
rect 68523 36688 68524 36728
rect 68564 36688 68565 36728
rect 68523 36679 68565 36688
rect 68619 36728 68661 36737
rect 68619 36688 68620 36728
rect 68660 36688 68661 36728
rect 68619 36679 68661 36688
rect 69099 36728 69141 36737
rect 69099 36688 69100 36728
rect 69140 36688 69141 36728
rect 69099 36679 69141 36688
rect 69291 36728 69333 36737
rect 69291 36688 69292 36728
rect 69332 36688 69333 36728
rect 69291 36679 69333 36688
rect 69379 36728 69437 36729
rect 69379 36688 69388 36728
rect 69428 36688 69437 36728
rect 69379 36687 69437 36688
rect 69579 36728 69621 36737
rect 69579 36688 69580 36728
rect 69620 36688 69621 36728
rect 69579 36679 69621 36688
rect 69763 36728 69821 36729
rect 69763 36688 69772 36728
rect 69812 36688 69821 36728
rect 69763 36687 69821 36688
rect 72067 36728 72125 36729
rect 72067 36688 72076 36728
rect 72116 36688 72125 36728
rect 72067 36687 72125 36688
rect 72931 36728 72989 36729
rect 72931 36688 72940 36728
rect 72980 36688 72989 36728
rect 72931 36687 72989 36688
rect 73891 36728 73949 36729
rect 73891 36688 73900 36728
rect 73940 36688 73949 36728
rect 73891 36687 73949 36688
rect 74755 36728 74813 36729
rect 74755 36688 74764 36728
rect 74804 36688 74813 36728
rect 74755 36687 74813 36688
rect 76107 36728 76149 36737
rect 76107 36688 76108 36728
rect 76148 36688 76149 36728
rect 76107 36679 76149 36688
rect 76299 36728 76341 36737
rect 76299 36688 76300 36728
rect 76340 36688 76341 36728
rect 76299 36679 76341 36688
rect 76387 36728 76445 36729
rect 76387 36688 76396 36728
rect 76436 36688 76445 36728
rect 76387 36687 76445 36688
rect 76587 36728 76629 36737
rect 76587 36688 76588 36728
rect 76628 36688 76629 36728
rect 76587 36679 76629 36688
rect 76779 36728 76821 36737
rect 76779 36688 76780 36728
rect 76820 36688 76821 36728
rect 76779 36679 76821 36688
rect 76867 36728 76925 36729
rect 76867 36688 76876 36728
rect 76916 36688 76925 36728
rect 76867 36687 76925 36688
rect 77067 36728 77109 36737
rect 77067 36688 77068 36728
rect 77108 36688 77109 36728
rect 77067 36679 77109 36688
rect 77443 36728 77501 36729
rect 77443 36688 77452 36728
rect 77492 36688 77501 36728
rect 77443 36687 77501 36688
rect 78307 36728 78365 36729
rect 78307 36688 78316 36728
rect 78356 36688 78365 36728
rect 78307 36687 78365 36688
rect 67747 36644 67805 36645
rect 67747 36604 67756 36644
rect 67796 36604 67805 36644
rect 67747 36603 67805 36604
rect 52491 36560 52533 36569
rect 52491 36520 52492 36560
rect 52532 36520 52533 36560
rect 52491 36511 52533 36520
rect 57291 36560 57333 36569
rect 57291 36520 57292 36560
rect 57332 36520 57333 36560
rect 57291 36511 57333 36520
rect 63619 36560 63677 36561
rect 63619 36520 63628 36560
rect 63668 36520 63677 36560
rect 63619 36519 63677 36520
rect 67179 36560 67221 36569
rect 67179 36520 67180 36560
rect 67220 36520 67221 36560
rect 67179 36511 67221 36520
rect 68899 36560 68957 36561
rect 68899 36520 68908 36560
rect 68948 36520 68957 36560
rect 68899 36519 68957 36520
rect 69675 36560 69717 36569
rect 69675 36520 69676 36560
rect 69716 36520 69717 36560
rect 69675 36511 69717 36520
rect 76107 36560 76149 36569
rect 76107 36520 76108 36560
rect 76148 36520 76149 36560
rect 76107 36511 76149 36520
rect 76587 36560 76629 36569
rect 76587 36520 76588 36560
rect 76628 36520 76629 36560
rect 76587 36511 76629 36520
rect 57091 36476 57149 36477
rect 57091 36436 57100 36476
rect 57140 36436 57149 36476
rect 57091 36435 57149 36436
rect 58147 36476 58205 36477
rect 58147 36436 58156 36476
rect 58196 36436 58205 36476
rect 58147 36435 58205 36436
rect 61507 36476 61565 36477
rect 61507 36436 61516 36476
rect 61556 36436 61565 36476
rect 61507 36435 61565 36436
rect 66507 36476 66549 36485
rect 66507 36436 66508 36476
rect 66548 36436 66549 36476
rect 66507 36427 66549 36436
rect 67947 36476 67989 36485
rect 67947 36436 67948 36476
rect 67988 36436 67989 36476
rect 67947 36427 67989 36436
rect 69099 36476 69141 36485
rect 69099 36436 69100 36476
rect 69140 36436 69141 36476
rect 69099 36427 69141 36436
rect 70915 36476 70973 36477
rect 70915 36436 70924 36476
rect 70964 36436 70973 36476
rect 70915 36435 70973 36436
rect 75907 36476 75965 36477
rect 75907 36436 75916 36476
rect 75956 36436 75965 36476
rect 75907 36435 75965 36436
rect 576 36308 79584 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79584 36308
rect 576 36244 79584 36268
rect 62283 36140 62325 36149
rect 62283 36100 62284 36140
rect 62324 36100 62325 36140
rect 62283 36091 62325 36100
rect 73803 36140 73845 36149
rect 73803 36100 73804 36140
rect 73844 36100 73845 36140
rect 73803 36091 73845 36100
rect 77547 36140 77589 36149
rect 77547 36100 77548 36140
rect 77588 36100 77589 36140
rect 77547 36091 77589 36100
rect 49227 36056 49269 36065
rect 49227 36016 49228 36056
rect 49268 36016 49269 36056
rect 49227 36007 49269 36016
rect 60363 36056 60405 36065
rect 60363 36016 60364 36056
rect 60404 36016 60405 36056
rect 60363 36007 60405 36016
rect 69483 36056 69525 36065
rect 69483 36016 69484 36056
rect 69524 36016 69525 36056
rect 69483 36007 69525 36016
rect 73507 36056 73565 36057
rect 73507 36016 73516 36056
rect 73556 36016 73565 36056
rect 73507 36015 73565 36016
rect 74091 36056 74133 36065
rect 74091 36016 74092 36056
rect 74132 36016 74133 36056
rect 74091 36007 74133 36016
rect 77835 36056 77877 36065
rect 77835 36016 77836 36056
rect 77876 36016 77877 36056
rect 77835 36007 77877 36016
rect 50947 35972 51005 35973
rect 50947 35932 50956 35972
rect 50996 35932 51005 35972
rect 50947 35931 51005 35932
rect 57091 35972 57149 35973
rect 57091 35932 57100 35972
rect 57140 35932 57149 35972
rect 57091 35931 57149 35932
rect 51339 35888 51381 35897
rect 51339 35848 51340 35888
rect 51380 35848 51381 35888
rect 51339 35839 51381 35848
rect 51523 35888 51581 35889
rect 51523 35848 51532 35888
rect 51572 35848 51581 35888
rect 51523 35847 51581 35848
rect 52387 35888 52445 35889
rect 52387 35848 52396 35888
rect 52436 35848 52445 35888
rect 52387 35847 52445 35848
rect 53276 35888 53334 35889
rect 53276 35848 53285 35888
rect 53325 35848 53334 35888
rect 53276 35847 53334 35848
rect 55555 35888 55613 35889
rect 55555 35848 55564 35888
rect 55604 35848 55613 35888
rect 55555 35847 55613 35848
rect 55659 35888 55701 35897
rect 55659 35848 55660 35888
rect 55700 35848 55701 35888
rect 55659 35839 55701 35848
rect 55851 35888 55893 35897
rect 55851 35848 55852 35888
rect 55892 35848 55893 35888
rect 55851 35839 55893 35848
rect 56043 35888 56085 35897
rect 56043 35848 56044 35888
rect 56084 35848 56085 35888
rect 56043 35839 56085 35848
rect 56139 35888 56181 35897
rect 56139 35848 56140 35888
rect 56180 35848 56181 35888
rect 56139 35839 56181 35848
rect 56235 35888 56277 35897
rect 56235 35848 56236 35888
rect 56276 35848 56277 35888
rect 56235 35839 56277 35848
rect 56331 35888 56373 35897
rect 56331 35848 56332 35888
rect 56372 35848 56373 35888
rect 56331 35839 56373 35848
rect 56515 35888 56573 35889
rect 56515 35848 56524 35888
rect 56564 35848 56573 35888
rect 56515 35847 56573 35848
rect 56619 35888 56661 35897
rect 56619 35848 56620 35888
rect 56660 35848 56661 35888
rect 56619 35839 56661 35848
rect 56715 35888 56757 35897
rect 56715 35848 56716 35888
rect 56756 35848 56757 35888
rect 56715 35839 56757 35848
rect 58539 35888 58581 35897
rect 58539 35848 58540 35888
rect 58580 35848 58581 35888
rect 58539 35839 58581 35848
rect 58635 35888 58677 35897
rect 58635 35848 58636 35888
rect 58676 35848 58677 35888
rect 58635 35839 58677 35848
rect 58723 35888 58781 35889
rect 58723 35848 58732 35888
rect 58772 35848 58781 35888
rect 58723 35847 58781 35848
rect 58923 35888 58965 35897
rect 58923 35848 58924 35888
rect 58964 35848 58965 35888
rect 58923 35839 58965 35848
rect 59115 35888 59157 35897
rect 59115 35848 59116 35888
rect 59156 35848 59157 35888
rect 59115 35839 59157 35848
rect 59203 35888 59261 35889
rect 59203 35848 59212 35888
rect 59252 35848 59261 35888
rect 59203 35847 59261 35848
rect 59395 35888 59453 35889
rect 59395 35848 59404 35888
rect 59444 35848 59453 35888
rect 59395 35847 59453 35848
rect 59595 35888 59637 35897
rect 59595 35848 59596 35888
rect 59636 35848 59637 35888
rect 59595 35839 59637 35848
rect 61987 35888 62045 35889
rect 61987 35848 61996 35888
rect 62036 35848 62045 35888
rect 61987 35847 62045 35848
rect 62091 35888 62133 35897
rect 62091 35848 62092 35888
rect 62132 35848 62133 35888
rect 62091 35839 62133 35848
rect 62283 35888 62325 35897
rect 62283 35848 62284 35888
rect 62324 35848 62325 35888
rect 62283 35839 62325 35848
rect 64395 35888 64437 35897
rect 64395 35848 64396 35888
rect 64436 35848 64437 35888
rect 64395 35839 64437 35848
rect 64771 35888 64829 35889
rect 64771 35848 64780 35888
rect 64820 35848 64829 35888
rect 64771 35847 64829 35848
rect 65635 35888 65693 35889
rect 65635 35848 65644 35888
rect 65684 35848 65693 35888
rect 65635 35847 65693 35848
rect 66987 35888 67029 35897
rect 66987 35848 66988 35888
rect 67028 35848 67029 35888
rect 66987 35839 67029 35848
rect 67083 35888 67125 35897
rect 67083 35848 67084 35888
rect 67124 35848 67125 35888
rect 67083 35839 67125 35848
rect 67179 35888 67221 35897
rect 67179 35848 67180 35888
rect 67220 35848 67221 35888
rect 67179 35839 67221 35848
rect 67275 35888 67317 35897
rect 67275 35848 67276 35888
rect 67316 35848 67317 35888
rect 67275 35839 67317 35848
rect 69675 35888 69717 35897
rect 69675 35848 69676 35888
rect 69716 35848 69717 35888
rect 69675 35839 69717 35848
rect 69867 35888 69909 35897
rect 69867 35848 69868 35888
rect 69908 35848 69909 35888
rect 69867 35839 69909 35848
rect 69955 35888 70013 35889
rect 69955 35848 69964 35888
rect 70004 35848 70013 35888
rect 69955 35847 70013 35848
rect 71499 35888 71541 35897
rect 71499 35848 71500 35888
rect 71540 35848 71541 35888
rect 71499 35839 71541 35848
rect 71683 35888 71741 35889
rect 71683 35848 71692 35888
rect 71732 35848 71741 35888
rect 71683 35847 71741 35848
rect 71883 35888 71925 35897
rect 71883 35848 71884 35888
rect 71924 35848 71925 35888
rect 71883 35839 71925 35848
rect 72075 35888 72117 35897
rect 72075 35848 72076 35888
rect 72116 35848 72117 35888
rect 72075 35839 72117 35848
rect 72163 35888 72221 35889
rect 72163 35848 72172 35888
rect 72212 35848 72221 35888
rect 72163 35847 72221 35848
rect 72835 35888 72893 35889
rect 72835 35848 72844 35888
rect 72884 35848 72893 35888
rect 72835 35847 72893 35848
rect 73131 35888 73173 35897
rect 73131 35848 73132 35888
rect 73172 35848 73173 35888
rect 73131 35839 73173 35848
rect 73227 35888 73269 35897
rect 73227 35848 73228 35888
rect 73268 35848 73269 35888
rect 73227 35839 73269 35848
rect 73699 35888 73757 35889
rect 73699 35848 73708 35888
rect 73748 35848 73757 35888
rect 73699 35847 73757 35848
rect 73899 35888 73941 35897
rect 73899 35848 73900 35888
rect 73940 35848 73941 35888
rect 73899 35839 73941 35848
rect 76203 35888 76245 35897
rect 76203 35848 76204 35888
rect 76244 35848 76245 35888
rect 76203 35839 76245 35848
rect 76395 35888 76437 35897
rect 76395 35848 76396 35888
rect 76436 35848 76437 35888
rect 76395 35839 76437 35848
rect 76483 35888 76541 35889
rect 76483 35848 76492 35888
rect 76532 35848 76541 35888
rect 76483 35847 76541 35848
rect 77059 35888 77117 35889
rect 77059 35848 77068 35888
rect 77108 35848 77117 35888
rect 77059 35847 77117 35848
rect 77259 35888 77301 35897
rect 77259 35848 77260 35888
rect 77300 35848 77301 35888
rect 77259 35839 77301 35848
rect 77443 35888 77501 35889
rect 77443 35848 77452 35888
rect 77492 35848 77501 35888
rect 77443 35847 77501 35848
rect 77643 35888 77685 35897
rect 77643 35848 77644 35888
rect 77684 35848 77685 35888
rect 77643 35839 77685 35848
rect 51435 35804 51477 35813
rect 51435 35764 51436 35804
rect 51476 35764 51477 35804
rect 51435 35755 51477 35764
rect 52011 35804 52053 35813
rect 52011 35764 52012 35804
rect 52052 35764 52053 35804
rect 52011 35755 52053 35764
rect 59019 35804 59061 35813
rect 59019 35764 59020 35804
rect 59060 35764 59061 35804
rect 59019 35755 59061 35764
rect 59499 35804 59541 35813
rect 59499 35764 59500 35804
rect 59540 35764 59541 35804
rect 59499 35755 59541 35764
rect 69771 35804 69813 35813
rect 69771 35764 69772 35804
rect 69812 35764 69813 35804
rect 69771 35755 69813 35764
rect 71595 35804 71637 35813
rect 71595 35764 71596 35804
rect 71636 35764 71637 35804
rect 71595 35755 71637 35764
rect 76299 35804 76341 35813
rect 76299 35764 76300 35804
rect 76340 35764 76341 35804
rect 76299 35755 76341 35764
rect 77163 35804 77205 35813
rect 77163 35764 77164 35804
rect 77204 35764 77205 35804
rect 77163 35755 77205 35764
rect 50763 35720 50805 35729
rect 50763 35680 50764 35720
rect 50804 35680 50805 35720
rect 50763 35671 50805 35680
rect 54403 35720 54461 35721
rect 54403 35680 54412 35720
rect 54452 35680 54461 35720
rect 54403 35679 54461 35680
rect 55747 35720 55805 35721
rect 55747 35680 55756 35720
rect 55796 35680 55805 35720
rect 55747 35679 55805 35680
rect 56907 35720 56949 35729
rect 56907 35680 56908 35720
rect 56948 35680 56949 35720
rect 56907 35671 56949 35680
rect 66787 35720 66845 35721
rect 66787 35680 66796 35720
rect 66836 35680 66845 35720
rect 66787 35679 66845 35680
rect 71971 35720 72029 35721
rect 71971 35680 71980 35720
rect 72020 35680 72029 35720
rect 71971 35679 72029 35680
rect 576 35552 79584 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79584 35552
rect 576 35488 79584 35512
rect 52195 35384 52253 35385
rect 52195 35344 52204 35384
rect 52244 35344 52253 35384
rect 52195 35343 52253 35344
rect 76579 35384 76637 35385
rect 76579 35344 76588 35384
rect 76628 35344 76637 35384
rect 76579 35343 76637 35344
rect 52683 35300 52725 35309
rect 52683 35260 52684 35300
rect 52724 35260 52725 35300
rect 52683 35251 52725 35260
rect 54891 35300 54933 35309
rect 54891 35260 54892 35300
rect 54932 35260 54933 35300
rect 54891 35251 54933 35260
rect 55179 35300 55221 35309
rect 55179 35260 55180 35300
rect 55220 35260 55221 35300
rect 55179 35251 55221 35260
rect 66027 35300 66069 35309
rect 66027 35260 66028 35300
rect 66068 35260 66069 35300
rect 66027 35251 66069 35260
rect 71307 35300 71349 35309
rect 71307 35260 71308 35300
rect 71348 35260 71349 35300
rect 71307 35251 71349 35260
rect 73419 35300 73461 35309
rect 73419 35260 73420 35300
rect 73460 35260 73461 35300
rect 73419 35251 73461 35260
rect 49699 35216 49757 35217
rect 49699 35176 49708 35216
rect 49748 35176 49757 35216
rect 49699 35175 49757 35176
rect 50563 35216 50621 35217
rect 50563 35176 50572 35216
rect 50612 35176 50621 35216
rect 50563 35175 50621 35176
rect 50955 35216 50997 35225
rect 50955 35176 50956 35216
rect 50996 35176 50997 35216
rect 50955 35167 50997 35176
rect 51435 35216 51477 35225
rect 51435 35176 51436 35216
rect 51476 35176 51477 35216
rect 51435 35167 51477 35176
rect 51531 35216 51573 35225
rect 51531 35176 51532 35216
rect 51572 35176 51573 35216
rect 51531 35167 51573 35176
rect 51811 35216 51869 35217
rect 51811 35176 51820 35216
rect 51860 35176 51869 35216
rect 51811 35175 51869 35176
rect 52107 35216 52149 35225
rect 52107 35176 52108 35216
rect 52148 35176 52149 35216
rect 52107 35167 52149 35176
rect 52299 35216 52341 35225
rect 52299 35176 52300 35216
rect 52340 35176 52341 35216
rect 52299 35167 52341 35176
rect 52387 35216 52445 35217
rect 52387 35176 52396 35216
rect 52436 35176 52445 35216
rect 52387 35175 52445 35176
rect 52579 35216 52637 35217
rect 52579 35176 52588 35216
rect 52628 35176 52637 35216
rect 52579 35175 52637 35176
rect 52779 35216 52821 35225
rect 52779 35176 52780 35216
rect 52820 35176 52821 35216
rect 52779 35167 52821 35176
rect 54787 35216 54845 35217
rect 54787 35176 54796 35216
rect 54836 35176 54845 35216
rect 54787 35175 54845 35176
rect 54987 35216 55029 35225
rect 54987 35176 54988 35216
rect 55028 35176 55029 35216
rect 54987 35167 55029 35176
rect 55555 35216 55613 35217
rect 55555 35176 55564 35216
rect 55604 35176 55613 35216
rect 55555 35175 55613 35176
rect 56419 35216 56477 35217
rect 56419 35176 56428 35216
rect 56468 35176 56477 35216
rect 56419 35175 56477 35176
rect 57771 35216 57813 35225
rect 57771 35176 57772 35216
rect 57812 35176 57813 35216
rect 57771 35167 57813 35176
rect 57963 35216 58005 35225
rect 57963 35176 57964 35216
rect 58004 35176 58005 35216
rect 57963 35167 58005 35176
rect 58051 35216 58109 35217
rect 58051 35176 58060 35216
rect 58100 35176 58109 35216
rect 58051 35175 58109 35176
rect 59883 35216 59925 35225
rect 59883 35176 59884 35216
rect 59924 35176 59925 35216
rect 59883 35167 59925 35176
rect 60259 35216 60317 35217
rect 60259 35176 60268 35216
rect 60308 35176 60317 35216
rect 60259 35175 60317 35176
rect 61123 35216 61181 35217
rect 61123 35176 61132 35216
rect 61172 35176 61181 35216
rect 61123 35175 61181 35176
rect 62763 35216 62805 35225
rect 62763 35176 62764 35216
rect 62804 35176 62805 35216
rect 62763 35167 62805 35176
rect 62859 35216 62901 35225
rect 62859 35176 62860 35216
rect 62900 35176 62901 35216
rect 62859 35167 62901 35176
rect 63139 35216 63197 35217
rect 63139 35176 63148 35216
rect 63188 35176 63197 35216
rect 63139 35175 63197 35176
rect 65923 35216 65981 35217
rect 65923 35176 65932 35216
rect 65972 35176 65981 35216
rect 65923 35175 65981 35176
rect 66123 35216 66165 35225
rect 66123 35176 66124 35216
rect 66164 35176 66165 35216
rect 66123 35167 66165 35176
rect 66603 35216 66645 35225
rect 66603 35176 66604 35216
rect 66644 35176 66645 35216
rect 66603 35167 66645 35176
rect 66699 35216 66741 35225
rect 66699 35176 66700 35216
rect 66740 35176 66741 35216
rect 66699 35167 66741 35176
rect 66979 35216 67037 35217
rect 66979 35176 66988 35216
rect 67028 35176 67037 35216
rect 66979 35175 67037 35176
rect 67275 35216 67317 35225
rect 67275 35176 67276 35216
rect 67316 35176 67317 35216
rect 67275 35167 67317 35176
rect 67651 35216 67709 35217
rect 67651 35176 67660 35216
rect 67700 35176 67709 35216
rect 67651 35175 67709 35176
rect 68515 35216 68573 35217
rect 68515 35176 68524 35216
rect 68564 35176 68573 35216
rect 68515 35175 68573 35176
rect 70347 35216 70389 35225
rect 70347 35176 70348 35216
rect 70388 35176 70389 35216
rect 70347 35167 70389 35176
rect 70443 35216 70485 35225
rect 70443 35176 70444 35216
rect 70484 35176 70485 35216
rect 70443 35167 70485 35176
rect 70539 35216 70581 35225
rect 70539 35176 70540 35216
rect 70580 35176 70581 35216
rect 70539 35167 70581 35176
rect 70635 35216 70677 35225
rect 70635 35176 70636 35216
rect 70676 35176 70677 35216
rect 70635 35167 70677 35176
rect 70915 35216 70973 35217
rect 70915 35176 70924 35216
rect 70964 35176 70973 35216
rect 70915 35175 70973 35176
rect 71211 35216 71253 35225
rect 71211 35176 71212 35216
rect 71252 35176 71253 35216
rect 71211 35167 71253 35176
rect 71787 35216 71829 35225
rect 71787 35176 71788 35216
rect 71828 35176 71829 35216
rect 71787 35167 71829 35176
rect 71979 35216 72021 35225
rect 71979 35176 71980 35216
rect 72020 35176 72021 35216
rect 71979 35167 72021 35176
rect 72067 35216 72125 35217
rect 72067 35176 72076 35216
rect 72116 35176 72125 35216
rect 72067 35175 72125 35176
rect 73315 35216 73373 35217
rect 73315 35176 73324 35216
rect 73364 35176 73373 35216
rect 73315 35175 73373 35176
rect 73515 35216 73557 35225
rect 73515 35176 73516 35216
rect 73556 35176 73557 35216
rect 73515 35167 73557 35176
rect 74187 35216 74229 35225
rect 74187 35176 74188 35216
rect 74228 35176 74229 35216
rect 74187 35167 74229 35176
rect 74563 35216 74621 35217
rect 74563 35176 74572 35216
rect 74612 35176 74621 35216
rect 74563 35175 74621 35176
rect 75427 35216 75485 35217
rect 75427 35176 75436 35216
rect 75476 35176 75485 35216
rect 75427 35175 75485 35176
rect 77067 35216 77109 35225
rect 77067 35176 77068 35216
rect 77108 35176 77109 35216
rect 77067 35167 77109 35176
rect 77443 35216 77501 35217
rect 77443 35176 77452 35216
rect 77492 35176 77501 35216
rect 77443 35175 77501 35176
rect 78307 35216 78365 35217
rect 78307 35176 78316 35216
rect 78356 35176 78365 35216
rect 78307 35175 78365 35176
rect 47115 35048 47157 35057
rect 47115 35008 47116 35048
rect 47156 35008 47157 35048
rect 47115 34999 47157 35008
rect 51139 35048 51197 35049
rect 51139 35008 51148 35048
rect 51188 35008 51197 35048
rect 51139 35007 51197 35008
rect 58443 35048 58485 35057
rect 58443 35008 58444 35048
rect 58484 35008 58485 35048
rect 58443 34999 58485 35008
rect 63627 35048 63669 35057
rect 63627 35008 63628 35048
rect 63668 35008 63669 35048
rect 63627 34999 63669 35008
rect 64875 35048 64917 35057
rect 64875 35008 64876 35048
rect 64916 35008 64917 35048
rect 64875 34999 64917 35008
rect 66307 35048 66365 35049
rect 66307 35008 66316 35048
rect 66356 35008 66365 35048
rect 66307 35007 66365 35008
rect 71587 35048 71645 35049
rect 71587 35008 71596 35048
rect 71636 35008 71645 35048
rect 71587 35007 71645 35008
rect 72555 35048 72597 35057
rect 72555 35008 72556 35048
rect 72596 35008 72597 35048
rect 72555 34999 72597 35008
rect 48547 34964 48605 34965
rect 48547 34924 48556 34964
rect 48596 34924 48605 34964
rect 48547 34923 48605 34924
rect 57571 34964 57629 34965
rect 57571 34924 57580 34964
rect 57620 34924 57629 34964
rect 57571 34923 57629 34924
rect 57771 34964 57813 34973
rect 57771 34924 57772 34964
rect 57812 34924 57813 34964
rect 57771 34915 57813 34924
rect 62275 34964 62333 34965
rect 62275 34924 62284 34964
rect 62324 34924 62333 34964
rect 62275 34923 62333 34924
rect 62467 34964 62525 34965
rect 62467 34924 62476 34964
rect 62516 34924 62525 34964
rect 62467 34923 62525 34924
rect 69667 34964 69725 34965
rect 69667 34924 69676 34964
rect 69716 34924 69725 34964
rect 69667 34923 69725 34924
rect 71787 34964 71829 34973
rect 71787 34924 71788 34964
rect 71828 34924 71829 34964
rect 71787 34915 71829 34924
rect 76579 34964 76637 34965
rect 76579 34924 76588 34964
rect 76628 34924 76637 34964
rect 76579 34923 76637 34924
rect 79459 34964 79517 34965
rect 79459 34924 79468 34964
rect 79508 34924 79517 34964
rect 79459 34923 79517 34924
rect 576 34796 79584 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79584 34796
rect 576 34732 79584 34756
rect 50955 34628 50997 34637
rect 50955 34588 50956 34628
rect 50996 34588 50997 34628
rect 50955 34579 50997 34588
rect 56515 34628 56573 34629
rect 56515 34588 56524 34628
rect 56564 34588 56573 34628
rect 56515 34587 56573 34588
rect 66891 34628 66933 34637
rect 66891 34588 66892 34628
rect 66932 34588 66933 34628
rect 66891 34579 66933 34588
rect 68803 34628 68861 34629
rect 68803 34588 68812 34628
rect 68852 34588 68861 34628
rect 68803 34587 68861 34588
rect 77251 34628 77309 34629
rect 77251 34588 77260 34628
rect 77300 34588 77309 34628
rect 77251 34587 77309 34588
rect 46443 34544 46485 34553
rect 46443 34504 46444 34544
rect 46484 34504 46485 34544
rect 46443 34495 46485 34504
rect 49227 34544 49269 34553
rect 49227 34504 49228 34544
rect 49268 34504 49269 34544
rect 49227 34495 49269 34504
rect 52011 34544 52053 34553
rect 52011 34504 52012 34544
rect 52052 34504 52053 34544
rect 52011 34495 52053 34504
rect 52203 34544 52245 34553
rect 52203 34504 52204 34544
rect 52244 34504 52245 34544
rect 52203 34495 52245 34504
rect 55563 34544 55605 34553
rect 55563 34504 55564 34544
rect 55604 34504 55605 34544
rect 55563 34495 55605 34504
rect 57771 34544 57813 34553
rect 57771 34504 57772 34544
rect 57812 34504 57813 34544
rect 57771 34495 57813 34504
rect 61995 34544 62037 34553
rect 61995 34504 61996 34544
rect 62036 34504 62037 34544
rect 61995 34495 62037 34504
rect 67467 34544 67509 34553
rect 67467 34504 67468 34544
rect 67508 34504 67509 34544
rect 67467 34495 67509 34504
rect 67755 34544 67797 34553
rect 67755 34504 67756 34544
rect 67796 34504 67797 34544
rect 67755 34495 67797 34504
rect 71883 34544 71925 34553
rect 71883 34504 71884 34544
rect 71924 34504 71925 34544
rect 71883 34495 71925 34504
rect 74667 34544 74709 34553
rect 74667 34504 74668 34544
rect 74708 34504 74709 34544
rect 74667 34495 74709 34504
rect 76011 34544 76053 34553
rect 76011 34504 76012 34544
rect 76052 34504 76053 34544
rect 76011 34495 76053 34504
rect 77451 34544 77493 34553
rect 77451 34504 77452 34544
rect 77492 34504 77493 34544
rect 77451 34495 77493 34504
rect 46147 34376 46205 34377
rect 46147 34336 46156 34376
rect 46196 34336 46205 34376
rect 46147 34335 46205 34336
rect 46251 34376 46293 34385
rect 46251 34336 46252 34376
rect 46292 34336 46293 34376
rect 46251 34327 46293 34336
rect 46443 34376 46485 34385
rect 46443 34336 46444 34376
rect 46484 34336 46485 34376
rect 46443 34327 46485 34336
rect 46635 34376 46677 34385
rect 46635 34336 46636 34376
rect 46676 34336 46677 34376
rect 46635 34327 46677 34336
rect 47011 34376 47069 34377
rect 47011 34336 47020 34376
rect 47060 34336 47069 34376
rect 47011 34335 47069 34336
rect 47875 34376 47933 34377
rect 47875 34336 47884 34376
rect 47924 34336 47933 34376
rect 47875 34335 47933 34336
rect 49227 34376 49269 34385
rect 49227 34336 49228 34376
rect 49268 34336 49269 34376
rect 49227 34327 49269 34336
rect 49419 34376 49461 34385
rect 49419 34336 49420 34376
rect 49460 34336 49461 34376
rect 49419 34327 49461 34336
rect 49507 34376 49565 34377
rect 49507 34336 49516 34376
rect 49556 34336 49565 34376
rect 49507 34335 49565 34336
rect 50475 34376 50517 34385
rect 50475 34336 50476 34376
rect 50516 34336 50517 34376
rect 50475 34327 50517 34336
rect 50571 34376 50613 34385
rect 50571 34336 50572 34376
rect 50612 34336 50613 34376
rect 50571 34327 50613 34336
rect 50667 34376 50709 34385
rect 50667 34336 50668 34376
rect 50708 34336 50709 34376
rect 50667 34327 50709 34336
rect 50763 34376 50805 34385
rect 50763 34336 50764 34376
rect 50804 34336 50805 34376
rect 50763 34327 50805 34336
rect 50955 34376 50997 34385
rect 50955 34336 50956 34376
rect 50996 34336 50997 34376
rect 50955 34327 50997 34336
rect 51147 34376 51189 34385
rect 51147 34336 51148 34376
rect 51188 34336 51189 34376
rect 51147 34327 51189 34336
rect 51235 34376 51293 34377
rect 51235 34336 51244 34376
rect 51284 34336 51293 34376
rect 51235 34335 51293 34336
rect 52203 34376 52245 34385
rect 52203 34336 52204 34376
rect 52244 34336 52245 34376
rect 52203 34327 52245 34336
rect 52395 34376 52437 34385
rect 52395 34336 52396 34376
rect 52436 34336 52437 34376
rect 52395 34327 52437 34336
rect 52483 34376 52541 34377
rect 52483 34336 52492 34376
rect 52532 34336 52541 34376
rect 52483 34335 52541 34336
rect 53835 34376 53877 34385
rect 53835 34336 53836 34376
rect 53876 34336 53877 34376
rect 53835 34327 53877 34336
rect 54027 34376 54069 34385
rect 54027 34336 54028 34376
rect 54068 34336 54069 34376
rect 54027 34327 54069 34336
rect 54115 34376 54173 34377
rect 54115 34336 54124 34376
rect 54164 34336 54173 34376
rect 54115 34335 54173 34336
rect 55843 34376 55901 34377
rect 55843 34336 55852 34376
rect 55892 34336 55901 34376
rect 55843 34335 55901 34336
rect 56139 34376 56181 34385
rect 56139 34336 56140 34376
rect 56180 34336 56181 34376
rect 56139 34327 56181 34336
rect 57475 34376 57533 34377
rect 57475 34336 57484 34376
rect 57524 34336 57533 34376
rect 57475 34335 57533 34336
rect 57579 34376 57621 34385
rect 57579 34336 57580 34376
rect 57620 34336 57621 34376
rect 57579 34327 57621 34336
rect 57771 34376 57813 34385
rect 57771 34336 57772 34376
rect 57812 34336 57813 34376
rect 57771 34327 57813 34336
rect 57963 34376 58005 34385
rect 57963 34336 57964 34376
rect 58004 34336 58005 34376
rect 57963 34327 58005 34336
rect 58339 34376 58397 34377
rect 58339 34336 58348 34376
rect 58388 34336 58397 34376
rect 58339 34335 58397 34336
rect 59203 34376 59261 34377
rect 59203 34336 59212 34376
rect 59252 34336 59261 34376
rect 59203 34335 59261 34336
rect 61515 34376 61557 34385
rect 61515 34336 61516 34376
rect 61556 34336 61557 34376
rect 61515 34327 61557 34336
rect 61611 34376 61653 34385
rect 61611 34336 61612 34376
rect 61652 34336 61653 34376
rect 61611 34327 61653 34336
rect 61707 34376 61749 34385
rect 61707 34336 61708 34376
rect 61748 34336 61749 34376
rect 61707 34327 61749 34336
rect 61803 34376 61845 34385
rect 61803 34336 61804 34376
rect 61844 34336 61845 34376
rect 61803 34327 61845 34336
rect 61995 34376 62037 34385
rect 61995 34336 61996 34376
rect 62036 34336 62037 34376
rect 61995 34327 62037 34336
rect 62187 34376 62229 34385
rect 62187 34336 62188 34376
rect 62228 34336 62229 34376
rect 62187 34327 62229 34336
rect 62275 34376 62333 34377
rect 62275 34336 62284 34376
rect 62324 34336 62333 34376
rect 62275 34335 62333 34336
rect 62667 34376 62709 34385
rect 62667 34336 62668 34376
rect 62708 34336 62709 34376
rect 62667 34327 62709 34336
rect 62859 34376 62901 34385
rect 62859 34336 62860 34376
rect 62900 34336 62901 34376
rect 62859 34327 62901 34336
rect 62947 34376 63005 34377
rect 62947 34336 62956 34376
rect 62996 34336 63005 34376
rect 62947 34335 63005 34336
rect 63523 34376 63581 34377
rect 63523 34336 63532 34376
rect 63572 34336 63581 34376
rect 63523 34335 63581 34336
rect 64387 34376 64445 34377
rect 64387 34336 64396 34376
rect 64436 34336 64445 34376
rect 64387 34335 64445 34336
rect 66123 34376 66165 34385
rect 66123 34336 66124 34376
rect 66164 34336 66165 34376
rect 66123 34327 66165 34336
rect 66315 34376 66357 34385
rect 66315 34336 66316 34376
rect 66356 34336 66357 34376
rect 66315 34327 66357 34336
rect 66403 34376 66461 34377
rect 66403 34336 66412 34376
rect 66452 34336 66461 34376
rect 66403 34335 66461 34336
rect 66891 34376 66933 34385
rect 66891 34336 66892 34376
rect 66932 34336 66933 34376
rect 66891 34327 66933 34336
rect 67083 34376 67125 34385
rect 67083 34336 67084 34376
rect 67124 34336 67125 34376
rect 67083 34327 67125 34336
rect 67171 34376 67229 34377
rect 67171 34336 67180 34376
rect 67220 34336 67229 34376
rect 67171 34335 67229 34336
rect 67363 34376 67421 34377
rect 67363 34336 67372 34376
rect 67412 34336 67421 34376
rect 67363 34335 67421 34336
rect 67563 34376 67605 34385
rect 67563 34336 67564 34376
rect 67604 34336 67605 34376
rect 67563 34327 67605 34336
rect 69955 34376 70013 34377
rect 69955 34336 69964 34376
rect 70004 34336 70013 34376
rect 69955 34335 70013 34336
rect 70819 34376 70877 34377
rect 70819 34336 70828 34376
rect 70868 34336 70877 34376
rect 70819 34335 70877 34336
rect 71211 34376 71253 34385
rect 71211 34336 71212 34376
rect 71252 34336 71253 34376
rect 71211 34327 71253 34336
rect 71587 34376 71645 34377
rect 71587 34336 71596 34376
rect 71636 34336 71645 34376
rect 71587 34335 71645 34336
rect 71691 34376 71733 34385
rect 71691 34336 71692 34376
rect 71732 34336 71733 34376
rect 71691 34327 71733 34336
rect 71883 34376 71925 34385
rect 71883 34336 71884 34376
rect 71924 34336 71925 34376
rect 71883 34327 71925 34336
rect 72075 34376 72117 34385
rect 72075 34336 72076 34376
rect 72116 34336 72117 34376
rect 72075 34327 72117 34336
rect 72451 34376 72509 34377
rect 72451 34336 72460 34376
rect 72500 34336 72509 34376
rect 72451 34335 72509 34336
rect 73315 34376 73373 34377
rect 73315 34336 73324 34376
rect 73364 34336 73373 34376
rect 73315 34335 73373 34336
rect 75627 34376 75669 34385
rect 75627 34336 75628 34376
rect 75668 34336 75669 34376
rect 75627 34327 75669 34336
rect 75723 34376 75765 34385
rect 75723 34336 75724 34376
rect 75764 34336 75765 34376
rect 75723 34327 75765 34336
rect 75819 34376 75861 34385
rect 75819 34336 75820 34376
rect 75860 34336 75861 34376
rect 75819 34327 75861 34336
rect 76011 34376 76053 34385
rect 76011 34336 76012 34376
rect 76052 34336 76053 34376
rect 76011 34327 76053 34336
rect 76203 34376 76245 34385
rect 76203 34336 76204 34376
rect 76244 34336 76245 34376
rect 76203 34327 76245 34336
rect 76291 34376 76349 34377
rect 76291 34336 76300 34376
rect 76340 34336 76349 34376
rect 76291 34335 76349 34336
rect 76579 34376 76637 34377
rect 76579 34336 76588 34376
rect 76628 34336 76637 34376
rect 76579 34335 76637 34336
rect 76875 34376 76917 34385
rect 76875 34336 76876 34376
rect 76916 34336 76917 34376
rect 76875 34327 76917 34336
rect 76971 34376 77013 34385
rect 76971 34336 76972 34376
rect 77012 34336 77013 34376
rect 76971 34327 77013 34336
rect 77451 34376 77493 34385
rect 77451 34336 77452 34376
rect 77492 34336 77493 34376
rect 77451 34327 77493 34336
rect 77643 34376 77685 34385
rect 77643 34336 77644 34376
rect 77684 34336 77685 34376
rect 77643 34327 77685 34336
rect 77731 34376 77789 34377
rect 77731 34336 77740 34376
rect 77780 34336 77789 34376
rect 77731 34335 77789 34336
rect 77923 34376 77981 34377
rect 77923 34336 77932 34376
rect 77972 34336 77981 34376
rect 77923 34335 77981 34336
rect 78123 34376 78165 34385
rect 78123 34336 78124 34376
rect 78164 34336 78165 34376
rect 78123 34327 78165 34336
rect 56235 34292 56277 34301
rect 56235 34252 56236 34292
rect 56276 34252 56277 34292
rect 56235 34243 56277 34252
rect 62763 34292 62805 34301
rect 62763 34252 62764 34292
rect 62804 34252 62805 34292
rect 62763 34243 62805 34252
rect 63147 34292 63189 34301
rect 63147 34252 63148 34292
rect 63188 34252 63189 34292
rect 63147 34243 63189 34252
rect 78027 34292 78069 34301
rect 78027 34252 78028 34292
rect 78068 34252 78069 34292
rect 78027 34243 78069 34252
rect 49027 34208 49085 34209
rect 49027 34168 49036 34208
rect 49076 34168 49085 34208
rect 49027 34167 49085 34168
rect 53923 34208 53981 34209
rect 53923 34168 53932 34208
rect 53972 34168 53981 34208
rect 53923 34167 53981 34168
rect 60355 34208 60413 34209
rect 60355 34168 60364 34208
rect 60404 34168 60413 34208
rect 60355 34167 60413 34168
rect 65539 34208 65597 34209
rect 65539 34168 65548 34208
rect 65588 34168 65597 34208
rect 65539 34167 65597 34168
rect 66211 34208 66269 34209
rect 66211 34168 66220 34208
rect 66260 34168 66269 34208
rect 66211 34167 66269 34168
rect 74467 34208 74525 34209
rect 74467 34168 74476 34208
rect 74516 34168 74525 34208
rect 74467 34167 74525 34168
rect 75523 34208 75581 34209
rect 75523 34168 75532 34208
rect 75572 34168 75581 34208
rect 75523 34167 75581 34168
rect 576 34040 79584 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79584 34040
rect 576 33976 79584 34000
rect 46723 33872 46781 33873
rect 46723 33832 46732 33872
rect 46772 33832 46781 33872
rect 46723 33831 46781 33832
rect 58339 33872 58397 33873
rect 58339 33832 58348 33872
rect 58388 33832 58397 33872
rect 58339 33831 58397 33832
rect 62275 33872 62333 33873
rect 62275 33832 62284 33872
rect 62324 33832 62333 33872
rect 62275 33831 62333 33832
rect 51627 33788 51669 33797
rect 51627 33748 51628 33788
rect 51668 33748 51669 33788
rect 51627 33739 51669 33748
rect 62763 33788 62805 33797
rect 62763 33748 62764 33788
rect 62804 33748 62805 33788
rect 62763 33739 62805 33748
rect 63147 33788 63189 33797
rect 63147 33748 63148 33788
rect 63188 33748 63189 33788
rect 63147 33739 63189 33748
rect 66219 33788 66261 33797
rect 66219 33748 66220 33788
rect 66260 33748 66261 33788
rect 66219 33739 66261 33748
rect 71691 33788 71733 33797
rect 71691 33748 71692 33788
rect 71732 33748 71733 33788
rect 71691 33739 71733 33748
rect 46827 33704 46869 33713
rect 46827 33664 46828 33704
rect 46868 33664 46869 33704
rect 46827 33655 46869 33664
rect 46923 33704 46965 33713
rect 46923 33664 46924 33704
rect 46964 33664 46965 33704
rect 46923 33655 46965 33664
rect 47019 33704 47061 33713
rect 47019 33664 47020 33704
rect 47060 33664 47061 33704
rect 47019 33655 47061 33664
rect 49227 33704 49269 33713
rect 49227 33664 49228 33704
rect 49268 33664 49269 33704
rect 49227 33655 49269 33664
rect 49419 33704 49461 33713
rect 49419 33664 49420 33704
rect 49460 33664 49461 33704
rect 49419 33655 49461 33664
rect 49507 33704 49565 33705
rect 49507 33664 49516 33704
rect 49556 33664 49565 33704
rect 49507 33663 49565 33664
rect 52003 33704 52061 33705
rect 52003 33664 52012 33704
rect 52052 33664 52061 33704
rect 52003 33663 52061 33664
rect 52867 33704 52925 33705
rect 52867 33664 52876 33704
rect 52916 33664 52925 33704
rect 52867 33663 52925 33664
rect 54307 33704 54365 33705
rect 54307 33664 54316 33704
rect 54356 33664 54365 33704
rect 54307 33663 54365 33664
rect 54603 33704 54645 33713
rect 54603 33664 54604 33704
rect 54644 33664 54645 33704
rect 54603 33655 54645 33664
rect 54699 33704 54741 33713
rect 54699 33664 54700 33704
rect 54740 33664 54741 33704
rect 54699 33655 54741 33664
rect 55171 33704 55229 33705
rect 55171 33664 55180 33704
rect 55220 33664 55229 33704
rect 55171 33663 55229 33664
rect 55275 33704 55317 33713
rect 55275 33664 55276 33704
rect 55316 33664 55317 33704
rect 55275 33655 55317 33664
rect 55371 33704 55413 33713
rect 55371 33664 55372 33704
rect 55412 33664 55413 33704
rect 55371 33655 55413 33664
rect 58443 33704 58485 33713
rect 58443 33664 58444 33704
rect 58484 33664 58485 33704
rect 58443 33655 58485 33664
rect 58539 33704 58581 33713
rect 58539 33664 58540 33704
rect 58580 33664 58581 33704
rect 58539 33655 58581 33664
rect 58635 33704 58677 33713
rect 58635 33664 58636 33704
rect 58676 33664 58677 33704
rect 58635 33655 58677 33664
rect 58819 33704 58877 33705
rect 58819 33664 58828 33704
rect 58868 33664 58877 33704
rect 58819 33663 58877 33664
rect 59019 33704 59061 33713
rect 59019 33664 59020 33704
rect 59060 33664 59061 33704
rect 59019 33655 59061 33664
rect 62187 33704 62229 33713
rect 62187 33664 62188 33704
rect 62228 33664 62229 33704
rect 62187 33655 62229 33664
rect 62379 33704 62421 33713
rect 62379 33664 62380 33704
rect 62420 33664 62421 33704
rect 62379 33655 62421 33664
rect 62467 33704 62525 33705
rect 62467 33664 62476 33704
rect 62516 33664 62525 33704
rect 62467 33663 62525 33664
rect 62667 33704 62709 33713
rect 62667 33664 62668 33704
rect 62708 33664 62709 33704
rect 62667 33655 62709 33664
rect 62851 33704 62909 33705
rect 62851 33664 62860 33704
rect 62900 33664 62909 33704
rect 62851 33663 62909 33664
rect 63043 33704 63101 33705
rect 63043 33664 63052 33704
rect 63092 33664 63101 33704
rect 63043 33663 63101 33664
rect 63243 33704 63285 33713
rect 63243 33664 63244 33704
rect 63284 33664 63285 33704
rect 63243 33655 63285 33664
rect 66123 33704 66165 33713
rect 66123 33664 66124 33704
rect 66164 33664 66165 33704
rect 66123 33655 66165 33664
rect 66315 33704 66357 33713
rect 66315 33664 66316 33704
rect 66356 33664 66357 33704
rect 66315 33655 66357 33664
rect 66403 33704 66461 33705
rect 66403 33664 66412 33704
rect 66452 33664 66461 33704
rect 66403 33663 66461 33664
rect 66595 33704 66653 33705
rect 66595 33664 66604 33704
rect 66644 33664 66653 33704
rect 66595 33663 66653 33664
rect 66795 33704 66837 33713
rect 66795 33664 66796 33704
rect 66836 33664 66837 33704
rect 66795 33655 66837 33664
rect 71587 33704 71645 33705
rect 71587 33664 71596 33704
rect 71636 33664 71645 33704
rect 71587 33663 71645 33664
rect 71787 33704 71829 33713
rect 71787 33664 71788 33704
rect 71828 33664 71829 33704
rect 71787 33655 71829 33664
rect 71979 33704 72021 33713
rect 71979 33664 71980 33704
rect 72020 33664 72021 33704
rect 71979 33655 72021 33664
rect 72171 33704 72213 33713
rect 72171 33664 72172 33704
rect 72212 33664 72213 33704
rect 72171 33655 72213 33664
rect 72259 33704 72317 33705
rect 72259 33664 72268 33704
rect 72308 33664 72317 33704
rect 72259 33663 72317 33664
rect 72459 33704 72501 33713
rect 72459 33664 72460 33704
rect 72500 33664 72501 33704
rect 72459 33655 72501 33664
rect 72555 33704 72597 33713
rect 72555 33664 72556 33704
rect 72596 33664 72597 33704
rect 72555 33655 72597 33664
rect 72643 33704 72701 33705
rect 72643 33664 72652 33704
rect 72692 33664 72701 33704
rect 72643 33663 72701 33664
rect 75715 33704 75773 33705
rect 75715 33664 75724 33704
rect 75764 33664 75773 33704
rect 75715 33663 75773 33664
rect 75819 33704 75861 33713
rect 75819 33664 75820 33704
rect 75860 33664 75861 33704
rect 75819 33655 75861 33664
rect 76011 33704 76053 33713
rect 76011 33664 76012 33704
rect 76052 33664 76053 33704
rect 76011 33655 76053 33664
rect 76203 33704 76245 33713
rect 76203 33664 76204 33704
rect 76244 33664 76245 33704
rect 76203 33655 76245 33664
rect 76299 33704 76341 33713
rect 76299 33664 76300 33704
rect 76340 33664 76341 33704
rect 76299 33655 76341 33664
rect 76395 33704 76437 33713
rect 76395 33664 76396 33704
rect 76436 33664 76437 33704
rect 76395 33655 76437 33664
rect 76491 33704 76533 33713
rect 76491 33664 76492 33704
rect 76532 33664 76533 33704
rect 76491 33655 76533 33664
rect 76683 33704 76725 33713
rect 76683 33664 76684 33704
rect 76724 33664 76725 33704
rect 76683 33655 76725 33664
rect 76875 33704 76917 33713
rect 76875 33664 76876 33704
rect 76916 33664 76917 33704
rect 76875 33655 76917 33664
rect 76963 33704 77021 33705
rect 76963 33664 76972 33704
rect 77012 33664 77021 33704
rect 76963 33663 77021 33664
rect 77259 33704 77301 33713
rect 77259 33664 77260 33704
rect 77300 33664 77301 33704
rect 77259 33655 77301 33664
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77451 33655 77493 33664
rect 77539 33704 77597 33705
rect 77539 33664 77548 33704
rect 77588 33664 77597 33704
rect 77539 33663 77597 33664
rect 54027 33620 54069 33629
rect 54027 33580 54028 33620
rect 54068 33580 54069 33620
rect 54027 33571 54069 33580
rect 48843 33536 48885 33545
rect 48843 33496 48844 33536
rect 48884 33496 48885 33536
rect 48843 33487 48885 33496
rect 54979 33536 55037 33537
rect 54979 33496 54988 33536
rect 55028 33496 55037 33536
rect 54979 33495 55037 33496
rect 55851 33536 55893 33545
rect 55851 33496 55852 33536
rect 55892 33496 55893 33536
rect 55851 33487 55893 33496
rect 59211 33536 59253 33545
rect 59211 33496 59212 33536
rect 59252 33496 59253 33536
rect 59211 33487 59253 33496
rect 63723 33536 63765 33545
rect 63723 33496 63724 33536
rect 63764 33496 63765 33536
rect 63723 33487 63765 33496
rect 66987 33536 67029 33545
rect 66987 33496 66988 33536
rect 67028 33496 67029 33536
rect 66987 33487 67029 33496
rect 69867 33536 69909 33545
rect 69867 33496 69868 33536
rect 69908 33496 69909 33536
rect 69867 33487 69909 33496
rect 72843 33536 72885 33545
rect 72843 33496 72844 33536
rect 72884 33496 72885 33536
rect 72843 33487 72885 33496
rect 75147 33536 75189 33545
rect 75147 33496 75148 33536
rect 75188 33496 75189 33536
rect 75147 33487 75189 33496
rect 77835 33536 77877 33545
rect 77835 33496 77836 33536
rect 77876 33496 77877 33536
rect 77835 33487 77877 33496
rect 49227 33452 49269 33461
rect 49227 33412 49228 33452
rect 49268 33412 49269 33452
rect 49227 33403 49269 33412
rect 58923 33452 58965 33461
rect 58923 33412 58924 33452
rect 58964 33412 58965 33452
rect 58923 33403 58965 33412
rect 66699 33452 66741 33461
rect 66699 33412 66700 33452
rect 66740 33412 66741 33452
rect 66699 33403 66741 33412
rect 71979 33452 72021 33461
rect 71979 33412 71980 33452
rect 72020 33412 72021 33452
rect 71979 33403 72021 33412
rect 76011 33452 76053 33461
rect 76011 33412 76012 33452
rect 76052 33412 76053 33452
rect 76011 33403 76053 33412
rect 76683 33452 76725 33461
rect 76683 33412 76684 33452
rect 76724 33412 76725 33452
rect 76683 33403 76725 33412
rect 77259 33452 77301 33461
rect 77259 33412 77260 33452
rect 77300 33412 77301 33452
rect 77259 33403 77301 33412
rect 576 33284 79584 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79584 33284
rect 576 33220 79584 33244
rect 60931 33116 60989 33117
rect 60931 33076 60940 33116
rect 60980 33076 60989 33116
rect 60931 33075 60989 33076
rect 77155 33116 77213 33117
rect 77155 33076 77164 33116
rect 77204 33076 77213 33116
rect 77155 33075 77213 33076
rect 78411 33116 78453 33125
rect 78411 33076 78412 33116
rect 78452 33076 78453 33116
rect 78411 33067 78453 33076
rect 43851 33032 43893 33041
rect 43851 32992 43852 33032
rect 43892 32992 43893 33032
rect 43851 32983 43893 32992
rect 47107 33032 47165 33033
rect 47107 32992 47116 33032
rect 47156 32992 47165 33032
rect 47107 32991 47165 32992
rect 47307 33032 47349 33041
rect 47307 32992 47308 33032
rect 47348 32992 47349 33032
rect 47307 32983 47349 32992
rect 52299 33032 52341 33041
rect 52299 32992 52300 33032
rect 52340 32992 52341 33032
rect 52299 32983 52341 32992
rect 55083 33032 55125 33041
rect 55083 32992 55084 33032
rect 55124 32992 55125 33032
rect 55083 32983 55125 32992
rect 61131 33032 61173 33041
rect 61131 32992 61132 33032
rect 61172 32992 61173 33032
rect 61131 32983 61173 32992
rect 78115 33032 78173 33033
rect 78115 32992 78124 33032
rect 78164 32992 78173 33032
rect 78115 32991 78173 32992
rect 42691 32948 42749 32949
rect 42691 32908 42700 32948
rect 42740 32908 42749 32948
rect 42691 32907 42749 32908
rect 47787 32948 47829 32957
rect 47787 32908 47788 32948
rect 47828 32908 47829 32948
rect 47787 32899 47829 32908
rect 69195 32875 69237 32884
rect 45867 32864 45909 32873
rect 45867 32824 45868 32864
rect 45908 32824 45909 32864
rect 45867 32815 45909 32824
rect 46059 32864 46101 32873
rect 46059 32824 46060 32864
rect 46100 32824 46101 32864
rect 46059 32815 46101 32824
rect 46147 32864 46205 32865
rect 46147 32824 46156 32864
rect 46196 32824 46205 32864
rect 46147 32823 46205 32824
rect 46435 32864 46493 32865
rect 46435 32824 46444 32864
rect 46484 32824 46493 32864
rect 46435 32823 46493 32824
rect 46731 32864 46773 32873
rect 46731 32824 46732 32864
rect 46772 32824 46773 32864
rect 46731 32815 46773 32824
rect 46827 32864 46869 32873
rect 46827 32824 46828 32864
rect 46868 32824 46869 32864
rect 46827 32815 46869 32824
rect 47683 32864 47741 32865
rect 47683 32824 47692 32864
rect 47732 32824 47741 32864
rect 47683 32823 47741 32824
rect 47883 32864 47925 32873
rect 47883 32824 47884 32864
rect 47924 32824 47925 32864
rect 47883 32815 47925 32824
rect 48459 32864 48501 32873
rect 48459 32824 48460 32864
rect 48500 32824 48501 32864
rect 48459 32815 48501 32824
rect 48835 32864 48893 32865
rect 48835 32824 48844 32864
rect 48884 32824 48893 32864
rect 48835 32823 48893 32824
rect 49699 32864 49757 32865
rect 49699 32824 49708 32864
rect 49748 32824 49757 32864
rect 49699 32823 49757 32824
rect 51051 32864 51093 32873
rect 51051 32824 51052 32864
rect 51092 32824 51093 32864
rect 51051 32815 51093 32824
rect 51235 32864 51293 32865
rect 51235 32824 51244 32864
rect 51284 32824 51293 32864
rect 51235 32823 51293 32824
rect 52579 32864 52637 32865
rect 52579 32824 52588 32864
rect 52628 32824 52637 32864
rect 52579 32823 52637 32824
rect 53451 32864 53493 32873
rect 53451 32824 53452 32864
rect 53492 32824 53493 32864
rect 53451 32815 53493 32824
rect 53547 32864 53589 32873
rect 53547 32824 53548 32864
rect 53588 32824 53589 32864
rect 53547 32815 53589 32824
rect 53643 32864 53685 32873
rect 53643 32824 53644 32864
rect 53684 32824 53685 32864
rect 53643 32815 53685 32824
rect 53739 32864 53781 32873
rect 53739 32824 53740 32864
rect 53780 32824 53781 32864
rect 53739 32815 53781 32824
rect 54403 32864 54461 32865
rect 54403 32824 54412 32864
rect 54452 32824 54461 32864
rect 54403 32823 54461 32824
rect 54507 32864 54549 32873
rect 54507 32824 54508 32864
rect 54548 32824 54549 32864
rect 54507 32815 54549 32824
rect 54603 32864 54645 32873
rect 54603 32824 54604 32864
rect 54644 32824 54645 32864
rect 54603 32815 54645 32824
rect 54787 32864 54845 32865
rect 54787 32824 54796 32864
rect 54836 32824 54845 32864
rect 54787 32823 54845 32824
rect 54891 32864 54933 32873
rect 54891 32824 54892 32864
rect 54932 32824 54933 32864
rect 54891 32815 54933 32824
rect 55083 32864 55125 32873
rect 55083 32824 55084 32864
rect 55124 32824 55125 32864
rect 55083 32815 55125 32824
rect 55275 32864 55317 32873
rect 55275 32824 55276 32864
rect 55316 32824 55317 32864
rect 55275 32815 55317 32824
rect 55651 32864 55709 32865
rect 55651 32824 55660 32864
rect 55700 32824 55709 32864
rect 55651 32823 55709 32824
rect 56515 32864 56573 32865
rect 56515 32824 56524 32864
rect 56564 32824 56573 32864
rect 56515 32823 56573 32824
rect 58059 32864 58101 32873
rect 58059 32824 58060 32864
rect 58100 32824 58101 32864
rect 58059 32815 58101 32824
rect 58251 32864 58293 32873
rect 58251 32824 58252 32864
rect 58292 32824 58293 32864
rect 58251 32815 58293 32824
rect 58339 32864 58397 32865
rect 58339 32824 58348 32864
rect 58388 32824 58397 32864
rect 58339 32823 58397 32824
rect 58915 32864 58973 32865
rect 58915 32824 58924 32864
rect 58964 32824 58973 32864
rect 58915 32823 58973 32824
rect 59779 32864 59837 32865
rect 59779 32824 59788 32864
rect 59828 32824 59837 32864
rect 59779 32823 59837 32824
rect 62475 32864 62517 32873
rect 62475 32824 62476 32864
rect 62516 32824 62517 32864
rect 62475 32815 62517 32824
rect 62571 32864 62613 32873
rect 62571 32824 62572 32864
rect 62612 32824 62613 32864
rect 62571 32815 62613 32824
rect 62667 32864 62709 32873
rect 62667 32824 62668 32864
rect 62708 32824 62709 32864
rect 62667 32815 62709 32824
rect 62859 32864 62901 32873
rect 62859 32824 62860 32864
rect 62900 32824 62901 32864
rect 62859 32815 62901 32824
rect 63043 32864 63101 32865
rect 63043 32824 63052 32864
rect 63092 32824 63101 32864
rect 63043 32823 63101 32824
rect 63619 32864 63677 32865
rect 63619 32824 63628 32864
rect 63668 32824 63677 32864
rect 63619 32823 63677 32824
rect 64483 32864 64541 32865
rect 64483 32824 64492 32864
rect 64532 32824 64541 32864
rect 64483 32823 64541 32824
rect 65835 32864 65877 32873
rect 65835 32824 65836 32864
rect 65876 32824 65877 32864
rect 65835 32815 65877 32824
rect 65931 32864 65973 32873
rect 65931 32824 65932 32864
rect 65972 32824 65973 32864
rect 65931 32815 65973 32824
rect 66027 32864 66069 32873
rect 66027 32824 66028 32864
rect 66068 32824 66069 32864
rect 66027 32815 66069 32824
rect 66123 32864 66165 32873
rect 66123 32824 66124 32864
rect 66164 32824 66165 32864
rect 66123 32815 66165 32824
rect 66315 32864 66357 32873
rect 66315 32824 66316 32864
rect 66356 32824 66357 32864
rect 66315 32815 66357 32824
rect 66691 32864 66749 32865
rect 66691 32824 66700 32864
rect 66740 32824 66749 32864
rect 66691 32823 66749 32824
rect 67555 32864 67613 32865
rect 67555 32824 67564 32864
rect 67604 32824 67613 32864
rect 67555 32823 67613 32824
rect 68899 32864 68957 32865
rect 68899 32824 68908 32864
rect 68948 32824 68957 32864
rect 68899 32823 68957 32824
rect 69003 32864 69045 32873
rect 69003 32824 69004 32864
rect 69044 32824 69045 32864
rect 69195 32835 69196 32875
rect 69236 32835 69237 32875
rect 69195 32826 69237 32835
rect 69763 32864 69821 32865
rect 69003 32815 69045 32824
rect 69763 32824 69772 32864
rect 69812 32824 69821 32864
rect 69763 32823 69821 32824
rect 70627 32864 70685 32865
rect 70627 32824 70636 32864
rect 70676 32824 70685 32864
rect 70627 32823 70685 32824
rect 72171 32864 72213 32873
rect 72171 32824 72172 32864
rect 72212 32824 72213 32864
rect 72171 32815 72213 32824
rect 72547 32864 72605 32865
rect 72547 32824 72556 32864
rect 72596 32824 72605 32864
rect 72547 32823 72605 32824
rect 73411 32864 73469 32865
rect 73411 32824 73420 32864
rect 73460 32824 73469 32864
rect 73411 32823 73469 32824
rect 74763 32864 74805 32873
rect 74763 32824 74764 32864
rect 74804 32824 74805 32864
rect 74763 32815 74805 32824
rect 75139 32864 75197 32865
rect 75139 32824 75148 32864
rect 75188 32824 75197 32864
rect 75139 32823 75197 32824
rect 76003 32864 76061 32865
rect 76003 32824 76012 32864
rect 76052 32824 76061 32864
rect 76003 32823 76061 32824
rect 77443 32864 77501 32865
rect 77443 32824 77452 32864
rect 77492 32824 77501 32864
rect 77443 32823 77501 32824
rect 77739 32864 77781 32873
rect 77739 32824 77740 32864
rect 77780 32824 77781 32864
rect 77739 32815 77781 32824
rect 77835 32864 77877 32873
rect 77835 32824 77836 32864
rect 77876 32824 77877 32864
rect 77835 32815 77877 32824
rect 78307 32864 78365 32865
rect 78307 32824 78316 32864
rect 78356 32824 78365 32864
rect 78307 32823 78365 32824
rect 78507 32864 78549 32873
rect 78507 32824 78508 32864
rect 78548 32824 78549 32864
rect 78507 32815 78549 32824
rect 51147 32780 51189 32789
rect 51147 32740 51148 32780
rect 51188 32740 51189 32780
rect 51147 32731 51189 32740
rect 58155 32780 58197 32789
rect 58155 32740 58156 32780
rect 58196 32740 58197 32780
rect 58155 32731 58197 32740
rect 58539 32780 58581 32789
rect 58539 32740 58540 32780
rect 58580 32740 58581 32780
rect 58539 32731 58581 32740
rect 62955 32780 62997 32789
rect 62955 32740 62956 32780
rect 62996 32740 62997 32780
rect 62955 32731 62997 32740
rect 63243 32780 63285 32789
rect 63243 32740 63244 32780
rect 63284 32740 63285 32780
rect 63243 32731 63285 32740
rect 69387 32780 69429 32789
rect 69387 32740 69388 32780
rect 69428 32740 69429 32780
rect 69387 32731 69429 32740
rect 42891 32696 42933 32705
rect 42891 32656 42892 32696
rect 42932 32656 42933 32696
rect 42891 32647 42933 32656
rect 45955 32696 46013 32697
rect 45955 32656 45964 32696
rect 46004 32656 46013 32696
rect 45955 32655 46013 32656
rect 50851 32696 50909 32697
rect 50851 32656 50860 32696
rect 50900 32656 50909 32696
rect 50851 32655 50909 32656
rect 57667 32696 57725 32697
rect 57667 32656 57676 32696
rect 57716 32656 57725 32696
rect 57667 32655 57725 32656
rect 60931 32696 60989 32697
rect 60931 32656 60940 32696
rect 60980 32656 60989 32696
rect 60931 32655 60989 32656
rect 62371 32696 62429 32697
rect 62371 32656 62380 32696
rect 62420 32656 62429 32696
rect 62371 32655 62429 32656
rect 65635 32696 65693 32697
rect 65635 32656 65644 32696
rect 65684 32656 65693 32696
rect 65635 32655 65693 32656
rect 68707 32696 68765 32697
rect 68707 32656 68716 32696
rect 68756 32656 68765 32696
rect 68707 32655 68765 32656
rect 69091 32696 69149 32697
rect 69091 32656 69100 32696
rect 69140 32656 69149 32696
rect 69091 32655 69149 32656
rect 71779 32696 71837 32697
rect 71779 32656 71788 32696
rect 71828 32656 71837 32696
rect 71779 32655 71837 32656
rect 74563 32696 74621 32697
rect 74563 32656 74572 32696
rect 74612 32656 74621 32696
rect 74563 32655 74621 32656
rect 576 32528 79584 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79584 32528
rect 576 32464 79584 32488
rect 66507 32402 66549 32411
rect 48643 32360 48701 32361
rect 48643 32320 48652 32360
rect 48692 32320 48701 32360
rect 48643 32319 48701 32320
rect 49611 32360 49653 32369
rect 66507 32362 66508 32402
rect 66548 32362 66549 32402
rect 49611 32320 49612 32360
rect 49652 32320 49653 32360
rect 49611 32311 49653 32320
rect 53539 32360 53597 32361
rect 53539 32320 53548 32360
rect 53588 32320 53597 32360
rect 53539 32319 53597 32320
rect 62755 32360 62813 32361
rect 62755 32320 62764 32360
rect 62804 32320 62813 32360
rect 62755 32319 62813 32320
rect 64003 32360 64061 32361
rect 64003 32320 64012 32360
rect 64052 32320 64061 32360
rect 66507 32353 66549 32362
rect 75907 32360 75965 32361
rect 64003 32319 64061 32320
rect 75907 32320 75916 32360
rect 75956 32320 75965 32360
rect 75907 32319 75965 32320
rect 46059 32276 46101 32285
rect 46059 32236 46060 32276
rect 46100 32236 46101 32276
rect 46059 32227 46101 32236
rect 50475 32276 50517 32285
rect 50475 32236 50476 32276
rect 50516 32236 50517 32276
rect 50475 32227 50517 32236
rect 58731 32276 58773 32285
rect 58731 32236 58732 32276
rect 58772 32236 58773 32276
rect 58731 32227 58773 32236
rect 66219 32276 66261 32285
rect 66219 32236 66220 32276
rect 66260 32236 66261 32276
rect 63339 32219 63381 32228
rect 66219 32227 66261 32236
rect 72075 32276 72117 32285
rect 72075 32236 72076 32276
rect 72116 32236 72117 32276
rect 72075 32227 72117 32236
rect 77067 32276 77109 32285
rect 77067 32236 77068 32276
rect 77108 32236 77109 32276
rect 77067 32227 77109 32236
rect 42315 32192 42357 32201
rect 42315 32152 42316 32192
rect 42356 32152 42357 32192
rect 42315 32143 42357 32152
rect 42411 32192 42453 32201
rect 42411 32152 42412 32192
rect 42452 32152 42453 32192
rect 42411 32143 42453 32152
rect 42507 32192 42549 32201
rect 42507 32152 42508 32192
rect 42548 32152 42549 32192
rect 42507 32143 42549 32152
rect 42603 32192 42645 32201
rect 42603 32152 42604 32192
rect 42644 32152 42645 32192
rect 42603 32143 42645 32152
rect 42891 32192 42933 32201
rect 42891 32152 42892 32192
rect 42932 32152 42933 32192
rect 42891 32143 42933 32152
rect 43075 32192 43133 32193
rect 43075 32152 43084 32192
rect 43124 32152 43133 32192
rect 43075 32151 43133 32152
rect 43371 32192 43413 32201
rect 43371 32152 43372 32192
rect 43412 32152 43413 32192
rect 43371 32143 43413 32152
rect 43747 32192 43805 32193
rect 43747 32152 43756 32192
rect 43796 32152 43805 32192
rect 43747 32151 43805 32152
rect 44611 32192 44669 32193
rect 44611 32152 44620 32192
rect 44660 32152 44669 32192
rect 44611 32151 44669 32152
rect 46435 32192 46493 32193
rect 46435 32152 46444 32192
rect 46484 32152 46493 32192
rect 46435 32151 46493 32152
rect 47299 32192 47357 32193
rect 47299 32152 47308 32192
rect 47348 32152 47357 32192
rect 47299 32151 47357 32152
rect 48747 32192 48789 32201
rect 48747 32152 48748 32192
rect 48788 32152 48789 32192
rect 48747 32143 48789 32152
rect 48843 32192 48885 32201
rect 48843 32152 48844 32192
rect 48884 32152 48885 32192
rect 48843 32143 48885 32152
rect 48939 32192 48981 32201
rect 48939 32152 48940 32192
rect 48980 32152 48981 32192
rect 48939 32143 48981 32152
rect 49123 32192 49181 32193
rect 49123 32152 49132 32192
rect 49172 32152 49181 32192
rect 49123 32151 49181 32152
rect 50083 32192 50141 32193
rect 50083 32152 50092 32192
rect 50132 32152 50141 32192
rect 50083 32151 50141 32152
rect 50379 32192 50421 32201
rect 50379 32152 50380 32192
rect 50420 32152 50421 32192
rect 50379 32143 50421 32152
rect 50563 32192 50621 32193
rect 50563 32152 50572 32192
rect 50612 32152 50621 32192
rect 50563 32151 50621 32152
rect 51147 32192 51189 32201
rect 51147 32152 51148 32192
rect 51188 32152 51189 32192
rect 51147 32143 51189 32152
rect 51523 32192 51581 32193
rect 51523 32152 51532 32192
rect 51572 32152 51581 32192
rect 51523 32151 51581 32152
rect 52387 32192 52445 32193
rect 52387 32152 52396 32192
rect 52436 32152 52445 32192
rect 52387 32151 52445 32152
rect 54219 32192 54261 32201
rect 54219 32152 54220 32192
rect 54260 32152 54261 32192
rect 54219 32143 54261 32152
rect 54411 32192 54453 32201
rect 54411 32152 54412 32192
rect 54452 32152 54453 32192
rect 54411 32143 54453 32152
rect 54499 32192 54557 32193
rect 54499 32152 54508 32192
rect 54548 32152 54557 32192
rect 54499 32151 54557 32152
rect 54699 32192 54741 32201
rect 54699 32152 54700 32192
rect 54740 32152 54741 32192
rect 54699 32143 54741 32152
rect 54795 32192 54837 32201
rect 54795 32152 54796 32192
rect 54836 32152 54837 32192
rect 54795 32143 54837 32152
rect 54891 32192 54933 32201
rect 54891 32152 54892 32192
rect 54932 32152 54933 32192
rect 54891 32143 54933 32152
rect 54987 32192 55029 32201
rect 54987 32152 54988 32192
rect 55028 32152 55029 32192
rect 54987 32143 55029 32152
rect 55651 32192 55709 32193
rect 55651 32152 55660 32192
rect 55700 32152 55709 32192
rect 55651 32151 55709 32152
rect 55851 32192 55893 32201
rect 55851 32152 55852 32192
rect 55892 32152 55893 32192
rect 55851 32143 55893 32152
rect 58339 32192 58397 32193
rect 58339 32152 58348 32192
rect 58388 32152 58397 32192
rect 58339 32151 58397 32152
rect 58635 32192 58677 32201
rect 58635 32152 58636 32192
rect 58676 32152 58677 32192
rect 58635 32143 58677 32152
rect 59211 32192 59253 32201
rect 59211 32152 59212 32192
rect 59252 32152 59253 32192
rect 59211 32143 59253 32152
rect 59395 32192 59453 32193
rect 59395 32152 59404 32192
rect 59444 32152 59453 32192
rect 59395 32151 59453 32152
rect 59587 32192 59645 32193
rect 59587 32152 59596 32192
rect 59636 32152 59645 32192
rect 59587 32151 59645 32152
rect 59691 32192 59733 32201
rect 59691 32152 59692 32192
rect 59732 32152 59733 32192
rect 59691 32143 59733 32152
rect 59883 32192 59925 32201
rect 59883 32152 59884 32192
rect 59924 32152 59925 32192
rect 59883 32143 59925 32152
rect 60363 32192 60405 32201
rect 60363 32152 60364 32192
rect 60404 32152 60405 32192
rect 60363 32143 60405 32152
rect 60739 32192 60797 32193
rect 60739 32152 60748 32192
rect 60788 32152 60797 32192
rect 60739 32151 60797 32152
rect 61603 32192 61661 32193
rect 61603 32152 61612 32192
rect 61652 32152 61661 32192
rect 61603 32151 61661 32152
rect 63243 32192 63285 32201
rect 63243 32152 63244 32192
rect 63284 32152 63285 32192
rect 63339 32179 63340 32219
rect 63380 32179 63381 32219
rect 63339 32170 63381 32179
rect 63619 32192 63677 32193
rect 63243 32143 63285 32152
rect 63619 32152 63628 32192
rect 63668 32152 63677 32192
rect 63619 32151 63677 32152
rect 63915 32192 63957 32201
rect 63915 32152 63916 32192
rect 63956 32152 63957 32192
rect 63915 32143 63957 32152
rect 64107 32192 64149 32201
rect 64107 32152 64108 32192
rect 64148 32152 64149 32192
rect 64107 32143 64149 32152
rect 64195 32192 64253 32193
rect 64195 32152 64204 32192
rect 64244 32152 64253 32192
rect 64195 32151 64253 32152
rect 64387 32192 64445 32193
rect 64387 32152 64396 32192
rect 64436 32152 64445 32192
rect 64387 32151 64445 32152
rect 64587 32192 64629 32201
rect 64587 32152 64588 32192
rect 64628 32152 64629 32192
rect 64587 32143 64629 32152
rect 65827 32192 65885 32193
rect 65827 32152 65836 32192
rect 65876 32152 65885 32192
rect 65827 32151 65885 32152
rect 66123 32192 66165 32201
rect 66123 32152 66124 32192
rect 66164 32152 66165 32192
rect 66123 32143 66165 32152
rect 66699 32192 66741 32201
rect 66699 32152 66700 32192
rect 66740 32152 66741 32192
rect 66699 32143 66741 32152
rect 67075 32192 67133 32193
rect 67075 32152 67084 32192
rect 67124 32152 67133 32192
rect 67075 32151 67133 32152
rect 67939 32192 67997 32193
rect 67939 32152 67948 32192
rect 67988 32152 67997 32192
rect 67939 32151 67997 32152
rect 69763 32192 69821 32193
rect 69763 32152 69772 32192
rect 69812 32152 69821 32192
rect 69763 32151 69821 32152
rect 69867 32192 69909 32201
rect 69867 32152 69868 32192
rect 69908 32152 69909 32192
rect 69867 32143 69909 32152
rect 70059 32192 70101 32201
rect 70059 32152 70060 32192
rect 70100 32152 70101 32192
rect 70059 32143 70101 32152
rect 70251 32192 70293 32201
rect 70251 32152 70252 32192
rect 70292 32152 70293 32192
rect 70251 32143 70293 32152
rect 70347 32192 70389 32201
rect 70347 32152 70348 32192
rect 70388 32152 70389 32192
rect 70347 32143 70389 32152
rect 70443 32192 70485 32201
rect 70443 32152 70444 32192
rect 70484 32152 70485 32192
rect 70443 32143 70485 32152
rect 70539 32192 70581 32201
rect 70539 32152 70540 32192
rect 70580 32152 70581 32192
rect 70539 32143 70581 32152
rect 70731 32192 70773 32201
rect 70731 32152 70732 32192
rect 70772 32152 70773 32192
rect 70731 32143 70773 32152
rect 70923 32192 70965 32201
rect 70923 32152 70924 32192
rect 70964 32152 70965 32192
rect 70923 32143 70965 32152
rect 71011 32192 71069 32193
rect 71011 32152 71020 32192
rect 71060 32152 71069 32192
rect 71011 32151 71069 32152
rect 71683 32192 71741 32193
rect 71683 32152 71692 32192
rect 71732 32152 71741 32192
rect 71683 32151 71741 32152
rect 71979 32192 72021 32201
rect 71979 32152 71980 32192
rect 72020 32152 72021 32192
rect 71979 32143 72021 32152
rect 72547 32192 72605 32193
rect 72547 32152 72556 32192
rect 72596 32152 72605 32192
rect 72547 32151 72605 32152
rect 72747 32192 72789 32201
rect 72747 32152 72748 32192
rect 72788 32152 72789 32192
rect 72747 32143 72789 32152
rect 75819 32192 75861 32201
rect 75819 32152 75820 32192
rect 75860 32152 75861 32192
rect 75819 32143 75861 32152
rect 76011 32192 76053 32201
rect 76011 32152 76012 32192
rect 76052 32152 76053 32192
rect 76011 32143 76053 32152
rect 76099 32192 76157 32193
rect 76099 32152 76108 32192
rect 76148 32152 76157 32192
rect 76099 32151 76157 32152
rect 77443 32192 77501 32193
rect 77443 32152 77452 32192
rect 77492 32152 77501 32192
rect 77443 32151 77501 32152
rect 78307 32192 78365 32193
rect 78307 32152 78316 32192
rect 78356 32152 78365 32192
rect 78307 32151 78365 32152
rect 40683 32024 40725 32033
rect 40683 31984 40684 32024
rect 40724 31984 40725 32024
rect 40683 31975 40725 31984
rect 54219 32024 54261 32033
rect 54219 31984 54220 32024
rect 54260 31984 54261 32024
rect 54219 31975 54261 31984
rect 59011 32024 59069 32025
rect 59011 31984 59020 32024
rect 59060 31984 59069 32024
rect 59011 31983 59069 31984
rect 59307 32024 59349 32033
rect 59307 31984 59308 32024
rect 59348 31984 59349 32024
rect 59307 31975 59349 31984
rect 62947 32024 63005 32025
rect 62947 31984 62956 32024
rect 62996 31984 63005 32024
rect 62947 31983 63005 31984
rect 64491 32024 64533 32033
rect 64491 31984 64492 32024
rect 64532 31984 64533 32024
rect 64491 31975 64533 31984
rect 70059 32024 70101 32033
rect 70059 31984 70060 32024
rect 70100 31984 70101 32024
rect 70059 31975 70101 31984
rect 72355 32024 72413 32025
rect 72355 31984 72364 32024
rect 72404 31984 72413 32024
rect 72355 31983 72413 31984
rect 74091 32024 74133 32033
rect 74091 31984 74092 32024
rect 74132 31984 74133 32024
rect 74091 31975 74133 31984
rect 42987 31940 43029 31949
rect 42987 31900 42988 31940
rect 43028 31900 43029 31940
rect 42987 31891 43029 31900
rect 45763 31940 45821 31941
rect 45763 31900 45772 31940
rect 45812 31900 45821 31940
rect 45763 31899 45821 31900
rect 48451 31940 48509 31941
rect 48451 31900 48460 31940
rect 48500 31900 48509 31940
rect 48451 31899 48509 31900
rect 53539 31940 53597 31941
rect 53539 31900 53548 31940
rect 53588 31900 53597 31940
rect 53539 31899 53597 31900
rect 55755 31940 55797 31949
rect 55755 31900 55756 31940
rect 55796 31900 55797 31940
rect 55755 31891 55797 31900
rect 59883 31940 59925 31949
rect 59883 31900 59884 31940
rect 59924 31900 59925 31940
rect 59883 31891 59925 31900
rect 69091 31940 69149 31941
rect 69091 31900 69100 31940
rect 69140 31900 69149 31940
rect 69091 31899 69149 31900
rect 70731 31940 70773 31949
rect 70731 31900 70732 31940
rect 70772 31900 70773 31940
rect 70731 31891 70773 31900
rect 72651 31940 72693 31949
rect 72651 31900 72652 31940
rect 72692 31900 72693 31940
rect 72651 31891 72693 31900
rect 79459 31940 79517 31941
rect 79459 31900 79468 31940
rect 79508 31900 79517 31940
rect 79459 31899 79517 31900
rect 576 31772 79584 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79584 31772
rect 576 31708 79584 31732
rect 42787 31604 42845 31605
rect 42787 31564 42796 31604
rect 42836 31564 42845 31604
rect 42787 31563 42845 31564
rect 44043 31604 44085 31613
rect 44043 31564 44044 31604
rect 44084 31564 44085 31604
rect 44043 31555 44085 31564
rect 46731 31604 46773 31613
rect 46731 31564 46732 31604
rect 46772 31564 46773 31604
rect 46731 31555 46773 31564
rect 49227 31604 49269 31613
rect 49227 31564 49228 31604
rect 49268 31564 49269 31604
rect 49227 31555 49269 31564
rect 50179 31604 50237 31605
rect 50179 31564 50188 31604
rect 50228 31564 50237 31604
rect 50179 31563 50237 31564
rect 51435 31604 51477 31613
rect 51435 31564 51436 31604
rect 51476 31564 51477 31604
rect 51435 31555 51477 31564
rect 55267 31604 55325 31605
rect 55267 31564 55276 31604
rect 55316 31564 55325 31604
rect 55267 31563 55325 31564
rect 60267 31604 60309 31613
rect 60267 31564 60268 31604
rect 60308 31564 60309 31604
rect 60267 31555 60309 31564
rect 60843 31604 60885 31613
rect 60843 31564 60844 31604
rect 60884 31564 60885 31604
rect 60843 31555 60885 31564
rect 66315 31604 66357 31613
rect 66315 31564 66316 31604
rect 66356 31564 66357 31604
rect 66315 31555 66357 31564
rect 71403 31604 71445 31613
rect 71403 31564 71404 31604
rect 71444 31564 71445 31604
rect 71403 31555 71445 31564
rect 72075 31604 72117 31613
rect 72075 31564 72076 31604
rect 72116 31564 72117 31604
rect 72075 31555 72117 31564
rect 76003 31604 76061 31605
rect 76003 31564 76012 31604
rect 76052 31564 76061 31604
rect 76003 31563 76061 31564
rect 77931 31604 77973 31613
rect 77931 31564 77932 31604
rect 77972 31564 77973 31604
rect 77931 31555 77973 31564
rect 51627 31520 51669 31529
rect 51627 31480 51628 31520
rect 51668 31480 51669 31520
rect 51627 31471 51669 31480
rect 63051 31520 63093 31529
rect 63051 31480 63052 31520
rect 63092 31480 63093 31520
rect 63051 31471 63093 31480
rect 63531 31520 63573 31529
rect 63531 31480 63532 31520
rect 63572 31480 63573 31520
rect 63531 31471 63573 31480
rect 66891 31520 66933 31529
rect 66891 31480 66892 31520
rect 66932 31480 66933 31520
rect 66891 31471 66933 31480
rect 67179 31520 67221 31529
rect 67179 31480 67180 31520
rect 67220 31480 67221 31520
rect 67179 31471 67221 31480
rect 68715 31520 68757 31529
rect 68715 31480 68716 31520
rect 68756 31480 68757 31520
rect 68715 31471 68757 31480
rect 71115 31520 71157 31529
rect 71115 31480 71116 31520
rect 71156 31480 71157 31520
rect 71115 31471 71157 31480
rect 72267 31520 72309 31529
rect 72267 31480 72268 31520
rect 72308 31480 72309 31520
rect 72267 31471 72309 31480
rect 60067 31436 60125 31437
rect 60067 31396 60076 31436
rect 60116 31396 60125 31436
rect 60067 31395 60125 31396
rect 60643 31436 60701 31437
rect 60643 31396 60652 31436
rect 60692 31396 60701 31436
rect 60643 31395 60701 31396
rect 71875 31436 71933 31437
rect 71875 31396 71884 31436
rect 71924 31396 71933 31436
rect 71875 31395 71933 31396
rect 40579 31352 40637 31353
rect 40579 31312 40588 31352
rect 40628 31312 40637 31352
rect 40579 31311 40637 31312
rect 41443 31352 41501 31353
rect 41443 31312 41452 31352
rect 41492 31312 41501 31352
rect 43459 31352 43517 31353
rect 41443 31311 41501 31312
rect 43179 31325 43221 31334
rect 43179 31285 43180 31325
rect 43220 31285 43221 31325
rect 43459 31312 43468 31352
rect 43508 31312 43517 31352
rect 43459 31311 43517 31312
rect 43747 31352 43805 31353
rect 43747 31312 43756 31352
rect 43796 31312 43805 31352
rect 43747 31311 43805 31312
rect 43851 31352 43893 31361
rect 43851 31312 43852 31352
rect 43892 31312 43893 31352
rect 43851 31303 43893 31312
rect 44043 31352 44085 31361
rect 44043 31312 44044 31352
rect 44084 31312 44085 31352
rect 44043 31303 44085 31312
rect 46627 31352 46685 31353
rect 46627 31312 46636 31352
rect 46676 31312 46685 31352
rect 46627 31311 46685 31312
rect 46827 31352 46869 31361
rect 46827 31312 46828 31352
rect 46868 31312 46869 31352
rect 46827 31303 46869 31312
rect 48547 31352 48605 31353
rect 48547 31312 48556 31352
rect 48596 31312 48605 31352
rect 48547 31311 48605 31312
rect 48931 31352 48989 31353
rect 48931 31312 48940 31352
rect 48980 31312 48989 31352
rect 48931 31311 48989 31312
rect 49035 31352 49077 31361
rect 49035 31312 49036 31352
rect 49076 31312 49077 31352
rect 49035 31303 49077 31312
rect 49227 31352 49269 31361
rect 49227 31312 49228 31352
rect 49268 31312 49269 31352
rect 49227 31303 49269 31312
rect 49707 31352 49749 31361
rect 49707 31312 49708 31352
rect 49748 31312 49749 31352
rect 49707 31303 49749 31312
rect 49899 31352 49941 31361
rect 49899 31312 49900 31352
rect 49940 31312 49941 31352
rect 49899 31303 49941 31312
rect 49987 31352 50045 31353
rect 49987 31312 49996 31352
rect 50036 31312 50045 31352
rect 49987 31311 50045 31312
rect 50475 31352 50517 31361
rect 50475 31312 50476 31352
rect 50516 31312 50517 31352
rect 50475 31303 50517 31312
rect 50571 31352 50613 31361
rect 50571 31312 50572 31352
rect 50612 31312 50613 31352
rect 50571 31303 50613 31312
rect 50851 31352 50909 31353
rect 50851 31312 50860 31352
rect 50900 31312 50909 31352
rect 50851 31311 50909 31312
rect 51139 31352 51197 31353
rect 51139 31312 51148 31352
rect 51188 31312 51197 31352
rect 51139 31311 51197 31312
rect 51243 31352 51285 31361
rect 51243 31312 51244 31352
rect 51284 31312 51285 31352
rect 51243 31303 51285 31312
rect 51435 31352 51477 31361
rect 51435 31312 51436 31352
rect 51476 31312 51477 31352
rect 54115 31352 54173 31353
rect 51435 31303 51477 31312
rect 53251 31339 53309 31340
rect 53251 31299 53260 31339
rect 53300 31299 53309 31339
rect 54115 31312 54124 31352
rect 54164 31312 54173 31352
rect 54115 31311 54173 31312
rect 55659 31352 55701 31361
rect 55659 31312 55660 31352
rect 55700 31312 55701 31352
rect 55659 31303 55701 31312
rect 55851 31352 55893 31361
rect 55851 31312 55852 31352
rect 55892 31312 55893 31352
rect 55851 31303 55893 31312
rect 55939 31352 55997 31353
rect 55939 31312 55948 31352
rect 55988 31312 55997 31352
rect 55939 31311 55997 31312
rect 56515 31352 56573 31353
rect 56515 31312 56524 31352
rect 56564 31312 56573 31352
rect 56515 31311 56573 31312
rect 57379 31352 57437 31353
rect 57379 31312 57388 31352
rect 57428 31312 57437 31352
rect 57379 31311 57437 31312
rect 59595 31352 59637 31361
rect 59595 31312 59596 31352
rect 59636 31312 59637 31352
rect 59595 31303 59637 31312
rect 59691 31352 59733 31361
rect 59691 31312 59692 31352
rect 59732 31312 59733 31352
rect 59691 31303 59733 31312
rect 59787 31352 59829 31361
rect 59787 31312 59788 31352
rect 59828 31312 59829 31352
rect 59787 31303 59829 31312
rect 62475 31352 62517 31361
rect 62475 31312 62476 31352
rect 62516 31312 62517 31352
rect 62475 31303 62517 31312
rect 62667 31352 62709 31361
rect 62667 31312 62668 31352
rect 62708 31312 62709 31352
rect 62667 31303 62709 31312
rect 62755 31352 62813 31353
rect 62755 31312 62764 31352
rect 62804 31312 62813 31352
rect 63243 31352 63285 31361
rect 62755 31311 62813 31312
rect 63051 31314 63093 31323
rect 53251 31298 53309 31299
rect 40203 31268 40245 31277
rect 40203 31228 40204 31268
rect 40244 31228 40245 31268
rect 40203 31219 40245 31228
rect 43083 31268 43125 31277
rect 43179 31276 43221 31285
rect 43083 31228 43084 31268
rect 43124 31228 43125 31268
rect 43083 31219 43125 31228
rect 52875 31268 52917 31277
rect 52875 31228 52876 31268
rect 52916 31228 52917 31268
rect 52875 31219 52917 31228
rect 56139 31268 56181 31277
rect 56139 31228 56140 31268
rect 56180 31228 56181 31268
rect 56139 31219 56181 31228
rect 62571 31268 62613 31277
rect 62571 31228 62572 31268
rect 62612 31228 62613 31268
rect 63051 31274 63052 31314
rect 63092 31274 63093 31314
rect 63243 31312 63244 31352
rect 63284 31312 63285 31352
rect 66315 31352 66357 31361
rect 63243 31303 63285 31312
rect 63331 31337 63389 31338
rect 63331 31297 63340 31337
rect 63380 31297 63389 31337
rect 66315 31312 66316 31352
rect 66356 31312 66357 31352
rect 66315 31303 66357 31312
rect 66507 31352 66549 31361
rect 66507 31312 66508 31352
rect 66548 31312 66549 31352
rect 66507 31303 66549 31312
rect 66595 31352 66653 31353
rect 66595 31312 66604 31352
rect 66644 31312 66653 31352
rect 66595 31311 66653 31312
rect 66787 31352 66845 31353
rect 66787 31312 66796 31352
rect 66836 31312 66845 31352
rect 66787 31311 66845 31312
rect 66987 31352 67029 31361
rect 66987 31312 66988 31352
rect 67028 31312 67029 31352
rect 66987 31303 67029 31312
rect 70539 31352 70581 31361
rect 70539 31312 70540 31352
rect 70580 31312 70581 31352
rect 70539 31303 70581 31312
rect 70731 31352 70773 31361
rect 70731 31312 70732 31352
rect 70772 31312 70773 31352
rect 70731 31303 70773 31312
rect 70819 31352 70877 31353
rect 70819 31312 70828 31352
rect 70868 31312 70877 31352
rect 70819 31311 70877 31312
rect 71019 31352 71061 31361
rect 71019 31312 71020 31352
rect 71060 31312 71061 31352
rect 71019 31303 71061 31312
rect 71203 31352 71261 31353
rect 71203 31312 71212 31352
rect 71252 31312 71261 31352
rect 71203 31311 71261 31312
rect 71403 31352 71445 31361
rect 71403 31312 71404 31352
rect 71444 31312 71445 31352
rect 71403 31303 71445 31312
rect 71595 31352 71637 31361
rect 71595 31312 71596 31352
rect 71636 31312 71637 31352
rect 73987 31352 74045 31353
rect 71595 31303 71637 31312
rect 71683 31337 71741 31338
rect 63331 31296 63389 31297
rect 71683 31297 71692 31337
rect 71732 31297 71741 31337
rect 73987 31312 73996 31352
rect 74036 31312 74045 31352
rect 73987 31311 74045 31312
rect 74851 31352 74909 31353
rect 74851 31312 74860 31352
rect 74900 31312 74909 31352
rect 74851 31311 74909 31312
rect 76971 31352 77013 31361
rect 76971 31312 76972 31352
rect 77012 31312 77013 31352
rect 76971 31303 77013 31312
rect 77155 31352 77213 31353
rect 77155 31312 77164 31352
rect 77204 31312 77213 31352
rect 77155 31311 77213 31312
rect 77443 31352 77501 31353
rect 77443 31312 77452 31352
rect 77492 31312 77501 31352
rect 77443 31311 77501 31312
rect 77643 31352 77685 31361
rect 77643 31312 77644 31352
rect 77684 31312 77685 31352
rect 77643 31303 77685 31312
rect 77827 31352 77885 31353
rect 77827 31312 77836 31352
rect 77876 31312 77885 31352
rect 77827 31311 77885 31312
rect 78027 31352 78069 31361
rect 78027 31312 78028 31352
rect 78068 31312 78069 31352
rect 78027 31303 78069 31312
rect 71683 31296 71741 31297
rect 63051 31265 63093 31274
rect 73611 31268 73653 31277
rect 62571 31219 62613 31228
rect 73611 31228 73612 31268
rect 73652 31228 73653 31268
rect 73611 31219 73653 31228
rect 77067 31268 77109 31277
rect 77067 31228 77068 31268
rect 77108 31228 77109 31268
rect 77067 31219 77109 31228
rect 77547 31268 77589 31277
rect 77547 31228 77548 31268
rect 77588 31228 77589 31268
rect 77547 31219 77589 31228
rect 42595 31184 42653 31185
rect 42595 31144 42604 31184
rect 42644 31144 42653 31184
rect 42595 31143 42653 31144
rect 49795 31184 49853 31185
rect 49795 31144 49804 31184
rect 49844 31144 49853 31184
rect 49795 31143 49853 31144
rect 55267 31184 55325 31185
rect 55267 31144 55276 31184
rect 55316 31144 55325 31184
rect 55267 31143 55325 31144
rect 55747 31184 55805 31185
rect 55747 31144 55756 31184
rect 55796 31144 55805 31184
rect 55747 31143 55805 31144
rect 58531 31184 58589 31185
rect 58531 31144 58540 31184
rect 58580 31144 58589 31184
rect 58531 31143 58589 31144
rect 59875 31184 59933 31185
rect 59875 31144 59884 31184
rect 59924 31144 59933 31184
rect 59875 31143 59933 31144
rect 60267 31184 60309 31193
rect 60267 31144 60268 31184
rect 60308 31144 60309 31184
rect 60267 31135 60309 31144
rect 60843 31184 60885 31193
rect 60843 31144 60844 31184
rect 60884 31144 60885 31184
rect 60843 31135 60885 31144
rect 70627 31184 70685 31185
rect 70627 31144 70636 31184
rect 70676 31144 70685 31184
rect 70627 31143 70685 31144
rect 76003 31184 76061 31185
rect 76003 31144 76012 31184
rect 76052 31144 76061 31184
rect 76003 31143 76061 31144
rect 576 31016 79584 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79584 31016
rect 576 30952 79584 30976
rect 76875 30890 76917 30899
rect 42507 30848 42549 30857
rect 42507 30808 42508 30848
rect 42548 30808 42549 30848
rect 42507 30799 42549 30808
rect 42787 30848 42845 30849
rect 42787 30808 42796 30848
rect 42836 30808 42845 30848
rect 42787 30807 42845 30808
rect 49227 30848 49269 30857
rect 49227 30808 49228 30848
rect 49268 30808 49269 30848
rect 49227 30799 49269 30808
rect 50379 30848 50421 30857
rect 50379 30808 50380 30848
rect 50420 30808 50421 30848
rect 50379 30799 50421 30808
rect 51531 30848 51573 30857
rect 51531 30808 51532 30848
rect 51572 30808 51573 30848
rect 51531 30799 51573 30808
rect 57955 30848 58013 30849
rect 57955 30808 57964 30848
rect 58004 30808 58013 30848
rect 57955 30807 58013 30808
rect 70819 30848 70877 30849
rect 70819 30808 70828 30848
rect 70868 30808 70877 30848
rect 70819 30807 70877 30808
rect 71499 30848 71541 30857
rect 76875 30850 76876 30890
rect 76916 30850 76917 30890
rect 71499 30808 71500 30848
rect 71540 30808 71541 30848
rect 71499 30799 71541 30808
rect 74851 30848 74909 30849
rect 74851 30808 74860 30848
rect 74900 30808 74909 30848
rect 74851 30807 74909 30808
rect 75427 30848 75485 30849
rect 75427 30808 75436 30848
rect 75476 30808 75485 30848
rect 76875 30841 76917 30850
rect 79459 30848 79517 30849
rect 75427 30807 75485 30808
rect 79459 30808 79468 30848
rect 79508 30808 79517 30848
rect 79459 30807 79517 30808
rect 43275 30764 43317 30773
rect 43275 30724 43276 30764
rect 43316 30724 43317 30764
rect 43275 30715 43317 30724
rect 55563 30764 55605 30773
rect 55563 30724 55564 30764
rect 55604 30724 55605 30764
rect 55563 30715 55605 30724
rect 56139 30764 56181 30773
rect 56139 30724 56140 30764
rect 56180 30724 56181 30764
rect 56139 30715 56181 30724
rect 68235 30764 68277 30773
rect 68235 30724 68236 30764
rect 68276 30724 68277 30764
rect 68235 30715 68277 30724
rect 71691 30764 71733 30773
rect 71691 30724 71692 30764
rect 71732 30724 71733 30764
rect 71691 30715 71733 30724
rect 43170 30701 43228 30702
rect 41451 30680 41493 30689
rect 41451 30640 41452 30680
rect 41492 30640 41493 30680
rect 41451 30631 41493 30640
rect 41643 30680 41685 30689
rect 41643 30640 41644 30680
rect 41684 30640 41685 30680
rect 41643 30631 41685 30640
rect 41731 30680 41789 30681
rect 41731 30640 41740 30680
rect 41780 30640 41789 30680
rect 41731 30639 41789 30640
rect 42699 30680 42741 30689
rect 42699 30640 42700 30680
rect 42740 30640 42741 30680
rect 42699 30631 42741 30640
rect 42891 30680 42933 30689
rect 42891 30640 42892 30680
rect 42932 30640 42933 30680
rect 42891 30631 42933 30640
rect 42979 30680 43037 30681
rect 42979 30640 42988 30680
rect 43028 30640 43037 30680
rect 43170 30661 43179 30701
rect 43219 30661 43228 30701
rect 51158 30701 51200 30710
rect 43170 30660 43228 30661
rect 43363 30680 43421 30681
rect 42979 30639 43037 30640
rect 43363 30640 43372 30680
rect 43412 30640 43421 30680
rect 43363 30639 43421 30640
rect 43755 30680 43797 30689
rect 43755 30640 43756 30680
rect 43796 30640 43797 30680
rect 43755 30631 43797 30640
rect 43947 30680 43989 30689
rect 43947 30640 43948 30680
rect 43988 30640 43989 30680
rect 43947 30631 43989 30640
rect 44035 30680 44093 30681
rect 44035 30640 44044 30680
rect 44084 30640 44093 30680
rect 44035 30639 44093 30640
rect 44619 30680 44661 30689
rect 44619 30640 44620 30680
rect 44660 30640 44661 30680
rect 44619 30631 44661 30640
rect 44715 30680 44757 30689
rect 44715 30640 44716 30680
rect 44756 30640 44757 30680
rect 44715 30631 44757 30640
rect 44811 30680 44853 30689
rect 44811 30640 44812 30680
rect 44852 30640 44853 30680
rect 44811 30631 44853 30640
rect 44907 30680 44949 30689
rect 44907 30640 44908 30680
rect 44948 30640 44949 30680
rect 44907 30631 44949 30640
rect 46059 30680 46101 30689
rect 46059 30640 46060 30680
rect 46100 30640 46101 30680
rect 46059 30631 46101 30640
rect 46251 30680 46293 30689
rect 46251 30640 46252 30680
rect 46292 30640 46293 30680
rect 46251 30631 46293 30640
rect 46339 30680 46397 30681
rect 46339 30640 46348 30680
rect 46388 30640 46397 30680
rect 46339 30639 46397 30640
rect 49611 30680 49653 30689
rect 49611 30640 49612 30680
rect 49652 30640 49653 30680
rect 49611 30631 49653 30640
rect 49707 30680 49749 30689
rect 49707 30640 49708 30680
rect 49748 30640 49749 30680
rect 49707 30631 49749 30640
rect 49803 30680 49845 30689
rect 49803 30640 49804 30680
rect 49844 30640 49845 30680
rect 49803 30631 49845 30640
rect 49899 30680 49941 30689
rect 49899 30640 49900 30680
rect 49940 30640 49941 30680
rect 49899 30631 49941 30640
rect 50563 30680 50621 30681
rect 50563 30640 50572 30680
rect 50612 30640 50621 30680
rect 50563 30639 50621 30640
rect 50763 30680 50805 30689
rect 50763 30640 50764 30680
rect 50804 30640 50805 30680
rect 50763 30631 50805 30640
rect 50955 30680 50997 30689
rect 50955 30640 50956 30680
rect 50996 30640 50997 30680
rect 51158 30661 51159 30701
rect 51199 30661 51200 30701
rect 65635 30701 65693 30702
rect 51158 30652 51200 30661
rect 54603 30680 54645 30689
rect 50955 30631 50997 30640
rect 54603 30640 54604 30680
rect 54644 30640 54645 30680
rect 54603 30631 54645 30640
rect 54795 30680 54837 30689
rect 54795 30640 54796 30680
rect 54836 30640 54837 30680
rect 54795 30631 54837 30640
rect 54883 30680 54941 30681
rect 54883 30640 54892 30680
rect 54932 30640 54941 30680
rect 54883 30639 54941 30640
rect 55171 30680 55229 30681
rect 55171 30640 55180 30680
rect 55220 30640 55229 30680
rect 55171 30639 55229 30640
rect 55467 30680 55509 30689
rect 55467 30640 55468 30680
rect 55508 30640 55509 30680
rect 56235 30680 56277 30689
rect 55467 30631 55509 30640
rect 56035 30657 56093 30658
rect 56035 30617 56044 30657
rect 56084 30617 56093 30657
rect 56235 30640 56236 30680
rect 56276 30640 56277 30680
rect 56235 30631 56277 30640
rect 59107 30680 59165 30681
rect 59107 30640 59116 30680
rect 59156 30640 59165 30680
rect 59107 30639 59165 30640
rect 59971 30680 60029 30681
rect 59971 30640 59980 30680
rect 60020 30640 60029 30680
rect 59971 30639 60029 30640
rect 60363 30680 60405 30689
rect 60363 30640 60364 30680
rect 60404 30640 60405 30680
rect 60363 30631 60405 30640
rect 60555 30680 60597 30689
rect 60555 30640 60556 30680
rect 60596 30640 60597 30680
rect 60555 30631 60597 30640
rect 60747 30680 60789 30689
rect 60747 30640 60748 30680
rect 60788 30640 60789 30680
rect 60747 30631 60789 30640
rect 60835 30680 60893 30681
rect 60835 30640 60844 30680
rect 60884 30640 60893 30680
rect 60835 30639 60893 30640
rect 61027 30680 61085 30681
rect 61027 30640 61036 30680
rect 61076 30640 61085 30680
rect 61027 30639 61085 30640
rect 61227 30680 61269 30689
rect 61227 30640 61228 30680
rect 61268 30640 61269 30680
rect 61227 30631 61269 30640
rect 63051 30680 63093 30689
rect 63051 30640 63052 30680
rect 63092 30640 63093 30680
rect 63051 30631 63093 30640
rect 63427 30680 63485 30681
rect 63427 30640 63436 30680
rect 63476 30640 63485 30680
rect 63427 30639 63485 30640
rect 64291 30680 64349 30681
rect 64291 30640 64300 30680
rect 64340 30640 64349 30680
rect 65635 30661 65644 30701
rect 65684 30661 65693 30701
rect 65635 30660 65693 30661
rect 65835 30680 65877 30689
rect 64291 30639 64349 30640
rect 65835 30640 65836 30680
rect 65876 30640 65877 30680
rect 65835 30631 65877 30640
rect 66019 30680 66077 30681
rect 66019 30640 66028 30680
rect 66068 30640 66077 30680
rect 66019 30639 66077 30640
rect 66219 30680 66261 30689
rect 66219 30640 66220 30680
rect 66260 30640 66261 30680
rect 66219 30631 66261 30640
rect 68611 30680 68669 30681
rect 68611 30640 68620 30680
rect 68660 30640 68669 30680
rect 68611 30639 68669 30640
rect 69475 30680 69533 30681
rect 69475 30640 69484 30680
rect 69524 30640 69533 30680
rect 69475 30639 69533 30640
rect 70923 30680 70965 30689
rect 70923 30640 70924 30680
rect 70964 30640 70965 30680
rect 70923 30631 70965 30640
rect 71019 30680 71061 30689
rect 71019 30640 71020 30680
rect 71060 30640 71061 30680
rect 71019 30631 71061 30640
rect 71115 30680 71157 30689
rect 71115 30640 71116 30680
rect 71156 30640 71157 30680
rect 71115 30631 71157 30640
rect 72067 30680 72125 30681
rect 72067 30640 72076 30680
rect 72116 30640 72125 30680
rect 72067 30639 72125 30640
rect 72931 30680 72989 30681
rect 72931 30640 72940 30680
rect 72980 30640 72989 30680
rect 72931 30639 72989 30640
rect 74955 30680 74997 30689
rect 74955 30640 74956 30680
rect 74996 30640 74997 30680
rect 74955 30631 74997 30640
rect 75051 30680 75093 30689
rect 75051 30640 75052 30680
rect 75092 30640 75093 30680
rect 75051 30631 75093 30640
rect 75147 30680 75189 30689
rect 75147 30640 75148 30680
rect 75188 30640 75189 30680
rect 75147 30631 75189 30640
rect 75339 30680 75381 30689
rect 75339 30640 75340 30680
rect 75380 30640 75381 30680
rect 75339 30631 75381 30640
rect 75531 30680 75573 30689
rect 75531 30640 75532 30680
rect 75572 30640 75573 30680
rect 75531 30631 75573 30640
rect 75619 30680 75677 30681
rect 75619 30640 75628 30680
rect 75668 30640 75677 30680
rect 75619 30639 75677 30640
rect 76195 30680 76253 30681
rect 76195 30640 76204 30680
rect 76244 30640 76253 30680
rect 76195 30639 76253 30640
rect 76491 30680 76533 30689
rect 76491 30640 76492 30680
rect 76532 30640 76533 30680
rect 76491 30631 76533 30640
rect 76587 30680 76629 30689
rect 76587 30640 76588 30680
rect 76628 30640 76629 30680
rect 76587 30631 76629 30640
rect 77067 30680 77109 30689
rect 77067 30640 77068 30680
rect 77108 30640 77109 30680
rect 77067 30631 77109 30640
rect 77443 30680 77501 30681
rect 77443 30640 77452 30680
rect 77492 30640 77501 30680
rect 77443 30639 77501 30640
rect 78307 30680 78365 30681
rect 78307 30640 78316 30680
rect 78356 30640 78365 30680
rect 78307 30639 78365 30640
rect 56035 30616 56093 30617
rect 40867 30596 40925 30597
rect 40867 30556 40876 30596
rect 40916 30556 40925 30596
rect 40867 30555 40925 30556
rect 42307 30596 42365 30597
rect 42307 30556 42316 30596
rect 42356 30556 42365 30596
rect 42307 30555 42365 30556
rect 49411 30596 49469 30597
rect 49411 30556 49420 30596
rect 49460 30556 49469 30596
rect 49411 30555 49469 30556
rect 50179 30596 50237 30597
rect 50179 30556 50188 30596
rect 50228 30556 50237 30596
rect 50179 30555 50237 30556
rect 51331 30596 51389 30597
rect 51331 30556 51340 30596
rect 51380 30556 51389 30596
rect 51331 30555 51389 30556
rect 71299 30596 71357 30597
rect 71299 30556 71308 30596
rect 71348 30556 71357 30596
rect 71299 30555 71357 30556
rect 43755 30512 43797 30521
rect 43755 30472 43756 30512
rect 43796 30472 43797 30512
rect 43755 30463 43797 30472
rect 44235 30512 44277 30521
rect 44235 30472 44236 30512
rect 44276 30472 44277 30512
rect 44235 30463 44277 30472
rect 46827 30512 46869 30521
rect 46827 30472 46828 30512
rect 46868 30472 46869 30512
rect 46827 30463 46869 30472
rect 48267 30512 48309 30521
rect 48267 30472 48268 30512
rect 48308 30472 48309 30512
rect 48267 30463 48309 30472
rect 51723 30512 51765 30521
rect 51723 30472 51724 30512
rect 51764 30472 51765 30512
rect 51723 30463 51765 30472
rect 53355 30512 53397 30521
rect 53355 30472 53356 30512
rect 53396 30472 53397 30512
rect 53355 30463 53397 30472
rect 54603 30512 54645 30521
rect 54603 30472 54604 30512
rect 54644 30472 54645 30512
rect 54603 30463 54645 30472
rect 55843 30512 55901 30513
rect 55843 30472 55852 30512
rect 55892 30472 55901 30512
rect 55843 30471 55901 30472
rect 56619 30512 56661 30521
rect 56619 30472 56620 30512
rect 56660 30472 56661 30512
rect 56619 30463 56661 30472
rect 60555 30512 60597 30521
rect 60555 30472 60556 30512
rect 60596 30472 60597 30512
rect 60555 30463 60597 30472
rect 61419 30512 61461 30521
rect 61419 30472 61420 30512
rect 61460 30472 61461 30512
rect 61419 30463 61461 30472
rect 66507 30512 66549 30521
rect 66507 30472 66508 30512
rect 66548 30472 66549 30512
rect 66507 30463 66549 30472
rect 40683 30428 40725 30437
rect 40683 30388 40684 30428
rect 40724 30388 40725 30428
rect 40683 30379 40725 30388
rect 41451 30428 41493 30437
rect 41451 30388 41452 30428
rect 41492 30388 41493 30428
rect 41451 30379 41493 30388
rect 42507 30428 42549 30437
rect 42507 30388 42508 30428
rect 42548 30388 42549 30428
rect 42507 30379 42549 30388
rect 46059 30428 46101 30437
rect 46059 30388 46060 30428
rect 46100 30388 46101 30428
rect 46059 30379 46101 30388
rect 50379 30428 50421 30437
rect 50379 30388 50380 30428
rect 50420 30388 50421 30428
rect 50379 30379 50421 30388
rect 50667 30428 50709 30437
rect 50667 30388 50668 30428
rect 50708 30388 50709 30428
rect 50667 30379 50709 30388
rect 51051 30428 51093 30437
rect 51051 30388 51052 30428
rect 51092 30388 51093 30428
rect 51051 30379 51093 30388
rect 61131 30428 61173 30437
rect 61131 30388 61132 30428
rect 61172 30388 61173 30428
rect 61131 30379 61173 30388
rect 65443 30428 65501 30429
rect 65443 30388 65452 30428
rect 65492 30388 65501 30428
rect 65443 30387 65501 30388
rect 65739 30428 65781 30437
rect 65739 30388 65740 30428
rect 65780 30388 65781 30428
rect 65739 30379 65781 30388
rect 66123 30428 66165 30437
rect 66123 30388 66124 30428
rect 66164 30388 66165 30428
rect 66123 30379 66165 30388
rect 70627 30428 70685 30429
rect 70627 30388 70636 30428
rect 70676 30388 70685 30428
rect 70627 30387 70685 30388
rect 71499 30428 71541 30437
rect 71499 30388 71500 30428
rect 71540 30388 71541 30428
rect 71499 30379 71541 30388
rect 74083 30428 74141 30429
rect 74083 30388 74092 30428
rect 74132 30388 74141 30428
rect 74083 30387 74141 30388
rect 576 30260 79584 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79584 30260
rect 576 30196 79584 30220
rect 40203 30092 40245 30101
rect 40203 30052 40204 30092
rect 40244 30052 40245 30092
rect 40203 30043 40245 30052
rect 45859 30092 45917 30093
rect 45859 30052 45868 30092
rect 45908 30052 45917 30092
rect 45859 30051 45917 30052
rect 47115 30092 47157 30101
rect 47115 30052 47116 30092
rect 47156 30052 47157 30092
rect 47115 30043 47157 30052
rect 50179 30092 50237 30093
rect 50179 30052 50188 30092
rect 50228 30052 50237 30092
rect 50179 30051 50237 30052
rect 54891 30092 54933 30101
rect 54891 30052 54892 30092
rect 54932 30052 54933 30092
rect 54891 30043 54933 30052
rect 62947 30092 63005 30093
rect 62947 30052 62956 30092
rect 62996 30052 63005 30092
rect 62947 30051 63005 30052
rect 63627 30092 63669 30101
rect 63627 30052 63628 30092
rect 63668 30052 63669 30092
rect 63627 30043 63669 30052
rect 65827 30092 65885 30093
rect 65827 30052 65836 30092
rect 65876 30052 65885 30092
rect 65827 30051 65885 30052
rect 69291 30092 69333 30101
rect 69291 30052 69292 30092
rect 69332 30052 69333 30092
rect 69291 30043 69333 30052
rect 70723 30092 70781 30093
rect 70723 30052 70732 30092
rect 70772 30052 70781 30092
rect 70723 30051 70781 30052
rect 71691 30092 71733 30101
rect 71691 30052 71692 30092
rect 71732 30052 71733 30092
rect 71691 30043 71733 30052
rect 72171 30092 72213 30101
rect 72171 30052 72172 30092
rect 72212 30052 72213 30092
rect 72171 30043 72213 30052
rect 75723 30092 75765 30101
rect 75723 30052 75724 30092
rect 75764 30052 75765 30092
rect 75723 30043 75765 30052
rect 77067 30092 77109 30101
rect 77067 30052 77068 30092
rect 77108 30052 77109 30092
rect 77067 30043 77109 30052
rect 38859 30008 38901 30017
rect 38859 29968 38860 30008
rect 38900 29968 38901 30008
rect 38859 29959 38901 29968
rect 40011 30008 40053 30017
rect 40011 29968 40012 30008
rect 40052 29968 40053 30008
rect 40011 29959 40053 29968
rect 46051 30008 46109 30009
rect 46051 29968 46060 30008
rect 46100 29968 46109 30008
rect 46051 29967 46109 29968
rect 54699 30008 54741 30017
rect 54699 29968 54700 30008
rect 54740 29968 54741 30008
rect 54699 29959 54741 29968
rect 55563 30008 55605 30017
rect 55563 29968 55564 30008
rect 55604 29968 55605 30008
rect 55563 29959 55605 29968
rect 58635 30008 58677 30017
rect 58635 29968 58636 30008
rect 58676 29968 58677 30008
rect 58635 29959 58677 29968
rect 58827 30008 58869 30017
rect 58827 29968 58828 30008
rect 58868 29968 58869 30008
rect 58827 29959 58869 29968
rect 60355 30008 60413 30009
rect 60355 29968 60364 30008
rect 60404 29968 60413 30008
rect 60355 29967 60413 29968
rect 73899 30008 73941 30017
rect 73899 29968 73900 30008
rect 73940 29968 73941 30008
rect 73899 29959 73941 29968
rect 77643 30008 77685 30017
rect 77643 29968 77644 30008
rect 77684 29968 77685 30008
rect 77643 29959 77685 29968
rect 39811 29924 39869 29925
rect 39811 29884 39820 29924
rect 39860 29884 39869 29924
rect 39811 29883 39869 29884
rect 40387 29924 40445 29925
rect 40387 29884 40396 29924
rect 40436 29884 40445 29924
rect 40387 29883 40445 29884
rect 50371 29924 50429 29925
rect 50371 29884 50380 29924
rect 50420 29884 50429 29924
rect 50371 29883 50429 29884
rect 54499 29924 54557 29925
rect 54499 29884 54508 29924
rect 54548 29884 54557 29924
rect 54499 29883 54557 29884
rect 59011 29924 59069 29925
rect 59011 29884 59020 29924
rect 59060 29884 59069 29924
rect 59011 29883 59069 29884
rect 59395 29924 59453 29925
rect 59395 29884 59404 29924
rect 59444 29884 59453 29924
rect 59395 29883 59453 29884
rect 69091 29924 69149 29925
rect 69091 29884 69100 29924
rect 69140 29884 69149 29924
rect 69091 29883 69149 29884
rect 71875 29924 71933 29925
rect 71875 29884 71884 29924
rect 71924 29884 71933 29924
rect 71875 29883 71933 29884
rect 75043 29924 75101 29925
rect 75043 29884 75052 29924
rect 75092 29884 75101 29924
rect 75043 29883 75101 29884
rect 40587 29840 40629 29849
rect 40587 29800 40588 29840
rect 40628 29800 40629 29840
rect 40587 29791 40629 29800
rect 40683 29840 40725 29849
rect 40683 29800 40684 29840
rect 40724 29800 40725 29840
rect 40683 29791 40725 29800
rect 40779 29840 40821 29849
rect 40779 29800 40780 29840
rect 40820 29800 40821 29840
rect 40779 29791 40821 29800
rect 41347 29840 41405 29841
rect 41347 29800 41356 29840
rect 41396 29800 41405 29840
rect 41347 29799 41405 29800
rect 41547 29840 41589 29849
rect 41547 29800 41548 29840
rect 41588 29800 41589 29840
rect 41547 29791 41589 29800
rect 43843 29840 43901 29841
rect 43843 29800 43852 29840
rect 43892 29800 43901 29840
rect 43843 29799 43901 29800
rect 44707 29840 44765 29841
rect 44707 29800 44716 29840
rect 44756 29800 44765 29840
rect 44707 29799 44765 29800
rect 46347 29840 46389 29849
rect 46347 29800 46348 29840
rect 46388 29800 46389 29840
rect 46347 29791 46389 29800
rect 46443 29840 46485 29849
rect 46443 29800 46444 29840
rect 46484 29800 46485 29840
rect 46443 29791 46485 29800
rect 46723 29840 46781 29841
rect 46723 29800 46732 29840
rect 46772 29800 46781 29840
rect 46723 29799 46781 29800
rect 47011 29840 47069 29841
rect 47011 29800 47020 29840
rect 47060 29800 47069 29840
rect 48163 29840 48221 29841
rect 47011 29799 47069 29800
rect 47211 29827 47253 29836
rect 47211 29787 47212 29827
rect 47252 29787 47253 29827
rect 48163 29800 48172 29840
rect 48212 29800 48221 29840
rect 48163 29799 48221 29800
rect 49027 29840 49085 29841
rect 49027 29800 49036 29840
rect 49076 29800 49085 29840
rect 49027 29799 49085 29800
rect 50755 29840 50813 29841
rect 50755 29800 50764 29840
rect 50804 29800 50813 29840
rect 51051 29840 51093 29849
rect 50755 29799 50813 29800
rect 47211 29778 47253 29787
rect 50859 29798 50901 29807
rect 41451 29756 41493 29765
rect 41451 29716 41452 29756
rect 41492 29716 41493 29756
rect 41451 29707 41493 29716
rect 43467 29756 43509 29765
rect 43467 29716 43468 29756
rect 43508 29716 43509 29756
rect 43467 29707 43509 29716
rect 47787 29756 47829 29765
rect 47787 29716 47788 29756
rect 47828 29716 47829 29756
rect 50859 29758 50860 29798
rect 50900 29758 50901 29798
rect 51051 29800 51052 29840
rect 51092 29800 51093 29840
rect 51051 29791 51093 29800
rect 51619 29840 51677 29841
rect 51619 29800 51628 29840
rect 51668 29800 51677 29840
rect 51619 29799 51677 29800
rect 52483 29840 52541 29841
rect 52483 29800 52492 29840
rect 52532 29800 52541 29840
rect 52483 29799 52541 29800
rect 54891 29840 54933 29849
rect 54891 29800 54892 29840
rect 54932 29800 54933 29840
rect 54891 29791 54933 29800
rect 55083 29840 55125 29849
rect 55083 29800 55084 29840
rect 55124 29800 55125 29840
rect 55083 29791 55125 29800
rect 55171 29840 55229 29841
rect 55171 29800 55180 29840
rect 55220 29800 55229 29840
rect 55171 29799 55229 29800
rect 55467 29840 55509 29849
rect 55467 29800 55468 29840
rect 55508 29800 55509 29840
rect 55467 29791 55509 29800
rect 55651 29840 55709 29841
rect 55651 29800 55660 29840
rect 55700 29800 55709 29840
rect 55651 29799 55709 29800
rect 55851 29840 55893 29849
rect 55851 29800 55852 29840
rect 55892 29800 55893 29840
rect 55851 29791 55893 29800
rect 56043 29840 56085 29849
rect 56043 29800 56044 29840
rect 56084 29800 56085 29840
rect 56043 29791 56085 29800
rect 56131 29840 56189 29841
rect 56131 29800 56140 29840
rect 56180 29800 56189 29840
rect 56131 29799 56189 29800
rect 59683 29840 59741 29841
rect 59683 29800 59692 29840
rect 59732 29800 59741 29840
rect 59683 29799 59741 29800
rect 59979 29840 60021 29849
rect 59979 29800 59980 29840
rect 60020 29800 60021 29840
rect 59979 29791 60021 29800
rect 60075 29840 60117 29849
rect 60075 29800 60076 29840
rect 60116 29800 60117 29840
rect 60075 29791 60117 29800
rect 60931 29840 60989 29841
rect 60931 29800 60940 29840
rect 60980 29800 60989 29840
rect 60931 29799 60989 29800
rect 61795 29840 61853 29841
rect 61795 29800 61804 29840
rect 61844 29800 61853 29840
rect 61795 29799 61853 29800
rect 63243 29840 63285 29849
rect 63243 29800 63244 29840
rect 63284 29800 63285 29840
rect 63435 29840 63477 29849
rect 63243 29791 63285 29800
rect 63339 29819 63381 29828
rect 63339 29779 63340 29819
rect 63380 29779 63381 29819
rect 63435 29800 63436 29840
rect 63476 29800 63477 29840
rect 63435 29791 63477 29800
rect 63627 29840 63669 29849
rect 63627 29800 63628 29840
rect 63668 29800 63669 29840
rect 63627 29791 63669 29800
rect 63819 29840 63861 29849
rect 63819 29800 63820 29840
rect 63860 29800 63861 29840
rect 63819 29791 63861 29800
rect 63907 29840 63965 29841
rect 63907 29800 63916 29840
rect 63956 29800 63965 29840
rect 63907 29799 63965 29800
rect 65155 29840 65213 29841
rect 65155 29800 65164 29840
rect 65204 29800 65213 29840
rect 65155 29799 65213 29800
rect 65451 29840 65493 29849
rect 65451 29800 65452 29840
rect 65492 29800 65493 29840
rect 65451 29791 65493 29800
rect 65547 29840 65589 29849
rect 65547 29800 65548 29840
rect 65588 29800 65589 29840
rect 65547 29791 65589 29800
rect 66403 29840 66461 29841
rect 66403 29800 66412 29840
rect 66452 29800 66461 29840
rect 66403 29799 66461 29800
rect 67267 29840 67325 29841
rect 67267 29800 67276 29840
rect 67316 29800 67325 29840
rect 67267 29799 67325 29800
rect 69483 29840 69525 29849
rect 69483 29800 69484 29840
rect 69524 29800 69525 29840
rect 69483 29791 69525 29800
rect 69675 29840 69717 29849
rect 69675 29800 69676 29840
rect 69716 29800 69717 29840
rect 69675 29791 69717 29800
rect 69763 29840 69821 29841
rect 69763 29800 69772 29840
rect 69812 29800 69821 29840
rect 69763 29799 69821 29800
rect 69955 29840 70013 29841
rect 69955 29800 69964 29840
rect 70004 29800 70013 29840
rect 69955 29799 70013 29800
rect 70059 29840 70101 29849
rect 70059 29800 70060 29840
rect 70100 29800 70101 29840
rect 70059 29791 70101 29800
rect 70251 29840 70293 29849
rect 70251 29800 70252 29840
rect 70292 29800 70293 29840
rect 70251 29791 70293 29800
rect 71019 29840 71061 29849
rect 71019 29800 71020 29840
rect 71060 29800 71061 29840
rect 71019 29791 71061 29800
rect 71115 29840 71157 29849
rect 71115 29800 71116 29840
rect 71156 29800 71157 29840
rect 71115 29791 71157 29800
rect 71395 29840 71453 29841
rect 71395 29800 71404 29840
rect 71444 29800 71453 29840
rect 71395 29799 71453 29800
rect 72067 29840 72125 29841
rect 72067 29800 72076 29840
rect 72116 29800 72125 29840
rect 72067 29799 72125 29800
rect 72267 29840 72309 29849
rect 72267 29800 72268 29840
rect 72308 29800 72309 29840
rect 72267 29791 72309 29800
rect 75339 29840 75381 29849
rect 75339 29800 75340 29840
rect 75380 29800 75381 29840
rect 75339 29791 75381 29800
rect 75435 29840 75477 29849
rect 75435 29800 75436 29840
rect 75476 29800 75477 29840
rect 75435 29791 75477 29800
rect 75531 29840 75573 29849
rect 75531 29800 75532 29840
rect 75572 29800 75573 29840
rect 75531 29791 75573 29800
rect 75723 29840 75765 29849
rect 75723 29800 75724 29840
rect 75764 29800 75765 29840
rect 75723 29791 75765 29800
rect 75915 29840 75957 29849
rect 75915 29800 75916 29840
rect 75956 29800 75957 29840
rect 75915 29791 75957 29800
rect 76003 29840 76061 29841
rect 76003 29800 76012 29840
rect 76052 29800 76061 29840
rect 76003 29799 76061 29800
rect 76483 29840 76541 29841
rect 76483 29800 76492 29840
rect 76532 29800 76541 29840
rect 76483 29799 76541 29800
rect 76683 29840 76725 29849
rect 76683 29800 76684 29840
rect 76724 29800 76725 29840
rect 76683 29791 76725 29800
rect 77067 29840 77109 29849
rect 77067 29800 77068 29840
rect 77108 29800 77109 29840
rect 77067 29791 77109 29800
rect 77259 29840 77301 29849
rect 77259 29800 77260 29840
rect 77300 29800 77301 29840
rect 77259 29791 77301 29800
rect 77347 29840 77405 29841
rect 77347 29800 77356 29840
rect 77396 29800 77405 29840
rect 77347 29799 77405 29800
rect 63339 29770 63381 29779
rect 50859 29749 50901 29758
rect 51243 29756 51285 29765
rect 47787 29707 47829 29716
rect 51243 29716 51244 29756
rect 51284 29716 51285 29756
rect 51243 29707 51285 29716
rect 60555 29756 60597 29765
rect 60555 29716 60556 29756
rect 60596 29716 60597 29756
rect 60555 29707 60597 29716
rect 63147 29756 63189 29765
rect 63147 29716 63148 29756
rect 63188 29716 63189 29756
rect 63147 29707 63189 29716
rect 66027 29756 66069 29765
rect 66027 29716 66028 29756
rect 66068 29716 66069 29756
rect 66027 29707 66069 29716
rect 69579 29756 69621 29765
rect 69579 29716 69580 29756
rect 69620 29716 69621 29756
rect 69579 29707 69621 29716
rect 76587 29756 76629 29765
rect 76587 29716 76588 29756
rect 76628 29716 76629 29756
rect 76587 29707 76629 29716
rect 40867 29672 40925 29673
rect 40867 29632 40876 29672
rect 40916 29632 40925 29672
rect 40867 29631 40925 29632
rect 50179 29672 50237 29673
rect 50179 29632 50188 29672
rect 50228 29632 50237 29672
rect 50179 29631 50237 29632
rect 50571 29672 50613 29681
rect 50571 29632 50572 29672
rect 50612 29632 50613 29672
rect 50571 29623 50613 29632
rect 50947 29672 51005 29673
rect 50947 29632 50956 29672
rect 50996 29632 51005 29672
rect 50947 29631 51005 29632
rect 53635 29672 53693 29673
rect 53635 29632 53644 29672
rect 53684 29632 53693 29672
rect 53635 29631 53693 29632
rect 55939 29672 55997 29673
rect 55939 29632 55948 29672
rect 55988 29632 55997 29672
rect 55939 29631 55997 29632
rect 59211 29672 59253 29681
rect 59211 29632 59212 29672
rect 59252 29632 59253 29672
rect 59211 29623 59253 29632
rect 62947 29672 63005 29673
rect 62947 29632 62956 29672
rect 62996 29632 63005 29672
rect 62947 29631 63005 29632
rect 68419 29672 68477 29673
rect 68419 29632 68428 29672
rect 68468 29632 68477 29672
rect 68419 29631 68477 29632
rect 70147 29672 70205 29673
rect 70147 29632 70156 29672
rect 70196 29632 70205 29672
rect 70147 29631 70205 29632
rect 74859 29672 74901 29681
rect 74859 29632 74860 29672
rect 74900 29632 74901 29672
rect 74859 29623 74901 29632
rect 75235 29672 75293 29673
rect 75235 29632 75244 29672
rect 75284 29632 75293 29672
rect 75235 29631 75293 29632
rect 576 29504 79584 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79584 29504
rect 576 29440 79584 29464
rect 44995 29336 45053 29337
rect 44995 29296 45004 29336
rect 45044 29296 45053 29336
rect 44995 29295 45053 29296
rect 55363 29336 55421 29337
rect 55363 29296 55372 29336
rect 55412 29296 55421 29336
rect 55363 29295 55421 29296
rect 59307 29336 59349 29345
rect 59307 29296 59308 29336
rect 59348 29296 59349 29336
rect 59307 29287 59349 29296
rect 60451 29336 60509 29337
rect 60451 29296 60460 29336
rect 60500 29296 60509 29336
rect 60451 29295 60509 29296
rect 61131 29336 61173 29345
rect 61131 29296 61132 29336
rect 61172 29296 61173 29336
rect 61131 29287 61173 29296
rect 63427 29336 63485 29337
rect 63427 29296 63436 29336
rect 63476 29296 63485 29336
rect 63427 29295 63485 29296
rect 70339 29336 70397 29337
rect 70339 29296 70348 29336
rect 70388 29296 70397 29336
rect 70339 29295 70397 29296
rect 70827 29336 70869 29345
rect 70827 29296 70828 29336
rect 70868 29296 70869 29336
rect 70827 29287 70869 29296
rect 71691 29336 71733 29345
rect 71691 29296 71692 29336
rect 71732 29296 71733 29336
rect 71691 29287 71733 29296
rect 75811 29336 75869 29337
rect 75811 29296 75820 29336
rect 75860 29296 75869 29336
rect 75811 29295 75869 29296
rect 46059 29252 46101 29261
rect 46059 29212 46060 29252
rect 46100 29212 46101 29252
rect 46059 29203 46101 29212
rect 46347 29252 46389 29261
rect 46347 29212 46348 29252
rect 46388 29212 46389 29252
rect 46347 29203 46389 29212
rect 50475 29252 50517 29261
rect 50475 29212 50476 29252
rect 50516 29212 50517 29252
rect 50475 29203 50517 29212
rect 56331 29252 56373 29261
rect 56331 29212 56332 29252
rect 56372 29212 56373 29252
rect 56331 29203 56373 29212
rect 60843 29252 60885 29261
rect 60843 29212 60844 29252
rect 60884 29212 60885 29252
rect 60843 29203 60885 29212
rect 65739 29252 65781 29261
rect 65739 29212 65740 29252
rect 65780 29212 65781 29252
rect 65739 29203 65781 29212
rect 67755 29252 67797 29261
rect 67755 29212 67756 29252
rect 67796 29212 67797 29252
rect 67755 29203 67797 29212
rect 76491 29252 76533 29261
rect 76491 29212 76492 29252
rect 76532 29212 76533 29252
rect 76491 29203 76533 29212
rect 38379 29168 38421 29177
rect 38379 29128 38380 29168
rect 38420 29128 38421 29168
rect 38379 29119 38421 29128
rect 38755 29168 38813 29169
rect 38755 29128 38764 29168
rect 38804 29128 38813 29168
rect 38755 29127 38813 29128
rect 39619 29168 39677 29169
rect 39619 29128 39628 29168
rect 39668 29128 39677 29168
rect 39619 29127 39677 29128
rect 41059 29168 41117 29169
rect 41059 29128 41068 29168
rect 41108 29128 41117 29168
rect 41059 29127 41117 29128
rect 41355 29168 41397 29177
rect 41355 29128 41356 29168
rect 41396 29128 41397 29168
rect 41355 29119 41397 29128
rect 41451 29168 41493 29177
rect 41451 29128 41452 29168
rect 41492 29128 41493 29168
rect 41451 29119 41493 29128
rect 41923 29168 41981 29169
rect 41923 29128 41932 29168
rect 41972 29128 41981 29168
rect 41923 29127 41981 29128
rect 42027 29168 42069 29177
rect 42027 29128 42028 29168
rect 42068 29128 42069 29168
rect 42027 29119 42069 29128
rect 42219 29168 42261 29177
rect 42219 29128 42220 29168
rect 42260 29128 42261 29168
rect 42219 29119 42261 29128
rect 44907 29168 44949 29177
rect 44907 29128 44908 29168
rect 44948 29128 44949 29168
rect 44907 29119 44949 29128
rect 45099 29168 45141 29177
rect 45099 29128 45100 29168
rect 45140 29128 45141 29168
rect 45099 29119 45141 29128
rect 45187 29168 45245 29169
rect 45187 29128 45196 29168
rect 45236 29128 45245 29168
rect 45187 29127 45245 29128
rect 45963 29168 46005 29177
rect 45963 29128 45964 29168
rect 46004 29128 46005 29168
rect 45963 29119 46005 29128
rect 46147 29168 46205 29169
rect 46147 29128 46156 29168
rect 46196 29128 46205 29168
rect 46147 29127 46205 29128
rect 46723 29168 46781 29169
rect 46723 29128 46732 29168
rect 46772 29128 46781 29168
rect 46723 29127 46781 29128
rect 47587 29168 47645 29169
rect 47587 29128 47596 29168
rect 47636 29128 47645 29168
rect 47587 29127 47645 29128
rect 49515 29168 49557 29177
rect 49515 29128 49516 29168
rect 49556 29128 49557 29168
rect 49515 29119 49557 29128
rect 49707 29168 49749 29177
rect 49707 29128 49708 29168
rect 49748 29128 49749 29168
rect 49707 29119 49749 29128
rect 49795 29168 49853 29169
rect 49795 29128 49804 29168
rect 49844 29128 49853 29168
rect 49795 29127 49853 29128
rect 50083 29168 50141 29169
rect 50083 29128 50092 29168
rect 50132 29128 50141 29168
rect 50083 29127 50141 29128
rect 50379 29168 50421 29177
rect 50379 29128 50380 29168
rect 50420 29128 50421 29168
rect 50379 29119 50421 29128
rect 51811 29168 51869 29169
rect 51811 29128 51820 29168
rect 51860 29128 51869 29168
rect 51811 29127 51869 29128
rect 52971 29168 53013 29177
rect 52971 29128 52972 29168
rect 53012 29128 53013 29168
rect 52971 29119 53013 29128
rect 53347 29168 53405 29169
rect 53347 29128 53356 29168
rect 53396 29128 53405 29168
rect 53347 29127 53405 29128
rect 54211 29168 54269 29169
rect 54211 29128 54220 29168
rect 54260 29128 54269 29168
rect 54211 29127 54269 29128
rect 55563 29168 55605 29177
rect 55563 29128 55564 29168
rect 55604 29128 55605 29168
rect 55563 29119 55605 29128
rect 55659 29168 55701 29177
rect 55659 29128 55660 29168
rect 55700 29128 55701 29168
rect 55659 29119 55701 29128
rect 55755 29168 55797 29177
rect 55755 29128 55756 29168
rect 55796 29128 55797 29168
rect 55755 29119 55797 29128
rect 55851 29168 55893 29177
rect 55851 29128 55852 29168
rect 55892 29128 55893 29168
rect 55851 29119 55893 29128
rect 56707 29168 56765 29169
rect 56707 29128 56716 29168
rect 56756 29128 56765 29168
rect 56707 29127 56765 29128
rect 57571 29168 57629 29169
rect 57571 29128 57580 29168
rect 57620 29128 57629 29168
rect 57571 29127 57629 29128
rect 59499 29168 59541 29177
rect 59499 29128 59500 29168
rect 59540 29128 59541 29168
rect 59499 29119 59541 29128
rect 59691 29168 59733 29177
rect 59691 29128 59692 29168
rect 59732 29128 59733 29168
rect 59691 29119 59733 29128
rect 59779 29168 59837 29169
rect 59779 29128 59788 29168
rect 59828 29128 59837 29168
rect 59779 29127 59837 29128
rect 60259 29168 60317 29169
rect 60259 29128 60268 29168
rect 60308 29128 60317 29168
rect 60259 29127 60317 29128
rect 60363 29168 60405 29177
rect 60363 29128 60364 29168
rect 60404 29128 60405 29168
rect 60363 29119 60405 29128
rect 60555 29168 60597 29177
rect 60555 29128 60556 29168
rect 60596 29128 60597 29168
rect 60555 29119 60597 29128
rect 60747 29168 60789 29177
rect 60747 29128 60748 29168
rect 60788 29128 60789 29168
rect 60747 29119 60789 29128
rect 60931 29168 60989 29169
rect 60931 29128 60940 29168
rect 60980 29128 60989 29168
rect 63531 29168 63573 29177
rect 60931 29127 60989 29128
rect 63339 29157 63381 29166
rect 63339 29117 63340 29157
rect 63380 29117 63381 29157
rect 63531 29128 63532 29168
rect 63572 29128 63573 29168
rect 63531 29119 63573 29128
rect 63619 29168 63677 29169
rect 63619 29128 63628 29168
rect 63668 29128 63677 29168
rect 63619 29127 63677 29128
rect 63819 29168 63861 29177
rect 63819 29128 63820 29168
rect 63860 29128 63861 29168
rect 63819 29119 63861 29128
rect 63915 29168 63957 29177
rect 63915 29128 63916 29168
rect 63956 29128 63957 29168
rect 63915 29119 63957 29128
rect 64011 29168 64053 29177
rect 64011 29128 64012 29168
rect 64052 29128 64053 29168
rect 64011 29119 64053 29128
rect 64107 29168 64149 29177
rect 64107 29128 64108 29168
rect 64148 29128 64149 29168
rect 64107 29119 64149 29128
rect 64963 29168 65021 29169
rect 64963 29128 64972 29168
rect 65012 29128 65021 29168
rect 64963 29127 65021 29128
rect 65163 29168 65205 29177
rect 65163 29128 65164 29168
rect 65204 29128 65205 29168
rect 65163 29119 65205 29128
rect 65643 29168 65685 29177
rect 65643 29128 65644 29168
rect 65684 29128 65685 29168
rect 65643 29119 65685 29128
rect 65835 29168 65877 29177
rect 65835 29128 65836 29168
rect 65876 29128 65877 29168
rect 65835 29119 65877 29128
rect 65923 29168 65981 29169
rect 65923 29128 65932 29168
rect 65972 29128 65981 29168
rect 65923 29127 65981 29128
rect 68131 29168 68189 29169
rect 68131 29128 68140 29168
rect 68180 29128 68189 29168
rect 68131 29127 68189 29128
rect 68995 29168 69053 29169
rect 68995 29128 69004 29168
rect 69044 29128 69053 29168
rect 68995 29127 69053 29128
rect 70443 29168 70485 29177
rect 70443 29128 70444 29168
rect 70484 29128 70485 29168
rect 70443 29119 70485 29128
rect 70539 29168 70581 29177
rect 70539 29128 70540 29168
rect 70580 29128 70581 29168
rect 70539 29119 70581 29128
rect 70635 29168 70677 29177
rect 70635 29128 70636 29168
rect 70676 29128 70677 29168
rect 70635 29119 70677 29128
rect 71299 29168 71357 29169
rect 71299 29128 71308 29168
rect 71348 29128 71357 29168
rect 71299 29127 71357 29128
rect 71499 29168 71541 29177
rect 71499 29128 71500 29168
rect 71540 29128 71541 29168
rect 73795 29168 73853 29169
rect 71499 29119 71541 29128
rect 73419 29126 73461 29135
rect 73795 29128 73804 29168
rect 73844 29128 73853 29168
rect 73795 29127 73853 29128
rect 74659 29168 74717 29169
rect 74659 29128 74668 29168
rect 74708 29128 74717 29168
rect 74659 29127 74717 29128
rect 76099 29168 76157 29169
rect 76099 29128 76108 29168
rect 76148 29128 76157 29168
rect 76099 29127 76157 29128
rect 76395 29168 76437 29177
rect 76395 29128 76396 29168
rect 76436 29128 76437 29168
rect 63339 29108 63381 29117
rect 51139 29084 51197 29085
rect 51139 29044 51148 29084
rect 51188 29044 51197 29084
rect 51139 29043 51197 29044
rect 51523 29084 51581 29085
rect 51523 29044 51532 29084
rect 51572 29044 51581 29084
rect 51523 29043 51581 29044
rect 59107 29084 59165 29085
rect 59107 29044 59116 29084
rect 59156 29044 59165 29084
rect 59107 29043 59165 29044
rect 61315 29084 61373 29085
rect 61315 29044 61324 29084
rect 61364 29044 61373 29084
rect 61315 29043 61373 29044
rect 70155 29084 70197 29093
rect 73419 29086 73420 29126
rect 73460 29086 73461 29126
rect 76395 29119 76437 29128
rect 77067 29168 77109 29177
rect 77067 29128 77068 29168
rect 77108 29128 77109 29168
rect 77067 29119 77109 29128
rect 77443 29168 77501 29169
rect 77443 29128 77452 29168
rect 77492 29128 77501 29168
rect 77443 29127 77501 29128
rect 78307 29168 78365 29169
rect 78307 29128 78316 29168
rect 78356 29128 78365 29168
rect 78307 29127 78365 29128
rect 70155 29044 70156 29084
rect 70196 29044 70197 29084
rect 70155 29035 70197 29044
rect 71011 29084 71069 29085
rect 71011 29044 71020 29084
rect 71060 29044 71069 29084
rect 71011 29043 71069 29044
rect 71875 29084 71933 29085
rect 71875 29044 71884 29084
rect 71924 29044 71933 29084
rect 73419 29077 73461 29086
rect 71875 29043 71933 29044
rect 41731 29000 41789 29001
rect 41731 28960 41740 29000
rect 41780 28960 41789 29000
rect 41731 28959 41789 28960
rect 42411 29000 42453 29009
rect 42411 28960 42412 29000
rect 42452 28960 42453 29000
rect 42411 28951 42453 28960
rect 49515 29000 49557 29009
rect 49515 28960 49516 29000
rect 49556 28960 49557 29000
rect 49515 28951 49557 28960
rect 50755 29000 50813 29001
rect 50755 28960 50764 29000
rect 50804 28960 50813 29000
rect 50755 28959 50813 28960
rect 62379 29000 62421 29009
rect 62379 28960 62380 29000
rect 62420 28960 62421 29000
rect 62379 28951 62421 28960
rect 76771 29000 76829 29001
rect 76771 28960 76780 29000
rect 76820 28960 76829 29000
rect 76771 28959 76829 28960
rect 40771 28916 40829 28917
rect 40771 28876 40780 28916
rect 40820 28876 40829 28916
rect 40771 28875 40829 28876
rect 42219 28916 42261 28925
rect 42219 28876 42220 28916
rect 42260 28876 42261 28916
rect 42219 28867 42261 28876
rect 48739 28916 48797 28917
rect 48739 28876 48748 28916
rect 48788 28876 48797 28916
rect 48739 28875 48797 28876
rect 50955 28916 50997 28925
rect 50955 28876 50956 28916
rect 50996 28876 50997 28916
rect 50955 28867 50997 28876
rect 51339 28916 51381 28925
rect 51339 28876 51340 28916
rect 51380 28876 51381 28916
rect 51339 28867 51381 28876
rect 58723 28916 58781 28917
rect 58723 28876 58732 28916
rect 58772 28876 58781 28916
rect 58723 28875 58781 28876
rect 59499 28916 59541 28925
rect 59499 28876 59500 28916
rect 59540 28876 59541 28916
rect 59499 28867 59541 28876
rect 65067 28916 65109 28925
rect 65067 28876 65068 28916
rect 65108 28876 65109 28916
rect 65067 28867 65109 28876
rect 70827 28916 70869 28925
rect 70827 28876 70828 28916
rect 70868 28876 70869 28916
rect 70827 28867 70869 28876
rect 71403 28916 71445 28925
rect 71403 28876 71404 28916
rect 71444 28876 71445 28916
rect 71403 28867 71445 28876
rect 71691 28916 71733 28925
rect 71691 28876 71692 28916
rect 71732 28876 71733 28916
rect 71691 28867 71733 28876
rect 79459 28916 79517 28917
rect 79459 28876 79468 28916
rect 79508 28876 79517 28916
rect 79459 28875 79517 28876
rect 576 28748 79584 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79584 28748
rect 576 28684 79584 28708
rect 39627 28580 39669 28589
rect 39627 28540 39628 28580
rect 39668 28540 39669 28580
rect 39627 28531 39669 28540
rect 41451 28580 41493 28589
rect 41451 28540 41452 28580
rect 41492 28540 41493 28580
rect 41451 28531 41493 28540
rect 45291 28580 45333 28589
rect 45291 28540 45292 28580
rect 45332 28540 45333 28580
rect 45291 28531 45333 28540
rect 51243 28580 51285 28589
rect 51243 28540 51244 28580
rect 51284 28540 51285 28580
rect 51243 28531 51285 28540
rect 55267 28580 55325 28581
rect 55267 28540 55276 28580
rect 55316 28540 55325 28580
rect 55267 28539 55325 28540
rect 59019 28580 59061 28589
rect 59019 28540 59020 28580
rect 59060 28540 59061 28580
rect 59019 28531 59061 28540
rect 65251 28580 65309 28581
rect 65251 28540 65260 28580
rect 65300 28540 65309 28580
rect 65251 28539 65309 28540
rect 73795 28580 73853 28581
rect 73795 28540 73804 28580
rect 73844 28540 73853 28580
rect 73795 28539 73853 28540
rect 76683 28580 76725 28589
rect 76683 28540 76684 28580
rect 76724 28540 76725 28580
rect 76683 28531 76725 28540
rect 38187 28496 38229 28505
rect 38187 28456 38188 28496
rect 38228 28456 38229 28496
rect 38187 28447 38229 28456
rect 44331 28496 44373 28505
rect 44331 28456 44332 28496
rect 44372 28456 44373 28496
rect 44331 28447 44373 28456
rect 47499 28496 47541 28505
rect 47499 28456 47500 28496
rect 47540 28456 47541 28496
rect 47499 28447 47541 28456
rect 49227 28496 49269 28505
rect 49227 28456 49228 28496
rect 49268 28456 49269 28496
rect 49227 28447 49269 28456
rect 52491 28496 52533 28505
rect 52491 28456 52492 28496
rect 52532 28456 52533 28496
rect 52491 28447 52533 28456
rect 56811 28496 56853 28505
rect 56811 28456 56812 28496
rect 56852 28456 56853 28496
rect 56811 28447 56853 28456
rect 58635 28496 58677 28505
rect 58635 28456 58636 28496
rect 58676 28456 58677 28496
rect 58635 28447 58677 28456
rect 59787 28496 59829 28505
rect 59787 28456 59788 28496
rect 59828 28456 59829 28496
rect 59787 28447 59829 28456
rect 68331 28496 68373 28505
rect 68331 28456 68332 28496
rect 68372 28456 68373 28496
rect 68331 28447 68373 28456
rect 71011 28496 71069 28497
rect 71011 28456 71020 28496
rect 71060 28456 71069 28496
rect 71011 28455 71069 28456
rect 77547 28496 77589 28505
rect 77547 28456 77548 28496
rect 77588 28456 77589 28496
rect 77547 28447 77589 28456
rect 39427 28412 39485 28413
rect 39427 28372 39436 28412
rect 39476 28372 39485 28412
rect 39427 28371 39485 28372
rect 40003 28412 40061 28413
rect 40003 28372 40012 28412
rect 40052 28372 40061 28412
rect 40003 28371 40061 28372
rect 51043 28412 51101 28413
rect 51043 28372 51052 28412
rect 51092 28372 51101 28412
rect 51043 28371 51101 28372
rect 54403 28412 54461 28413
rect 54403 28372 54412 28412
rect 54452 28372 54461 28412
rect 54403 28371 54461 28372
rect 58435 28412 58493 28413
rect 58435 28372 58444 28412
rect 58484 28372 58493 28412
rect 58435 28371 58493 28372
rect 58819 28412 58877 28413
rect 58819 28372 58828 28412
rect 58868 28372 58877 28412
rect 58819 28371 58877 28372
rect 60931 28412 60989 28413
rect 60931 28372 60940 28412
rect 60980 28372 60989 28412
rect 60931 28371 60989 28372
rect 70051 28412 70109 28413
rect 70051 28372 70060 28412
rect 70100 28372 70109 28412
rect 70051 28371 70109 28372
rect 40203 28328 40245 28337
rect 40203 28288 40204 28328
rect 40244 28288 40245 28328
rect 40203 28279 40245 28288
rect 40395 28328 40437 28337
rect 40395 28288 40396 28328
rect 40436 28288 40437 28328
rect 40395 28279 40437 28288
rect 40483 28328 40541 28329
rect 40483 28288 40492 28328
rect 40532 28288 40541 28328
rect 40483 28287 40541 28288
rect 40875 28328 40917 28337
rect 40875 28288 40876 28328
rect 40916 28288 40917 28328
rect 40875 28279 40917 28288
rect 41067 28328 41109 28337
rect 41067 28288 41068 28328
rect 41108 28288 41109 28328
rect 41067 28279 41109 28288
rect 41155 28328 41213 28329
rect 41155 28288 41164 28328
rect 41204 28288 41213 28328
rect 41155 28287 41213 28288
rect 41355 28328 41397 28337
rect 41355 28288 41356 28328
rect 41396 28288 41397 28328
rect 41355 28279 41397 28288
rect 41539 28328 41597 28329
rect 41539 28288 41548 28328
rect 41588 28288 41597 28328
rect 41539 28287 41597 28288
rect 41739 28328 41781 28337
rect 41739 28288 41740 28328
rect 41780 28288 41781 28328
rect 41739 28279 41781 28288
rect 42115 28328 42173 28329
rect 42115 28288 42124 28328
rect 42164 28288 42173 28328
rect 42115 28287 42173 28288
rect 42979 28328 43037 28329
rect 42979 28288 42988 28328
rect 43028 28288 43037 28328
rect 42979 28287 43037 28288
rect 44995 28328 45053 28329
rect 44995 28288 45004 28328
rect 45044 28288 45053 28328
rect 44995 28287 45053 28288
rect 45099 28328 45141 28337
rect 45099 28288 45100 28328
rect 45140 28288 45141 28328
rect 45099 28279 45141 28288
rect 45291 28328 45333 28337
rect 45291 28288 45292 28328
rect 45332 28288 45333 28328
rect 45291 28279 45333 28288
rect 45483 28328 45525 28337
rect 45483 28288 45484 28328
rect 45524 28288 45525 28328
rect 45483 28279 45525 28288
rect 45675 28328 45717 28337
rect 45675 28288 45676 28328
rect 45716 28288 45717 28328
rect 45675 28279 45717 28288
rect 45763 28328 45821 28329
rect 45763 28288 45772 28328
rect 45812 28288 45821 28328
rect 45763 28287 45821 28288
rect 49419 28328 49461 28337
rect 49419 28288 49420 28328
rect 49460 28288 49461 28328
rect 49419 28279 49461 28288
rect 49611 28328 49653 28337
rect 49611 28288 49612 28328
rect 49652 28288 49653 28328
rect 49611 28279 49653 28288
rect 49699 28328 49757 28329
rect 49699 28288 49708 28328
rect 49748 28288 49757 28328
rect 49699 28287 49757 28288
rect 49891 28328 49949 28329
rect 49891 28288 49900 28328
rect 49940 28288 49949 28328
rect 49891 28287 49949 28288
rect 49995 28328 50037 28337
rect 49995 28288 49996 28328
rect 50036 28288 50037 28328
rect 49995 28279 50037 28288
rect 50187 28328 50229 28337
rect 50187 28288 50188 28328
rect 50228 28288 50229 28328
rect 50187 28279 50229 28288
rect 50475 28328 50517 28337
rect 50475 28288 50476 28328
rect 50516 28288 50517 28328
rect 50475 28279 50517 28288
rect 50571 28328 50613 28337
rect 50571 28288 50572 28328
rect 50612 28288 50613 28328
rect 50571 28279 50613 28288
rect 50667 28328 50709 28337
rect 50667 28288 50668 28328
rect 50708 28288 50709 28328
rect 50667 28279 50709 28288
rect 51715 28328 51773 28329
rect 51715 28288 51724 28328
rect 51764 28288 51773 28328
rect 51715 28287 51773 28288
rect 51819 28328 51861 28337
rect 51819 28288 51820 28328
rect 51860 28288 51861 28328
rect 51819 28279 51861 28288
rect 51915 28328 51957 28337
rect 51915 28288 51916 28328
rect 51956 28288 51957 28328
rect 51915 28279 51957 28288
rect 52099 28328 52157 28329
rect 52099 28288 52108 28328
rect 52148 28288 52157 28328
rect 52099 28287 52157 28288
rect 52299 28328 52341 28337
rect 52299 28288 52300 28328
rect 52340 28288 52341 28328
rect 52299 28279 52341 28288
rect 53059 28328 53117 28329
rect 53059 28288 53068 28328
rect 53108 28288 53117 28328
rect 53059 28287 53117 28288
rect 55563 28328 55605 28337
rect 55563 28288 55564 28328
rect 55604 28288 55605 28328
rect 55563 28279 55605 28288
rect 55659 28328 55701 28337
rect 55659 28288 55660 28328
rect 55700 28288 55701 28328
rect 55659 28279 55701 28288
rect 55939 28328 55997 28329
rect 55939 28288 55948 28328
rect 55988 28288 55997 28328
rect 55939 28287 55997 28288
rect 56227 28328 56285 28329
rect 56227 28288 56236 28328
rect 56276 28288 56285 28328
rect 56227 28287 56285 28288
rect 56427 28328 56469 28337
rect 56427 28288 56428 28328
rect 56468 28288 56469 28328
rect 56427 28279 56469 28288
rect 59211 28328 59253 28337
rect 59211 28288 59212 28328
rect 59252 28288 59253 28328
rect 59211 28279 59253 28288
rect 59403 28328 59445 28337
rect 59403 28288 59404 28328
rect 59444 28288 59445 28328
rect 59403 28279 59445 28288
rect 59491 28328 59549 28329
rect 59491 28288 59500 28328
rect 59540 28288 59549 28328
rect 59491 28287 59549 28288
rect 59691 28328 59733 28337
rect 59691 28288 59692 28328
rect 59732 28288 59733 28328
rect 59691 28279 59733 28288
rect 59875 28328 59933 28329
rect 59875 28288 59884 28328
rect 59924 28288 59933 28328
rect 59875 28287 59933 28288
rect 60075 28328 60117 28337
rect 60075 28288 60076 28328
rect 60116 28288 60117 28328
rect 60075 28279 60117 28288
rect 60267 28328 60309 28337
rect 60267 28288 60268 28328
rect 60308 28288 60309 28328
rect 60267 28279 60309 28288
rect 60355 28328 60413 28329
rect 60355 28288 60364 28328
rect 60404 28288 60413 28328
rect 60355 28287 60413 28288
rect 60547 28328 60605 28329
rect 60547 28288 60556 28328
rect 60596 28288 60605 28328
rect 60547 28287 60605 28288
rect 60651 28328 60693 28337
rect 60651 28288 60652 28328
rect 60692 28288 60693 28328
rect 60651 28279 60693 28288
rect 60747 28328 60789 28337
rect 60747 28288 60748 28328
rect 60788 28288 60789 28328
rect 60747 28279 60789 28288
rect 62275 28328 62333 28329
rect 62275 28288 62284 28328
rect 62324 28288 62333 28328
rect 62275 28287 62333 28288
rect 63139 28328 63197 28329
rect 63139 28288 63148 28328
rect 63188 28288 63197 28328
rect 63139 28287 63197 28288
rect 64579 28328 64637 28329
rect 64579 28288 64588 28328
rect 64628 28288 64637 28328
rect 64579 28287 64637 28288
rect 64875 28328 64917 28337
rect 64875 28288 64876 28328
rect 64916 28288 64917 28328
rect 64875 28279 64917 28288
rect 66115 28328 66173 28329
rect 66115 28288 66124 28328
rect 66164 28288 66173 28328
rect 66115 28287 66173 28288
rect 66979 28328 67037 28329
rect 66979 28288 66988 28328
rect 67028 28288 67037 28328
rect 66979 28287 67037 28288
rect 70339 28328 70397 28329
rect 70339 28288 70348 28328
rect 70388 28288 70397 28328
rect 70339 28287 70397 28288
rect 70635 28328 70677 28337
rect 70635 28288 70636 28328
rect 70676 28288 70677 28328
rect 70635 28279 70677 28288
rect 70731 28328 70773 28337
rect 70731 28288 70732 28328
rect 70772 28288 70773 28328
rect 70731 28279 70773 28288
rect 71779 28328 71837 28329
rect 71779 28288 71788 28328
rect 71828 28288 71837 28328
rect 71779 28287 71837 28288
rect 72643 28328 72701 28329
rect 72643 28288 72652 28328
rect 72692 28288 72701 28328
rect 72643 28287 72701 28288
rect 75243 28328 75285 28337
rect 75243 28288 75244 28328
rect 75284 28288 75285 28328
rect 75243 28279 75285 28288
rect 75435 28328 75477 28337
rect 75435 28288 75436 28328
rect 75476 28288 75477 28328
rect 75435 28279 75477 28288
rect 75523 28328 75581 28329
rect 75523 28288 75532 28328
rect 75572 28288 75581 28328
rect 75523 28287 75581 28288
rect 76683 28328 76725 28337
rect 76683 28288 76684 28328
rect 76724 28288 76725 28328
rect 76683 28279 76725 28288
rect 76875 28328 76917 28337
rect 76875 28288 76876 28328
rect 76916 28288 76917 28328
rect 76875 28279 76917 28288
rect 76963 28328 77021 28329
rect 76963 28288 76972 28328
rect 77012 28288 77021 28328
rect 76963 28287 77021 28288
rect 77155 28328 77213 28329
rect 77155 28288 77164 28328
rect 77204 28288 77213 28328
rect 77155 28287 77213 28288
rect 77355 28328 77397 28337
rect 77355 28288 77356 28328
rect 77396 28288 77397 28328
rect 77355 28279 77397 28288
rect 40971 28244 41013 28253
rect 40971 28204 40972 28244
rect 41012 28204 41013 28244
rect 40971 28195 41013 28204
rect 52203 28244 52245 28253
rect 52203 28204 52204 28244
rect 52244 28204 52245 28244
rect 52203 28195 52245 28204
rect 56331 28244 56373 28253
rect 56331 28204 56332 28244
rect 56372 28204 56373 28244
rect 56331 28195 56373 28204
rect 61899 28244 61941 28253
rect 61899 28204 61900 28244
rect 61940 28204 61941 28244
rect 61899 28195 61941 28204
rect 64971 28244 65013 28253
rect 64971 28204 64972 28244
rect 65012 28204 65013 28244
rect 64971 28195 65013 28204
rect 65739 28244 65781 28253
rect 65739 28204 65740 28244
rect 65780 28204 65781 28244
rect 65739 28195 65781 28204
rect 71403 28244 71445 28253
rect 71403 28204 71404 28244
rect 71444 28204 71445 28244
rect 71403 28195 71445 28204
rect 75339 28244 75381 28253
rect 75339 28204 75340 28244
rect 75380 28204 75381 28244
rect 75339 28195 75381 28204
rect 77259 28244 77301 28253
rect 77259 28204 77260 28244
rect 77300 28204 77301 28244
rect 77259 28195 77301 28204
rect 39819 28160 39861 28169
rect 39819 28120 39820 28160
rect 39860 28120 39861 28160
rect 39819 28111 39861 28120
rect 40291 28160 40349 28161
rect 40291 28120 40300 28160
rect 40340 28120 40349 28160
rect 40291 28119 40349 28120
rect 44131 28160 44189 28161
rect 44131 28120 44140 28160
rect 44180 28120 44189 28160
rect 44131 28119 44189 28120
rect 45571 28160 45629 28161
rect 45571 28120 45580 28160
rect 45620 28120 45629 28160
rect 45571 28119 45629 28120
rect 49507 28160 49565 28161
rect 49507 28120 49516 28160
rect 49556 28120 49565 28160
rect 49507 28119 49565 28120
rect 50083 28160 50141 28161
rect 50083 28120 50092 28160
rect 50132 28120 50141 28160
rect 50083 28119 50141 28120
rect 50371 28160 50429 28161
rect 50371 28120 50380 28160
rect 50420 28120 50429 28160
rect 50371 28119 50429 28120
rect 51243 28160 51285 28169
rect 51243 28120 51244 28160
rect 51284 28120 51285 28160
rect 51243 28111 51285 28120
rect 59019 28160 59061 28169
rect 59019 28120 59020 28160
rect 59060 28120 59061 28160
rect 59019 28111 59061 28120
rect 59299 28160 59357 28161
rect 59299 28120 59308 28160
rect 59348 28120 59357 28160
rect 59299 28119 59357 28120
rect 60163 28160 60221 28161
rect 60163 28120 60172 28160
rect 60212 28120 60221 28160
rect 60163 28119 60221 28120
rect 61131 28160 61173 28169
rect 61131 28120 61132 28160
rect 61172 28120 61173 28160
rect 61131 28111 61173 28120
rect 64291 28160 64349 28161
rect 64291 28120 64300 28160
rect 64340 28120 64349 28160
rect 64291 28119 64349 28120
rect 68131 28160 68189 28161
rect 68131 28120 68140 28160
rect 68180 28120 68189 28160
rect 68131 28119 68189 28120
rect 69867 28160 69909 28169
rect 69867 28120 69868 28160
rect 69908 28120 69909 28160
rect 69867 28111 69909 28120
rect 73795 28160 73853 28161
rect 73795 28120 73804 28160
rect 73844 28120 73853 28160
rect 73795 28119 73853 28120
rect 576 27992 79584 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79584 27992
rect 576 27928 79584 27952
rect 45955 27824 46013 27825
rect 45955 27784 45964 27824
rect 46004 27784 46013 27824
rect 45955 27783 46013 27784
rect 51235 27824 51293 27825
rect 51235 27784 51244 27824
rect 51284 27784 51293 27824
rect 51235 27783 51293 27784
rect 54499 27824 54557 27825
rect 54499 27784 54508 27824
rect 54548 27784 54557 27824
rect 54499 27783 54557 27784
rect 54787 27824 54845 27825
rect 54787 27784 54796 27824
rect 54836 27784 54845 27824
rect 54787 27783 54845 27784
rect 59683 27824 59741 27825
rect 59683 27784 59692 27824
rect 59732 27784 59741 27824
rect 59683 27783 59741 27784
rect 64003 27824 64061 27825
rect 64003 27784 64012 27824
rect 64052 27784 64061 27824
rect 64003 27783 64061 27784
rect 68619 27824 68661 27833
rect 68619 27784 68620 27824
rect 68660 27784 68661 27824
rect 68619 27775 68661 27784
rect 75523 27824 75581 27825
rect 75523 27784 75532 27824
rect 75572 27784 75581 27824
rect 75523 27783 75581 27784
rect 37707 27740 37749 27749
rect 37707 27700 37708 27740
rect 37748 27700 37749 27740
rect 37707 27691 37749 27700
rect 40395 27740 40437 27749
rect 40395 27700 40396 27740
rect 40436 27700 40437 27740
rect 40395 27691 40437 27700
rect 43563 27740 43605 27749
rect 43563 27700 43564 27740
rect 43604 27700 43605 27740
rect 43563 27691 43605 27700
rect 46443 27740 46485 27749
rect 46443 27700 46444 27740
rect 46484 27700 46485 27740
rect 46443 27691 46485 27700
rect 48843 27740 48885 27749
rect 48843 27700 48844 27740
rect 48884 27700 48885 27740
rect 48843 27691 48885 27700
rect 51723 27740 51765 27749
rect 51723 27700 51724 27740
rect 51764 27700 51765 27740
rect 51723 27691 51765 27700
rect 52107 27740 52149 27749
rect 52107 27700 52108 27740
rect 52148 27700 52149 27740
rect 52107 27691 52149 27700
rect 57099 27740 57141 27749
rect 57099 27700 57100 27740
rect 57140 27700 57141 27740
rect 57099 27691 57141 27700
rect 60459 27740 60501 27749
rect 60459 27700 60460 27740
rect 60500 27700 60501 27740
rect 60459 27691 60501 27700
rect 65259 27740 65301 27749
rect 65259 27700 65260 27740
rect 65300 27700 65301 27740
rect 65259 27691 65301 27700
rect 70731 27740 70773 27749
rect 70731 27700 70732 27740
rect 70772 27700 70773 27740
rect 70731 27691 70773 27700
rect 71115 27740 71157 27749
rect 71115 27700 71116 27740
rect 71156 27700 71157 27740
rect 71115 27691 71157 27700
rect 38083 27656 38141 27657
rect 38083 27616 38092 27656
rect 38132 27616 38141 27656
rect 38083 27615 38141 27616
rect 38947 27656 39005 27657
rect 38947 27616 38956 27656
rect 38996 27616 39005 27656
rect 38947 27615 39005 27616
rect 40299 27656 40341 27665
rect 40299 27616 40300 27656
rect 40340 27616 40341 27656
rect 40299 27607 40341 27616
rect 40491 27656 40533 27665
rect 40491 27616 40492 27656
rect 40532 27616 40533 27656
rect 40491 27607 40533 27616
rect 40579 27656 40637 27657
rect 40579 27616 40588 27656
rect 40628 27616 40637 27656
rect 40579 27615 40637 27616
rect 40963 27656 41021 27657
rect 40963 27616 40972 27656
rect 41012 27616 41021 27656
rect 40963 27615 41021 27616
rect 41163 27656 41205 27665
rect 41163 27616 41164 27656
rect 41204 27616 41205 27656
rect 41163 27607 41205 27616
rect 43939 27656 43997 27657
rect 43939 27616 43948 27656
rect 43988 27616 43997 27656
rect 43939 27615 43997 27616
rect 44803 27656 44861 27657
rect 44803 27616 44812 27656
rect 44852 27616 44861 27656
rect 44803 27615 44861 27616
rect 46539 27656 46581 27665
rect 46539 27616 46540 27656
rect 46580 27616 46581 27656
rect 46539 27607 46581 27616
rect 46819 27656 46877 27657
rect 46819 27616 46828 27656
rect 46868 27616 46877 27656
rect 46819 27615 46877 27616
rect 47115 27656 47157 27665
rect 47115 27616 47116 27656
rect 47156 27616 47157 27656
rect 47115 27607 47157 27616
rect 47307 27656 47349 27665
rect 47307 27616 47308 27656
rect 47348 27616 47349 27656
rect 47307 27607 47349 27616
rect 47395 27656 47453 27657
rect 47395 27616 47404 27656
rect 47444 27616 47453 27656
rect 47395 27615 47453 27616
rect 47587 27656 47645 27657
rect 47587 27616 47596 27656
rect 47636 27616 47645 27656
rect 47587 27615 47645 27616
rect 47691 27656 47733 27665
rect 47691 27616 47692 27656
rect 47732 27616 47733 27656
rect 47691 27607 47733 27616
rect 47787 27656 47829 27665
rect 47787 27616 47788 27656
rect 47828 27616 47829 27656
rect 47787 27607 47829 27616
rect 49219 27656 49277 27657
rect 49219 27616 49228 27656
rect 49268 27616 49277 27656
rect 49219 27615 49277 27616
rect 50083 27656 50141 27657
rect 50083 27616 50092 27656
rect 50132 27616 50141 27656
rect 50083 27615 50141 27616
rect 51627 27656 51669 27665
rect 51627 27616 51628 27656
rect 51668 27616 51669 27656
rect 51627 27607 51669 27616
rect 51819 27656 51861 27665
rect 51819 27616 51820 27656
rect 51860 27616 51861 27656
rect 51819 27607 51861 27616
rect 51907 27656 51965 27657
rect 51907 27616 51916 27656
rect 51956 27616 51965 27656
rect 51907 27615 51965 27616
rect 52483 27656 52541 27657
rect 52483 27616 52492 27656
rect 52532 27616 52541 27656
rect 52483 27615 52541 27616
rect 53347 27656 53405 27657
rect 53347 27616 53356 27656
rect 53396 27616 53405 27656
rect 53347 27615 53405 27616
rect 54699 27656 54741 27665
rect 54699 27616 54700 27656
rect 54740 27616 54741 27656
rect 54699 27607 54741 27616
rect 54891 27656 54933 27665
rect 54891 27616 54892 27656
rect 54932 27616 54933 27656
rect 54891 27607 54933 27616
rect 54979 27656 55037 27657
rect 54979 27616 54988 27656
rect 55028 27616 55037 27656
rect 54979 27615 55037 27616
rect 55179 27656 55221 27665
rect 55179 27616 55180 27656
rect 55220 27616 55221 27656
rect 55179 27607 55221 27616
rect 55371 27656 55413 27665
rect 55371 27616 55372 27656
rect 55412 27616 55413 27656
rect 55371 27607 55413 27616
rect 55459 27656 55517 27657
rect 55459 27616 55468 27656
rect 55508 27616 55517 27656
rect 55459 27615 55517 27616
rect 55659 27656 55701 27665
rect 55659 27616 55660 27656
rect 55700 27616 55701 27656
rect 55659 27607 55701 27616
rect 55755 27656 55797 27665
rect 55755 27616 55756 27656
rect 55796 27616 55797 27656
rect 55755 27607 55797 27616
rect 55851 27656 55893 27665
rect 55851 27616 55852 27656
rect 55892 27616 55893 27656
rect 55851 27607 55893 27616
rect 55947 27656 55989 27665
rect 55947 27616 55948 27656
rect 55988 27616 55989 27656
rect 55947 27607 55989 27616
rect 57475 27656 57533 27657
rect 57475 27616 57484 27656
rect 57524 27616 57533 27656
rect 57475 27615 57533 27616
rect 58339 27656 58397 27657
rect 58339 27616 58348 27656
rect 58388 27616 58397 27656
rect 58339 27615 58397 27616
rect 59787 27656 59829 27665
rect 59787 27616 59788 27656
rect 59828 27616 59829 27656
rect 59787 27607 59829 27616
rect 59883 27656 59925 27665
rect 59883 27616 59884 27656
rect 59924 27616 59925 27656
rect 59883 27607 59925 27616
rect 59979 27656 60021 27665
rect 59979 27616 59980 27656
rect 60020 27616 60021 27656
rect 59979 27607 60021 27616
rect 60835 27656 60893 27657
rect 60835 27616 60844 27656
rect 60884 27616 60893 27656
rect 60835 27615 60893 27616
rect 61699 27656 61757 27657
rect 61699 27616 61708 27656
rect 61748 27616 61757 27656
rect 61699 27615 61757 27616
rect 63811 27656 63869 27657
rect 63811 27616 63820 27656
rect 63860 27616 63869 27656
rect 63811 27615 63869 27616
rect 63915 27656 63957 27665
rect 63915 27616 63916 27656
rect 63956 27616 63957 27656
rect 63915 27607 63957 27616
rect 64107 27656 64149 27665
rect 64107 27616 64108 27656
rect 64148 27616 64149 27656
rect 64107 27607 64149 27616
rect 65163 27656 65205 27665
rect 65163 27616 65164 27656
rect 65204 27616 65205 27656
rect 65163 27607 65205 27616
rect 65355 27656 65397 27665
rect 65355 27616 65356 27656
rect 65396 27616 65397 27656
rect 65355 27607 65397 27616
rect 65443 27656 65501 27657
rect 65443 27616 65452 27656
rect 65492 27616 65501 27656
rect 65443 27615 65501 27616
rect 65635 27656 65693 27657
rect 65635 27616 65644 27656
rect 65684 27616 65693 27656
rect 65635 27615 65693 27616
rect 65835 27656 65877 27665
rect 65835 27616 65836 27656
rect 65876 27616 65877 27656
rect 65835 27607 65877 27616
rect 69579 27656 69621 27665
rect 69579 27616 69580 27656
rect 69620 27616 69621 27656
rect 69579 27607 69621 27616
rect 69771 27656 69813 27665
rect 69771 27616 69772 27656
rect 69812 27616 69813 27656
rect 69771 27607 69813 27616
rect 69859 27656 69917 27657
rect 69859 27616 69868 27656
rect 69908 27616 69917 27656
rect 69859 27615 69917 27616
rect 70059 27656 70101 27665
rect 70059 27616 70060 27656
rect 70100 27616 70101 27656
rect 70059 27607 70101 27616
rect 70251 27656 70293 27665
rect 70251 27616 70252 27656
rect 70292 27616 70293 27656
rect 70251 27607 70293 27616
rect 70339 27656 70397 27657
rect 70339 27616 70348 27656
rect 70388 27616 70397 27656
rect 70339 27615 70397 27616
rect 70627 27656 70685 27657
rect 70627 27616 70636 27656
rect 70676 27616 70685 27656
rect 70627 27615 70685 27616
rect 70827 27656 70869 27665
rect 70827 27616 70828 27656
rect 70868 27616 70869 27656
rect 70827 27607 70869 27616
rect 71019 27656 71061 27665
rect 71019 27616 71020 27656
rect 71060 27616 71061 27656
rect 71019 27607 71061 27616
rect 71211 27656 71253 27665
rect 71211 27616 71212 27656
rect 71252 27616 71253 27656
rect 71211 27607 71253 27616
rect 71299 27656 71357 27657
rect 71299 27616 71308 27656
rect 71348 27616 71357 27656
rect 71299 27615 71357 27616
rect 74859 27656 74901 27665
rect 74859 27616 74860 27656
rect 74900 27616 74901 27656
rect 74859 27607 74901 27616
rect 75051 27656 75093 27665
rect 75051 27616 75052 27656
rect 75092 27616 75093 27656
rect 75051 27607 75093 27616
rect 75139 27656 75197 27657
rect 75139 27616 75148 27656
rect 75188 27616 75197 27656
rect 75139 27615 75197 27616
rect 75435 27656 75477 27665
rect 75435 27616 75436 27656
rect 75476 27616 75477 27656
rect 75435 27607 75477 27616
rect 75627 27656 75669 27665
rect 75627 27616 75628 27656
rect 75668 27616 75669 27656
rect 75627 27607 75669 27616
rect 75715 27656 75773 27657
rect 75715 27616 75724 27656
rect 75764 27616 75773 27656
rect 75715 27615 75773 27616
rect 76771 27656 76829 27657
rect 76771 27616 76780 27656
rect 76820 27616 76829 27656
rect 76771 27615 76829 27616
rect 76875 27656 76917 27665
rect 76875 27616 76876 27656
rect 76916 27616 76917 27656
rect 76875 27607 76917 27616
rect 76971 27656 77013 27665
rect 76971 27616 76972 27656
rect 77012 27616 77013 27656
rect 76971 27607 77013 27616
rect 77155 27656 77213 27657
rect 77155 27616 77164 27656
rect 77204 27616 77213 27656
rect 77155 27615 77213 27616
rect 77355 27656 77397 27665
rect 77355 27616 77356 27656
rect 77396 27616 77397 27656
rect 77355 27607 77397 27616
rect 41539 27572 41597 27573
rect 41539 27532 41548 27572
rect 41588 27532 41597 27572
rect 41539 27531 41597 27532
rect 65739 27572 65781 27581
rect 65739 27532 65740 27572
rect 65780 27532 65781 27572
rect 65739 27523 65781 27532
rect 67555 27572 67613 27573
rect 67555 27532 67564 27572
rect 67604 27532 67613 27572
rect 67555 27531 67613 27532
rect 68419 27572 68477 27573
rect 68419 27532 68428 27572
rect 68468 27532 68477 27572
rect 68419 27531 68477 27532
rect 36459 27488 36501 27497
rect 36459 27448 36460 27488
rect 36500 27448 36501 27488
rect 36459 27439 36501 27448
rect 41355 27488 41397 27497
rect 41355 27448 41356 27488
rect 41396 27448 41397 27488
rect 41355 27439 41397 27448
rect 55179 27488 55221 27497
rect 55179 27448 55180 27488
rect 55220 27448 55221 27488
rect 55179 27439 55221 27448
rect 66219 27488 66261 27497
rect 66219 27448 66220 27488
rect 66260 27448 66261 27488
rect 66219 27439 66261 27448
rect 69387 27488 69429 27497
rect 69387 27448 69388 27488
rect 69428 27448 69429 27488
rect 69387 27439 69429 27448
rect 70059 27488 70101 27497
rect 70059 27448 70060 27488
rect 70100 27448 70101 27488
rect 70059 27439 70101 27448
rect 71883 27488 71925 27497
rect 71883 27448 71884 27488
rect 71924 27448 71925 27488
rect 71883 27439 71925 27448
rect 73515 27488 73557 27497
rect 73515 27448 73516 27488
rect 73556 27448 73557 27488
rect 73515 27439 73557 27448
rect 77547 27488 77589 27497
rect 77547 27448 77548 27488
rect 77588 27448 77589 27488
rect 77547 27439 77589 27448
rect 40099 27404 40157 27405
rect 40099 27364 40108 27404
rect 40148 27364 40157 27404
rect 40099 27363 40157 27364
rect 41067 27404 41109 27413
rect 41067 27364 41068 27404
rect 41108 27364 41109 27404
rect 41067 27355 41109 27364
rect 46147 27404 46205 27405
rect 46147 27364 46156 27404
rect 46196 27364 46205 27404
rect 46147 27363 46205 27364
rect 47115 27404 47157 27413
rect 47115 27364 47116 27404
rect 47156 27364 47157 27404
rect 47115 27355 47157 27364
rect 51235 27404 51293 27405
rect 51235 27364 51244 27404
rect 51284 27364 51293 27404
rect 51235 27363 51293 27364
rect 59491 27404 59549 27405
rect 59491 27364 59500 27404
rect 59540 27364 59549 27404
rect 59491 27363 59549 27364
rect 62851 27404 62909 27405
rect 62851 27364 62860 27404
rect 62900 27364 62909 27404
rect 62851 27363 62909 27364
rect 67371 27404 67413 27413
rect 67371 27364 67372 27404
rect 67412 27364 67413 27404
rect 67371 27355 67413 27364
rect 69579 27404 69621 27413
rect 69579 27364 69580 27404
rect 69620 27364 69621 27404
rect 69579 27355 69621 27364
rect 74859 27404 74901 27413
rect 74859 27364 74860 27404
rect 74900 27364 74901 27404
rect 74859 27355 74901 27364
rect 77259 27404 77301 27413
rect 77259 27364 77260 27404
rect 77300 27364 77301 27404
rect 77259 27355 77301 27364
rect 576 27236 79584 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79584 27236
rect 576 27172 79584 27196
rect 41059 27068 41117 27069
rect 41059 27028 41068 27068
rect 41108 27028 41117 27068
rect 41059 27027 41117 27028
rect 44907 27068 44949 27077
rect 44907 27028 44908 27068
rect 44948 27028 44949 27068
rect 44907 27019 44949 27028
rect 45867 27068 45909 27077
rect 45867 27028 45868 27068
rect 45908 27028 45909 27068
rect 45867 27019 45909 27028
rect 46347 27068 46389 27077
rect 46347 27028 46348 27068
rect 46388 27028 46389 27068
rect 46347 27019 46389 27028
rect 49411 27068 49469 27069
rect 49411 27028 49420 27068
rect 49460 27028 49469 27068
rect 49411 27027 49469 27028
rect 51907 27068 51965 27069
rect 51907 27028 51916 27068
rect 51956 27028 51965 27068
rect 51907 27027 51965 27028
rect 54211 27068 54269 27069
rect 54211 27028 54220 27068
rect 54260 27028 54269 27068
rect 54211 27027 54269 27028
rect 58443 27068 58485 27077
rect 58443 27028 58444 27068
rect 58484 27028 58485 27068
rect 58443 27019 58485 27028
rect 59395 27068 59453 27069
rect 59395 27028 59404 27068
rect 59444 27028 59453 27068
rect 59395 27027 59453 27028
rect 60747 27068 60789 27077
rect 60747 27028 60748 27068
rect 60788 27028 60789 27068
rect 60747 27019 60789 27028
rect 63819 27068 63861 27077
rect 63819 27028 63820 27068
rect 63860 27028 63861 27068
rect 63819 27019 63861 27028
rect 71883 27068 71925 27077
rect 71883 27028 71884 27068
rect 71924 27028 71925 27068
rect 71883 27019 71925 27028
rect 72075 27068 72117 27077
rect 72075 27028 72076 27068
rect 72116 27028 72117 27068
rect 72075 27019 72117 27028
rect 76867 27068 76925 27069
rect 76867 27028 76876 27068
rect 76916 27028 76925 27068
rect 76867 27027 76925 27028
rect 33003 26984 33045 26993
rect 33003 26944 33004 26984
rect 33044 26944 33045 26984
rect 33003 26935 33045 26944
rect 35307 26984 35349 26993
rect 35307 26944 35308 26984
rect 35348 26944 35349 26984
rect 35307 26935 35349 26944
rect 38859 26984 38901 26993
rect 38859 26944 38860 26984
rect 38900 26944 38901 26984
rect 38859 26935 38901 26944
rect 53451 26984 53493 26993
rect 53451 26944 53452 26984
rect 53492 26944 53493 26984
rect 53451 26935 53493 26944
rect 57579 26984 57621 26993
rect 57579 26944 57580 26984
rect 57620 26944 57621 26984
rect 57579 26935 57621 26944
rect 61131 26984 61173 26993
rect 61131 26944 61132 26984
rect 61172 26944 61173 26984
rect 61131 26935 61173 26944
rect 62091 26984 62133 26993
rect 62091 26944 62092 26984
rect 62132 26944 62133 26984
rect 62091 26935 62133 26944
rect 35587 26900 35645 26901
rect 35587 26860 35596 26900
rect 35636 26860 35645 26900
rect 35587 26859 35645 26860
rect 38659 26900 38717 26901
rect 38659 26860 38668 26900
rect 38708 26860 38717 26900
rect 38659 26859 38717 26860
rect 39043 26900 39101 26901
rect 39043 26860 39052 26900
rect 39092 26860 39101 26900
rect 39043 26859 39101 26860
rect 39427 26900 39485 26901
rect 39427 26860 39436 26900
rect 39476 26860 39485 26900
rect 39427 26859 39485 26860
rect 44707 26900 44765 26901
rect 44707 26860 44716 26900
rect 44756 26860 44765 26900
rect 44707 26859 44765 26860
rect 52099 26900 52157 26901
rect 52099 26860 52108 26900
rect 52148 26860 52157 26900
rect 52099 26859 52157 26860
rect 58243 26900 58301 26901
rect 58243 26860 58252 26900
rect 58292 26860 58301 26900
rect 58243 26859 58301 26860
rect 59011 26900 59069 26901
rect 59011 26860 59020 26900
rect 59060 26860 59069 26900
rect 59011 26859 59069 26860
rect 60355 26900 60413 26901
rect 60355 26860 60364 26900
rect 60404 26860 60413 26900
rect 60355 26859 60413 26860
rect 60931 26900 60989 26901
rect 60931 26860 60940 26900
rect 60980 26860 60989 26900
rect 60931 26859 60989 26860
rect 71683 26900 71741 26901
rect 71683 26860 71692 26900
rect 71732 26860 71741 26900
rect 71683 26859 71741 26860
rect 72259 26900 72317 26901
rect 72259 26860 72268 26900
rect 72308 26860 72317 26900
rect 72259 26859 72317 26860
rect 75435 26900 75477 26909
rect 75435 26860 75436 26900
rect 75476 26860 75477 26900
rect 73411 26852 73469 26853
rect 4291 26816 4349 26817
rect 4291 26776 4300 26816
rect 4340 26776 4349 26816
rect 4291 26775 4349 26776
rect 35203 26816 35261 26817
rect 35203 26776 35212 26816
rect 35252 26776 35261 26816
rect 35203 26775 35261 26776
rect 35403 26816 35445 26825
rect 35403 26776 35404 26816
rect 35444 26776 35445 26816
rect 35403 26767 35445 26776
rect 36355 26816 36413 26817
rect 36355 26776 36364 26816
rect 36404 26776 36413 26816
rect 36355 26775 36413 26776
rect 37219 26816 37277 26817
rect 37219 26776 37228 26816
rect 37268 26776 37277 26816
rect 37219 26775 37277 26776
rect 39819 26816 39861 26825
rect 39819 26776 39820 26816
rect 39860 26776 39861 26816
rect 39819 26767 39861 26776
rect 39915 26816 39957 26825
rect 39915 26776 39916 26816
rect 39956 26776 39957 26816
rect 39915 26767 39957 26776
rect 40011 26816 40053 26825
rect 40011 26776 40012 26816
rect 40052 26776 40053 26816
rect 40011 26767 40053 26776
rect 40107 26816 40149 26825
rect 40107 26776 40108 26816
rect 40148 26776 40149 26816
rect 40107 26767 40149 26776
rect 40387 26816 40445 26817
rect 40387 26776 40396 26816
rect 40436 26776 40445 26816
rect 40387 26775 40445 26776
rect 40683 26816 40725 26825
rect 40683 26776 40684 26816
rect 40724 26776 40725 26816
rect 40683 26767 40725 26776
rect 40779 26816 40821 26825
rect 40779 26776 40780 26816
rect 40820 26776 40821 26816
rect 40779 26767 40821 26776
rect 41251 26816 41309 26817
rect 41251 26776 41260 26816
rect 41300 26776 41309 26816
rect 41251 26775 41309 26776
rect 41355 26816 41397 26825
rect 41355 26776 41356 26816
rect 41396 26776 41397 26816
rect 41355 26767 41397 26776
rect 41451 26816 41493 26825
rect 41451 26776 41452 26816
rect 41492 26776 41493 26816
rect 41451 26767 41493 26776
rect 42019 26816 42077 26817
rect 42019 26776 42028 26816
rect 42068 26776 42077 26816
rect 42019 26775 42077 26776
rect 42883 26816 42941 26817
rect 42883 26776 42892 26816
rect 42932 26776 42941 26816
rect 42883 26775 42941 26776
rect 45099 26816 45141 26825
rect 45099 26776 45100 26816
rect 45140 26776 45141 26816
rect 45099 26767 45141 26776
rect 45195 26816 45237 26825
rect 45195 26776 45196 26816
rect 45236 26776 45237 26816
rect 45195 26767 45237 26776
rect 45291 26816 45333 26825
rect 45291 26776 45292 26816
rect 45332 26776 45333 26816
rect 45291 26767 45333 26776
rect 45387 26816 45429 26825
rect 45387 26776 45388 26816
rect 45428 26776 45429 26816
rect 45387 26767 45429 26776
rect 45571 26816 45629 26817
rect 45571 26776 45580 26816
rect 45620 26776 45629 26816
rect 45571 26775 45629 26776
rect 45675 26816 45717 26825
rect 45675 26776 45676 26816
rect 45716 26776 45717 26816
rect 45675 26767 45717 26776
rect 45867 26816 45909 26825
rect 45867 26776 45868 26816
rect 45908 26776 45909 26816
rect 46435 26816 46493 26817
rect 45867 26767 45909 26776
rect 46242 26803 46284 26812
rect 46242 26763 46243 26803
rect 46283 26763 46284 26803
rect 46435 26776 46444 26816
rect 46484 26776 46493 26816
rect 46435 26775 46493 26776
rect 46627 26816 46685 26817
rect 46627 26776 46636 26816
rect 46676 26776 46685 26816
rect 46627 26775 46685 26776
rect 46827 26816 46869 26825
rect 46827 26776 46828 26816
rect 46868 26776 46869 26816
rect 46827 26767 46869 26776
rect 47019 26816 47061 26825
rect 47019 26776 47020 26816
rect 47060 26776 47061 26816
rect 47019 26767 47061 26776
rect 47395 26816 47453 26817
rect 47395 26776 47404 26816
rect 47444 26776 47453 26816
rect 47395 26775 47453 26776
rect 48259 26816 48317 26817
rect 48259 26776 48268 26816
rect 48308 26776 48317 26816
rect 48259 26775 48317 26776
rect 50091 26816 50133 26825
rect 50091 26776 50092 26816
rect 50132 26776 50133 26816
rect 50091 26767 50133 26776
rect 50283 26816 50325 26825
rect 50283 26776 50284 26816
rect 50324 26776 50325 26816
rect 50283 26767 50325 26776
rect 50371 26816 50429 26817
rect 50371 26776 50380 26816
rect 50420 26776 50429 26816
rect 50371 26775 50429 26776
rect 50563 26816 50621 26817
rect 50563 26776 50572 26816
rect 50612 26776 50621 26816
rect 50563 26775 50621 26776
rect 50667 26816 50709 26825
rect 50667 26776 50668 26816
rect 50708 26776 50709 26816
rect 50667 26767 50709 26776
rect 50859 26816 50901 26825
rect 50859 26776 50860 26816
rect 50900 26776 50901 26816
rect 50859 26767 50901 26776
rect 51235 26816 51293 26817
rect 51235 26776 51244 26816
rect 51284 26776 51293 26816
rect 51235 26775 51293 26776
rect 51531 26816 51573 26825
rect 51531 26776 51532 26816
rect 51572 26776 51573 26816
rect 51531 26767 51573 26776
rect 51627 26816 51669 26825
rect 51627 26776 51628 26816
rect 51668 26776 51669 26816
rect 51627 26767 51669 26776
rect 55363 26816 55421 26817
rect 55363 26776 55372 26816
rect 55412 26776 55421 26816
rect 55363 26775 55421 26776
rect 56227 26816 56285 26817
rect 56227 26776 56236 26816
rect 56276 26776 56285 26816
rect 56227 26775 56285 26776
rect 59787 26816 59829 26825
rect 59787 26776 59788 26816
rect 59828 26776 59829 26816
rect 59787 26767 59829 26776
rect 60067 26816 60125 26817
rect 60067 26776 60076 26816
rect 60116 26776 60125 26816
rect 60067 26775 60125 26776
rect 63819 26816 63861 26825
rect 63819 26776 63820 26816
rect 63860 26776 63861 26816
rect 63819 26767 63861 26776
rect 64011 26816 64053 26825
rect 64011 26776 64012 26816
rect 64052 26776 64053 26816
rect 64011 26767 64053 26776
rect 64099 26816 64157 26817
rect 64099 26776 64108 26816
rect 64148 26776 64157 26816
rect 64099 26775 64157 26776
rect 66883 26816 66941 26817
rect 66883 26776 66892 26816
rect 66932 26776 66941 26816
rect 66883 26775 66941 26776
rect 67747 26816 67805 26817
rect 67747 26776 67756 26816
rect 67796 26776 67805 26816
rect 67747 26775 67805 26776
rect 68331 26816 68373 26825
rect 68331 26776 68332 26816
rect 68372 26776 68373 26816
rect 68331 26767 68373 26776
rect 68523 26816 68565 26825
rect 68523 26776 68524 26816
rect 68564 26776 68565 26816
rect 68523 26767 68565 26776
rect 68611 26816 68669 26817
rect 68611 26776 68620 26816
rect 68660 26776 68669 26816
rect 68611 26775 68669 26776
rect 69099 26816 69141 26825
rect 69099 26776 69100 26816
rect 69140 26776 69141 26816
rect 69099 26767 69141 26776
rect 69475 26816 69533 26817
rect 69475 26776 69484 26816
rect 69524 26776 69533 26816
rect 69475 26775 69533 26776
rect 70339 26816 70397 26817
rect 70339 26776 70348 26816
rect 70388 26776 70397 26816
rect 70339 26775 70397 26776
rect 73035 26816 73077 26825
rect 73035 26776 73036 26816
rect 73076 26776 73077 26816
rect 73411 26812 73420 26852
rect 73460 26812 73469 26852
rect 75435 26851 75477 26860
rect 73411 26811 73469 26812
rect 74275 26816 74333 26817
rect 73035 26767 73077 26776
rect 74275 26776 74284 26816
rect 74324 26776 74333 26816
rect 74275 26775 74333 26776
rect 75627 26816 75669 26825
rect 75627 26776 75628 26816
rect 75668 26776 75669 26816
rect 75627 26767 75669 26776
rect 75723 26816 75765 26825
rect 75723 26776 75724 26816
rect 75764 26776 75765 26816
rect 75915 26816 75957 26825
rect 75723 26767 75765 26776
rect 75819 26795 75861 26804
rect 46242 26754 46284 26763
rect 75819 26755 75820 26795
rect 75860 26755 75861 26795
rect 75915 26776 75916 26816
rect 75956 26776 75957 26816
rect 75915 26767 75957 26776
rect 76195 26816 76253 26817
rect 76195 26776 76204 26816
rect 76244 26776 76253 26816
rect 76195 26775 76253 26776
rect 76491 26816 76533 26825
rect 76491 26776 76492 26816
rect 76532 26776 76533 26816
rect 76491 26767 76533 26776
rect 76587 26816 76629 26825
rect 76587 26776 76588 26816
rect 76628 26776 76629 26816
rect 76587 26767 76629 26776
rect 77443 26816 77501 26817
rect 77443 26776 77452 26816
rect 77492 26776 77501 26816
rect 77443 26775 77501 26776
rect 78307 26816 78365 26817
rect 78307 26776 78316 26816
rect 78356 26776 78365 26816
rect 78307 26775 78365 26776
rect 75819 26746 75861 26755
rect 35979 26732 36021 26741
rect 35979 26692 35980 26732
rect 36020 26692 36021 26732
rect 35979 26683 36021 26692
rect 41643 26732 41685 26741
rect 41643 26692 41644 26732
rect 41684 26692 41685 26732
rect 41643 26683 41685 26692
rect 46731 26732 46773 26741
rect 46731 26692 46732 26732
rect 46772 26692 46773 26732
rect 46731 26683 46773 26692
rect 50187 26732 50229 26741
rect 50187 26692 50188 26732
rect 50228 26692 50229 26732
rect 50187 26683 50229 26692
rect 56619 26732 56661 26741
rect 56619 26692 56620 26732
rect 56660 26692 56661 26732
rect 56619 26683 56661 26692
rect 59691 26732 59733 26741
rect 59691 26692 59692 26732
rect 59732 26692 59733 26732
rect 59691 26683 59733 26692
rect 68139 26732 68181 26741
rect 68139 26692 68140 26732
rect 68180 26692 68181 26732
rect 68139 26683 68181 26692
rect 77067 26732 77109 26741
rect 77067 26692 77068 26732
rect 77108 26692 77109 26732
rect 77067 26683 77109 26692
rect 4203 26648 4245 26657
rect 4203 26608 4204 26648
rect 4244 26608 4245 26648
rect 4203 26599 4245 26608
rect 35787 26648 35829 26657
rect 35787 26608 35788 26648
rect 35828 26608 35829 26648
rect 35787 26599 35829 26608
rect 38371 26648 38429 26649
rect 38371 26608 38380 26648
rect 38420 26608 38429 26648
rect 38371 26607 38429 26608
rect 39243 26648 39285 26657
rect 39243 26608 39244 26648
rect 39284 26608 39285 26648
rect 39243 26599 39285 26608
rect 39627 26648 39669 26657
rect 39627 26608 39628 26648
rect 39668 26608 39669 26648
rect 39627 26599 39669 26608
rect 44035 26648 44093 26649
rect 44035 26608 44044 26648
rect 44084 26608 44093 26648
rect 44035 26607 44093 26608
rect 44907 26648 44949 26657
rect 44907 26608 44908 26648
rect 44948 26608 44949 26648
rect 44907 26599 44949 26608
rect 49411 26648 49469 26649
rect 49411 26608 49420 26648
rect 49460 26608 49469 26648
rect 49411 26607 49469 26608
rect 50755 26648 50813 26649
rect 50755 26608 50764 26648
rect 50804 26608 50813 26648
rect 50755 26607 50813 26608
rect 52299 26648 52341 26657
rect 52299 26608 52300 26648
rect 52340 26608 52341 26648
rect 52299 26599 52341 26608
rect 58827 26648 58869 26657
rect 58827 26608 58828 26648
rect 58868 26608 58869 26648
rect 58827 26599 58869 26608
rect 60555 26648 60597 26657
rect 60555 26608 60556 26648
rect 60596 26608 60597 26648
rect 60555 26599 60597 26608
rect 60747 26648 60789 26657
rect 60747 26608 60748 26648
rect 60788 26608 60789 26648
rect 60747 26599 60789 26608
rect 65731 26648 65789 26649
rect 65731 26608 65740 26648
rect 65780 26608 65789 26648
rect 65731 26607 65789 26608
rect 68419 26648 68477 26649
rect 68419 26608 68428 26648
rect 68468 26608 68477 26648
rect 68419 26607 68477 26608
rect 71491 26648 71549 26649
rect 71491 26608 71500 26648
rect 71540 26608 71549 26648
rect 71491 26607 71549 26608
rect 71883 26648 71925 26657
rect 71883 26608 71884 26648
rect 71924 26608 71925 26648
rect 71883 26599 71925 26608
rect 79459 26648 79517 26649
rect 79459 26608 79468 26648
rect 79508 26608 79517 26648
rect 79459 26607 79517 26608
rect 576 26480 79584 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79584 26480
rect 576 26416 79584 26440
rect 35875 26312 35933 26313
rect 35875 26272 35884 26312
rect 35924 26272 35933 26312
rect 35875 26271 35933 26272
rect 39147 26312 39189 26321
rect 39147 26272 39148 26312
rect 39188 26272 39189 26312
rect 39147 26263 39189 26272
rect 56419 26312 56477 26313
rect 56419 26272 56428 26312
rect 56468 26272 56477 26312
rect 56419 26271 56477 26272
rect 57675 26312 57717 26321
rect 57675 26272 57676 26312
rect 57716 26272 57717 26312
rect 57675 26263 57717 26272
rect 61227 26312 61269 26321
rect 61227 26272 61228 26312
rect 61268 26272 61269 26312
rect 61227 26263 61269 26272
rect 67747 26312 67805 26313
rect 67747 26272 67756 26312
rect 67796 26272 67805 26312
rect 67747 26271 67805 26272
rect 69571 26312 69629 26313
rect 69571 26272 69580 26312
rect 69620 26272 69629 26312
rect 69571 26271 69629 26272
rect 75235 26312 75293 26313
rect 75235 26272 75244 26312
rect 75284 26272 75293 26312
rect 75235 26271 75293 26272
rect 76963 26312 77021 26313
rect 76963 26272 76972 26312
rect 77012 26272 77021 26312
rect 76963 26271 77021 26272
rect 36363 26228 36405 26237
rect 36363 26188 36364 26228
rect 36404 26188 36405 26228
rect 48747 26228 48789 26237
rect 36363 26179 36405 26188
rect 39819 26186 39861 26195
rect 33379 26144 33437 26145
rect 33379 26104 33388 26144
rect 33428 26104 33437 26144
rect 33379 26103 33437 26104
rect 34243 26144 34301 26145
rect 34243 26104 34252 26144
rect 34292 26104 34301 26144
rect 34243 26103 34301 26104
rect 34635 26144 34677 26153
rect 34635 26104 34636 26144
rect 34676 26104 34677 26144
rect 34635 26095 34677 26104
rect 34915 26144 34973 26145
rect 34915 26104 34924 26144
rect 34964 26104 34973 26144
rect 34915 26103 34973 26104
rect 35211 26144 35253 26153
rect 35211 26104 35212 26144
rect 35252 26104 35253 26144
rect 35211 26095 35253 26104
rect 35307 26144 35349 26153
rect 35307 26104 35308 26144
rect 35348 26104 35349 26144
rect 35307 26095 35349 26104
rect 35787 26144 35829 26153
rect 35787 26104 35788 26144
rect 35828 26104 35829 26144
rect 35787 26095 35829 26104
rect 35979 26144 36021 26153
rect 35979 26104 35980 26144
rect 36020 26104 36021 26144
rect 35979 26095 36021 26104
rect 36067 26144 36125 26145
rect 36067 26104 36076 26144
rect 36116 26104 36125 26144
rect 36067 26103 36125 26104
rect 36259 26144 36317 26145
rect 36259 26104 36268 26144
rect 36308 26104 36317 26144
rect 36259 26103 36317 26104
rect 36459 26144 36501 26153
rect 36459 26104 36460 26144
rect 36500 26104 36501 26144
rect 36459 26095 36501 26104
rect 39339 26144 39381 26153
rect 39339 26104 39340 26144
rect 39380 26104 39381 26144
rect 39339 26095 39381 26104
rect 39531 26144 39573 26153
rect 39819 26146 39820 26186
rect 39860 26146 39861 26186
rect 48747 26188 48748 26228
rect 48788 26188 48789 26228
rect 48747 26179 48789 26188
rect 52107 26228 52149 26237
rect 52107 26188 52108 26228
rect 52148 26188 52149 26228
rect 52107 26179 52149 26188
rect 55851 26228 55893 26237
rect 55851 26188 55852 26228
rect 55892 26188 55893 26228
rect 55851 26179 55893 26188
rect 61611 26228 61653 26237
rect 61611 26188 61612 26228
rect 61652 26188 61653 26228
rect 61611 26179 61653 26188
rect 64779 26228 64821 26237
rect 64779 26188 64780 26228
rect 64820 26188 64821 26228
rect 64779 26179 64821 26188
rect 71307 26228 71349 26237
rect 71307 26188 71308 26228
rect 71348 26188 71349 26228
rect 71307 26179 71349 26188
rect 71883 26228 71925 26237
rect 71883 26188 71884 26228
rect 71924 26188 71925 26228
rect 71883 26179 71925 26188
rect 39531 26104 39532 26144
rect 39572 26104 39573 26144
rect 39531 26095 39573 26104
rect 39619 26144 39677 26145
rect 39619 26104 39628 26144
rect 39668 26104 39677 26144
rect 39819 26137 39861 26146
rect 40099 26144 40157 26145
rect 39619 26103 39677 26104
rect 40003 26130 40061 26131
rect 40003 26090 40012 26130
rect 40052 26090 40061 26130
rect 40099 26104 40108 26144
rect 40148 26104 40157 26144
rect 40099 26103 40157 26104
rect 41155 26144 41213 26145
rect 41155 26104 41164 26144
rect 41204 26104 41213 26144
rect 41155 26103 41213 26104
rect 41259 26144 41301 26153
rect 41259 26104 41260 26144
rect 41300 26104 41301 26144
rect 41259 26095 41301 26104
rect 41451 26144 41493 26153
rect 41451 26104 41452 26144
rect 41492 26104 41493 26144
rect 41451 26095 41493 26104
rect 43659 26144 43701 26153
rect 43659 26104 43660 26144
rect 43700 26104 43701 26144
rect 43659 26095 43701 26104
rect 44035 26144 44093 26145
rect 44035 26104 44044 26144
rect 44084 26104 44093 26144
rect 44035 26103 44093 26104
rect 44899 26144 44957 26145
rect 44899 26104 44908 26144
rect 44948 26104 44957 26144
rect 44899 26103 44957 26104
rect 47211 26144 47253 26153
rect 47211 26104 47212 26144
rect 47252 26104 47253 26144
rect 47211 26095 47253 26104
rect 47971 26144 48029 26145
rect 47971 26104 47980 26144
rect 48020 26104 48029 26144
rect 47971 26103 48029 26104
rect 48171 26144 48213 26153
rect 48171 26104 48172 26144
rect 48212 26104 48213 26144
rect 48171 26095 48213 26104
rect 49123 26144 49181 26145
rect 49123 26104 49132 26144
rect 49172 26104 49181 26144
rect 49123 26103 49181 26104
rect 49987 26144 50045 26145
rect 49987 26104 49996 26144
rect 50036 26104 50045 26144
rect 49987 26103 50045 26104
rect 52003 26144 52061 26145
rect 52003 26104 52012 26144
rect 52052 26104 52061 26144
rect 52003 26103 52061 26104
rect 52203 26144 52245 26153
rect 52203 26104 52204 26144
rect 52244 26104 52245 26144
rect 52203 26095 52245 26104
rect 52387 26144 52445 26145
rect 52387 26104 52396 26144
rect 52436 26104 52445 26144
rect 52387 26103 52445 26104
rect 52587 26144 52629 26153
rect 52587 26104 52588 26144
rect 52628 26104 52629 26144
rect 52587 26095 52629 26104
rect 55459 26144 55517 26145
rect 55459 26104 55468 26144
rect 55508 26104 55517 26144
rect 55459 26103 55517 26104
rect 55755 26144 55797 26153
rect 55755 26104 55756 26144
rect 55796 26104 55797 26144
rect 55755 26095 55797 26104
rect 56331 26144 56373 26153
rect 56331 26104 56332 26144
rect 56372 26104 56373 26144
rect 56331 26095 56373 26104
rect 56523 26144 56565 26153
rect 56523 26104 56524 26144
rect 56564 26104 56565 26144
rect 56523 26095 56565 26104
rect 56611 26144 56669 26145
rect 56611 26104 56620 26144
rect 56660 26104 56669 26144
rect 56611 26103 56669 26104
rect 56811 26144 56853 26153
rect 56811 26104 56812 26144
rect 56852 26104 56853 26144
rect 56811 26095 56853 26104
rect 57003 26144 57045 26153
rect 57003 26104 57004 26144
rect 57044 26104 57045 26144
rect 57003 26095 57045 26104
rect 57091 26144 57149 26145
rect 57091 26104 57100 26144
rect 57140 26104 57149 26144
rect 57091 26103 57149 26104
rect 58347 26144 58389 26153
rect 58347 26104 58348 26144
rect 58388 26104 58389 26144
rect 58347 26095 58389 26104
rect 58539 26144 58581 26153
rect 58539 26104 58540 26144
rect 58580 26104 58581 26144
rect 58539 26095 58581 26104
rect 58627 26144 58685 26145
rect 58627 26104 58636 26144
rect 58676 26104 58685 26144
rect 58627 26103 58685 26104
rect 58827 26144 58869 26153
rect 58827 26104 58828 26144
rect 58868 26104 58869 26144
rect 58827 26095 58869 26104
rect 59019 26144 59061 26153
rect 59019 26104 59020 26144
rect 59060 26104 59061 26144
rect 59019 26095 59061 26104
rect 59107 26144 59165 26145
rect 59107 26104 59116 26144
rect 59156 26104 59165 26144
rect 59107 26103 59165 26104
rect 59395 26144 59453 26145
rect 59395 26104 59404 26144
rect 59444 26104 59453 26144
rect 59395 26103 59453 26104
rect 59499 26144 59541 26153
rect 59499 26104 59500 26144
rect 59540 26104 59541 26144
rect 59499 26095 59541 26104
rect 59595 26144 59637 26153
rect 59595 26104 59596 26144
rect 59636 26104 59637 26144
rect 59595 26095 59637 26104
rect 59779 26144 59837 26145
rect 59779 26104 59788 26144
rect 59828 26104 59837 26144
rect 59779 26103 59837 26104
rect 59883 26144 59925 26153
rect 59883 26104 59884 26144
rect 59924 26104 59925 26144
rect 59883 26095 59925 26104
rect 60075 26144 60117 26153
rect 60075 26104 60076 26144
rect 60116 26104 60117 26144
rect 60075 26095 60117 26104
rect 61987 26144 62045 26145
rect 61987 26104 61996 26144
rect 62036 26104 62045 26144
rect 61987 26103 62045 26104
rect 62851 26144 62909 26145
rect 62851 26104 62860 26144
rect 62900 26104 62909 26144
rect 62851 26103 62909 26104
rect 64203 26144 64245 26153
rect 64203 26104 64204 26144
rect 64244 26104 64245 26144
rect 64203 26095 64245 26104
rect 64299 26144 64341 26153
rect 64299 26104 64300 26144
rect 64340 26104 64341 26144
rect 64299 26095 64341 26104
rect 64395 26144 64437 26153
rect 64395 26104 64396 26144
rect 64436 26104 64437 26144
rect 64395 26095 64437 26104
rect 64491 26144 64533 26153
rect 64491 26104 64492 26144
rect 64532 26104 64533 26144
rect 64875 26144 64917 26153
rect 64491 26095 64533 26104
rect 64683 26133 64725 26142
rect 40003 26089 40061 26090
rect 64683 26093 64684 26133
rect 64724 26093 64725 26133
rect 64875 26104 64876 26144
rect 64916 26104 64917 26144
rect 64875 26095 64917 26104
rect 64963 26144 65021 26145
rect 64963 26104 64972 26144
rect 65012 26104 65021 26144
rect 64963 26103 65021 26104
rect 65451 26144 65493 26153
rect 65451 26104 65452 26144
rect 65492 26104 65493 26144
rect 65451 26095 65493 26104
rect 65643 26144 65685 26153
rect 65643 26104 65644 26144
rect 65684 26104 65685 26144
rect 65643 26095 65685 26104
rect 65731 26144 65789 26145
rect 65731 26104 65740 26144
rect 65780 26104 65789 26144
rect 65731 26103 65789 26104
rect 67179 26144 67221 26153
rect 67179 26104 67180 26144
rect 67220 26104 67221 26144
rect 67179 26095 67221 26104
rect 67275 26144 67317 26153
rect 67275 26104 67276 26144
rect 67316 26104 67317 26144
rect 67275 26095 67317 26104
rect 67371 26144 67413 26153
rect 67371 26104 67372 26144
rect 67412 26104 67413 26144
rect 67371 26095 67413 26104
rect 67467 26144 67509 26153
rect 67467 26104 67468 26144
rect 67508 26104 67509 26144
rect 67467 26095 67509 26104
rect 67659 26144 67701 26153
rect 67659 26104 67660 26144
rect 67700 26104 67701 26144
rect 67659 26095 67701 26104
rect 67851 26144 67893 26153
rect 67851 26104 67852 26144
rect 67892 26104 67893 26144
rect 67851 26095 67893 26104
rect 67939 26144 67997 26145
rect 67939 26104 67948 26144
rect 67988 26104 67997 26144
rect 67939 26103 67997 26104
rect 68131 26144 68189 26145
rect 68131 26104 68140 26144
rect 68180 26104 68189 26144
rect 68131 26103 68189 26104
rect 68331 26144 68373 26153
rect 68331 26104 68332 26144
rect 68372 26104 68373 26144
rect 68331 26095 68373 26104
rect 69291 26144 69333 26153
rect 69291 26104 69292 26144
rect 69332 26104 69333 26144
rect 69291 26095 69333 26104
rect 69387 26144 69429 26153
rect 69387 26104 69388 26144
rect 69428 26104 69429 26144
rect 69387 26095 69429 26104
rect 69483 26144 69525 26153
rect 69483 26104 69484 26144
rect 69524 26104 69525 26144
rect 69483 26095 69525 26104
rect 70915 26144 70973 26145
rect 70915 26104 70924 26144
rect 70964 26104 70973 26144
rect 70915 26103 70973 26104
rect 71211 26144 71253 26153
rect 71211 26104 71212 26144
rect 71252 26104 71253 26144
rect 71211 26095 71253 26104
rect 71787 26144 71829 26153
rect 71787 26104 71788 26144
rect 71828 26104 71829 26144
rect 71787 26095 71829 26104
rect 71971 26144 72029 26145
rect 71971 26104 71980 26144
rect 72020 26104 72029 26144
rect 71971 26103 72029 26104
rect 74179 26144 74237 26145
rect 74179 26104 74188 26144
rect 74228 26104 74237 26144
rect 74179 26103 74237 26104
rect 74283 26144 74325 26153
rect 74283 26104 74284 26144
rect 74324 26104 74325 26144
rect 74283 26095 74325 26104
rect 74475 26144 74517 26153
rect 74475 26104 74476 26144
rect 74516 26104 74517 26144
rect 74475 26095 74517 26104
rect 74667 26144 74709 26153
rect 74667 26104 74668 26144
rect 74708 26104 74709 26144
rect 74667 26095 74709 26104
rect 74763 26144 74805 26153
rect 74763 26104 74764 26144
rect 74804 26104 74805 26144
rect 74763 26095 74805 26104
rect 74859 26144 74901 26153
rect 74859 26104 74860 26144
rect 74900 26104 74901 26144
rect 74859 26095 74901 26104
rect 74955 26144 74997 26153
rect 74955 26104 74956 26144
rect 74996 26104 74997 26144
rect 74955 26095 74997 26104
rect 75147 26144 75189 26153
rect 75147 26104 75148 26144
rect 75188 26104 75189 26144
rect 75147 26095 75189 26104
rect 75339 26144 75381 26153
rect 75339 26104 75340 26144
rect 75380 26104 75381 26144
rect 75339 26095 75381 26104
rect 75427 26144 75485 26145
rect 75427 26104 75436 26144
rect 75476 26104 75485 26144
rect 75427 26103 75485 26104
rect 76875 26144 76917 26153
rect 76875 26104 76876 26144
rect 76916 26104 76917 26144
rect 76875 26095 76917 26104
rect 77067 26144 77109 26153
rect 77067 26104 77068 26144
rect 77108 26104 77109 26144
rect 77067 26095 77109 26104
rect 77155 26144 77213 26145
rect 77155 26104 77164 26144
rect 77204 26104 77213 26144
rect 77155 26103 77213 26104
rect 64683 26084 64725 26093
rect 643 26060 701 26061
rect 643 26020 652 26060
rect 692 26020 701 26060
rect 643 26019 701 26020
rect 38947 26060 39005 26061
rect 38947 26020 38956 26060
rect 38996 26020 39005 26060
rect 38947 26019 39005 26020
rect 40483 26060 40541 26061
rect 40483 26020 40492 26060
rect 40532 26020 40541 26060
rect 40483 26019 40541 26020
rect 48075 26060 48117 26069
rect 48075 26020 48076 26060
rect 48116 26020 48117 26060
rect 48075 26011 48117 26020
rect 51523 26060 51581 26061
rect 51523 26020 51532 26060
rect 51572 26020 51581 26060
rect 51523 26019 51581 26020
rect 57475 26060 57533 26061
rect 57475 26020 57484 26060
rect 57524 26020 57533 26060
rect 57475 26019 57533 26020
rect 60259 26060 60317 26061
rect 60259 26020 60268 26060
rect 60308 26020 60317 26060
rect 60259 26019 60317 26020
rect 60643 26060 60701 26061
rect 60643 26020 60652 26060
rect 60692 26020 60701 26060
rect 60643 26019 60701 26020
rect 61027 26060 61085 26061
rect 61027 26020 61036 26060
rect 61076 26020 61085 26060
rect 61027 26019 61085 26020
rect 68803 26060 68861 26061
rect 68803 26020 68812 26060
rect 68852 26020 68861 26060
rect 68803 26019 68861 26020
rect 70435 26060 70493 26061
rect 70435 26020 70444 26060
rect 70484 26020 70493 26060
rect 70435 26019 70493 26020
rect 843 25976 885 25985
rect 843 25936 844 25976
rect 884 25936 885 25976
rect 843 25927 885 25936
rect 32227 25976 32285 25977
rect 32227 25936 32236 25976
rect 32276 25936 32285 25976
rect 32227 25935 32285 25936
rect 35587 25976 35645 25977
rect 35587 25936 35596 25976
rect 35636 25936 35645 25976
rect 35587 25935 35645 25936
rect 39819 25976 39861 25985
rect 39819 25936 39820 25976
rect 39860 25936 39861 25976
rect 39819 25927 39861 25936
rect 40683 25976 40725 25985
rect 40683 25936 40684 25976
rect 40724 25936 40725 25976
rect 40683 25927 40725 25936
rect 41451 25976 41493 25985
rect 41451 25936 41452 25976
rect 41492 25936 41493 25976
rect 41451 25927 41493 25936
rect 42123 25976 42165 25985
rect 42123 25936 42124 25976
rect 42164 25936 42165 25976
rect 42123 25927 42165 25936
rect 47019 25976 47061 25985
rect 47019 25936 47020 25976
rect 47060 25936 47061 25976
rect 47019 25927 47061 25936
rect 47595 25976 47637 25985
rect 47595 25936 47596 25976
rect 47636 25936 47637 25976
rect 47595 25927 47637 25936
rect 48555 25976 48597 25985
rect 48555 25936 48556 25976
rect 48596 25936 48597 25976
rect 48555 25927 48597 25936
rect 51723 25976 51765 25985
rect 51723 25936 51724 25976
rect 51764 25936 51765 25976
rect 51723 25927 51765 25936
rect 52779 25976 52821 25985
rect 52779 25936 52780 25976
rect 52820 25936 52821 25976
rect 52779 25927 52821 25936
rect 54891 25976 54933 25985
rect 54891 25936 54892 25976
rect 54932 25936 54933 25976
rect 54891 25927 54933 25936
rect 56811 25976 56853 25985
rect 56811 25936 56812 25976
rect 56852 25936 56853 25976
rect 56811 25927 56853 25936
rect 57867 25976 57909 25985
rect 57867 25936 57868 25976
rect 57908 25936 57909 25976
rect 57867 25927 57909 25936
rect 58347 25976 58389 25985
rect 58347 25936 58348 25976
rect 58388 25936 58389 25976
rect 58347 25927 58389 25936
rect 58827 25976 58869 25985
rect 58827 25936 58828 25976
rect 58868 25936 58869 25976
rect 58827 25927 58869 25936
rect 60459 25976 60501 25985
rect 60459 25936 60460 25976
rect 60500 25936 60501 25976
rect 60459 25927 60501 25936
rect 60843 25976 60885 25985
rect 60843 25936 60844 25976
rect 60884 25936 60885 25976
rect 60843 25927 60885 25936
rect 65451 25976 65493 25985
rect 65451 25936 65452 25976
rect 65492 25936 65493 25976
rect 65451 25927 65493 25936
rect 66411 25976 66453 25985
rect 66411 25936 66412 25976
rect 66452 25936 66453 25976
rect 66411 25927 66453 25936
rect 68619 25976 68661 25985
rect 68619 25936 68620 25976
rect 68660 25936 68661 25976
rect 68619 25927 68661 25936
rect 71587 25976 71645 25977
rect 71587 25936 71596 25976
rect 71636 25936 71645 25976
rect 74475 25976 74517 25985
rect 71587 25935 71645 25936
rect 73419 25934 73461 25943
rect 39147 25892 39189 25901
rect 39147 25852 39148 25892
rect 39188 25852 39189 25892
rect 39147 25843 39189 25852
rect 39339 25892 39381 25901
rect 39339 25852 39340 25892
rect 39380 25852 39381 25892
rect 39339 25843 39381 25852
rect 46051 25892 46109 25893
rect 46051 25852 46060 25892
rect 46100 25852 46109 25892
rect 46051 25851 46109 25852
rect 51139 25892 51197 25893
rect 51139 25852 51148 25892
rect 51188 25852 51197 25892
rect 51139 25851 51197 25852
rect 52491 25892 52533 25901
rect 52491 25852 52492 25892
rect 52532 25852 52533 25892
rect 52491 25843 52533 25852
rect 56131 25892 56189 25893
rect 56131 25852 56140 25892
rect 56180 25852 56189 25892
rect 56131 25851 56189 25852
rect 60075 25892 60117 25901
rect 60075 25852 60076 25892
rect 60116 25852 60117 25892
rect 60075 25843 60117 25852
rect 64003 25892 64061 25893
rect 64003 25852 64012 25892
rect 64052 25852 64061 25892
rect 64003 25851 64061 25852
rect 68235 25892 68277 25901
rect 68235 25852 68236 25892
rect 68276 25852 68277 25892
rect 68235 25843 68277 25852
rect 70635 25892 70677 25901
rect 70635 25852 70636 25892
rect 70676 25852 70677 25892
rect 73419 25894 73420 25934
rect 73460 25894 73461 25934
rect 74475 25936 74476 25976
rect 74516 25936 74517 25976
rect 74475 25927 74517 25936
rect 73419 25885 73461 25894
rect 70635 25843 70677 25852
rect 576 25724 79584 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79584 25724
rect 576 25660 79584 25684
rect 34923 25556 34965 25565
rect 34923 25516 34924 25556
rect 34964 25516 34965 25556
rect 34923 25507 34965 25516
rect 40395 25556 40437 25565
rect 40395 25516 40396 25556
rect 40436 25516 40437 25556
rect 40395 25507 40437 25516
rect 45099 25556 45141 25565
rect 45099 25516 45100 25556
rect 45140 25516 45141 25556
rect 45099 25507 45141 25516
rect 46819 25556 46877 25557
rect 46819 25516 46828 25556
rect 46868 25516 46877 25556
rect 46819 25515 46877 25516
rect 52099 25556 52157 25557
rect 52099 25516 52108 25556
rect 52148 25516 52157 25556
rect 52099 25515 52157 25516
rect 56235 25556 56277 25565
rect 56235 25516 56236 25556
rect 56276 25516 56277 25556
rect 56235 25507 56277 25516
rect 67747 25556 67805 25557
rect 67747 25516 67756 25556
rect 67796 25516 67805 25556
rect 67747 25515 67805 25516
rect 75619 25556 75677 25557
rect 75619 25516 75628 25556
rect 75668 25516 75677 25556
rect 75619 25515 75677 25516
rect 75915 25556 75957 25565
rect 75915 25516 75916 25556
rect 75956 25516 75957 25556
rect 75915 25507 75957 25516
rect 35691 25472 35733 25481
rect 35691 25432 35692 25472
rect 35732 25432 35733 25472
rect 35691 25423 35733 25432
rect 44139 25472 44181 25481
rect 44139 25432 44140 25472
rect 44180 25432 44181 25472
rect 44139 25423 44181 25432
rect 55755 25472 55797 25481
rect 55755 25432 55756 25472
rect 55796 25432 55797 25472
rect 55755 25423 55797 25432
rect 63811 25472 63869 25473
rect 63811 25432 63820 25472
rect 63860 25432 63869 25472
rect 63811 25431 63869 25432
rect 76491 25472 76533 25481
rect 76491 25432 76492 25472
rect 76532 25432 76533 25472
rect 76491 25423 76533 25432
rect 643 25388 701 25389
rect 54699 25388 54741 25397
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 40579 25387 40637 25388
rect 40579 25347 40588 25387
rect 40628 25347 40637 25387
rect 40579 25346 40637 25347
rect 54699 25348 54700 25388
rect 54740 25348 54741 25388
rect 54699 25339 54741 25348
rect 76004 25319 76046 25328
rect 30115 25304 30173 25305
rect 30115 25264 30124 25304
rect 30164 25264 30173 25304
rect 30115 25263 30173 25264
rect 30979 25304 31037 25305
rect 30979 25264 30988 25304
rect 31028 25264 31037 25304
rect 30979 25263 31037 25264
rect 32803 25304 32861 25305
rect 32803 25264 32812 25304
rect 32852 25264 32861 25304
rect 33291 25304 33333 25313
rect 32803 25263 32861 25264
rect 33099 25262 33141 25271
rect 29739 25220 29781 25229
rect 29739 25180 29740 25220
rect 29780 25180 29781 25220
rect 33099 25222 33100 25262
rect 33140 25222 33141 25262
rect 33291 25264 33292 25304
rect 33332 25264 33333 25304
rect 33291 25255 33333 25264
rect 33379 25304 33437 25305
rect 33379 25264 33388 25304
rect 33428 25264 33437 25304
rect 33379 25263 33437 25264
rect 34443 25304 34485 25313
rect 34443 25264 34444 25304
rect 34484 25264 34485 25304
rect 34443 25255 34485 25264
rect 34539 25304 34581 25313
rect 34539 25264 34540 25304
rect 34580 25264 34581 25304
rect 34539 25255 34581 25264
rect 34635 25304 34677 25313
rect 34635 25264 34636 25304
rect 34676 25264 34677 25304
rect 34635 25255 34677 25264
rect 34731 25304 34773 25313
rect 34731 25264 34732 25304
rect 34772 25264 34773 25304
rect 34731 25255 34773 25264
rect 34923 25304 34965 25313
rect 34923 25264 34924 25304
rect 34964 25264 34965 25304
rect 34923 25255 34965 25264
rect 35115 25304 35157 25313
rect 35115 25264 35116 25304
rect 35156 25264 35157 25304
rect 35115 25255 35157 25264
rect 35203 25304 35261 25305
rect 35203 25264 35212 25304
rect 35252 25264 35261 25304
rect 35203 25263 35261 25264
rect 35691 25304 35733 25313
rect 35691 25264 35692 25304
rect 35732 25264 35733 25304
rect 35691 25255 35733 25264
rect 35883 25304 35925 25313
rect 35883 25264 35884 25304
rect 35924 25264 35925 25304
rect 35883 25255 35925 25264
rect 35971 25304 36029 25305
rect 35971 25264 35980 25304
rect 36020 25264 36029 25304
rect 35971 25263 36029 25264
rect 37227 25304 37269 25313
rect 37227 25264 37228 25304
rect 37268 25264 37269 25304
rect 37227 25255 37269 25264
rect 37603 25304 37661 25305
rect 37603 25264 37612 25304
rect 37652 25264 37661 25304
rect 37603 25263 37661 25264
rect 38467 25304 38525 25305
rect 38467 25264 38476 25304
rect 38516 25264 38525 25304
rect 38467 25263 38525 25264
rect 39819 25304 39861 25313
rect 39819 25264 39820 25304
rect 39860 25264 39861 25304
rect 39819 25255 39861 25264
rect 39915 25304 39957 25313
rect 39915 25264 39916 25304
rect 39956 25264 39957 25304
rect 39915 25255 39957 25264
rect 40011 25304 40053 25313
rect 40011 25264 40012 25304
rect 40052 25264 40053 25304
rect 40011 25255 40053 25264
rect 40107 25304 40149 25313
rect 40107 25264 40108 25304
rect 40148 25264 40149 25304
rect 40107 25255 40149 25264
rect 41251 25304 41309 25305
rect 41251 25264 41260 25304
rect 41300 25264 41309 25304
rect 41251 25263 41309 25264
rect 42115 25304 42173 25305
rect 42115 25264 42124 25304
rect 42164 25264 42173 25304
rect 42115 25263 42173 25264
rect 44803 25304 44861 25305
rect 44803 25264 44812 25304
rect 44852 25264 44861 25304
rect 44803 25263 44861 25264
rect 44907 25304 44949 25313
rect 44907 25264 44908 25304
rect 44948 25264 44949 25304
rect 44907 25255 44949 25264
rect 45099 25304 45141 25313
rect 45099 25264 45100 25304
rect 45140 25264 45141 25304
rect 45099 25255 45141 25264
rect 45291 25304 45333 25313
rect 45291 25264 45292 25304
rect 45332 25264 45333 25304
rect 45291 25255 45333 25264
rect 45387 25304 45429 25313
rect 45387 25264 45388 25304
rect 45428 25264 45429 25304
rect 45387 25255 45429 25264
rect 45483 25304 45525 25313
rect 45483 25264 45484 25304
rect 45524 25264 45525 25304
rect 45483 25255 45525 25264
rect 45579 25304 45621 25313
rect 45579 25264 45580 25304
rect 45620 25264 45621 25304
rect 45579 25255 45621 25264
rect 45763 25304 45821 25305
rect 45763 25264 45772 25304
rect 45812 25264 45821 25304
rect 45763 25263 45821 25264
rect 46147 25304 46205 25305
rect 46147 25264 46156 25304
rect 46196 25264 46205 25304
rect 46147 25263 46205 25264
rect 46443 25304 46485 25313
rect 46443 25264 46444 25304
rect 46484 25264 46485 25304
rect 46443 25255 46485 25264
rect 46539 25304 46581 25313
rect 46539 25264 46540 25304
rect 46580 25264 46581 25304
rect 46539 25255 46581 25264
rect 47395 25304 47453 25305
rect 47395 25264 47404 25304
rect 47444 25264 47453 25304
rect 47395 25263 47453 25264
rect 48259 25304 48317 25305
rect 48259 25264 48268 25304
rect 48308 25264 48317 25304
rect 48259 25263 48317 25264
rect 50571 25304 50613 25313
rect 50571 25264 50572 25304
rect 50612 25264 50613 25304
rect 50571 25255 50613 25264
rect 50667 25304 50709 25313
rect 50667 25264 50668 25304
rect 50708 25264 50709 25304
rect 50667 25255 50709 25264
rect 50763 25304 50805 25313
rect 50763 25264 50764 25304
rect 50804 25264 50805 25304
rect 50763 25255 50805 25264
rect 50859 25304 50901 25313
rect 50859 25264 50860 25304
rect 50900 25264 50901 25304
rect 50859 25255 50901 25264
rect 51427 25304 51485 25305
rect 51427 25264 51436 25304
rect 51476 25264 51485 25304
rect 51427 25263 51485 25264
rect 51723 25304 51765 25313
rect 51723 25264 51724 25304
rect 51764 25264 51765 25304
rect 51723 25255 51765 25264
rect 52675 25304 52733 25305
rect 52675 25264 52684 25304
rect 52724 25264 52733 25304
rect 52675 25263 52733 25264
rect 53539 25304 53597 25305
rect 53539 25264 53548 25304
rect 53588 25264 53597 25304
rect 53539 25263 53597 25264
rect 55275 25304 55317 25313
rect 55275 25264 55276 25304
rect 55316 25264 55317 25304
rect 55275 25255 55317 25264
rect 55467 25304 55509 25313
rect 55467 25264 55468 25304
rect 55508 25264 55509 25304
rect 55467 25255 55509 25264
rect 55555 25304 55613 25305
rect 55555 25264 55564 25304
rect 55604 25264 55613 25304
rect 55555 25263 55613 25264
rect 56139 25304 56181 25313
rect 56139 25264 56140 25304
rect 56180 25264 56181 25304
rect 56139 25255 56181 25264
rect 56323 25304 56381 25305
rect 56323 25264 56332 25304
rect 56372 25264 56381 25304
rect 56323 25263 56381 25264
rect 57387 25304 57429 25313
rect 57387 25264 57388 25304
rect 57428 25264 57429 25304
rect 57387 25255 57429 25264
rect 57763 25304 57821 25305
rect 57763 25264 57772 25304
rect 57812 25264 57821 25304
rect 57763 25263 57821 25264
rect 58627 25304 58685 25305
rect 58627 25264 58636 25304
rect 58676 25264 58685 25304
rect 58627 25263 58685 25264
rect 60267 25304 60309 25313
rect 60267 25264 60268 25304
rect 60308 25264 60309 25304
rect 60267 25255 60309 25264
rect 60643 25304 60701 25305
rect 60643 25264 60652 25304
rect 60692 25264 60701 25304
rect 60643 25263 60701 25264
rect 61507 25304 61565 25305
rect 61507 25264 61516 25304
rect 61556 25264 61565 25304
rect 61507 25263 61565 25264
rect 63139 25304 63197 25305
rect 63139 25264 63148 25304
rect 63188 25264 63197 25304
rect 63139 25263 63197 25264
rect 63435 25304 63477 25313
rect 63435 25264 63436 25304
rect 63476 25264 63477 25304
rect 63435 25255 63477 25264
rect 63531 25304 63573 25313
rect 63531 25264 63532 25304
rect 63572 25264 63573 25304
rect 63531 25255 63573 25264
rect 64387 25304 64445 25305
rect 64387 25264 64396 25304
rect 64436 25264 64445 25304
rect 64387 25263 64445 25264
rect 65251 25304 65309 25305
rect 65251 25264 65260 25304
rect 65300 25264 65309 25304
rect 65251 25263 65309 25264
rect 67075 25304 67133 25305
rect 67075 25264 67084 25304
rect 67124 25264 67133 25304
rect 67075 25263 67133 25264
rect 67371 25304 67413 25313
rect 67371 25264 67372 25304
rect 67412 25264 67413 25304
rect 67371 25255 67413 25264
rect 67467 25304 67509 25313
rect 67467 25264 67468 25304
rect 67508 25264 67509 25304
rect 67467 25255 67509 25264
rect 68323 25304 68381 25305
rect 68323 25264 68332 25304
rect 68372 25264 68381 25304
rect 68323 25263 68381 25264
rect 69187 25304 69245 25305
rect 69187 25264 69196 25304
rect 69236 25264 69245 25304
rect 69187 25263 69245 25264
rect 71011 25304 71069 25305
rect 71011 25264 71020 25304
rect 71060 25264 71069 25304
rect 71011 25263 71069 25264
rect 71875 25304 71933 25305
rect 71875 25264 71884 25304
rect 71924 25264 71933 25304
rect 71875 25263 71933 25264
rect 73227 25304 73269 25313
rect 73227 25264 73228 25304
rect 73268 25264 73269 25304
rect 73227 25255 73269 25264
rect 73603 25304 73661 25305
rect 73603 25264 73612 25304
rect 73652 25264 73661 25304
rect 73603 25263 73661 25264
rect 74467 25304 74525 25305
rect 74467 25264 74476 25304
rect 74516 25264 74525 25304
rect 74467 25263 74525 25264
rect 75811 25304 75869 25305
rect 75811 25264 75820 25304
rect 75860 25264 75869 25304
rect 76004 25279 76005 25319
rect 76045 25279 76046 25319
rect 76004 25270 76046 25279
rect 76195 25304 76253 25305
rect 75811 25263 75869 25264
rect 76195 25264 76204 25304
rect 76244 25264 76253 25304
rect 76195 25263 76253 25264
rect 76299 25304 76341 25313
rect 76299 25264 76300 25304
rect 76340 25264 76341 25304
rect 76299 25255 76341 25264
rect 76491 25304 76533 25313
rect 76491 25264 76492 25304
rect 76532 25264 76533 25304
rect 76491 25255 76533 25264
rect 76683 25304 76725 25313
rect 76683 25264 76684 25304
rect 76724 25264 76725 25304
rect 76683 25255 76725 25264
rect 77059 25304 77117 25305
rect 77059 25264 77068 25304
rect 77108 25264 77117 25304
rect 77059 25263 77117 25264
rect 77923 25304 77981 25305
rect 77923 25264 77932 25304
rect 77972 25264 77981 25304
rect 77923 25263 77981 25264
rect 33099 25213 33141 25222
rect 40875 25220 40917 25229
rect 29739 25171 29781 25180
rect 40875 25180 40876 25220
rect 40916 25180 40917 25220
rect 40875 25171 40917 25180
rect 47019 25220 47061 25229
rect 47019 25180 47020 25220
rect 47060 25180 47061 25220
rect 47019 25171 47061 25180
rect 51819 25220 51861 25229
rect 51819 25180 51820 25220
rect 51860 25180 51861 25220
rect 51819 25171 51861 25180
rect 52299 25220 52341 25229
rect 52299 25180 52300 25220
rect 52340 25180 52341 25220
rect 52299 25171 52341 25180
rect 64011 25220 64053 25229
rect 64011 25180 64012 25220
rect 64052 25180 64053 25220
rect 64011 25171 64053 25180
rect 67947 25220 67989 25229
rect 67947 25180 67948 25220
rect 67988 25180 67989 25220
rect 67947 25171 67989 25180
rect 70635 25220 70677 25229
rect 70635 25180 70636 25220
rect 70676 25180 70677 25220
rect 70635 25171 70677 25180
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 32131 25136 32189 25137
rect 32131 25096 32140 25136
rect 32180 25096 32189 25136
rect 32131 25095 32189 25096
rect 33187 25136 33245 25137
rect 33187 25096 33196 25136
rect 33236 25096 33245 25136
rect 33187 25095 33245 25096
rect 39619 25136 39677 25137
rect 39619 25096 39628 25136
rect 39668 25096 39677 25136
rect 39619 25095 39677 25096
rect 43267 25136 43325 25137
rect 43267 25096 43276 25136
rect 43316 25096 43325 25136
rect 43267 25095 43325 25096
rect 49411 25136 49469 25137
rect 49411 25096 49420 25136
rect 49460 25096 49469 25136
rect 49411 25095 49469 25096
rect 55363 25136 55421 25137
rect 55363 25096 55372 25136
rect 55412 25096 55421 25136
rect 55363 25095 55421 25096
rect 59779 25136 59837 25137
rect 59779 25096 59788 25136
rect 59828 25096 59837 25136
rect 59779 25095 59837 25096
rect 62659 25136 62717 25137
rect 62659 25096 62668 25136
rect 62708 25096 62717 25136
rect 62659 25095 62717 25096
rect 66403 25136 66461 25137
rect 66403 25096 66412 25136
rect 66452 25096 66461 25136
rect 66403 25095 66461 25096
rect 70339 25136 70397 25137
rect 70339 25096 70348 25136
rect 70388 25096 70397 25136
rect 70339 25095 70397 25096
rect 73027 25136 73085 25137
rect 73027 25096 73036 25136
rect 73076 25096 73085 25136
rect 73027 25095 73085 25096
rect 75619 25136 75677 25137
rect 75619 25096 75628 25136
rect 75668 25096 75677 25136
rect 75619 25095 75677 25096
rect 79075 25136 79133 25137
rect 79075 25096 79084 25136
rect 79124 25096 79133 25136
rect 79075 25095 79133 25096
rect 576 24968 79584 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79584 24968
rect 576 24904 79584 24928
rect 32227 24800 32285 24801
rect 32227 24760 32236 24800
rect 32276 24760 32285 24800
rect 32227 24759 32285 24760
rect 39147 24800 39189 24809
rect 39147 24760 39148 24800
rect 39188 24760 39189 24800
rect 39147 24751 39189 24760
rect 40579 24800 40637 24801
rect 40579 24760 40588 24800
rect 40628 24760 40637 24800
rect 40579 24759 40637 24760
rect 44995 24800 45053 24801
rect 44995 24760 45004 24800
rect 45044 24760 45053 24800
rect 44995 24759 45053 24760
rect 46819 24800 46877 24801
rect 46819 24760 46828 24800
rect 46868 24760 46877 24800
rect 46819 24759 46877 24760
rect 50187 24800 50229 24809
rect 50187 24760 50188 24800
rect 50228 24760 50229 24800
rect 50187 24751 50229 24760
rect 51435 24800 51477 24809
rect 51435 24760 51436 24800
rect 51476 24760 51477 24800
rect 51435 24751 51477 24760
rect 52195 24800 52253 24801
rect 52195 24760 52204 24800
rect 52244 24760 52253 24800
rect 52195 24759 52253 24760
rect 58339 24800 58397 24801
rect 58339 24760 58348 24800
rect 58388 24760 58397 24800
rect 58339 24759 58397 24760
rect 59019 24800 59061 24809
rect 59019 24760 59020 24800
rect 59060 24760 59061 24800
rect 59019 24751 59061 24760
rect 64003 24800 64061 24801
rect 64003 24760 64012 24800
rect 64052 24760 64061 24800
rect 64003 24759 64061 24760
rect 67747 24800 67805 24801
rect 67747 24760 67756 24800
rect 67796 24760 67805 24800
rect 67747 24759 67805 24760
rect 74371 24800 74429 24801
rect 74371 24760 74380 24800
rect 74420 24760 74429 24800
rect 74371 24759 74429 24760
rect 34923 24716 34965 24725
rect 34923 24676 34924 24716
rect 34964 24676 34965 24716
rect 34923 24667 34965 24676
rect 40011 24716 40053 24725
rect 40011 24676 40012 24716
rect 40052 24676 40053 24716
rect 40011 24667 40053 24676
rect 54891 24716 54933 24725
rect 54891 24676 54892 24716
rect 54932 24676 54933 24716
rect 54891 24667 54933 24676
rect 59499 24716 59541 24725
rect 59499 24676 59500 24716
rect 59540 24676 59541 24716
rect 59499 24667 59541 24676
rect 60267 24716 60309 24725
rect 60267 24676 60268 24716
rect 60308 24676 60309 24716
rect 60267 24667 60309 24676
rect 64491 24716 64533 24725
rect 64491 24676 64492 24716
rect 64532 24676 64533 24716
rect 64491 24667 64533 24676
rect 64875 24716 64917 24725
rect 64875 24676 64876 24716
rect 64916 24676 64917 24716
rect 64875 24667 64917 24676
rect 68235 24716 68277 24725
rect 68235 24676 68236 24716
rect 68276 24676 68277 24716
rect 68235 24667 68277 24676
rect 75819 24716 75861 24725
rect 75819 24676 75820 24716
rect 75860 24676 75861 24716
rect 75819 24667 75861 24676
rect 76491 24716 76533 24725
rect 76491 24676 76492 24716
rect 76532 24676 76533 24716
rect 76491 24667 76533 24676
rect 31659 24632 31701 24641
rect 31659 24592 31660 24632
rect 31700 24592 31701 24632
rect 31659 24583 31701 24592
rect 31755 24632 31797 24641
rect 31755 24592 31756 24632
rect 31796 24592 31797 24632
rect 31755 24583 31797 24592
rect 31851 24632 31893 24641
rect 31851 24592 31852 24632
rect 31892 24592 31893 24632
rect 31851 24583 31893 24592
rect 31947 24632 31989 24641
rect 31947 24592 31948 24632
rect 31988 24592 31989 24632
rect 31947 24583 31989 24592
rect 32139 24632 32181 24641
rect 32139 24592 32140 24632
rect 32180 24592 32181 24632
rect 32139 24583 32181 24592
rect 32331 24632 32373 24641
rect 32331 24592 32332 24632
rect 32372 24592 32373 24632
rect 32331 24583 32373 24592
rect 32419 24632 32477 24633
rect 32419 24592 32428 24632
rect 32468 24592 32477 24632
rect 32419 24591 32477 24592
rect 32715 24632 32757 24641
rect 32715 24592 32716 24632
rect 32756 24592 32757 24632
rect 32715 24583 32757 24592
rect 32899 24632 32957 24633
rect 32899 24592 32908 24632
rect 32948 24592 32957 24632
rect 32899 24591 32957 24592
rect 34147 24632 34205 24633
rect 34147 24592 34156 24632
rect 34196 24592 34205 24632
rect 34147 24591 34205 24592
rect 35299 24632 35357 24633
rect 35299 24592 35308 24632
rect 35348 24592 35357 24632
rect 35299 24591 35357 24592
rect 36163 24632 36221 24633
rect 36163 24592 36172 24632
rect 36212 24592 36221 24632
rect 36163 24591 36221 24592
rect 39619 24632 39677 24633
rect 39619 24592 39628 24632
rect 39668 24592 39677 24632
rect 39619 24591 39677 24592
rect 39915 24632 39957 24641
rect 39915 24592 39916 24632
rect 39956 24592 39957 24632
rect 39915 24583 39957 24592
rect 40491 24632 40533 24641
rect 40491 24592 40492 24632
rect 40532 24592 40533 24632
rect 40491 24583 40533 24592
rect 40683 24632 40725 24641
rect 40683 24592 40684 24632
rect 40724 24592 40725 24632
rect 40683 24583 40725 24592
rect 40771 24632 40829 24633
rect 40771 24592 40780 24632
rect 40820 24592 40829 24632
rect 40771 24591 40829 24592
rect 40963 24632 41021 24633
rect 40963 24592 40972 24632
rect 41012 24592 41021 24632
rect 40963 24591 41021 24592
rect 41163 24632 41205 24641
rect 41163 24592 41164 24632
rect 41204 24592 41205 24632
rect 41163 24583 41205 24592
rect 42315 24632 42357 24641
rect 42315 24592 42316 24632
rect 42356 24592 42357 24632
rect 42315 24583 42357 24592
rect 42691 24632 42749 24633
rect 42691 24592 42700 24632
rect 42740 24592 42749 24632
rect 42691 24591 42749 24592
rect 43555 24632 43613 24633
rect 43555 24592 43564 24632
rect 43604 24592 43613 24632
rect 43555 24591 43613 24592
rect 44907 24632 44949 24641
rect 44907 24592 44908 24632
rect 44948 24592 44949 24632
rect 44907 24583 44949 24592
rect 45099 24632 45141 24641
rect 45099 24592 45100 24632
rect 45140 24592 45141 24632
rect 45099 24583 45141 24592
rect 45187 24632 45245 24633
rect 45187 24592 45196 24632
rect 45236 24592 45245 24632
rect 45187 24591 45245 24592
rect 46731 24632 46773 24641
rect 46731 24592 46732 24632
rect 46772 24592 46773 24632
rect 46731 24583 46773 24592
rect 46923 24632 46965 24641
rect 46923 24592 46924 24632
rect 46964 24592 46965 24632
rect 46923 24583 46965 24592
rect 47011 24632 47069 24633
rect 47011 24592 47020 24632
rect 47060 24592 47069 24632
rect 47011 24591 47069 24592
rect 50379 24632 50421 24641
rect 50379 24592 50380 24632
rect 50420 24592 50421 24632
rect 50379 24583 50421 24592
rect 50571 24632 50613 24641
rect 50571 24592 50572 24632
rect 50612 24592 50613 24632
rect 50571 24583 50613 24592
rect 50659 24632 50717 24633
rect 50659 24592 50668 24632
rect 50708 24592 50717 24632
rect 50659 24591 50717 24592
rect 50851 24632 50909 24633
rect 50851 24592 50860 24632
rect 50900 24592 50909 24632
rect 50851 24591 50909 24592
rect 51051 24632 51093 24641
rect 51051 24592 51052 24632
rect 51092 24592 51093 24632
rect 51051 24583 51093 24592
rect 52107 24632 52149 24641
rect 52107 24592 52108 24632
rect 52148 24592 52149 24632
rect 52107 24583 52149 24592
rect 52299 24632 52341 24641
rect 52299 24592 52300 24632
rect 52340 24592 52341 24632
rect 52299 24583 52341 24592
rect 52387 24632 52445 24633
rect 52387 24592 52396 24632
rect 52436 24592 52445 24632
rect 52387 24591 52445 24592
rect 55267 24632 55325 24633
rect 55267 24592 55276 24632
rect 55316 24592 55325 24632
rect 55267 24591 55325 24592
rect 56131 24632 56189 24633
rect 56131 24592 56140 24632
rect 56180 24592 56189 24632
rect 56131 24591 56189 24592
rect 58059 24632 58101 24641
rect 58059 24592 58060 24632
rect 58100 24592 58101 24632
rect 58059 24583 58101 24592
rect 58155 24632 58197 24641
rect 58155 24592 58156 24632
rect 58196 24592 58197 24632
rect 58155 24583 58197 24592
rect 58251 24632 58293 24641
rect 58251 24592 58252 24632
rect 58292 24592 58293 24632
rect 58251 24583 58293 24592
rect 59595 24632 59637 24641
rect 59595 24592 59596 24632
rect 59636 24592 59637 24632
rect 59595 24583 59637 24592
rect 59875 24632 59933 24633
rect 59875 24592 59884 24632
rect 59924 24592 59933 24632
rect 59875 24591 59933 24592
rect 60163 24632 60221 24633
rect 60163 24592 60172 24632
rect 60212 24592 60221 24632
rect 60163 24591 60221 24592
rect 60363 24632 60405 24641
rect 60363 24592 60364 24632
rect 60404 24592 60405 24632
rect 60363 24583 60405 24592
rect 63915 24632 63957 24641
rect 63915 24592 63916 24632
rect 63956 24592 63957 24632
rect 63915 24583 63957 24592
rect 64107 24632 64149 24641
rect 64107 24592 64108 24632
rect 64148 24592 64149 24632
rect 64107 24583 64149 24592
rect 64195 24632 64253 24633
rect 64195 24592 64204 24632
rect 64244 24592 64253 24632
rect 64195 24591 64253 24592
rect 64387 24632 64445 24633
rect 64387 24592 64396 24632
rect 64436 24592 64445 24632
rect 64387 24591 64445 24592
rect 64587 24632 64629 24641
rect 64587 24592 64588 24632
rect 64628 24592 64629 24632
rect 64587 24583 64629 24592
rect 64779 24632 64821 24641
rect 64779 24592 64780 24632
rect 64820 24592 64821 24632
rect 64779 24583 64821 24592
rect 64963 24632 65021 24633
rect 64963 24592 64972 24632
rect 65012 24592 65021 24632
rect 64963 24591 65021 24592
rect 67659 24632 67701 24641
rect 67659 24592 67660 24632
rect 67700 24592 67701 24632
rect 67659 24583 67701 24592
rect 67851 24632 67893 24641
rect 67851 24592 67852 24632
rect 67892 24592 67893 24632
rect 67851 24583 67893 24592
rect 67939 24632 67997 24633
rect 67939 24592 67948 24632
rect 67988 24592 67997 24632
rect 67939 24591 67997 24592
rect 68131 24632 68189 24633
rect 68131 24592 68140 24632
rect 68180 24592 68189 24632
rect 68131 24591 68189 24592
rect 68331 24632 68373 24641
rect 68331 24592 68332 24632
rect 68372 24592 68373 24632
rect 68331 24583 68373 24592
rect 70731 24632 70773 24641
rect 70731 24592 70732 24632
rect 70772 24592 70773 24632
rect 70731 24583 70773 24592
rect 70923 24632 70965 24641
rect 70923 24592 70924 24632
rect 70964 24592 70965 24632
rect 70923 24583 70965 24592
rect 71011 24632 71069 24633
rect 71011 24592 71020 24632
rect 71060 24592 71069 24632
rect 71011 24591 71069 24592
rect 71203 24632 71261 24633
rect 71203 24592 71212 24632
rect 71252 24592 71261 24632
rect 71203 24591 71261 24592
rect 71307 24632 71349 24641
rect 71307 24592 71308 24632
rect 71348 24592 71349 24632
rect 71307 24583 71349 24592
rect 71403 24632 71445 24641
rect 71403 24592 71404 24632
rect 71444 24592 71445 24632
rect 71403 24583 71445 24592
rect 74283 24632 74325 24641
rect 74283 24592 74284 24632
rect 74324 24592 74325 24632
rect 74283 24583 74325 24592
rect 74475 24632 74517 24641
rect 74475 24592 74476 24632
rect 74516 24592 74517 24632
rect 74475 24583 74517 24592
rect 74563 24632 74621 24633
rect 74563 24592 74572 24632
rect 74612 24592 74621 24632
rect 74563 24591 74621 24592
rect 75427 24632 75485 24633
rect 75427 24592 75436 24632
rect 75476 24592 75485 24632
rect 75427 24591 75485 24592
rect 75723 24632 75765 24641
rect 75723 24592 75724 24632
rect 75764 24592 75765 24632
rect 75723 24583 75765 24592
rect 76387 24632 76445 24633
rect 76387 24592 76396 24632
rect 76436 24592 76445 24632
rect 76387 24591 76445 24592
rect 76587 24632 76629 24641
rect 76587 24592 76588 24632
rect 76628 24592 76629 24632
rect 76587 24583 76629 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 39331 24548 39389 24549
rect 39331 24508 39340 24548
rect 39380 24508 39389 24548
rect 39331 24507 39389 24508
rect 41067 24548 41109 24557
rect 41067 24508 41068 24548
rect 41108 24508 41109 24548
rect 41067 24499 41109 24508
rect 49987 24548 50045 24549
rect 49987 24508 49996 24548
rect 50036 24508 50045 24548
rect 49987 24507 50045 24508
rect 51235 24548 51293 24549
rect 51235 24508 51244 24548
rect 51284 24508 51293 24548
rect 51235 24507 51293 24508
rect 57291 24548 57333 24557
rect 57291 24508 57292 24548
rect 57332 24508 57333 24548
rect 57291 24499 57333 24508
rect 58819 24548 58877 24549
rect 58819 24508 58828 24548
rect 58868 24508 58877 24548
rect 58819 24507 58877 24508
rect 60739 24548 60797 24549
rect 60739 24508 60748 24548
rect 60788 24508 60797 24548
rect 60739 24507 60797 24508
rect 30219 24464 30261 24473
rect 30219 24424 30220 24464
rect 30260 24424 30261 24464
rect 30219 24415 30261 24424
rect 33867 24464 33909 24473
rect 33867 24424 33868 24464
rect 33908 24424 33909 24464
rect 33867 24415 33909 24424
rect 37707 24464 37749 24473
rect 37707 24424 37708 24464
rect 37748 24424 37749 24464
rect 37707 24415 37749 24424
rect 41355 24464 41397 24473
rect 41355 24424 41356 24464
rect 41396 24424 41397 24464
rect 41355 24415 41397 24424
rect 48555 24464 48597 24473
rect 48555 24424 48556 24464
rect 48596 24424 48597 24464
rect 48555 24415 48597 24424
rect 52587 24464 52629 24473
rect 52587 24424 52588 24464
rect 52628 24424 52629 24464
rect 52587 24415 52629 24424
rect 59203 24464 59261 24465
rect 59203 24424 59212 24464
rect 59252 24424 59261 24464
rect 59203 24423 59261 24424
rect 60939 24464 60981 24473
rect 60939 24424 60940 24464
rect 60980 24424 60981 24464
rect 60939 24415 60981 24424
rect 65163 24464 65205 24473
rect 65163 24424 65164 24464
rect 65204 24424 65205 24464
rect 65163 24415 65205 24424
rect 68523 24464 68565 24473
rect 68523 24424 68524 24464
rect 68564 24424 68565 24464
rect 68523 24415 68565 24424
rect 70731 24464 70773 24473
rect 70731 24424 70732 24464
rect 70772 24424 70773 24464
rect 70731 24415 70773 24424
rect 71595 24464 71637 24473
rect 71595 24424 71596 24464
rect 71636 24424 71637 24464
rect 71595 24415 71637 24424
rect 76099 24464 76157 24465
rect 76099 24424 76108 24464
rect 76148 24424 76157 24464
rect 76099 24423 76157 24424
rect 77163 24464 77205 24473
rect 77163 24424 77164 24464
rect 77204 24424 77205 24464
rect 77163 24415 77205 24424
rect 843 24380 885 24389
rect 843 24340 844 24380
rect 884 24340 885 24380
rect 843 24331 885 24340
rect 32811 24380 32853 24389
rect 32811 24340 32812 24380
rect 32852 24340 32853 24380
rect 32811 24331 32853 24340
rect 37315 24380 37373 24381
rect 37315 24340 37324 24380
rect 37364 24340 37373 24380
rect 37315 24339 37373 24340
rect 40291 24380 40349 24381
rect 40291 24340 40300 24380
rect 40340 24340 40349 24380
rect 40291 24339 40349 24340
rect 44707 24380 44765 24381
rect 44707 24340 44716 24380
rect 44756 24340 44765 24380
rect 44707 24339 44765 24340
rect 50187 24380 50229 24389
rect 50187 24340 50188 24380
rect 50228 24340 50229 24380
rect 50187 24331 50229 24340
rect 50379 24380 50421 24389
rect 50379 24340 50380 24380
rect 50420 24340 50421 24380
rect 50379 24331 50421 24340
rect 50955 24380 50997 24389
rect 50955 24340 50956 24380
rect 50996 24340 50997 24380
rect 50955 24331 50997 24340
rect 60555 24380 60597 24389
rect 60555 24340 60556 24380
rect 60596 24340 60597 24380
rect 60555 24331 60597 24340
rect 576 24212 79584 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 79584 24212
rect 576 24148 79584 24172
rect 36555 24044 36597 24053
rect 36555 24004 36556 24044
rect 36596 24004 36597 24044
rect 36555 23995 36597 24004
rect 40203 24044 40245 24053
rect 40203 24004 40204 24044
rect 40244 24004 40245 24044
rect 40203 23995 40245 24004
rect 41451 24044 41493 24053
rect 41451 24004 41452 24044
rect 41492 24004 41493 24044
rect 41451 23995 41493 24004
rect 44427 24044 44469 24053
rect 44427 24004 44428 24044
rect 44468 24004 44469 24044
rect 44427 23995 44469 24004
rect 55755 24044 55797 24053
rect 55755 24004 55756 24044
rect 55796 24004 55797 24044
rect 55755 23995 55797 24004
rect 28875 23960 28917 23969
rect 28875 23920 28876 23960
rect 28916 23920 28917 23960
rect 28875 23911 28917 23920
rect 32515 23960 32573 23961
rect 32515 23920 32524 23960
rect 32564 23920 32573 23960
rect 32515 23919 32573 23920
rect 35499 23960 35541 23969
rect 35499 23920 35500 23960
rect 35540 23920 35541 23960
rect 35499 23911 35541 23920
rect 40683 23960 40725 23969
rect 40683 23920 40684 23960
rect 40724 23920 40725 23960
rect 40683 23911 40725 23920
rect 42795 23960 42837 23969
rect 42795 23920 42796 23960
rect 42836 23920 42837 23960
rect 42795 23911 42837 23920
rect 45667 23960 45725 23961
rect 45667 23920 45676 23960
rect 45716 23920 45725 23960
rect 45667 23919 45725 23920
rect 46923 23960 46965 23969
rect 46923 23920 46924 23960
rect 46964 23920 46965 23960
rect 46923 23911 46965 23920
rect 51435 23960 51477 23969
rect 51435 23920 51436 23960
rect 51476 23920 51477 23960
rect 51435 23911 51477 23920
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 1795 23876 1853 23877
rect 1795 23836 1804 23876
rect 1844 23836 1853 23876
rect 1795 23835 1853 23836
rect 1987 23876 2045 23877
rect 1987 23836 1996 23876
rect 2036 23836 2045 23876
rect 1987 23835 2045 23836
rect 30883 23876 30941 23877
rect 30883 23836 30892 23876
rect 30932 23836 30941 23876
rect 30883 23835 30941 23836
rect 40483 23876 40541 23877
rect 40483 23836 40492 23876
rect 40532 23836 40541 23876
rect 40483 23835 40541 23836
rect 41251 23876 41309 23877
rect 41251 23836 41260 23876
rect 41300 23836 41309 23876
rect 41251 23835 41309 23836
rect 51235 23806 51293 23807
rect 31275 23792 31317 23801
rect 31275 23752 31276 23792
rect 31316 23752 31317 23792
rect 31275 23743 31317 23752
rect 31467 23792 31509 23801
rect 31467 23752 31468 23792
rect 31508 23752 31509 23792
rect 31467 23743 31509 23752
rect 31555 23792 31613 23793
rect 31555 23752 31564 23792
rect 31604 23752 31613 23792
rect 31555 23751 31613 23752
rect 31843 23792 31901 23793
rect 31843 23752 31852 23792
rect 31892 23752 31901 23792
rect 31843 23751 31901 23752
rect 32139 23792 32181 23801
rect 32139 23752 32140 23792
rect 32180 23752 32181 23792
rect 32139 23743 32181 23752
rect 32235 23792 32277 23801
rect 32235 23752 32236 23792
rect 32276 23752 32277 23792
rect 32235 23743 32277 23752
rect 33283 23792 33341 23793
rect 33283 23752 33292 23792
rect 33332 23752 33341 23792
rect 33283 23751 33341 23752
rect 34147 23792 34205 23793
rect 34147 23752 34156 23792
rect 34196 23752 34205 23792
rect 34147 23751 34205 23752
rect 36075 23792 36117 23801
rect 36075 23752 36076 23792
rect 36116 23752 36117 23792
rect 36075 23743 36117 23752
rect 36171 23792 36213 23801
rect 36171 23752 36172 23792
rect 36212 23752 36213 23792
rect 36171 23743 36213 23752
rect 36267 23792 36309 23801
rect 36267 23752 36268 23792
rect 36308 23752 36309 23792
rect 36267 23743 36309 23752
rect 36363 23792 36405 23801
rect 36363 23752 36364 23792
rect 36404 23752 36405 23792
rect 36363 23743 36405 23752
rect 36555 23792 36597 23801
rect 36555 23752 36556 23792
rect 36596 23752 36597 23792
rect 36555 23743 36597 23752
rect 36747 23792 36789 23801
rect 36747 23752 36748 23792
rect 36788 23752 36789 23792
rect 36747 23743 36789 23752
rect 36835 23792 36893 23793
rect 36835 23752 36844 23792
rect 36884 23752 36893 23792
rect 36835 23751 36893 23752
rect 38763 23792 38805 23801
rect 38763 23752 38764 23792
rect 38804 23752 38805 23792
rect 38763 23743 38805 23752
rect 38859 23792 38901 23801
rect 38859 23752 38860 23792
rect 38900 23752 38901 23792
rect 38859 23743 38901 23752
rect 38955 23792 38997 23801
rect 38955 23752 38956 23792
rect 38996 23752 38997 23792
rect 38955 23743 38997 23752
rect 39243 23792 39285 23801
rect 39243 23752 39244 23792
rect 39284 23752 39285 23792
rect 39243 23743 39285 23752
rect 39435 23792 39477 23801
rect 39435 23752 39436 23792
rect 39476 23752 39477 23792
rect 39435 23743 39477 23752
rect 39523 23792 39581 23793
rect 39523 23752 39532 23792
rect 39572 23752 39581 23792
rect 39523 23751 39581 23752
rect 40099 23792 40157 23793
rect 40099 23752 40108 23792
rect 40148 23752 40157 23792
rect 40099 23751 40157 23752
rect 40299 23792 40341 23801
rect 40299 23752 40300 23792
rect 40340 23752 40341 23792
rect 40299 23743 40341 23752
rect 40867 23792 40925 23793
rect 40867 23752 40876 23792
rect 40916 23752 40925 23792
rect 40867 23751 40925 23752
rect 41067 23792 41109 23801
rect 41067 23752 41068 23792
rect 41108 23752 41109 23792
rect 41067 23743 41109 23752
rect 44043 23792 44085 23801
rect 44043 23752 44044 23792
rect 44084 23752 44085 23792
rect 44043 23743 44085 23752
rect 44139 23792 44181 23801
rect 44139 23752 44140 23792
rect 44180 23752 44181 23792
rect 44139 23743 44181 23752
rect 44235 23792 44277 23801
rect 44235 23752 44236 23792
rect 44276 23752 44277 23792
rect 44235 23743 44277 23752
rect 44427 23792 44469 23801
rect 44427 23752 44428 23792
rect 44468 23752 44469 23792
rect 44427 23743 44469 23752
rect 44619 23792 44661 23801
rect 44619 23752 44620 23792
rect 44660 23752 44661 23792
rect 44619 23743 44661 23752
rect 44707 23792 44765 23793
rect 44707 23752 44716 23792
rect 44756 23752 44765 23792
rect 44707 23751 44765 23752
rect 44995 23792 45053 23793
rect 44995 23752 45004 23792
rect 45044 23752 45053 23792
rect 44995 23751 45053 23752
rect 45291 23792 45333 23801
rect 45291 23752 45292 23792
rect 45332 23752 45333 23792
rect 45291 23743 45333 23752
rect 45387 23792 45429 23801
rect 45387 23752 45388 23792
rect 45428 23752 45429 23792
rect 45387 23743 45429 23752
rect 45867 23792 45909 23801
rect 45867 23752 45868 23792
rect 45908 23752 45909 23792
rect 45867 23743 45909 23752
rect 45963 23792 46005 23801
rect 45963 23752 45964 23792
rect 46004 23752 46005 23792
rect 45963 23743 46005 23752
rect 46051 23792 46109 23793
rect 46051 23752 46060 23792
rect 46100 23752 46109 23792
rect 46051 23751 46109 23752
rect 48451 23792 48509 23793
rect 48451 23752 48460 23792
rect 48500 23752 48509 23792
rect 48451 23751 48509 23752
rect 49315 23792 49373 23793
rect 49315 23752 49324 23792
rect 49364 23752 49373 23792
rect 49315 23751 49373 23752
rect 50667 23792 50709 23801
rect 50667 23752 50668 23792
rect 50708 23752 50709 23792
rect 50667 23743 50709 23752
rect 50859 23792 50901 23801
rect 50859 23752 50860 23792
rect 50900 23752 50901 23792
rect 50859 23743 50901 23752
rect 50947 23792 51005 23793
rect 50947 23752 50956 23792
rect 50996 23752 51005 23792
rect 50947 23751 51005 23752
rect 51139 23792 51197 23793
rect 51139 23752 51148 23792
rect 51188 23752 51197 23792
rect 51235 23766 51244 23806
rect 51284 23766 51293 23806
rect 51235 23765 51293 23766
rect 51435 23792 51477 23801
rect 51139 23751 51197 23752
rect 51435 23752 51436 23792
rect 51476 23752 51477 23792
rect 51435 23743 51477 23752
rect 51723 23792 51765 23801
rect 51723 23752 51724 23792
rect 51764 23752 51765 23792
rect 51723 23743 51765 23752
rect 52099 23792 52157 23793
rect 52099 23752 52108 23792
rect 52148 23752 52157 23792
rect 52099 23751 52157 23752
rect 52963 23792 53021 23793
rect 52963 23752 52972 23792
rect 53012 23752 53021 23792
rect 52963 23751 53021 23752
rect 54787 23792 54845 23793
rect 54787 23752 54796 23792
rect 54836 23752 54845 23792
rect 54787 23751 54845 23752
rect 55171 23792 55229 23793
rect 55171 23752 55180 23792
rect 55220 23752 55229 23792
rect 55171 23751 55229 23752
rect 55651 23792 55709 23793
rect 55651 23752 55660 23792
rect 55700 23752 55709 23792
rect 55651 23751 55709 23752
rect 55851 23792 55893 23801
rect 55851 23752 55852 23792
rect 55892 23752 55893 23792
rect 55851 23743 55893 23752
rect 56131 23792 56189 23793
rect 56131 23752 56140 23792
rect 56180 23752 56189 23792
rect 56131 23751 56189 23752
rect 56419 23792 56477 23793
rect 56419 23752 56428 23792
rect 56468 23752 56477 23792
rect 56419 23751 56477 23752
rect 56611 23792 56669 23793
rect 56611 23752 56620 23792
rect 56660 23752 56669 23792
rect 56611 23751 56669 23752
rect 56899 23792 56957 23793
rect 56899 23752 56908 23792
rect 56948 23752 56957 23792
rect 56899 23751 56957 23752
rect 57283 23792 57341 23793
rect 57283 23752 57292 23792
rect 57332 23752 57341 23792
rect 57283 23751 57341 23752
rect 57667 23792 57725 23793
rect 57667 23752 57676 23792
rect 57716 23752 57725 23792
rect 57667 23751 57725 23752
rect 58051 23792 58109 23793
rect 58051 23752 58060 23792
rect 58100 23752 58109 23792
rect 58051 23751 58109 23752
rect 58435 23792 58493 23793
rect 58435 23752 58444 23792
rect 58484 23752 58493 23792
rect 58435 23751 58493 23752
rect 58819 23792 58877 23793
rect 58819 23752 58828 23792
rect 58868 23752 58877 23792
rect 58819 23751 58877 23752
rect 59299 23792 59357 23793
rect 59299 23752 59308 23792
rect 59348 23752 59357 23792
rect 59299 23751 59357 23752
rect 59683 23792 59741 23793
rect 59683 23752 59692 23792
rect 59732 23752 59741 23792
rect 59683 23751 59741 23752
rect 60067 23792 60125 23793
rect 60067 23752 60076 23792
rect 60116 23752 60125 23792
rect 60067 23751 60125 23752
rect 60451 23792 60509 23793
rect 60451 23752 60460 23792
rect 60500 23752 60509 23792
rect 60451 23751 60509 23752
rect 60835 23792 60893 23793
rect 60835 23752 60844 23792
rect 60884 23752 60893 23792
rect 60835 23751 60893 23752
rect 61315 23792 61373 23793
rect 61315 23752 61324 23792
rect 61364 23752 61373 23792
rect 61315 23751 61373 23752
rect 61699 23792 61757 23793
rect 61699 23752 61708 23792
rect 61748 23752 61757 23792
rect 61699 23751 61757 23752
rect 62083 23792 62141 23793
rect 62083 23752 62092 23792
rect 62132 23752 62141 23792
rect 62083 23751 62141 23752
rect 62467 23792 62525 23793
rect 62467 23752 62476 23792
rect 62516 23752 62525 23792
rect 62467 23751 62525 23752
rect 62851 23792 62909 23793
rect 62851 23752 62860 23792
rect 62900 23752 62909 23792
rect 62851 23751 62909 23752
rect 63235 23792 63293 23793
rect 63235 23752 63244 23792
rect 63284 23752 63293 23792
rect 63235 23751 63293 23752
rect 63619 23792 63677 23793
rect 63619 23752 63628 23792
rect 63668 23752 63677 23792
rect 63619 23751 63677 23752
rect 64099 23792 64157 23793
rect 64099 23752 64108 23792
rect 64148 23752 64157 23792
rect 64099 23751 64157 23752
rect 64483 23792 64541 23793
rect 64483 23752 64492 23792
rect 64532 23752 64541 23792
rect 64483 23751 64541 23752
rect 64867 23792 64925 23793
rect 64867 23752 64876 23792
rect 64916 23752 64925 23792
rect 64867 23751 64925 23752
rect 65251 23792 65309 23793
rect 65251 23752 65260 23792
rect 65300 23752 65309 23792
rect 65251 23751 65309 23752
rect 65731 23792 65789 23793
rect 65731 23752 65740 23792
rect 65780 23752 65789 23792
rect 65731 23751 65789 23752
rect 66115 23792 66173 23793
rect 66115 23752 66124 23792
rect 66164 23752 66173 23792
rect 66115 23751 66173 23752
rect 66499 23792 66557 23793
rect 66499 23752 66508 23792
rect 66548 23752 66557 23792
rect 66499 23751 66557 23752
rect 66883 23792 66941 23793
rect 66883 23752 66892 23792
rect 66932 23752 66941 23792
rect 66883 23751 66941 23752
rect 67267 23792 67325 23793
rect 67267 23752 67276 23792
rect 67316 23752 67325 23792
rect 67267 23751 67325 23752
rect 67651 23792 67709 23793
rect 67651 23752 67660 23792
rect 67700 23752 67709 23792
rect 67651 23751 67709 23752
rect 68131 23792 68189 23793
rect 68131 23752 68140 23792
rect 68180 23752 68189 23792
rect 68131 23751 68189 23752
rect 68515 23792 68573 23793
rect 68515 23752 68524 23792
rect 68564 23752 68573 23792
rect 68515 23751 68573 23752
rect 68899 23792 68957 23793
rect 68899 23752 68908 23792
rect 68948 23752 68957 23792
rect 68899 23751 68957 23752
rect 69283 23792 69341 23793
rect 69283 23752 69292 23792
rect 69332 23752 69341 23792
rect 69283 23751 69341 23752
rect 69667 23792 69725 23793
rect 69667 23752 69676 23792
rect 69716 23752 69725 23792
rect 69667 23751 69725 23752
rect 70147 23792 70205 23793
rect 70147 23752 70156 23792
rect 70196 23752 70205 23792
rect 70147 23751 70205 23752
rect 70531 23792 70589 23793
rect 70531 23752 70540 23792
rect 70580 23752 70589 23792
rect 70531 23751 70589 23752
rect 70915 23792 70973 23793
rect 70915 23752 70924 23792
rect 70964 23752 70973 23792
rect 70915 23751 70973 23752
rect 71299 23792 71357 23793
rect 71299 23752 71308 23792
rect 71348 23752 71357 23792
rect 71299 23751 71357 23752
rect 71683 23792 71741 23793
rect 71683 23752 71692 23792
rect 71732 23752 71741 23792
rect 71683 23751 71741 23752
rect 72067 23792 72125 23793
rect 72067 23752 72076 23792
rect 72116 23752 72125 23792
rect 72067 23751 72125 23752
rect 72451 23792 72509 23793
rect 72451 23752 72460 23792
rect 72500 23752 72509 23792
rect 72451 23751 72509 23752
rect 72835 23792 72893 23793
rect 72835 23752 72844 23792
rect 72884 23752 72893 23792
rect 72835 23751 72893 23752
rect 73315 23792 73373 23793
rect 73315 23752 73324 23792
rect 73364 23752 73373 23792
rect 73315 23751 73373 23752
rect 73699 23792 73757 23793
rect 73699 23752 73708 23792
rect 73748 23752 73757 23792
rect 73699 23751 73757 23752
rect 74083 23792 74141 23793
rect 74083 23752 74092 23792
rect 74132 23752 74141 23792
rect 74083 23751 74141 23752
rect 74467 23792 74525 23793
rect 74467 23752 74476 23792
rect 74516 23752 74525 23792
rect 74467 23751 74525 23752
rect 74851 23792 74909 23793
rect 74851 23752 74860 23792
rect 74900 23752 74909 23792
rect 74851 23751 74909 23752
rect 75235 23792 75293 23793
rect 75235 23752 75244 23792
rect 75284 23752 75293 23792
rect 75235 23751 75293 23752
rect 75619 23792 75677 23793
rect 75619 23752 75628 23792
rect 75668 23752 75677 23792
rect 75619 23751 75677 23752
rect 76099 23792 76157 23793
rect 76099 23752 76108 23792
rect 76148 23752 76157 23792
rect 76099 23751 76157 23752
rect 76963 23792 77021 23793
rect 76963 23752 76972 23792
rect 77012 23752 77021 23792
rect 76963 23751 77021 23752
rect 77251 23792 77309 23793
rect 77251 23752 77260 23792
rect 77300 23752 77309 23792
rect 77251 23751 77309 23752
rect 77539 23792 77597 23793
rect 77539 23752 77548 23792
rect 77588 23752 77597 23792
rect 77539 23751 77597 23752
rect 77731 23792 77789 23793
rect 77731 23752 77740 23792
rect 77780 23752 77789 23792
rect 77731 23751 77789 23752
rect 78115 23792 78173 23793
rect 78115 23752 78124 23792
rect 78164 23752 78173 23792
rect 78115 23751 78173 23752
rect 78499 23792 78557 23793
rect 78499 23752 78508 23792
rect 78548 23752 78557 23792
rect 78499 23751 78557 23752
rect 78787 23792 78845 23793
rect 78787 23752 78796 23792
rect 78836 23752 78845 23792
rect 78787 23751 78845 23752
rect 79075 23792 79133 23793
rect 79075 23752 79084 23792
rect 79124 23752 79133 23792
rect 79075 23751 79133 23752
rect 79363 23792 79421 23793
rect 79363 23752 79372 23792
rect 79412 23752 79421 23792
rect 79363 23751 79421 23752
rect 32907 23708 32949 23717
rect 32907 23668 32908 23708
rect 32948 23668 32949 23708
rect 32907 23659 32949 23668
rect 39051 23708 39093 23717
rect 39051 23668 39052 23708
rect 39092 23668 39093 23708
rect 39051 23659 39093 23668
rect 40971 23708 41013 23717
rect 40971 23668 40972 23708
rect 41012 23668 41013 23708
rect 40971 23659 41013 23668
rect 48075 23708 48117 23717
rect 48075 23668 48076 23708
rect 48116 23668 48117 23708
rect 48075 23659 48117 23668
rect 50763 23708 50805 23717
rect 50763 23668 50764 23708
rect 50804 23668 50805 23708
rect 50763 23659 50805 23668
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 1611 23624 1653 23633
rect 1611 23584 1612 23624
rect 1652 23584 1653 23624
rect 1611 23575 1653 23584
rect 2187 23624 2229 23633
rect 2187 23584 2188 23624
rect 2228 23584 2229 23624
rect 2187 23575 2229 23584
rect 31083 23624 31125 23633
rect 31083 23584 31084 23624
rect 31124 23584 31125 23624
rect 31083 23575 31125 23584
rect 31363 23624 31421 23625
rect 31363 23584 31372 23624
rect 31412 23584 31421 23624
rect 31363 23583 31421 23584
rect 35299 23624 35357 23625
rect 35299 23584 35308 23624
rect 35348 23584 35357 23624
rect 35299 23583 35357 23584
rect 39331 23624 39389 23625
rect 39331 23584 39340 23624
rect 39380 23584 39389 23624
rect 39331 23583 39389 23584
rect 41451 23624 41493 23633
rect 41451 23584 41452 23624
rect 41492 23584 41493 23624
rect 41451 23575 41493 23584
rect 43939 23624 43997 23625
rect 43939 23584 43948 23624
rect 43988 23584 43997 23624
rect 43939 23583 43997 23584
rect 50467 23624 50525 23625
rect 50467 23584 50476 23624
rect 50516 23584 50525 23624
rect 50467 23583 50525 23584
rect 54115 23624 54173 23625
rect 54115 23584 54124 23624
rect 54164 23584 54173 23624
rect 54115 23583 54173 23584
rect 54891 23624 54933 23633
rect 54891 23584 54892 23624
rect 54932 23584 54933 23624
rect 54891 23575 54933 23584
rect 55275 23624 55317 23633
rect 55275 23584 55276 23624
rect 55316 23584 55317 23624
rect 55275 23575 55317 23584
rect 56043 23624 56085 23633
rect 56043 23584 56044 23624
rect 56084 23584 56085 23624
rect 56043 23575 56085 23584
rect 56331 23624 56373 23633
rect 56331 23584 56332 23624
rect 56372 23584 56373 23624
rect 56331 23575 56373 23584
rect 56715 23624 56757 23633
rect 56715 23584 56716 23624
rect 56756 23584 56757 23624
rect 56715 23575 56757 23584
rect 57003 23624 57045 23633
rect 57003 23584 57004 23624
rect 57044 23584 57045 23624
rect 57003 23575 57045 23584
rect 57387 23624 57429 23633
rect 57387 23584 57388 23624
rect 57428 23584 57429 23624
rect 57387 23575 57429 23584
rect 57771 23624 57813 23633
rect 57771 23584 57772 23624
rect 57812 23584 57813 23624
rect 57771 23575 57813 23584
rect 58155 23624 58197 23633
rect 58155 23584 58156 23624
rect 58196 23584 58197 23624
rect 58155 23575 58197 23584
rect 58539 23624 58581 23633
rect 58539 23584 58540 23624
rect 58580 23584 58581 23624
rect 58539 23575 58581 23584
rect 58923 23624 58965 23633
rect 58923 23584 58924 23624
rect 58964 23584 58965 23624
rect 58923 23575 58965 23584
rect 59403 23624 59445 23633
rect 59403 23584 59404 23624
rect 59444 23584 59445 23624
rect 59403 23575 59445 23584
rect 59787 23624 59829 23633
rect 59787 23584 59788 23624
rect 59828 23584 59829 23624
rect 59787 23575 59829 23584
rect 60171 23624 60213 23633
rect 60171 23584 60172 23624
rect 60212 23584 60213 23624
rect 60171 23575 60213 23584
rect 60555 23624 60597 23633
rect 60555 23584 60556 23624
rect 60596 23584 60597 23624
rect 60555 23575 60597 23584
rect 60939 23624 60981 23633
rect 60939 23584 60940 23624
rect 60980 23584 60981 23624
rect 60939 23575 60981 23584
rect 61419 23624 61461 23633
rect 61419 23584 61420 23624
rect 61460 23584 61461 23624
rect 61419 23575 61461 23584
rect 61803 23624 61845 23633
rect 61803 23584 61804 23624
rect 61844 23584 61845 23624
rect 61803 23575 61845 23584
rect 62187 23624 62229 23633
rect 62187 23584 62188 23624
rect 62228 23584 62229 23624
rect 62187 23575 62229 23584
rect 62571 23624 62613 23633
rect 62571 23584 62572 23624
rect 62612 23584 62613 23624
rect 62571 23575 62613 23584
rect 62955 23624 62997 23633
rect 62955 23584 62956 23624
rect 62996 23584 62997 23624
rect 62955 23575 62997 23584
rect 63339 23624 63381 23633
rect 63339 23584 63340 23624
rect 63380 23584 63381 23624
rect 63339 23575 63381 23584
rect 63723 23624 63765 23633
rect 63723 23584 63724 23624
rect 63764 23584 63765 23624
rect 63723 23575 63765 23584
rect 64203 23624 64245 23633
rect 64203 23584 64204 23624
rect 64244 23584 64245 23624
rect 64203 23575 64245 23584
rect 64587 23624 64629 23633
rect 64587 23584 64588 23624
rect 64628 23584 64629 23624
rect 64587 23575 64629 23584
rect 64971 23624 65013 23633
rect 64971 23584 64972 23624
rect 65012 23584 65013 23624
rect 64971 23575 65013 23584
rect 65355 23624 65397 23633
rect 65355 23584 65356 23624
rect 65396 23584 65397 23624
rect 65355 23575 65397 23584
rect 65835 23624 65877 23633
rect 65835 23584 65836 23624
rect 65876 23584 65877 23624
rect 65835 23575 65877 23584
rect 66219 23624 66261 23633
rect 66219 23584 66220 23624
rect 66260 23584 66261 23624
rect 66219 23575 66261 23584
rect 66603 23624 66645 23633
rect 66603 23584 66604 23624
rect 66644 23584 66645 23624
rect 66603 23575 66645 23584
rect 66987 23624 67029 23633
rect 66987 23584 66988 23624
rect 67028 23584 67029 23624
rect 66987 23575 67029 23584
rect 67371 23624 67413 23633
rect 67371 23584 67372 23624
rect 67412 23584 67413 23624
rect 67371 23575 67413 23584
rect 67755 23624 67797 23633
rect 67755 23584 67756 23624
rect 67796 23584 67797 23624
rect 67755 23575 67797 23584
rect 68235 23624 68277 23633
rect 68235 23584 68236 23624
rect 68276 23584 68277 23624
rect 68235 23575 68277 23584
rect 68619 23624 68661 23633
rect 68619 23584 68620 23624
rect 68660 23584 68661 23624
rect 68619 23575 68661 23584
rect 69003 23624 69045 23633
rect 69003 23584 69004 23624
rect 69044 23584 69045 23624
rect 69003 23575 69045 23584
rect 69387 23624 69429 23633
rect 69387 23584 69388 23624
rect 69428 23584 69429 23624
rect 69387 23575 69429 23584
rect 69771 23624 69813 23633
rect 69771 23584 69772 23624
rect 69812 23584 69813 23624
rect 69771 23575 69813 23584
rect 70251 23624 70293 23633
rect 70251 23584 70252 23624
rect 70292 23584 70293 23624
rect 70251 23575 70293 23584
rect 70635 23624 70677 23633
rect 70635 23584 70636 23624
rect 70676 23584 70677 23624
rect 70635 23575 70677 23584
rect 71019 23624 71061 23633
rect 71019 23584 71020 23624
rect 71060 23584 71061 23624
rect 71019 23575 71061 23584
rect 71403 23624 71445 23633
rect 71403 23584 71404 23624
rect 71444 23584 71445 23624
rect 71403 23575 71445 23584
rect 71787 23624 71829 23633
rect 71787 23584 71788 23624
rect 71828 23584 71829 23624
rect 71787 23575 71829 23584
rect 72171 23624 72213 23633
rect 72171 23584 72172 23624
rect 72212 23584 72213 23624
rect 72171 23575 72213 23584
rect 72555 23624 72597 23633
rect 72555 23584 72556 23624
rect 72596 23584 72597 23624
rect 72555 23575 72597 23584
rect 72939 23624 72981 23633
rect 72939 23584 72940 23624
rect 72980 23584 72981 23624
rect 72939 23575 72981 23584
rect 73419 23624 73461 23633
rect 73419 23584 73420 23624
rect 73460 23584 73461 23624
rect 73419 23575 73461 23584
rect 73803 23624 73845 23633
rect 73803 23584 73804 23624
rect 73844 23584 73845 23624
rect 73803 23575 73845 23584
rect 74187 23624 74229 23633
rect 74187 23584 74188 23624
rect 74228 23584 74229 23624
rect 74187 23575 74229 23584
rect 74571 23624 74613 23633
rect 74571 23584 74572 23624
rect 74612 23584 74613 23624
rect 74571 23575 74613 23584
rect 74955 23624 74997 23633
rect 74955 23584 74956 23624
rect 74996 23584 74997 23624
rect 74955 23575 74997 23584
rect 75339 23624 75381 23633
rect 75339 23584 75340 23624
rect 75380 23584 75381 23624
rect 75339 23575 75381 23584
rect 75723 23624 75765 23633
rect 75723 23584 75724 23624
rect 75764 23584 75765 23624
rect 75723 23575 75765 23584
rect 76203 23624 76245 23633
rect 76203 23584 76204 23624
rect 76244 23584 76245 23624
rect 76203 23575 76245 23584
rect 76875 23624 76917 23633
rect 76875 23584 76876 23624
rect 76916 23584 76917 23624
rect 76875 23575 76917 23584
rect 77163 23624 77205 23633
rect 77163 23584 77164 23624
rect 77204 23584 77205 23624
rect 77163 23575 77205 23584
rect 77451 23624 77493 23633
rect 77451 23584 77452 23624
rect 77492 23584 77493 23624
rect 77451 23575 77493 23584
rect 77835 23624 77877 23633
rect 77835 23584 77836 23624
rect 77876 23584 77877 23624
rect 77835 23575 77877 23584
rect 78219 23624 78261 23633
rect 78219 23584 78220 23624
rect 78260 23584 78261 23624
rect 78219 23575 78261 23584
rect 78603 23624 78645 23633
rect 78603 23584 78604 23624
rect 78644 23584 78645 23624
rect 78603 23575 78645 23584
rect 78891 23624 78933 23633
rect 78891 23584 78892 23624
rect 78932 23584 78933 23624
rect 78891 23575 78933 23584
rect 79179 23624 79221 23633
rect 79179 23584 79180 23624
rect 79220 23584 79221 23624
rect 79179 23575 79221 23584
rect 79467 23624 79509 23633
rect 79467 23584 79468 23624
rect 79508 23584 79509 23624
rect 79467 23575 79509 23584
rect 576 23456 79584 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 79584 23456
rect 576 23392 79584 23416
rect 41067 23330 41109 23339
rect 41067 23290 41068 23330
rect 41108 23290 41109 23330
rect 51051 23330 51093 23339
rect 32611 23288 32669 23289
rect 32611 23248 32620 23288
rect 32660 23248 32669 23288
rect 32611 23247 32669 23248
rect 37891 23288 37949 23289
rect 37891 23248 37900 23288
rect 37940 23248 37949 23288
rect 37891 23247 37949 23248
rect 40867 23288 40925 23289
rect 40867 23248 40876 23288
rect 40916 23248 40925 23288
rect 41067 23281 41109 23290
rect 44707 23288 44765 23289
rect 40867 23247 40925 23248
rect 44707 23248 44716 23288
rect 44756 23248 44765 23288
rect 44707 23247 44765 23248
rect 48739 23288 48797 23289
rect 48739 23248 48748 23288
rect 48788 23248 48797 23288
rect 48739 23247 48797 23248
rect 49611 23288 49653 23297
rect 51051 23290 51052 23330
rect 51092 23290 51093 23330
rect 49611 23248 49612 23288
rect 49652 23248 49653 23288
rect 49611 23239 49653 23248
rect 50083 23288 50141 23289
rect 50083 23248 50092 23288
rect 50132 23248 50141 23288
rect 51051 23281 51093 23290
rect 50083 23247 50141 23248
rect 32235 23204 32277 23213
rect 32235 23164 32236 23204
rect 32276 23164 32277 23204
rect 32235 23155 32277 23164
rect 36651 23204 36693 23213
rect 36651 23164 36652 23204
rect 36692 23164 36693 23204
rect 36651 23155 36693 23164
rect 41355 23204 41397 23213
rect 41355 23164 41356 23204
rect 41396 23164 41397 23204
rect 41355 23155 41397 23164
rect 45579 23204 45621 23213
rect 45579 23164 45580 23204
rect 45620 23164 45621 23204
rect 45579 23155 45621 23164
rect 50763 23204 50805 23213
rect 50763 23164 50764 23204
rect 50804 23164 50805 23204
rect 50763 23155 50805 23164
rect 51339 23204 51381 23213
rect 51339 23164 51340 23204
rect 51380 23164 51381 23204
rect 51339 23155 51381 23164
rect 51235 23141 51293 23142
rect 1515 23120 1557 23129
rect 1515 23080 1516 23120
rect 1556 23080 1557 23120
rect 1515 23071 1557 23080
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 1941 23120
rect 1899 23071 1941 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 28395 23120 28437 23129
rect 28395 23080 28396 23120
rect 28436 23080 28437 23120
rect 28395 23071 28437 23080
rect 28771 23120 28829 23121
rect 28771 23080 28780 23120
rect 28820 23080 28829 23120
rect 28771 23079 28829 23080
rect 29635 23120 29693 23121
rect 29635 23080 29644 23120
rect 29684 23080 29693 23120
rect 29635 23079 29693 23080
rect 30987 23120 31029 23129
rect 30987 23080 30988 23120
rect 31028 23080 31029 23120
rect 30987 23071 31029 23080
rect 31179 23120 31221 23129
rect 31179 23080 31180 23120
rect 31220 23080 31221 23120
rect 31179 23071 31221 23080
rect 31267 23120 31325 23121
rect 31267 23080 31276 23120
rect 31316 23080 31325 23120
rect 31267 23079 31325 23080
rect 31747 23120 31805 23121
rect 31747 23080 31756 23120
rect 31796 23080 31805 23120
rect 31747 23079 31805 23080
rect 31947 23120 31989 23129
rect 31947 23080 31948 23120
rect 31988 23080 31989 23120
rect 31947 23071 31989 23080
rect 32131 23120 32189 23121
rect 32131 23080 32140 23120
rect 32180 23080 32189 23120
rect 32131 23079 32189 23080
rect 32331 23120 32373 23129
rect 32331 23080 32332 23120
rect 32372 23080 32373 23120
rect 32331 23071 32373 23080
rect 32523 23120 32565 23129
rect 32523 23080 32524 23120
rect 32564 23080 32565 23120
rect 32523 23071 32565 23080
rect 32715 23120 32757 23129
rect 32715 23080 32716 23120
rect 32756 23080 32757 23120
rect 32715 23071 32757 23080
rect 32803 23120 32861 23121
rect 32803 23080 32812 23120
rect 32852 23080 32861 23120
rect 32803 23079 32861 23080
rect 36259 23120 36317 23121
rect 36259 23080 36268 23120
rect 36308 23080 36317 23120
rect 36259 23079 36317 23080
rect 36555 23120 36597 23129
rect 36555 23080 36556 23120
rect 36596 23080 36597 23120
rect 36555 23071 36597 23080
rect 37131 23120 37173 23129
rect 37131 23080 37132 23120
rect 37172 23080 37173 23120
rect 37131 23071 37173 23080
rect 37227 23120 37269 23129
rect 37227 23080 37228 23120
rect 37268 23080 37269 23120
rect 37227 23071 37269 23080
rect 37315 23120 37373 23121
rect 37315 23080 37324 23120
rect 37364 23080 37373 23120
rect 37315 23079 37373 23080
rect 37803 23120 37845 23129
rect 37803 23080 37804 23120
rect 37844 23080 37845 23120
rect 37803 23071 37845 23080
rect 37995 23120 38037 23129
rect 37995 23080 37996 23120
rect 38036 23080 38037 23120
rect 37995 23071 38037 23080
rect 38083 23120 38141 23121
rect 38083 23080 38092 23120
rect 38132 23080 38141 23120
rect 38083 23079 38141 23080
rect 38475 23120 38517 23129
rect 38475 23080 38476 23120
rect 38516 23080 38517 23120
rect 38475 23071 38517 23080
rect 38851 23120 38909 23121
rect 38851 23080 38860 23120
rect 38900 23080 38909 23120
rect 38851 23079 38909 23080
rect 39715 23120 39773 23121
rect 39715 23080 39724 23120
rect 39764 23080 39773 23120
rect 39715 23079 39773 23080
rect 41451 23120 41493 23129
rect 41451 23080 41452 23120
rect 41492 23080 41493 23120
rect 41451 23071 41493 23080
rect 41731 23120 41789 23121
rect 41731 23080 41740 23120
rect 41780 23080 41789 23120
rect 41731 23079 41789 23080
rect 44619 23120 44661 23129
rect 44619 23080 44620 23120
rect 44660 23080 44661 23120
rect 44619 23071 44661 23080
rect 44811 23120 44853 23129
rect 44811 23080 44812 23120
rect 44852 23080 44853 23120
rect 44811 23071 44853 23080
rect 44899 23120 44957 23121
rect 44899 23080 44908 23120
rect 44948 23080 44957 23120
rect 44899 23079 44957 23080
rect 45483 23120 45525 23129
rect 45483 23080 45484 23120
rect 45524 23080 45525 23120
rect 45483 23071 45525 23080
rect 45667 23120 45725 23121
rect 45667 23080 45676 23120
rect 45716 23080 45725 23120
rect 45667 23079 45725 23080
rect 45859 23120 45917 23121
rect 45859 23080 45868 23120
rect 45908 23080 45917 23120
rect 45859 23079 45917 23080
rect 45963 23120 46005 23129
rect 45963 23080 45964 23120
rect 46004 23080 46005 23120
rect 45963 23071 46005 23080
rect 46155 23120 46197 23129
rect 46155 23080 46156 23120
rect 46196 23080 46197 23120
rect 46155 23071 46197 23080
rect 46347 23120 46389 23129
rect 46347 23080 46348 23120
rect 46388 23080 46389 23120
rect 46347 23071 46389 23080
rect 46723 23120 46781 23121
rect 46723 23080 46732 23120
rect 46772 23080 46781 23120
rect 46723 23079 46781 23080
rect 47587 23120 47645 23121
rect 47587 23080 47596 23120
rect 47636 23080 47645 23120
rect 49899 23120 49941 23129
rect 47587 23079 47645 23080
rect 49803 23075 49845 23084
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 49411 23036 49469 23037
rect 49411 22996 49420 23036
rect 49460 22996 49469 23036
rect 49803 23035 49804 23075
rect 49844 23035 49845 23075
rect 49899 23080 49900 23120
rect 49940 23080 49941 23120
rect 49899 23071 49941 23080
rect 49995 23120 50037 23129
rect 49995 23080 49996 23120
rect 50036 23080 50037 23120
rect 49995 23071 50037 23080
rect 50371 23120 50429 23121
rect 50371 23080 50380 23120
rect 50420 23080 50429 23120
rect 50371 23079 50429 23080
rect 50667 23120 50709 23129
rect 50667 23080 50668 23120
rect 50708 23080 50709 23120
rect 51235 23101 51244 23141
rect 51284 23101 51293 23141
rect 51235 23100 51293 23101
rect 51435 23120 51477 23129
rect 50667 23071 50709 23080
rect 51435 23080 51436 23120
rect 51476 23080 51477 23120
rect 51435 23071 51477 23080
rect 52491 23120 52533 23129
rect 52491 23080 52492 23120
rect 52532 23080 52533 23120
rect 52491 23071 52533 23080
rect 49803 23026 49845 23035
rect 51723 23036 51765 23045
rect 49411 22995 49469 22996
rect 51723 22996 51724 23036
rect 51764 22996 51765 23036
rect 51723 22987 51765 22996
rect 1515 22952 1557 22961
rect 1515 22912 1516 22952
rect 1556 22912 1557 22952
rect 1515 22903 1557 22912
rect 30987 22952 31029 22961
rect 30987 22912 30988 22952
rect 31028 22912 31029 22952
rect 30987 22903 31029 22912
rect 33387 22952 33429 22961
rect 33387 22912 33388 22952
rect 33428 22912 33429 22952
rect 33387 22903 33429 22912
rect 35979 22952 36021 22961
rect 35979 22912 35980 22952
rect 36020 22912 36021 22952
rect 35979 22903 36021 22912
rect 36931 22952 36989 22953
rect 36931 22912 36940 22952
rect 36980 22912 36989 22952
rect 36931 22911 36989 22912
rect 42027 22952 42069 22961
rect 42027 22912 42028 22952
rect 42068 22912 42069 22952
rect 42027 22903 42069 22912
rect 42891 22952 42933 22961
rect 42891 22912 42892 22952
rect 42932 22912 42933 22952
rect 42891 22903 42933 22912
rect 46155 22952 46197 22961
rect 46155 22912 46156 22952
rect 46196 22912 46197 22952
rect 46155 22903 46197 22912
rect 52299 22952 52341 22961
rect 52299 22912 52300 22952
rect 52340 22912 52341 22952
rect 52299 22903 52341 22912
rect 843 22868 885 22877
rect 843 22828 844 22868
rect 884 22828 885 22868
rect 843 22819 885 22828
rect 1707 22868 1749 22877
rect 1707 22828 1708 22868
rect 1748 22828 1749 22868
rect 1707 22819 1749 22828
rect 1899 22868 1941 22877
rect 1899 22828 1900 22868
rect 1940 22828 1941 22868
rect 1899 22819 1941 22828
rect 30787 22868 30845 22869
rect 30787 22828 30796 22868
rect 30836 22828 30845 22868
rect 30787 22827 30845 22828
rect 31851 22868 31893 22877
rect 31851 22828 31852 22868
rect 31892 22828 31893 22868
rect 31851 22819 31893 22828
rect 49611 22868 49653 22877
rect 49611 22828 49612 22868
rect 49652 22828 49653 22868
rect 49611 22819 49653 22828
rect 576 22700 52800 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 52800 22700
rect 576 22636 52800 22660
rect 28299 22532 28341 22541
rect 28299 22492 28300 22532
rect 28340 22492 28341 22532
rect 28299 22483 28341 22492
rect 31843 22532 31901 22533
rect 31843 22492 31852 22532
rect 31892 22492 31901 22532
rect 31843 22491 31901 22492
rect 35203 22532 35261 22533
rect 35203 22492 35212 22532
rect 35252 22492 35261 22532
rect 35203 22491 35261 22492
rect 39051 22532 39093 22541
rect 39051 22492 39052 22532
rect 39092 22492 39093 22532
rect 39051 22483 39093 22492
rect 43555 22532 43613 22533
rect 43555 22492 43564 22532
rect 43604 22492 43613 22532
rect 43555 22491 43613 22492
rect 50379 22532 50421 22541
rect 50379 22492 50380 22532
rect 50420 22492 50421 22532
rect 50379 22483 50421 22492
rect 52011 22532 52053 22541
rect 52011 22492 52012 22532
rect 52052 22492 52053 22532
rect 52011 22483 52053 22492
rect 52395 22532 52437 22541
rect 52395 22492 52396 22532
rect 52436 22492 52437 22532
rect 52395 22483 52437 22492
rect 52683 22532 52725 22541
rect 52683 22492 52684 22532
rect 52724 22492 52725 22532
rect 52683 22483 52725 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 27915 22448 27957 22457
rect 27915 22408 27916 22448
rect 27956 22408 27957 22448
rect 27915 22399 27957 22408
rect 38859 22448 38901 22457
rect 38859 22408 38860 22448
rect 38900 22408 38901 22448
rect 38859 22399 38901 22408
rect 40971 22448 41013 22457
rect 40971 22408 40972 22448
rect 41012 22408 41013 22448
rect 40971 22399 41013 22408
rect 44907 22448 44949 22457
rect 44907 22408 44908 22448
rect 44948 22408 44949 22448
rect 44907 22399 44949 22408
rect 46443 22448 46485 22457
rect 46443 22408 46444 22448
rect 46484 22408 46485 22448
rect 46443 22399 46485 22408
rect 48171 22448 48213 22457
rect 48171 22408 48172 22448
rect 48212 22408 48213 22448
rect 48171 22399 48213 22408
rect 27715 22364 27773 22365
rect 27715 22324 27724 22364
rect 27764 22324 27773 22364
rect 27715 22323 27773 22324
rect 28099 22364 28157 22365
rect 28099 22324 28108 22364
rect 28148 22324 28157 22364
rect 28099 22323 28157 22324
rect 50179 22364 50237 22365
rect 50179 22324 50188 22364
rect 50228 22324 50237 22364
rect 50179 22323 50237 22324
rect 28483 22280 28541 22281
rect 28483 22240 28492 22280
rect 28532 22240 28541 22280
rect 28483 22239 28541 22240
rect 28683 22280 28725 22289
rect 28683 22240 28684 22280
rect 28724 22240 28725 22280
rect 28683 22231 28725 22240
rect 28867 22280 28925 22281
rect 28867 22240 28876 22280
rect 28916 22240 28925 22280
rect 28867 22239 28925 22240
rect 29067 22280 29109 22289
rect 29067 22240 29068 22280
rect 29108 22240 29109 22280
rect 29067 22231 29109 22240
rect 29547 22280 29589 22289
rect 29547 22240 29548 22280
rect 29588 22240 29589 22280
rect 29547 22231 29589 22240
rect 29739 22280 29781 22289
rect 29739 22240 29740 22280
rect 29780 22240 29781 22280
rect 29739 22231 29781 22240
rect 29827 22280 29885 22281
rect 29827 22240 29836 22280
rect 29876 22240 29885 22280
rect 29827 22239 29885 22240
rect 30603 22280 30645 22289
rect 30603 22240 30604 22280
rect 30644 22240 30645 22280
rect 30603 22231 30645 22240
rect 30699 22280 30741 22289
rect 30699 22240 30700 22280
rect 30740 22240 30741 22280
rect 30699 22231 30741 22240
rect 30795 22280 30837 22289
rect 30795 22240 30796 22280
rect 30836 22240 30837 22280
rect 30795 22231 30837 22240
rect 30891 22280 30933 22289
rect 30891 22240 30892 22280
rect 30932 22240 30933 22280
rect 30891 22231 30933 22240
rect 31171 22280 31229 22281
rect 31171 22240 31180 22280
rect 31220 22240 31229 22280
rect 31171 22239 31229 22240
rect 31467 22280 31509 22289
rect 31467 22240 31468 22280
rect 31508 22240 31509 22280
rect 31467 22231 31509 22240
rect 31563 22280 31605 22289
rect 31563 22240 31564 22280
rect 31604 22240 31605 22280
rect 32331 22280 32373 22289
rect 31563 22231 31605 22240
rect 32139 22238 32181 22247
rect 28587 22196 28629 22205
rect 28587 22156 28588 22196
rect 28628 22156 28629 22196
rect 28587 22147 28629 22156
rect 28971 22196 29013 22205
rect 28971 22156 28972 22196
rect 29012 22156 29013 22196
rect 32139 22198 32140 22238
rect 32180 22198 32181 22238
rect 32331 22240 32332 22280
rect 32372 22240 32373 22280
rect 32331 22231 32373 22240
rect 32419 22280 32477 22281
rect 32419 22240 32428 22280
rect 32468 22240 32477 22280
rect 32419 22239 32477 22240
rect 33187 22280 33245 22281
rect 33187 22240 33196 22280
rect 33236 22240 33245 22280
rect 33187 22239 33245 22240
rect 34051 22280 34109 22281
rect 34051 22240 34060 22280
rect 34100 22240 34109 22280
rect 34051 22239 34109 22240
rect 36067 22280 36125 22281
rect 36067 22240 36076 22280
rect 36116 22240 36125 22280
rect 36067 22239 36125 22240
rect 36931 22280 36989 22281
rect 36931 22240 36940 22280
rect 36980 22240 36989 22280
rect 36931 22239 36989 22240
rect 39051 22280 39093 22289
rect 39051 22240 39052 22280
rect 39092 22240 39093 22280
rect 39051 22231 39093 22240
rect 39243 22280 39285 22289
rect 39243 22240 39244 22280
rect 39284 22240 39285 22280
rect 39243 22231 39285 22240
rect 39331 22280 39389 22281
rect 39331 22240 39340 22280
rect 39380 22240 39389 22280
rect 39331 22239 39389 22240
rect 40675 22280 40733 22281
rect 40675 22240 40684 22280
rect 40724 22240 40733 22280
rect 40675 22239 40733 22240
rect 40779 22280 40821 22289
rect 40779 22240 40780 22280
rect 40820 22240 40821 22280
rect 40779 22231 40821 22240
rect 40971 22280 41013 22289
rect 40971 22240 40972 22280
rect 41012 22240 41013 22280
rect 40971 22231 41013 22240
rect 41163 22280 41205 22289
rect 41163 22240 41164 22280
rect 41204 22240 41205 22280
rect 41163 22231 41205 22240
rect 41539 22280 41597 22281
rect 41539 22240 41548 22280
rect 41588 22240 41597 22280
rect 41539 22239 41597 22240
rect 42403 22280 42461 22281
rect 42403 22240 42412 22280
rect 42452 22240 42461 22280
rect 42403 22239 42461 22240
rect 44803 22280 44861 22281
rect 44803 22240 44812 22280
rect 44852 22240 44861 22280
rect 44803 22239 44861 22240
rect 45003 22280 45045 22289
rect 45003 22240 45004 22280
rect 45044 22240 45045 22280
rect 45003 22231 45045 22240
rect 45195 22280 45237 22289
rect 45195 22240 45196 22280
rect 45236 22240 45237 22280
rect 45195 22231 45237 22240
rect 45387 22280 45429 22289
rect 45387 22240 45388 22280
rect 45428 22240 45429 22280
rect 45387 22231 45429 22240
rect 45475 22280 45533 22281
rect 45475 22240 45484 22280
rect 45524 22240 45533 22280
rect 45475 22239 45533 22240
rect 45675 22280 45717 22289
rect 45675 22240 45676 22280
rect 45716 22240 45717 22280
rect 45675 22231 45717 22240
rect 45859 22280 45917 22281
rect 45859 22240 45868 22280
rect 45908 22240 45917 22280
rect 45859 22239 45917 22240
rect 48555 22280 48597 22289
rect 48555 22240 48556 22280
rect 48596 22240 48597 22280
rect 48555 22231 48597 22240
rect 48651 22280 48693 22289
rect 48651 22240 48652 22280
rect 48692 22240 48693 22280
rect 48651 22231 48693 22240
rect 48747 22280 48789 22289
rect 48747 22240 48748 22280
rect 48788 22240 48789 22280
rect 48747 22231 48789 22240
rect 49419 22280 49461 22289
rect 49419 22240 49420 22280
rect 49460 22240 49461 22280
rect 49419 22231 49461 22240
rect 49611 22280 49653 22289
rect 49611 22240 49612 22280
rect 49652 22240 49653 22280
rect 49611 22231 49653 22240
rect 49699 22280 49757 22281
rect 49699 22240 49708 22280
rect 49748 22240 49757 22280
rect 49699 22239 49757 22240
rect 50571 22280 50613 22289
rect 50571 22240 50572 22280
rect 50612 22240 50613 22280
rect 50571 22231 50613 22240
rect 50755 22280 50813 22281
rect 50755 22240 50764 22280
rect 50804 22240 50813 22280
rect 50755 22239 50813 22240
rect 51619 22280 51677 22281
rect 51619 22240 51628 22280
rect 51668 22240 51677 22280
rect 52291 22280 52349 22281
rect 51619 22239 51677 22240
rect 52099 22269 52157 22270
rect 52099 22229 52108 22269
rect 52148 22229 52157 22269
rect 52291 22240 52300 22280
rect 52340 22240 52349 22280
rect 52291 22239 52349 22240
rect 52579 22280 52637 22281
rect 52579 22240 52588 22280
rect 52628 22240 52637 22280
rect 52579 22239 52637 22240
rect 52099 22228 52157 22229
rect 32139 22189 32181 22198
rect 32235 22196 32277 22205
rect 28971 22147 29013 22156
rect 32235 22156 32236 22196
rect 32276 22156 32277 22196
rect 32235 22147 32277 22156
rect 32811 22196 32853 22205
rect 32811 22156 32812 22196
rect 32852 22156 32853 22196
rect 32811 22147 32853 22156
rect 35691 22196 35733 22205
rect 35691 22156 35692 22196
rect 35732 22156 35733 22196
rect 35691 22147 35733 22156
rect 45771 22196 45813 22205
rect 45771 22156 45772 22196
rect 45812 22156 45813 22196
rect 45771 22147 45813 22156
rect 50667 22196 50709 22205
rect 50667 22156 50668 22196
rect 50708 22156 50709 22196
rect 50667 22147 50709 22156
rect 28299 22112 28341 22121
rect 28299 22072 28300 22112
rect 28340 22072 28341 22112
rect 28299 22063 28341 22072
rect 29635 22112 29693 22113
rect 29635 22072 29644 22112
rect 29684 22072 29693 22112
rect 29635 22071 29693 22072
rect 35203 22112 35261 22113
rect 35203 22072 35212 22112
rect 35252 22072 35261 22112
rect 35203 22071 35261 22072
rect 38083 22112 38141 22113
rect 38083 22072 38092 22112
rect 38132 22072 38141 22112
rect 38083 22071 38141 22072
rect 43555 22112 43613 22113
rect 43555 22072 43564 22112
rect 43604 22072 43613 22112
rect 43555 22071 43613 22072
rect 45283 22112 45341 22113
rect 45283 22072 45292 22112
rect 45332 22072 45341 22112
rect 45283 22071 45341 22072
rect 48835 22112 48893 22113
rect 48835 22072 48844 22112
rect 48884 22072 48893 22112
rect 48835 22071 48893 22072
rect 49507 22112 49565 22113
rect 49507 22072 49516 22112
rect 49556 22072 49565 22112
rect 49507 22071 49565 22072
rect 576 21944 52800 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 52800 21944
rect 576 21880 52800 21904
rect 36163 21776 36221 21777
rect 36163 21736 36172 21776
rect 36212 21736 36221 21776
rect 36163 21735 36221 21736
rect 44803 21776 44861 21777
rect 44803 21736 44812 21776
rect 44852 21736 44861 21776
rect 44803 21735 44861 21736
rect 32427 21692 32469 21701
rect 32427 21652 32428 21692
rect 32468 21652 32469 21692
rect 32427 21643 32469 21652
rect 41259 21692 41301 21701
rect 41259 21652 41260 21692
rect 41300 21652 41301 21692
rect 41259 21643 41301 21652
rect 42411 21692 42453 21701
rect 42411 21652 42412 21692
rect 42452 21652 42453 21692
rect 42411 21643 42453 21652
rect 51051 21692 51093 21701
rect 51051 21652 51052 21692
rect 51092 21652 51093 21692
rect 51051 21643 51093 21652
rect 26659 21608 26717 21609
rect 26659 21568 26668 21608
rect 26708 21568 26717 21608
rect 26659 21567 26717 21568
rect 27523 21608 27581 21609
rect 27523 21568 27532 21608
rect 27572 21568 27581 21608
rect 27523 21567 27581 21568
rect 27915 21608 27957 21617
rect 27915 21568 27916 21608
rect 27956 21568 27957 21608
rect 27915 21559 27957 21568
rect 28195 21608 28253 21609
rect 28195 21568 28204 21608
rect 28244 21568 28253 21608
rect 28195 21567 28253 21568
rect 28491 21608 28533 21617
rect 28491 21568 28492 21608
rect 28532 21568 28533 21608
rect 28491 21559 28533 21568
rect 28587 21608 28629 21617
rect 28587 21568 28588 21608
rect 28628 21568 28629 21608
rect 28587 21559 28629 21568
rect 29355 21608 29397 21617
rect 29355 21568 29356 21608
rect 29396 21568 29397 21608
rect 29355 21559 29397 21568
rect 29731 21608 29789 21609
rect 29731 21568 29740 21608
rect 29780 21568 29789 21608
rect 29731 21567 29789 21568
rect 30595 21608 30653 21609
rect 30595 21568 30604 21608
rect 30644 21568 30653 21608
rect 30595 21567 30653 21568
rect 32331 21608 32373 21617
rect 32331 21568 32332 21608
rect 32372 21568 32373 21608
rect 32331 21559 32373 21568
rect 32515 21608 32573 21609
rect 32515 21568 32524 21608
rect 32564 21568 32573 21608
rect 32515 21567 32573 21568
rect 36075 21608 36117 21617
rect 36075 21568 36076 21608
rect 36116 21568 36117 21608
rect 36075 21559 36117 21568
rect 36267 21608 36309 21617
rect 36267 21568 36268 21608
rect 36308 21568 36309 21608
rect 36267 21559 36309 21568
rect 36355 21608 36413 21609
rect 36355 21568 36364 21608
rect 36404 21568 36413 21608
rect 36355 21567 36413 21568
rect 36547 21608 36605 21609
rect 36547 21568 36556 21608
rect 36596 21568 36605 21608
rect 36547 21567 36605 21568
rect 36747 21608 36789 21617
rect 36747 21568 36748 21608
rect 36788 21568 36789 21608
rect 36747 21559 36789 21568
rect 38955 21608 38997 21617
rect 38955 21568 38956 21608
rect 38996 21568 38997 21608
rect 38955 21559 38997 21568
rect 39051 21608 39093 21617
rect 39051 21568 39052 21608
rect 39092 21568 39093 21608
rect 39051 21559 39093 21568
rect 39147 21608 39189 21617
rect 39147 21568 39148 21608
rect 39188 21568 39189 21608
rect 39147 21559 39189 21568
rect 39243 21608 39285 21617
rect 39243 21568 39244 21608
rect 39284 21568 39285 21608
rect 39243 21559 39285 21568
rect 41155 21608 41213 21609
rect 41155 21568 41164 21608
rect 41204 21568 41213 21608
rect 41155 21567 41213 21568
rect 41355 21608 41397 21617
rect 41355 21568 41356 21608
rect 41396 21568 41397 21608
rect 41355 21559 41397 21568
rect 42787 21608 42845 21609
rect 42787 21568 42796 21608
rect 42836 21568 42845 21608
rect 42787 21567 42845 21568
rect 43651 21608 43709 21609
rect 43651 21568 43660 21608
rect 43700 21568 43709 21608
rect 43651 21567 43709 21568
rect 45291 21608 45333 21617
rect 45291 21568 45292 21608
rect 45332 21568 45333 21608
rect 45291 21559 45333 21568
rect 45387 21608 45429 21617
rect 45387 21568 45388 21608
rect 45428 21568 45429 21608
rect 45387 21559 45429 21568
rect 45667 21608 45725 21609
rect 45667 21568 45676 21608
rect 45716 21568 45725 21608
rect 45667 21567 45725 21568
rect 45963 21608 46005 21617
rect 45963 21568 45964 21608
rect 46004 21568 46005 21608
rect 45963 21559 46005 21568
rect 46339 21608 46397 21609
rect 46339 21568 46348 21608
rect 46388 21568 46397 21608
rect 46339 21567 46397 21568
rect 47203 21608 47261 21609
rect 47203 21568 47212 21608
rect 47252 21568 47261 21608
rect 47203 21567 47261 21568
rect 48843 21608 48885 21617
rect 48843 21568 48844 21608
rect 48884 21568 48885 21608
rect 48843 21559 48885 21568
rect 49035 21608 49077 21617
rect 49035 21568 49036 21608
rect 49076 21568 49077 21608
rect 49035 21559 49077 21568
rect 49123 21608 49181 21609
rect 49123 21568 49132 21608
rect 49172 21568 49181 21608
rect 49123 21567 49181 21568
rect 49507 21608 49565 21609
rect 49507 21568 49516 21608
rect 49556 21568 49565 21608
rect 49507 21567 49565 21568
rect 49611 21608 49653 21617
rect 49611 21568 49612 21608
rect 49652 21568 49653 21608
rect 49611 21559 49653 21568
rect 49707 21608 49749 21617
rect 49707 21568 49708 21608
rect 49748 21568 49749 21608
rect 49707 21559 49749 21568
rect 50187 21608 50229 21617
rect 50187 21568 50188 21608
rect 50228 21568 50229 21608
rect 50187 21559 50229 21568
rect 50283 21608 50325 21617
rect 50283 21568 50284 21608
rect 50324 21568 50325 21608
rect 50283 21559 50325 21568
rect 50563 21608 50621 21609
rect 50563 21568 50572 21608
rect 50612 21568 50621 21608
rect 50563 21567 50621 21568
rect 50851 21608 50909 21609
rect 50851 21568 50860 21608
rect 50900 21568 50909 21608
rect 50851 21567 50909 21568
rect 50955 21608 50997 21617
rect 50955 21568 50956 21608
rect 50996 21568 50997 21608
rect 50955 21559 50997 21568
rect 51147 21608 51189 21617
rect 51147 21568 51148 21608
rect 51188 21568 51189 21608
rect 51147 21559 51189 21568
rect 52291 21608 52349 21609
rect 52291 21568 52300 21608
rect 52340 21568 52349 21608
rect 52291 21567 52349 21568
rect 52395 21608 52437 21617
rect 52395 21568 52396 21608
rect 52436 21568 52437 21608
rect 52395 21559 52437 21568
rect 52579 21608 52637 21609
rect 52579 21568 52588 21608
rect 52628 21568 52637 21608
rect 52579 21567 52637 21568
rect 52683 21608 52725 21617
rect 52683 21568 52684 21608
rect 52724 21568 52725 21608
rect 52683 21559 52725 21568
rect 3043 21524 3101 21525
rect 3043 21484 3052 21524
rect 3092 21484 3101 21524
rect 3043 21483 3101 21484
rect 3619 21524 3677 21525
rect 3619 21484 3628 21524
rect 3668 21484 3677 21524
rect 3619 21483 3677 21484
rect 4003 21524 4061 21525
rect 4003 21484 4012 21524
rect 4052 21484 4061 21524
rect 4003 21483 4061 21484
rect 4195 21524 4253 21525
rect 4195 21484 4204 21524
rect 4244 21484 4253 21524
rect 4195 21483 4253 21484
rect 3243 21440 3285 21449
rect 3243 21400 3244 21440
rect 3284 21400 3285 21440
rect 3243 21391 3285 21400
rect 28867 21440 28925 21441
rect 28867 21400 28876 21440
rect 28916 21400 28925 21440
rect 28867 21399 28925 21400
rect 31747 21440 31805 21441
rect 31747 21400 31756 21440
rect 31796 21400 31805 21440
rect 31747 21399 31805 21400
rect 32715 21440 32757 21449
rect 32715 21400 32716 21440
rect 32756 21400 32757 21440
rect 32715 21391 32757 21400
rect 33291 21440 33333 21449
rect 33291 21400 33292 21440
rect 33332 21400 33333 21440
rect 33291 21391 33333 21400
rect 35691 21440 35733 21449
rect 35691 21400 35692 21440
rect 35732 21400 35733 21440
rect 35691 21391 35733 21400
rect 36651 21440 36693 21449
rect 36651 21400 36652 21440
rect 36692 21400 36693 21440
rect 36651 21391 36693 21400
rect 39435 21440 39477 21449
rect 39435 21400 39436 21440
rect 39476 21400 39477 21440
rect 39435 21391 39477 21400
rect 44995 21440 45053 21441
rect 44995 21400 45004 21440
rect 45044 21400 45053 21440
rect 44995 21399 45053 21400
rect 49891 21440 49949 21441
rect 49891 21400 49900 21440
rect 49940 21400 49949 21440
rect 49891 21399 49949 21400
rect 51339 21440 51381 21449
rect 51339 21400 51340 21440
rect 51380 21400 51381 21440
rect 51339 21391 51381 21400
rect 3435 21356 3477 21365
rect 3435 21316 3436 21356
rect 3476 21316 3477 21356
rect 3435 21307 3477 21316
rect 3819 21356 3861 21365
rect 3819 21316 3820 21356
rect 3860 21316 3861 21356
rect 3819 21307 3861 21316
rect 4395 21356 4437 21365
rect 4395 21316 4396 21356
rect 4436 21316 4437 21356
rect 4395 21307 4437 21316
rect 25507 21356 25565 21357
rect 25507 21316 25516 21356
rect 25556 21316 25565 21356
rect 25507 21315 25565 21316
rect 48355 21356 48413 21357
rect 48355 21316 48364 21356
rect 48404 21316 48413 21356
rect 48355 21315 48413 21316
rect 48843 21356 48885 21365
rect 48843 21316 48844 21356
rect 48884 21316 48885 21356
rect 48843 21307 48885 21316
rect 576 21188 52800 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 52800 21188
rect 576 21124 52800 21148
rect 26955 21020 26997 21029
rect 26955 20980 26956 21020
rect 26996 20980 26997 21020
rect 26955 20971 26997 20980
rect 28299 21020 28341 21029
rect 28299 20980 28300 21020
rect 28340 20980 28341 21020
rect 28299 20971 28341 20980
rect 29067 21020 29109 21029
rect 29067 20980 29068 21020
rect 29108 20980 29109 21020
rect 29067 20971 29109 20980
rect 43851 21020 43893 21029
rect 43851 20980 43852 21020
rect 43892 20980 43893 21020
rect 43851 20971 43893 20980
rect 46347 21020 46389 21029
rect 46347 20980 46348 21020
rect 46388 20980 46389 21020
rect 46347 20971 46389 20980
rect 50083 21020 50141 21021
rect 50083 20980 50092 21020
rect 50132 20980 50141 21020
rect 50083 20979 50141 20980
rect 52675 21020 52733 21021
rect 52675 20980 52684 21020
rect 52724 20980 52733 21020
rect 52675 20979 52733 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 26187 20936 26229 20945
rect 26187 20896 26188 20936
rect 26228 20896 26229 20936
rect 26187 20887 26229 20896
rect 29835 20936 29877 20945
rect 29835 20896 29836 20936
rect 29876 20896 29877 20936
rect 29835 20887 29877 20896
rect 38475 20936 38517 20945
rect 38475 20896 38476 20936
rect 38516 20896 38517 20936
rect 38475 20887 38517 20896
rect 41931 20936 41973 20945
rect 41931 20896 41932 20936
rect 41972 20896 41973 20936
rect 41931 20887 41973 20896
rect 5059 20852 5117 20853
rect 5059 20812 5068 20852
rect 5108 20812 5117 20852
rect 5059 20811 5117 20812
rect 23203 20852 23261 20853
rect 23203 20812 23212 20852
rect 23252 20812 23261 20852
rect 23203 20811 23261 20812
rect 26371 20852 26429 20853
rect 26371 20812 26380 20852
rect 26420 20812 26429 20852
rect 26371 20811 26429 20812
rect 26755 20852 26813 20853
rect 26755 20812 26764 20852
rect 26804 20812 26813 20852
rect 26755 20811 26813 20812
rect 27139 20852 27197 20853
rect 27139 20812 27148 20852
rect 27188 20812 27197 20852
rect 27139 20811 27197 20812
rect 42883 20852 42941 20853
rect 42883 20812 42892 20852
rect 42932 20812 42941 20852
rect 42883 20811 42941 20812
rect 43459 20852 43517 20853
rect 43459 20812 43468 20852
rect 43508 20812 43517 20852
rect 43459 20811 43517 20812
rect 43651 20852 43709 20853
rect 43651 20812 43660 20852
rect 43700 20812 43709 20852
rect 43651 20811 43709 20812
rect 44035 20852 44093 20853
rect 44035 20812 44044 20852
rect 44084 20812 44093 20852
rect 44035 20811 44093 20812
rect 44611 20852 44669 20853
rect 44611 20812 44620 20852
rect 44660 20812 44669 20852
rect 44611 20811 44669 20812
rect 3523 20768 3581 20769
rect 3523 20728 3532 20768
rect 3572 20728 3581 20768
rect 3523 20727 3581 20728
rect 3627 20768 3669 20777
rect 3627 20728 3628 20768
rect 3668 20728 3669 20768
rect 3627 20719 3669 20728
rect 3819 20768 3861 20777
rect 3819 20728 3820 20768
rect 3860 20728 3861 20768
rect 3819 20719 3861 20728
rect 27819 20768 27861 20777
rect 27819 20728 27820 20768
rect 27860 20728 27861 20768
rect 27819 20719 27861 20728
rect 27915 20768 27957 20777
rect 27915 20728 27916 20768
rect 27956 20728 27957 20768
rect 27915 20719 27957 20728
rect 28011 20768 28053 20777
rect 28011 20728 28012 20768
rect 28052 20728 28053 20768
rect 28011 20719 28053 20728
rect 28107 20768 28149 20777
rect 28107 20728 28108 20768
rect 28148 20728 28149 20768
rect 28107 20719 28149 20728
rect 28299 20768 28341 20777
rect 28299 20728 28300 20768
rect 28340 20728 28341 20768
rect 28299 20719 28341 20728
rect 28491 20768 28533 20777
rect 28491 20728 28492 20768
rect 28532 20728 28533 20768
rect 28491 20719 28533 20728
rect 28579 20768 28637 20769
rect 28579 20728 28588 20768
rect 28628 20728 28637 20768
rect 28579 20727 28637 20728
rect 28771 20768 28829 20769
rect 28771 20728 28780 20768
rect 28820 20728 28829 20768
rect 28771 20727 28829 20728
rect 28875 20768 28917 20777
rect 28875 20728 28876 20768
rect 28916 20728 28917 20768
rect 28875 20719 28917 20728
rect 29067 20768 29109 20777
rect 29067 20728 29068 20768
rect 29108 20728 29109 20768
rect 29067 20719 29109 20728
rect 32611 20768 32669 20769
rect 32611 20728 32620 20768
rect 32660 20728 32669 20768
rect 32611 20727 32669 20728
rect 33475 20768 33533 20769
rect 33475 20728 33484 20768
rect 33524 20728 33533 20768
rect 33475 20727 33533 20728
rect 35683 20768 35741 20769
rect 35683 20728 35692 20768
rect 35732 20728 35741 20768
rect 35683 20727 35741 20728
rect 36547 20768 36605 20769
rect 36547 20728 36556 20768
rect 36596 20728 36605 20768
rect 36547 20727 36605 20728
rect 38179 20768 38237 20769
rect 38179 20728 38188 20768
rect 38228 20728 38237 20768
rect 38179 20727 38237 20728
rect 38283 20768 38325 20777
rect 38283 20728 38284 20768
rect 38324 20728 38325 20768
rect 38283 20719 38325 20728
rect 38475 20768 38517 20777
rect 38475 20728 38476 20768
rect 38516 20728 38517 20768
rect 38475 20719 38517 20728
rect 38667 20768 38709 20777
rect 38667 20728 38668 20768
rect 38708 20728 38709 20768
rect 38667 20719 38709 20728
rect 39043 20768 39101 20769
rect 39043 20728 39052 20768
rect 39092 20728 39101 20768
rect 39043 20727 39101 20728
rect 39907 20768 39965 20769
rect 39907 20728 39916 20768
rect 39956 20728 39965 20768
rect 39907 20727 39965 20728
rect 42411 20768 42453 20777
rect 42411 20728 42412 20768
rect 42452 20728 42453 20768
rect 42411 20719 42453 20728
rect 42507 20768 42549 20777
rect 42507 20728 42508 20768
rect 42548 20728 42549 20768
rect 42507 20719 42549 20728
rect 42603 20768 42645 20777
rect 42603 20728 42604 20768
rect 42644 20728 42645 20768
rect 42603 20719 42645 20728
rect 44811 20768 44853 20777
rect 44811 20728 44812 20768
rect 44852 20728 44853 20768
rect 44811 20719 44853 20728
rect 44907 20768 44949 20777
rect 44907 20728 44908 20768
rect 44948 20728 44949 20768
rect 44907 20719 44949 20728
rect 45003 20768 45045 20777
rect 45003 20728 45004 20768
rect 45044 20728 45045 20768
rect 45003 20719 45045 20728
rect 45099 20768 45141 20777
rect 45099 20728 45100 20768
rect 45140 20728 45141 20768
rect 45099 20719 45141 20728
rect 45483 20768 45525 20777
rect 45483 20728 45484 20768
rect 45524 20728 45525 20768
rect 45483 20719 45525 20728
rect 45675 20768 45717 20777
rect 45675 20728 45676 20768
rect 45716 20728 45717 20768
rect 45675 20719 45717 20728
rect 45763 20768 45821 20769
rect 45763 20728 45772 20768
rect 45812 20728 45821 20768
rect 45763 20727 45821 20728
rect 46347 20768 46389 20777
rect 46347 20728 46348 20768
rect 46388 20728 46389 20768
rect 46347 20719 46389 20728
rect 46539 20768 46581 20777
rect 46539 20728 46540 20768
rect 46580 20728 46581 20768
rect 46539 20719 46581 20728
rect 46627 20768 46685 20769
rect 46627 20728 46636 20768
rect 46676 20728 46685 20768
rect 46627 20727 46685 20728
rect 47691 20768 47733 20777
rect 47691 20728 47692 20768
rect 47732 20728 47733 20768
rect 47691 20719 47733 20728
rect 48067 20768 48125 20769
rect 48067 20728 48076 20768
rect 48116 20728 48125 20768
rect 48067 20727 48125 20728
rect 48931 20768 48989 20769
rect 48931 20728 48940 20768
rect 48980 20728 48989 20768
rect 48931 20727 48989 20728
rect 50283 20768 50325 20777
rect 50283 20728 50284 20768
rect 50324 20728 50325 20768
rect 50283 20719 50325 20728
rect 50659 20768 50717 20769
rect 50659 20728 50668 20768
rect 50708 20728 50717 20768
rect 50659 20727 50717 20728
rect 51523 20768 51581 20769
rect 51523 20728 51532 20768
rect 51572 20728 51581 20768
rect 51523 20727 51581 20728
rect 32235 20684 32277 20693
rect 32235 20644 32236 20684
rect 32276 20644 32277 20684
rect 32235 20635 32277 20644
rect 35307 20684 35349 20693
rect 35307 20644 35308 20684
rect 35348 20644 35349 20684
rect 35307 20635 35349 20644
rect 3715 20600 3773 20601
rect 3715 20560 3724 20600
rect 3764 20560 3773 20600
rect 3715 20559 3773 20560
rect 5259 20600 5301 20609
rect 5259 20560 5260 20600
rect 5300 20560 5301 20600
rect 5259 20551 5301 20560
rect 23019 20600 23061 20609
rect 23019 20560 23020 20600
rect 23060 20560 23061 20600
rect 23019 20551 23061 20560
rect 26571 20600 26613 20609
rect 26571 20560 26572 20600
rect 26612 20560 26613 20600
rect 26571 20551 26613 20560
rect 26955 20600 26997 20609
rect 26955 20560 26956 20600
rect 26996 20560 26997 20600
rect 26955 20551 26997 20560
rect 27339 20600 27381 20609
rect 27339 20560 27340 20600
rect 27380 20560 27381 20600
rect 27339 20551 27381 20560
rect 34627 20600 34685 20601
rect 34627 20560 34636 20600
rect 34676 20560 34685 20600
rect 34627 20559 34685 20560
rect 37699 20600 37757 20601
rect 37699 20560 37708 20600
rect 37748 20560 37757 20600
rect 37699 20559 37757 20560
rect 41059 20600 41117 20601
rect 41059 20560 41068 20600
rect 41108 20560 41117 20600
rect 41059 20559 41117 20560
rect 42307 20600 42365 20601
rect 42307 20560 42316 20600
rect 42356 20560 42365 20600
rect 42307 20559 42365 20560
rect 43083 20600 43125 20609
rect 43083 20560 43084 20600
rect 43124 20560 43125 20600
rect 43083 20551 43125 20560
rect 43275 20600 43317 20609
rect 43275 20560 43276 20600
rect 43316 20560 43317 20600
rect 43275 20551 43317 20560
rect 44235 20600 44277 20609
rect 44235 20560 44236 20600
rect 44276 20560 44277 20600
rect 44235 20551 44277 20560
rect 44427 20600 44469 20609
rect 44427 20560 44428 20600
rect 44468 20560 44469 20600
rect 44427 20551 44469 20560
rect 45571 20600 45629 20601
rect 45571 20560 45580 20600
rect 45620 20560 45629 20600
rect 45571 20559 45629 20560
rect 576 20432 52800 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 52800 20432
rect 576 20368 52800 20392
rect 23499 20264 23541 20273
rect 23499 20224 23500 20264
rect 23540 20224 23541 20264
rect 23499 20215 23541 20224
rect 32323 20264 32381 20265
rect 32323 20224 32332 20264
rect 32372 20224 32381 20264
rect 32323 20223 32381 20224
rect 35683 20264 35741 20265
rect 35683 20224 35692 20264
rect 35732 20224 35741 20264
rect 35683 20223 35741 20224
rect 37987 20264 38045 20265
rect 37987 20224 37996 20264
rect 38036 20224 38045 20264
rect 37987 20223 38045 20224
rect 11019 20117 11061 20126
rect 4675 20096 4733 20097
rect 4675 20056 4684 20096
rect 4724 20056 4733 20096
rect 4675 20055 4733 20056
rect 10923 20096 10965 20105
rect 10923 20056 10924 20096
rect 10964 20056 10965 20096
rect 11019 20077 11020 20117
rect 11060 20077 11061 20117
rect 11019 20068 11061 20077
rect 11115 20096 11157 20105
rect 10923 20047 10965 20056
rect 11115 20056 11116 20096
rect 11156 20056 11157 20096
rect 11115 20047 11157 20056
rect 11211 20096 11253 20105
rect 11211 20056 11212 20096
rect 11252 20056 11253 20096
rect 11211 20047 11253 20056
rect 11403 20096 11445 20105
rect 11403 20056 11404 20096
rect 11444 20056 11445 20096
rect 11403 20047 11445 20056
rect 11595 20096 11637 20105
rect 11595 20056 11596 20096
rect 11636 20056 11637 20096
rect 11595 20047 11637 20056
rect 11683 20096 11741 20097
rect 11683 20056 11692 20096
rect 11732 20056 11741 20096
rect 11683 20055 11741 20056
rect 22539 20096 22581 20105
rect 22539 20056 22540 20096
rect 22580 20056 22581 20096
rect 22539 20047 22581 20056
rect 22731 20096 22773 20105
rect 22731 20056 22732 20096
rect 22772 20056 22773 20096
rect 22731 20047 22773 20056
rect 22819 20096 22877 20097
rect 22819 20056 22828 20096
rect 22868 20056 22877 20096
rect 22819 20055 22877 20056
rect 26475 20096 26517 20105
rect 26475 20056 26476 20096
rect 26516 20056 26517 20096
rect 26475 20047 26517 20056
rect 26667 20096 26709 20105
rect 26667 20056 26668 20096
rect 26708 20056 26709 20096
rect 26667 20047 26709 20056
rect 26755 20096 26813 20097
rect 26755 20056 26764 20096
rect 26804 20056 26813 20096
rect 26755 20055 26813 20056
rect 29931 20096 29973 20105
rect 29931 20056 29932 20096
rect 29972 20056 29973 20096
rect 29931 20047 29973 20056
rect 30027 20096 30069 20105
rect 30027 20056 30028 20096
rect 30068 20056 30069 20096
rect 30027 20047 30069 20056
rect 30123 20096 30165 20105
rect 30123 20056 30124 20096
rect 30164 20056 30165 20096
rect 30123 20047 30165 20056
rect 30219 20096 30261 20105
rect 30219 20056 30220 20096
rect 30260 20056 30261 20096
rect 30219 20047 30261 20056
rect 32131 20096 32189 20097
rect 32131 20056 32140 20096
rect 32180 20056 32189 20096
rect 32131 20055 32189 20056
rect 32235 20096 32277 20105
rect 32235 20056 32236 20096
rect 32276 20056 32277 20096
rect 32235 20047 32277 20056
rect 32427 20096 32469 20105
rect 32427 20056 32428 20096
rect 32468 20056 32469 20096
rect 32427 20047 32469 20056
rect 32619 20096 32661 20105
rect 32619 20056 32620 20096
rect 32660 20056 32661 20096
rect 32619 20047 32661 20056
rect 32715 20096 32757 20105
rect 32715 20056 32716 20096
rect 32756 20056 32757 20096
rect 32715 20047 32757 20056
rect 32811 20096 32853 20105
rect 32811 20056 32812 20096
rect 32852 20056 32853 20096
rect 32811 20047 32853 20056
rect 32907 20096 32949 20105
rect 32907 20056 32908 20096
rect 32948 20056 32949 20096
rect 32907 20047 32949 20056
rect 34819 20096 34877 20097
rect 34819 20056 34828 20096
rect 34868 20056 34877 20096
rect 34819 20055 34877 20056
rect 34923 20096 34965 20105
rect 34923 20056 34924 20096
rect 34964 20056 34965 20096
rect 34923 20047 34965 20056
rect 35115 20096 35157 20105
rect 35115 20056 35116 20096
rect 35156 20056 35157 20096
rect 35115 20047 35157 20056
rect 35491 20096 35549 20097
rect 35491 20056 35500 20096
rect 35540 20056 35549 20096
rect 35491 20055 35549 20056
rect 35595 20096 35637 20105
rect 35595 20056 35596 20096
rect 35636 20056 35637 20096
rect 35595 20047 35637 20056
rect 35787 20096 35829 20105
rect 35787 20056 35788 20096
rect 35828 20056 35829 20096
rect 35787 20047 35829 20056
rect 35979 20096 36021 20105
rect 35979 20056 35980 20096
rect 36020 20056 36021 20096
rect 35979 20047 36021 20056
rect 36075 20096 36117 20105
rect 36075 20056 36076 20096
rect 36116 20056 36117 20096
rect 36075 20047 36117 20056
rect 36171 20096 36213 20105
rect 36171 20056 36172 20096
rect 36212 20056 36213 20096
rect 36171 20047 36213 20056
rect 36267 20096 36309 20105
rect 36267 20056 36268 20096
rect 36308 20056 36309 20096
rect 36267 20047 36309 20056
rect 37795 20096 37853 20097
rect 37795 20056 37804 20096
rect 37844 20056 37853 20096
rect 37795 20055 37853 20056
rect 37899 20096 37941 20105
rect 37899 20056 37900 20096
rect 37940 20056 37941 20096
rect 37899 20047 37941 20056
rect 38091 20096 38133 20105
rect 38091 20056 38092 20096
rect 38132 20056 38133 20096
rect 38091 20047 38133 20056
rect 38275 20096 38333 20097
rect 38275 20056 38284 20096
rect 38324 20056 38333 20096
rect 38275 20055 38333 20056
rect 38475 20096 38517 20105
rect 38475 20056 38476 20096
rect 38516 20056 38517 20096
rect 38475 20047 38517 20056
rect 38659 20096 38717 20097
rect 38659 20056 38668 20096
rect 38708 20056 38717 20096
rect 38659 20055 38717 20056
rect 38859 20096 38901 20105
rect 38859 20056 38860 20096
rect 38900 20056 38901 20096
rect 38859 20047 38901 20056
rect 39139 20096 39197 20097
rect 39139 20056 39148 20096
rect 39188 20056 39197 20096
rect 39139 20055 39197 20056
rect 41451 20096 41493 20105
rect 41451 20056 41452 20096
rect 41492 20056 41493 20096
rect 41451 20047 41493 20056
rect 41827 20096 41885 20097
rect 41827 20056 41836 20096
rect 41876 20056 41885 20096
rect 41827 20055 41885 20056
rect 42691 20096 42749 20097
rect 42691 20056 42700 20096
rect 42740 20056 42749 20096
rect 42691 20055 42749 20056
rect 49131 20096 49173 20105
rect 49131 20056 49132 20096
rect 49172 20056 49173 20096
rect 49131 20047 49173 20056
rect 49315 20096 49373 20097
rect 49315 20056 49324 20096
rect 49364 20056 49373 20096
rect 49315 20055 49373 20056
rect 5059 20012 5117 20013
rect 5059 19972 5068 20012
rect 5108 19972 5117 20012
rect 5059 19971 5117 19972
rect 23683 20012 23741 20013
rect 23683 19972 23692 20012
rect 23732 19972 23741 20012
rect 23683 19971 23741 19972
rect 31747 20012 31805 20013
rect 31747 19972 31756 20012
rect 31796 19972 31805 20012
rect 31747 19971 31805 19972
rect 43851 20012 43893 20021
rect 43851 19972 43852 20012
rect 43892 19972 43893 20012
rect 43851 19963 43893 19972
rect 44515 20012 44573 20013
rect 44515 19972 44524 20012
rect 44564 19972 44573 20012
rect 44515 19971 44573 19972
rect 45283 20012 45341 20013
rect 45283 19972 45292 20012
rect 45332 19972 45341 20012
rect 45283 19971 45341 19972
rect 45667 20012 45725 20013
rect 45667 19972 45676 20012
rect 45716 19972 45725 20012
rect 45667 19971 45725 19972
rect 47491 20012 47549 20013
rect 47491 19972 47500 20012
rect 47540 19972 47549 20012
rect 47491 19971 47549 19972
rect 47875 20012 47933 20013
rect 47875 19972 47884 20012
rect 47924 19972 47933 20012
rect 47875 19971 47933 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 9579 19928 9621 19937
rect 9579 19888 9580 19928
rect 9620 19888 9621 19928
rect 9579 19879 9621 19888
rect 12747 19928 12789 19937
rect 12747 19888 12748 19928
rect 12788 19888 12789 19928
rect 12747 19879 12789 19888
rect 23115 19928 23157 19937
rect 23115 19888 23116 19928
rect 23156 19888 23157 19928
rect 23115 19879 23157 19888
rect 26475 19928 26517 19937
rect 26475 19888 26476 19928
rect 26516 19888 26517 19928
rect 26475 19879 26517 19888
rect 26955 19928 26997 19937
rect 26955 19888 26956 19928
rect 26996 19888 26997 19928
rect 26955 19879 26997 19888
rect 29739 19928 29781 19937
rect 29739 19888 29740 19928
rect 29780 19888 29781 19928
rect 29739 19879 29781 19888
rect 33387 19928 33429 19937
rect 33387 19888 33388 19928
rect 33428 19888 33429 19928
rect 33387 19879 33429 19888
rect 35115 19928 35157 19937
rect 35115 19888 35116 19928
rect 35156 19888 35157 19928
rect 35115 19879 35157 19888
rect 40779 19928 40821 19937
rect 40779 19888 40780 19928
rect 40820 19888 40821 19928
rect 40779 19879 40821 19888
rect 44715 19928 44757 19937
rect 44715 19888 44716 19928
rect 44756 19888 44757 19928
rect 44715 19879 44757 19888
rect 46731 19928 46773 19937
rect 46731 19888 46732 19928
rect 46772 19888 46773 19928
rect 46731 19879 46773 19888
rect 50091 19928 50133 19937
rect 50091 19888 50092 19928
rect 50132 19888 50133 19928
rect 50091 19879 50133 19888
rect 4587 19844 4629 19853
rect 4587 19804 4588 19844
rect 4628 19804 4629 19844
rect 4587 19795 4629 19804
rect 4875 19844 4917 19853
rect 4875 19804 4876 19844
rect 4916 19804 4917 19844
rect 4875 19795 4917 19804
rect 11403 19844 11445 19853
rect 11403 19804 11404 19844
rect 11444 19804 11445 19844
rect 11403 19795 11445 19804
rect 22539 19844 22581 19853
rect 22539 19804 22540 19844
rect 22580 19804 22581 19844
rect 22539 19795 22581 19804
rect 31947 19844 31989 19853
rect 31947 19804 31948 19844
rect 31988 19804 31989 19844
rect 31947 19795 31989 19804
rect 38379 19844 38421 19853
rect 38379 19804 38380 19844
rect 38420 19804 38421 19844
rect 38379 19795 38421 19804
rect 38763 19844 38805 19853
rect 38763 19804 38764 19844
rect 38804 19804 38805 19844
rect 38763 19795 38805 19804
rect 44331 19844 44373 19853
rect 44331 19804 44332 19844
rect 44372 19804 44373 19844
rect 44331 19795 44373 19804
rect 45099 19844 45141 19853
rect 45099 19804 45100 19844
rect 45140 19804 45141 19844
rect 45099 19795 45141 19804
rect 45483 19844 45525 19853
rect 45483 19804 45484 19844
rect 45524 19804 45525 19844
rect 45483 19795 45525 19804
rect 47307 19844 47349 19853
rect 47307 19804 47308 19844
rect 47348 19804 47349 19844
rect 47307 19795 47349 19804
rect 47691 19844 47733 19853
rect 47691 19804 47692 19844
rect 47732 19804 47733 19844
rect 47691 19795 47733 19804
rect 49227 19844 49269 19853
rect 49227 19804 49228 19844
rect 49268 19804 49269 19844
rect 49227 19795 49269 19804
rect 576 19676 52800 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 52800 19676
rect 576 19612 52800 19636
rect 14659 19508 14717 19509
rect 14659 19468 14668 19508
rect 14708 19468 14717 19508
rect 14659 19467 14717 19468
rect 32139 19508 32181 19517
rect 32139 19468 32140 19508
rect 32180 19468 32181 19508
rect 32139 19459 32181 19468
rect 35787 19508 35829 19517
rect 35787 19468 35788 19508
rect 35828 19468 35829 19508
rect 35787 19459 35829 19468
rect 39043 19508 39101 19509
rect 39043 19468 39052 19508
rect 39092 19468 39101 19508
rect 39043 19467 39101 19468
rect 40587 19508 40629 19517
rect 40587 19468 40588 19508
rect 40628 19468 40629 19508
rect 40587 19459 40629 19468
rect 48939 19508 48981 19517
rect 48939 19468 48940 19508
rect 48980 19468 48981 19508
rect 48939 19459 48981 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 29067 19424 29109 19433
rect 29067 19384 29068 19424
rect 29108 19384 29109 19424
rect 29067 19375 29109 19384
rect 33571 19424 33629 19425
rect 33571 19384 33580 19424
rect 33620 19384 33629 19424
rect 33571 19383 33629 19384
rect 36067 19424 36125 19425
rect 36067 19384 36076 19424
rect 36116 19384 36125 19424
rect 36067 19383 36125 19384
rect 37035 19424 37077 19433
rect 37035 19384 37036 19424
rect 37076 19384 37077 19424
rect 37035 19375 37077 19384
rect 38379 19424 38421 19433
rect 38379 19384 38380 19424
rect 38420 19384 38421 19424
rect 38379 19375 38421 19384
rect 40395 19424 40437 19433
rect 40395 19384 40396 19424
rect 40436 19384 40437 19424
rect 40395 19375 40437 19384
rect 41259 19424 41301 19433
rect 41259 19384 41260 19424
rect 41300 19384 41301 19424
rect 41259 19375 41301 19384
rect 43459 19424 43517 19425
rect 43459 19384 43468 19424
rect 43508 19384 43517 19424
rect 43459 19383 43517 19384
rect 40771 19351 40829 19352
rect 21763 19340 21821 19341
rect 21763 19300 21772 19340
rect 21812 19300 21821 19340
rect 21763 19299 21821 19300
rect 31659 19340 31701 19349
rect 31659 19300 31660 19340
rect 31700 19300 31701 19340
rect 23011 19292 23069 19293
rect 10051 19256 10109 19257
rect 10051 19216 10060 19256
rect 10100 19216 10109 19256
rect 10051 19215 10109 19216
rect 10915 19256 10973 19257
rect 10915 19216 10924 19256
rect 10964 19216 10973 19256
rect 10915 19215 10973 19216
rect 11307 19256 11349 19265
rect 11307 19216 11308 19256
rect 11348 19216 11349 19256
rect 11307 19207 11349 19216
rect 11787 19256 11829 19265
rect 11787 19216 11788 19256
rect 11828 19216 11829 19256
rect 11787 19207 11829 19216
rect 11979 19256 12021 19265
rect 11979 19216 11980 19256
rect 12020 19216 12021 19256
rect 11979 19207 12021 19216
rect 12067 19256 12125 19257
rect 12067 19216 12076 19256
rect 12116 19216 12125 19256
rect 12067 19215 12125 19216
rect 12643 19256 12701 19257
rect 12643 19216 12652 19256
rect 12692 19216 12701 19256
rect 12643 19215 12701 19216
rect 13507 19256 13565 19257
rect 13507 19216 13516 19256
rect 13556 19216 13565 19256
rect 13507 19215 13565 19216
rect 22155 19256 22197 19265
rect 22155 19216 22156 19256
rect 22196 19216 22197 19256
rect 22155 19207 22197 19216
rect 22251 19256 22293 19265
rect 22251 19216 22252 19256
rect 22292 19216 22293 19256
rect 22251 19207 22293 19216
rect 22347 19256 22389 19265
rect 22347 19216 22348 19256
rect 22388 19216 22389 19256
rect 22347 19207 22389 19216
rect 22443 19256 22485 19265
rect 22443 19216 22444 19256
rect 22484 19216 22485 19256
rect 22443 19207 22485 19216
rect 22635 19256 22677 19265
rect 22635 19216 22636 19256
rect 22676 19216 22677 19256
rect 23011 19252 23020 19292
rect 23060 19252 23069 19292
rect 31659 19291 31701 19300
rect 40195 19340 40253 19341
rect 40195 19300 40204 19340
rect 40244 19300 40253 19340
rect 40771 19311 40780 19351
rect 40820 19311 40829 19351
rect 40771 19310 40829 19311
rect 41539 19340 41597 19341
rect 40195 19299 40253 19300
rect 41539 19300 41548 19340
rect 41588 19300 41597 19340
rect 41539 19299 41597 19300
rect 43171 19298 43229 19299
rect 23011 19251 23069 19252
rect 23875 19256 23933 19257
rect 22635 19207 22677 19216
rect 23875 19216 23884 19256
rect 23924 19216 23933 19256
rect 23875 19215 23933 19216
rect 25219 19256 25277 19257
rect 25219 19216 25228 19256
rect 25268 19216 25277 19256
rect 25219 19215 25277 19216
rect 25323 19256 25365 19265
rect 25323 19216 25324 19256
rect 25364 19216 25365 19256
rect 25323 19207 25365 19216
rect 25515 19256 25557 19265
rect 25515 19216 25516 19256
rect 25556 19216 25557 19256
rect 25515 19207 25557 19216
rect 25803 19256 25845 19265
rect 25803 19216 25804 19256
rect 25844 19216 25845 19256
rect 25803 19207 25845 19216
rect 25899 19256 25941 19265
rect 25899 19216 25900 19256
rect 25940 19216 25941 19256
rect 25899 19207 25941 19216
rect 25995 19256 26037 19265
rect 25995 19216 25996 19256
rect 26036 19216 26037 19256
rect 25995 19207 26037 19216
rect 26563 19256 26621 19257
rect 26563 19216 26572 19256
rect 26612 19216 26621 19256
rect 26563 19215 26621 19216
rect 27427 19256 27485 19257
rect 27427 19216 27436 19256
rect 27476 19216 27485 19256
rect 27427 19215 27485 19216
rect 28771 19256 28829 19257
rect 28771 19216 28780 19256
rect 28820 19216 28829 19256
rect 28771 19215 28829 19216
rect 28875 19256 28917 19265
rect 28875 19216 28876 19256
rect 28916 19216 28917 19256
rect 28875 19207 28917 19216
rect 29067 19256 29109 19265
rect 29067 19216 29068 19256
rect 29108 19216 29109 19256
rect 29067 19207 29109 19216
rect 29259 19256 29301 19265
rect 29259 19216 29260 19256
rect 29300 19216 29301 19256
rect 29259 19207 29301 19216
rect 29635 19256 29693 19257
rect 29635 19216 29644 19256
rect 29684 19216 29693 19256
rect 29635 19215 29693 19216
rect 30499 19256 30557 19257
rect 30499 19216 30508 19256
rect 30548 19216 30557 19256
rect 30499 19215 30557 19216
rect 31843 19256 31901 19257
rect 31843 19216 31852 19256
rect 31892 19216 31901 19256
rect 31843 19215 31901 19216
rect 31947 19256 31989 19265
rect 31947 19216 31948 19256
rect 31988 19216 31989 19256
rect 31947 19207 31989 19216
rect 32139 19256 32181 19265
rect 32139 19216 32140 19256
rect 32180 19216 32181 19256
rect 32139 19207 32181 19216
rect 32899 19256 32957 19257
rect 32899 19216 32908 19256
rect 32948 19216 32957 19256
rect 32899 19215 32957 19216
rect 33195 19256 33237 19265
rect 33195 19216 33196 19256
rect 33236 19216 33237 19256
rect 33195 19207 33237 19216
rect 33291 19256 33333 19265
rect 33291 19216 33292 19256
rect 33332 19216 33333 19256
rect 33291 19207 33333 19216
rect 33771 19256 33813 19265
rect 33771 19216 33772 19256
rect 33812 19216 33813 19256
rect 33771 19207 33813 19216
rect 33955 19256 34013 19257
rect 33955 19216 33964 19256
rect 34004 19216 34013 19256
rect 33955 19215 34013 19216
rect 35683 19256 35741 19257
rect 35683 19216 35692 19256
rect 35732 19216 35741 19256
rect 35683 19215 35741 19216
rect 35883 19256 35925 19265
rect 35883 19216 35884 19256
rect 35924 19216 35925 19256
rect 35883 19207 35925 19216
rect 36363 19256 36405 19265
rect 36363 19216 36364 19256
rect 36404 19216 36405 19256
rect 36363 19207 36405 19216
rect 36459 19256 36501 19265
rect 36459 19216 36460 19256
rect 36500 19216 36501 19256
rect 36459 19207 36501 19216
rect 36739 19256 36797 19257
rect 36739 19216 36748 19256
rect 36788 19216 36797 19256
rect 36739 19215 36797 19216
rect 38571 19256 38613 19265
rect 38571 19216 38572 19256
rect 38612 19216 38613 19256
rect 38571 19207 38613 19216
rect 38763 19256 38805 19265
rect 38763 19216 38764 19256
rect 38804 19216 38805 19256
rect 38763 19207 38805 19216
rect 38851 19256 38909 19257
rect 38851 19216 38860 19256
rect 38900 19216 38909 19256
rect 38851 19215 38909 19216
rect 39339 19256 39381 19265
rect 39339 19216 39340 19256
rect 39380 19216 39381 19256
rect 39339 19207 39381 19216
rect 39435 19256 39477 19265
rect 39435 19216 39436 19256
rect 39476 19216 39477 19256
rect 39435 19207 39477 19216
rect 39715 19256 39773 19257
rect 39715 19216 39724 19256
rect 39764 19216 39773 19256
rect 39715 19215 39773 19216
rect 40963 19256 41021 19257
rect 40963 19216 40972 19256
rect 41012 19216 41021 19256
rect 40963 19215 41021 19216
rect 41067 19256 41109 19265
rect 41067 19216 41068 19256
rect 41108 19216 41109 19256
rect 41067 19207 41109 19216
rect 41259 19256 41301 19265
rect 41259 19216 41260 19256
rect 41300 19216 41301 19256
rect 41259 19207 41301 19216
rect 41923 19256 41981 19257
rect 41923 19216 41932 19256
rect 41972 19216 41981 19256
rect 41923 19215 41981 19216
rect 42027 19256 42069 19265
rect 42027 19216 42028 19256
rect 42068 19216 42069 19256
rect 42027 19207 42069 19216
rect 42219 19256 42261 19265
rect 42219 19216 42220 19256
rect 42260 19216 42261 19256
rect 42219 19207 42261 19216
rect 42787 19256 42845 19257
rect 42787 19216 42796 19256
rect 42836 19216 42845 19256
rect 42787 19215 42845 19216
rect 43083 19256 43125 19265
rect 43171 19258 43180 19298
rect 43220 19258 43229 19298
rect 43171 19257 43229 19258
rect 43083 19216 43084 19256
rect 43124 19216 43125 19256
rect 43083 19207 43125 19216
rect 44035 19256 44093 19257
rect 44035 19216 44044 19256
rect 44084 19216 44093 19256
rect 44035 19215 44093 19216
rect 44899 19256 44957 19257
rect 44899 19216 44908 19256
rect 44948 19216 44957 19256
rect 44899 19215 44957 19216
rect 46627 19256 46685 19257
rect 46627 19216 46636 19256
rect 46676 19216 46685 19256
rect 46627 19215 46685 19216
rect 47491 19256 47549 19257
rect 47491 19216 47500 19256
rect 47540 19216 47549 19256
rect 47491 19215 47549 19216
rect 48939 19256 48981 19265
rect 48939 19216 48940 19256
rect 48980 19216 48981 19256
rect 48939 19207 48981 19216
rect 49131 19256 49173 19265
rect 49131 19216 49132 19256
rect 49172 19216 49173 19256
rect 49131 19207 49173 19216
rect 49219 19256 49277 19257
rect 49219 19216 49228 19256
rect 49268 19216 49277 19256
rect 49219 19215 49277 19216
rect 49611 19256 49653 19265
rect 49611 19216 49612 19256
rect 49652 19216 49653 19256
rect 49611 19207 49653 19216
rect 49987 19256 50045 19257
rect 49987 19216 49996 19256
rect 50036 19216 50045 19256
rect 49987 19215 50045 19216
rect 50851 19256 50909 19257
rect 50851 19216 50860 19256
rect 50900 19216 50909 19256
rect 50851 19215 50909 19216
rect 11883 19172 11925 19181
rect 11883 19132 11884 19172
rect 11924 19132 11925 19172
rect 11883 19123 11925 19132
rect 12267 19172 12309 19181
rect 12267 19132 12268 19172
rect 12308 19132 12309 19172
rect 12267 19123 12309 19132
rect 26187 19172 26229 19181
rect 26187 19132 26188 19172
rect 26228 19132 26229 19172
rect 26187 19123 26229 19132
rect 33867 19172 33909 19181
rect 33867 19132 33868 19172
rect 33908 19132 33909 19172
rect 33867 19123 33909 19132
rect 42123 19172 42165 19181
rect 42123 19132 42124 19172
rect 42164 19132 42165 19172
rect 42123 19123 42165 19132
rect 43659 19172 43701 19181
rect 43659 19132 43660 19172
rect 43700 19132 43701 19172
rect 43659 19123 43701 19132
rect 46251 19172 46293 19181
rect 46251 19132 46252 19172
rect 46292 19132 46293 19172
rect 46251 19123 46293 19132
rect 8899 19088 8957 19089
rect 8899 19048 8908 19088
rect 8948 19048 8957 19088
rect 8899 19047 8957 19048
rect 14659 19088 14717 19089
rect 14659 19048 14668 19088
rect 14708 19048 14717 19088
rect 14659 19047 14717 19048
rect 21963 19088 22005 19097
rect 21963 19048 21964 19088
rect 22004 19048 22005 19088
rect 21963 19039 22005 19048
rect 25027 19088 25085 19089
rect 25027 19048 25036 19088
rect 25076 19048 25085 19088
rect 25027 19047 25085 19048
rect 25411 19088 25469 19089
rect 25411 19048 25420 19088
rect 25460 19048 25469 19088
rect 25411 19047 25469 19048
rect 25699 19088 25757 19089
rect 25699 19048 25708 19088
rect 25748 19048 25757 19088
rect 25699 19047 25757 19048
rect 28579 19088 28637 19089
rect 28579 19048 28588 19088
rect 28628 19048 28637 19088
rect 28579 19047 28637 19048
rect 38659 19088 38717 19089
rect 38659 19048 38668 19088
rect 38708 19048 38717 19088
rect 38659 19047 38717 19048
rect 41739 19088 41781 19097
rect 41739 19048 41740 19088
rect 41780 19048 41781 19088
rect 41739 19039 41781 19048
rect 46051 19088 46109 19089
rect 46051 19048 46060 19088
rect 46100 19048 46109 19088
rect 46051 19047 46109 19048
rect 48643 19088 48701 19089
rect 48643 19048 48652 19088
rect 48692 19048 48701 19088
rect 48643 19047 48701 19048
rect 52003 19088 52061 19089
rect 52003 19048 52012 19088
rect 52052 19048 52061 19088
rect 52003 19047 52061 19048
rect 576 18920 52800 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 52800 18920
rect 576 18856 52800 18880
rect 22539 18752 22581 18761
rect 22539 18712 22540 18752
rect 22580 18712 22581 18752
rect 22539 18703 22581 18712
rect 26275 18752 26333 18753
rect 26275 18712 26284 18752
rect 26324 18712 26333 18752
rect 26275 18711 26333 18712
rect 41155 18752 41213 18753
rect 41155 18712 41164 18752
rect 41204 18712 41213 18752
rect 41155 18711 41213 18712
rect 44035 18752 44093 18753
rect 44035 18712 44044 18752
rect 44084 18712 44093 18752
rect 44035 18711 44093 18712
rect 11019 18668 11061 18677
rect 11019 18628 11020 18668
rect 11060 18628 11061 18668
rect 11019 18619 11061 18628
rect 11595 18668 11637 18677
rect 11595 18628 11596 18668
rect 11636 18628 11637 18668
rect 11595 18619 11637 18628
rect 12171 18668 12213 18677
rect 12171 18628 12172 18668
rect 12212 18628 12213 18668
rect 12171 18619 12213 18628
rect 23019 18668 23061 18677
rect 23019 18628 23020 18668
rect 23060 18628 23061 18668
rect 23019 18619 23061 18628
rect 27243 18668 27285 18677
rect 27243 18628 27244 18668
rect 27284 18628 27285 18668
rect 27243 18619 27285 18628
rect 28875 18668 28917 18677
rect 28875 18628 28876 18668
rect 28916 18628 28917 18668
rect 28875 18619 28917 18628
rect 29739 18668 29781 18677
rect 29739 18628 29740 18668
rect 29780 18628 29781 18668
rect 29739 18619 29781 18628
rect 30315 18668 30357 18677
rect 30315 18628 30316 18668
rect 30356 18628 30357 18668
rect 30315 18619 30357 18628
rect 32523 18668 32565 18677
rect 32523 18628 32524 18668
rect 32564 18628 32565 18668
rect 32523 18619 32565 18628
rect 32907 18668 32949 18677
rect 32907 18628 32908 18668
rect 32948 18628 32949 18668
rect 32907 18619 32949 18628
rect 35787 18668 35829 18677
rect 35787 18628 35788 18668
rect 35828 18628 35829 18668
rect 35787 18619 35829 18628
rect 36171 18668 36213 18677
rect 36171 18628 36172 18668
rect 36212 18628 36213 18668
rect 36171 18619 36213 18628
rect 38763 18668 38805 18677
rect 38763 18628 38764 18668
rect 38804 18628 38805 18668
rect 38763 18619 38805 18628
rect 43659 18668 43701 18677
rect 43659 18628 43660 18668
rect 43700 18628 43701 18668
rect 43659 18619 43701 18628
rect 49323 18668 49365 18677
rect 49323 18628 49324 18668
rect 49364 18628 49365 18668
rect 49323 18619 49365 18628
rect 49219 18605 49277 18606
rect 10627 18584 10685 18585
rect 10627 18544 10636 18584
rect 10676 18544 10685 18584
rect 10627 18543 10685 18544
rect 10923 18584 10965 18593
rect 10923 18544 10924 18584
rect 10964 18544 10965 18584
rect 10923 18535 10965 18544
rect 11499 18584 11541 18593
rect 11499 18544 11500 18584
rect 11540 18544 11541 18584
rect 11499 18535 11541 18544
rect 11683 18584 11741 18585
rect 11683 18544 11692 18584
rect 11732 18544 11741 18584
rect 11683 18543 11741 18544
rect 12067 18584 12125 18585
rect 12067 18544 12076 18584
rect 12116 18544 12125 18584
rect 12067 18543 12125 18544
rect 12267 18584 12309 18593
rect 12267 18544 12268 18584
rect 12308 18544 12309 18584
rect 12267 18535 12309 18544
rect 23115 18584 23157 18593
rect 23115 18544 23116 18584
rect 23156 18544 23157 18584
rect 23115 18535 23157 18544
rect 23395 18584 23453 18585
rect 23395 18544 23404 18584
rect 23444 18544 23453 18584
rect 23395 18543 23453 18544
rect 26187 18584 26229 18593
rect 26187 18544 26188 18584
rect 26228 18544 26229 18584
rect 26187 18535 26229 18544
rect 26379 18584 26421 18593
rect 26379 18544 26380 18584
rect 26420 18544 26421 18584
rect 26379 18535 26421 18544
rect 26467 18584 26525 18585
rect 26467 18544 26476 18584
rect 26516 18544 26525 18584
rect 26467 18543 26525 18544
rect 26851 18584 26909 18585
rect 26851 18544 26860 18584
rect 26900 18544 26909 18584
rect 26851 18543 26909 18544
rect 27147 18584 27189 18593
rect 27147 18544 27148 18584
rect 27188 18544 27189 18584
rect 27147 18535 27189 18544
rect 27723 18584 27765 18593
rect 27723 18544 27724 18584
rect 27764 18544 27765 18584
rect 27723 18535 27765 18544
rect 27819 18584 27861 18593
rect 27819 18544 27820 18584
rect 27860 18544 27861 18584
rect 27819 18535 27861 18544
rect 27907 18584 27965 18585
rect 27907 18544 27916 18584
rect 27956 18544 27965 18584
rect 27907 18543 27965 18544
rect 28675 18584 28733 18585
rect 28675 18544 28684 18584
rect 28724 18544 28733 18584
rect 28675 18543 28733 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 28779 18535 28821 18544
rect 28971 18584 29013 18593
rect 28971 18544 28972 18584
rect 29012 18544 29013 18584
rect 28971 18535 29013 18544
rect 29635 18584 29693 18585
rect 29635 18544 29644 18584
rect 29684 18544 29693 18584
rect 29635 18543 29693 18544
rect 29835 18584 29877 18593
rect 29835 18544 29836 18584
rect 29876 18544 29877 18584
rect 29835 18535 29877 18544
rect 30411 18584 30453 18593
rect 30411 18544 30412 18584
rect 30452 18544 30453 18584
rect 30411 18535 30453 18544
rect 30691 18584 30749 18585
rect 30691 18544 30700 18584
rect 30740 18544 30749 18584
rect 30691 18543 30749 18544
rect 31179 18584 31221 18593
rect 31179 18544 31180 18584
rect 31220 18544 31221 18584
rect 31179 18535 31221 18544
rect 32427 18584 32469 18593
rect 32427 18544 32428 18584
rect 32468 18544 32469 18584
rect 32427 18535 32469 18544
rect 32619 18584 32661 18593
rect 32619 18544 32620 18584
rect 32660 18544 32661 18584
rect 32619 18535 32661 18544
rect 32707 18584 32765 18585
rect 32707 18544 32716 18584
rect 32756 18544 32765 18584
rect 32707 18543 32765 18544
rect 33283 18584 33341 18585
rect 33283 18544 33292 18584
rect 33332 18544 33341 18584
rect 33283 18543 33341 18544
rect 34147 18584 34205 18585
rect 34147 18544 34156 18584
rect 34196 18544 34205 18584
rect 34147 18543 34205 18544
rect 35691 18584 35733 18593
rect 35691 18544 35692 18584
rect 35732 18544 35733 18584
rect 35691 18535 35733 18544
rect 35883 18584 35925 18593
rect 35883 18544 35884 18584
rect 35924 18544 35925 18584
rect 35883 18535 35925 18544
rect 35971 18584 36029 18585
rect 35971 18544 35980 18584
rect 36020 18544 36029 18584
rect 35971 18543 36029 18544
rect 36547 18584 36605 18585
rect 36547 18544 36556 18584
rect 36596 18544 36605 18584
rect 36547 18543 36605 18544
rect 37411 18584 37469 18585
rect 37411 18544 37420 18584
rect 37460 18544 37469 18584
rect 37411 18543 37469 18544
rect 39139 18584 39197 18585
rect 39139 18544 39148 18584
rect 39188 18544 39197 18584
rect 39139 18543 39197 18544
rect 40003 18584 40061 18585
rect 40003 18544 40012 18584
rect 40052 18544 40061 18584
rect 40003 18543 40061 18544
rect 41931 18584 41973 18593
rect 41931 18544 41932 18584
rect 41972 18544 41973 18584
rect 41931 18535 41973 18544
rect 42123 18584 42165 18593
rect 42123 18544 42124 18584
rect 42164 18544 42165 18584
rect 42123 18535 42165 18544
rect 42211 18584 42269 18585
rect 42211 18544 42220 18584
rect 42260 18544 42269 18584
rect 42211 18543 42269 18544
rect 42411 18584 42453 18593
rect 42411 18544 42412 18584
rect 42452 18544 42453 18584
rect 42411 18535 42453 18544
rect 42603 18584 42645 18593
rect 42603 18544 42604 18584
rect 42644 18544 42645 18584
rect 42603 18535 42645 18544
rect 42691 18584 42749 18585
rect 42691 18544 42700 18584
rect 42740 18544 42749 18584
rect 42691 18543 42749 18544
rect 43563 18584 43605 18593
rect 43563 18544 43564 18584
rect 43604 18544 43605 18584
rect 43563 18535 43605 18544
rect 43747 18584 43805 18585
rect 43747 18544 43756 18584
rect 43796 18544 43805 18584
rect 43747 18543 43805 18544
rect 43947 18584 43989 18593
rect 43947 18544 43948 18584
rect 43988 18544 43989 18584
rect 43947 18535 43989 18544
rect 44139 18584 44181 18593
rect 44139 18544 44140 18584
rect 44180 18544 44181 18584
rect 44139 18535 44181 18544
rect 44227 18584 44285 18585
rect 44227 18544 44236 18584
rect 44276 18544 44285 18584
rect 44227 18543 44285 18544
rect 44419 18584 44477 18585
rect 44419 18544 44428 18584
rect 44468 18544 44477 18584
rect 44419 18543 44477 18544
rect 44619 18584 44661 18593
rect 44619 18544 44620 18584
rect 44660 18544 44661 18584
rect 44619 18535 44661 18544
rect 46723 18584 46781 18585
rect 46723 18544 46732 18584
rect 46772 18544 46781 18584
rect 46723 18543 46781 18544
rect 46827 18584 46869 18593
rect 46827 18544 46828 18584
rect 46868 18544 46869 18584
rect 46827 18535 46869 18544
rect 47019 18584 47061 18593
rect 47019 18544 47020 18584
rect 47060 18544 47061 18584
rect 47019 18535 47061 18544
rect 47403 18584 47445 18593
rect 47403 18544 47404 18584
rect 47444 18544 47445 18584
rect 47403 18535 47445 18544
rect 47499 18584 47541 18593
rect 47499 18544 47500 18584
rect 47540 18544 47541 18584
rect 47499 18535 47541 18544
rect 47595 18584 47637 18593
rect 47595 18544 47596 18584
rect 47636 18544 47637 18584
rect 47595 18535 47637 18544
rect 47691 18584 47733 18593
rect 47691 18544 47692 18584
rect 47732 18544 47733 18584
rect 47691 18535 47733 18544
rect 48355 18584 48413 18585
rect 48355 18544 48364 18584
rect 48404 18544 48413 18584
rect 48355 18543 48413 18544
rect 48651 18584 48693 18593
rect 48651 18544 48652 18584
rect 48692 18544 48693 18584
rect 48651 18535 48693 18544
rect 48747 18584 48789 18593
rect 48747 18544 48748 18584
rect 48788 18544 48789 18584
rect 49219 18565 49228 18605
rect 49268 18565 49277 18605
rect 49219 18564 49277 18565
rect 49419 18584 49461 18593
rect 48747 18535 48789 18544
rect 49419 18544 49420 18584
rect 49460 18544 49461 18584
rect 49419 18535 49461 18544
rect 52291 18584 52349 18585
rect 52291 18544 52300 18584
rect 52340 18544 52349 18584
rect 52291 18543 52349 18544
rect 52675 18584 52733 18585
rect 52675 18544 52684 18584
rect 52724 18544 52733 18584
rect 52675 18543 52733 18544
rect 1699 18500 1757 18501
rect 1699 18460 1708 18500
rect 1748 18460 1757 18500
rect 1699 18459 1757 18460
rect 21955 18500 22013 18501
rect 21955 18460 21964 18500
rect 22004 18460 22013 18500
rect 21955 18459 22013 18460
rect 22339 18500 22397 18501
rect 22339 18460 22348 18500
rect 22388 18460 22397 18500
rect 22339 18459 22397 18460
rect 23683 18500 23741 18501
rect 23683 18460 23692 18500
rect 23732 18460 23741 18500
rect 23683 18459 23741 18460
rect 24067 18500 24125 18501
rect 24067 18460 24076 18500
rect 24116 18460 24125 18500
rect 24067 18459 24125 18460
rect 24451 18500 24509 18501
rect 24451 18460 24460 18500
rect 24500 18460 24509 18500
rect 24451 18459 24509 18460
rect 24835 18500 24893 18501
rect 24835 18460 24844 18500
rect 24884 18460 24893 18500
rect 24835 18459 24893 18460
rect 25699 18500 25757 18501
rect 25699 18460 25708 18500
rect 25748 18460 25757 18500
rect 25699 18459 25757 18460
rect 35307 18500 35349 18509
rect 35307 18460 35308 18500
rect 35348 18460 35349 18500
rect 35307 18451 35349 18460
rect 41731 18500 41789 18501
rect 41731 18460 41740 18500
rect 41780 18460 41789 18500
rect 41731 18459 41789 18460
rect 43075 18500 43133 18501
rect 43075 18460 43084 18500
rect 43124 18460 43133 18500
rect 43075 18459 43133 18460
rect 49795 18500 49853 18501
rect 49795 18460 49804 18500
rect 49844 18460 49853 18500
rect 49795 18459 49853 18460
rect 50467 18500 50525 18501
rect 50467 18460 50476 18500
rect 50516 18460 50525 18500
rect 50467 18459 50525 18460
rect 51331 18500 51389 18501
rect 51331 18460 51340 18500
rect 51380 18460 51389 18500
rect 51331 18459 51389 18460
rect 51523 18500 51581 18501
rect 51523 18460 51532 18500
rect 51572 18460 51581 18500
rect 51523 18459 51581 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 11299 18416 11357 18417
rect 11299 18376 11308 18416
rect 11348 18376 11357 18416
rect 11299 18375 11357 18376
rect 22155 18416 22197 18425
rect 22155 18376 22156 18416
rect 22196 18376 22197 18416
rect 22155 18367 22197 18376
rect 25515 18416 25557 18425
rect 25515 18376 25516 18416
rect 25556 18376 25557 18416
rect 25515 18367 25557 18376
rect 27523 18416 27581 18417
rect 27523 18376 27532 18416
rect 27572 18376 27581 18416
rect 27523 18375 27581 18376
rect 30019 18416 30077 18417
rect 30019 18376 30028 18416
rect 30068 18376 30077 18416
rect 30019 18375 30077 18376
rect 41547 18416 41589 18425
rect 41547 18376 41548 18416
rect 41588 18376 41589 18416
rect 41547 18367 41589 18376
rect 44523 18416 44565 18425
rect 44523 18376 44524 18416
rect 44564 18376 44565 18416
rect 44523 18367 44565 18376
rect 47019 18416 47061 18425
rect 47019 18376 47020 18416
rect 47060 18376 47061 18416
rect 47019 18367 47061 18376
rect 49027 18416 49085 18417
rect 49027 18376 49036 18416
rect 49076 18376 49085 18416
rect 49027 18375 49085 18376
rect 50763 18416 50805 18425
rect 50763 18376 50764 18416
rect 50804 18376 50805 18416
rect 50763 18367 50805 18376
rect 1515 18332 1557 18341
rect 1515 18292 1516 18332
rect 1556 18292 1557 18332
rect 1515 18283 1557 18292
rect 22723 18332 22781 18333
rect 22723 18292 22732 18332
rect 22772 18292 22781 18332
rect 22723 18291 22781 18292
rect 23883 18332 23925 18341
rect 23883 18292 23884 18332
rect 23924 18292 23925 18332
rect 23883 18283 23925 18292
rect 24267 18332 24309 18341
rect 24267 18292 24268 18332
rect 24308 18292 24309 18332
rect 24267 18283 24309 18292
rect 24651 18332 24693 18341
rect 24651 18292 24652 18332
rect 24692 18292 24693 18332
rect 24651 18283 24693 18292
rect 25035 18332 25077 18341
rect 25035 18292 25036 18332
rect 25076 18292 25077 18332
rect 25035 18283 25077 18292
rect 31563 18332 31605 18341
rect 31563 18292 31564 18332
rect 31604 18292 31605 18332
rect 31563 18283 31605 18292
rect 38563 18332 38621 18333
rect 38563 18292 38572 18332
rect 38612 18292 38621 18332
rect 38563 18291 38621 18292
rect 41155 18332 41213 18333
rect 41155 18292 41164 18332
rect 41204 18292 41213 18332
rect 41155 18291 41213 18292
rect 41931 18332 41973 18341
rect 41931 18292 41932 18332
rect 41972 18292 41973 18332
rect 41931 18283 41973 18292
rect 42411 18332 42453 18341
rect 42411 18292 42412 18332
rect 42452 18292 42453 18332
rect 42411 18283 42453 18292
rect 42891 18332 42933 18341
rect 42891 18292 42892 18332
rect 42932 18292 42933 18332
rect 42891 18283 42933 18292
rect 49995 18332 50037 18341
rect 49995 18292 49996 18332
rect 50036 18292 50037 18332
rect 49995 18283 50037 18292
rect 50283 18332 50325 18341
rect 50283 18292 50284 18332
rect 50324 18292 50325 18332
rect 50283 18283 50325 18292
rect 51147 18332 51189 18341
rect 51147 18292 51148 18332
rect 51188 18292 51189 18332
rect 51147 18283 51189 18292
rect 51723 18332 51765 18341
rect 51723 18292 51724 18332
rect 51764 18292 51765 18332
rect 51723 18283 51765 18292
rect 52395 18332 52437 18341
rect 52395 18292 52396 18332
rect 52436 18292 52437 18332
rect 52395 18283 52437 18292
rect 52587 18332 52629 18341
rect 52587 18292 52588 18332
rect 52628 18292 52629 18332
rect 52587 18283 52629 18292
rect 576 18164 52800 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 52800 18164
rect 576 18100 52800 18124
rect 33387 17996 33429 18005
rect 33387 17956 33388 17996
rect 33428 17956 33429 17996
rect 33387 17947 33429 17956
rect 36555 17996 36597 18005
rect 36555 17956 36556 17996
rect 36596 17956 36597 17996
rect 36555 17947 36597 17956
rect 37035 17996 37077 18005
rect 37035 17956 37036 17996
rect 37076 17956 37077 17996
rect 37035 17947 37077 17956
rect 46443 17996 46485 18005
rect 46443 17956 46444 17996
rect 46484 17956 46485 17996
rect 46443 17947 46485 17956
rect 50091 17996 50133 18005
rect 50091 17956 50092 17996
rect 50132 17956 50133 17996
rect 50091 17947 50133 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 23211 17912 23253 17921
rect 23211 17872 23212 17912
rect 23252 17872 23253 17912
rect 23211 17863 23253 17872
rect 34827 17912 34869 17921
rect 34827 17872 34828 17912
rect 34868 17872 34869 17912
rect 34827 17863 34869 17872
rect 37899 17912 37941 17921
rect 37899 17872 37900 17912
rect 37940 17872 37941 17912
rect 37899 17863 37941 17872
rect 39435 17912 39477 17921
rect 39435 17872 39436 17912
rect 39476 17872 39477 17912
rect 39435 17863 39477 17872
rect 22635 17828 22677 17837
rect 22635 17788 22636 17828
rect 22676 17788 22677 17828
rect 22635 17779 22677 17788
rect 34339 17828 34397 17829
rect 34339 17788 34348 17828
rect 34388 17788 34397 17828
rect 34339 17787 34397 17788
rect 36835 17828 36893 17829
rect 36835 17788 36844 17828
rect 36884 17788 36893 17828
rect 36835 17787 36893 17788
rect 46819 17828 46877 17829
rect 46819 17788 46828 17828
rect 46868 17788 46877 17828
rect 46819 17787 46877 17788
rect 49515 17828 49557 17837
rect 49515 17788 49516 17828
rect 49556 17788 49557 17828
rect 49515 17779 49557 17788
rect 23011 17758 23069 17759
rect 22539 17744 22581 17753
rect 22539 17704 22540 17744
rect 22580 17704 22581 17744
rect 22539 17695 22581 17704
rect 22723 17744 22781 17745
rect 22723 17704 22732 17744
rect 22772 17704 22781 17744
rect 22723 17703 22781 17704
rect 22915 17744 22973 17745
rect 22915 17704 22924 17744
rect 22964 17704 22973 17744
rect 23011 17718 23020 17758
rect 23060 17718 23069 17758
rect 23011 17717 23069 17718
rect 23211 17744 23253 17753
rect 22915 17703 22973 17704
rect 23211 17704 23212 17744
rect 23252 17704 23253 17744
rect 23211 17695 23253 17704
rect 23403 17744 23445 17753
rect 23403 17704 23404 17744
rect 23444 17704 23445 17744
rect 23403 17695 23445 17704
rect 23779 17744 23837 17745
rect 23779 17704 23788 17744
rect 23828 17704 23837 17744
rect 23779 17703 23837 17704
rect 24643 17744 24701 17745
rect 24643 17704 24652 17744
rect 24692 17704 24701 17744
rect 24643 17703 24701 17704
rect 26667 17744 26709 17753
rect 26667 17704 26668 17744
rect 26708 17704 26709 17744
rect 26667 17695 26709 17704
rect 26859 17744 26901 17753
rect 26859 17704 26860 17744
rect 26900 17704 26901 17744
rect 26859 17695 26901 17704
rect 26947 17744 27005 17745
rect 26947 17704 26956 17744
rect 26996 17704 27005 17744
rect 26947 17703 27005 17704
rect 27523 17744 27581 17745
rect 27523 17704 27532 17744
rect 27572 17704 27581 17744
rect 27523 17703 27581 17704
rect 28387 17744 28445 17745
rect 28387 17704 28396 17744
rect 28436 17704 28445 17744
rect 28387 17703 28445 17704
rect 29835 17744 29877 17753
rect 29835 17704 29836 17744
rect 29876 17704 29877 17744
rect 29835 17695 29877 17704
rect 30027 17744 30069 17753
rect 30027 17704 30028 17744
rect 30068 17704 30069 17744
rect 30027 17695 30069 17704
rect 30115 17744 30173 17745
rect 30115 17704 30124 17744
rect 30164 17704 30173 17744
rect 30115 17703 30173 17704
rect 30691 17744 30749 17745
rect 30691 17704 30700 17744
rect 30740 17704 30749 17744
rect 30691 17703 30749 17704
rect 31555 17744 31613 17745
rect 31555 17704 31564 17744
rect 31604 17704 31613 17744
rect 31555 17703 31613 17704
rect 33283 17744 33341 17745
rect 33283 17704 33292 17744
rect 33332 17704 33341 17744
rect 33283 17703 33341 17704
rect 33483 17744 33525 17753
rect 33483 17704 33484 17744
rect 33524 17704 33525 17744
rect 33483 17695 33525 17704
rect 36451 17744 36509 17745
rect 36451 17704 36460 17744
rect 36500 17704 36509 17744
rect 36451 17703 36509 17704
rect 36651 17744 36693 17753
rect 36651 17704 36652 17744
rect 36692 17704 36693 17744
rect 36651 17695 36693 17704
rect 39819 17744 39861 17753
rect 39819 17704 39820 17744
rect 39860 17704 39861 17744
rect 39819 17695 39861 17704
rect 40195 17744 40253 17745
rect 40195 17704 40204 17744
rect 40244 17704 40253 17744
rect 40195 17703 40253 17704
rect 41059 17744 41117 17745
rect 41059 17704 41068 17744
rect 41108 17704 41117 17744
rect 41059 17703 41117 17704
rect 42603 17744 42645 17753
rect 42603 17704 42604 17744
rect 42644 17704 42645 17744
rect 42603 17695 42645 17704
rect 42795 17744 42837 17753
rect 42795 17704 42796 17744
rect 42836 17704 42837 17744
rect 42795 17695 42837 17704
rect 42883 17744 42941 17745
rect 42883 17704 42892 17744
rect 42932 17704 42941 17744
rect 42883 17703 42941 17704
rect 43459 17744 43517 17745
rect 43459 17704 43468 17744
rect 43508 17704 43517 17744
rect 43459 17703 43517 17704
rect 44323 17744 44381 17745
rect 44323 17704 44332 17744
rect 44372 17704 44381 17744
rect 44323 17703 44381 17704
rect 45771 17744 45813 17753
rect 45771 17704 45772 17744
rect 45812 17704 45813 17744
rect 45771 17695 45813 17704
rect 45955 17744 46013 17745
rect 45955 17704 45964 17744
rect 46004 17704 46013 17744
rect 45955 17703 46013 17704
rect 46147 17744 46205 17745
rect 46147 17704 46156 17744
rect 46196 17704 46205 17744
rect 46147 17703 46205 17704
rect 46251 17744 46293 17753
rect 46251 17704 46252 17744
rect 46292 17704 46293 17744
rect 46251 17695 46293 17704
rect 46443 17744 46485 17753
rect 46443 17704 46444 17744
rect 46484 17704 46485 17744
rect 46443 17695 46485 17704
rect 48643 17744 48701 17745
rect 48643 17704 48652 17744
rect 48692 17704 48701 17744
rect 48643 17703 48701 17704
rect 48747 17744 48789 17753
rect 48747 17704 48748 17744
rect 48788 17704 48789 17744
rect 48747 17695 48789 17704
rect 48939 17744 48981 17753
rect 48939 17704 48940 17744
rect 48980 17704 48981 17744
rect 48939 17695 48981 17704
rect 49419 17744 49461 17753
rect 49419 17704 49420 17744
rect 49460 17704 49461 17744
rect 49419 17695 49461 17704
rect 49603 17744 49661 17745
rect 49603 17704 49612 17744
rect 49652 17704 49661 17744
rect 49603 17703 49661 17704
rect 49795 17744 49853 17745
rect 49795 17704 49804 17744
rect 49844 17704 49853 17744
rect 49795 17703 49853 17704
rect 49899 17744 49941 17753
rect 49899 17704 49900 17744
rect 49940 17704 49941 17744
rect 49899 17695 49941 17704
rect 50091 17744 50133 17753
rect 50091 17704 50092 17744
rect 50132 17704 50133 17744
rect 50091 17695 50133 17704
rect 50283 17744 50325 17753
rect 50283 17704 50284 17744
rect 50324 17704 50325 17744
rect 50283 17695 50325 17704
rect 50659 17744 50717 17745
rect 50659 17704 50668 17744
rect 50708 17704 50717 17744
rect 50659 17703 50717 17704
rect 51523 17744 51581 17745
rect 51523 17704 51532 17744
rect 51572 17704 51581 17744
rect 51523 17703 51581 17704
rect 27147 17660 27189 17669
rect 27147 17620 27148 17660
rect 27188 17620 27189 17660
rect 27147 17611 27189 17620
rect 29931 17660 29973 17669
rect 29931 17620 29932 17660
rect 29972 17620 29973 17660
rect 29931 17611 29973 17620
rect 30315 17660 30357 17669
rect 30315 17620 30316 17660
rect 30356 17620 30357 17660
rect 30315 17611 30357 17620
rect 42699 17660 42741 17669
rect 42699 17620 42700 17660
rect 42740 17620 42741 17660
rect 42699 17611 42741 17620
rect 43083 17660 43125 17669
rect 43083 17620 43084 17660
rect 43124 17620 43125 17660
rect 43083 17611 43125 17620
rect 45867 17660 45909 17669
rect 45867 17620 45868 17660
rect 45908 17620 45909 17660
rect 45867 17611 45909 17620
rect 25795 17576 25853 17577
rect 25795 17536 25804 17576
rect 25844 17536 25853 17576
rect 25795 17535 25853 17536
rect 26755 17576 26813 17577
rect 26755 17536 26764 17576
rect 26804 17536 26813 17576
rect 26755 17535 26813 17536
rect 29539 17576 29597 17577
rect 29539 17536 29548 17576
rect 29588 17536 29597 17576
rect 29539 17535 29597 17536
rect 32707 17576 32765 17577
rect 32707 17536 32716 17576
rect 32756 17536 32765 17576
rect 32707 17535 32765 17536
rect 34155 17576 34197 17585
rect 34155 17536 34156 17576
rect 34196 17536 34197 17576
rect 34155 17527 34197 17536
rect 37035 17576 37077 17585
rect 37035 17536 37036 17576
rect 37076 17536 37077 17576
rect 37035 17527 37077 17536
rect 42211 17576 42269 17577
rect 42211 17536 42220 17576
rect 42260 17536 42269 17576
rect 42211 17535 42269 17536
rect 45475 17576 45533 17577
rect 45475 17536 45484 17576
rect 45524 17536 45533 17576
rect 45475 17535 45533 17536
rect 46635 17576 46677 17585
rect 46635 17536 46636 17576
rect 46676 17536 46677 17576
rect 46635 17527 46677 17536
rect 48835 17576 48893 17577
rect 48835 17536 48844 17576
rect 48884 17536 48893 17576
rect 48835 17535 48893 17536
rect 52675 17576 52733 17577
rect 52675 17536 52684 17576
rect 52724 17536 52733 17576
rect 52675 17535 52733 17536
rect 576 17408 52800 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 52800 17408
rect 576 17344 52800 17368
rect 23211 17240 23253 17249
rect 23211 17200 23212 17240
rect 23252 17200 23253 17240
rect 23211 17191 23253 17200
rect 41635 17240 41693 17241
rect 41635 17200 41644 17240
rect 41684 17200 41693 17240
rect 41635 17199 41693 17200
rect 51435 17240 51477 17249
rect 51435 17200 51436 17240
rect 51476 17200 51477 17240
rect 51435 17191 51477 17200
rect 52683 17240 52725 17249
rect 52683 17200 52684 17240
rect 52724 17200 52725 17240
rect 52683 17191 52725 17200
rect 23691 17156 23733 17165
rect 23691 17116 23692 17156
rect 23732 17116 23733 17156
rect 23691 17107 23733 17116
rect 27339 17156 27381 17165
rect 27339 17116 27340 17156
rect 27380 17116 27381 17156
rect 27339 17107 27381 17116
rect 30507 17156 30549 17165
rect 30507 17116 30508 17156
rect 30548 17116 30549 17156
rect 30507 17107 30549 17116
rect 42603 17156 42645 17165
rect 42603 17116 42604 17156
rect 42644 17116 42645 17156
rect 42603 17107 42645 17116
rect 44043 17156 44085 17165
rect 44043 17116 44044 17156
rect 44084 17116 44085 17156
rect 44043 17107 44085 17116
rect 45771 17156 45813 17165
rect 45771 17116 45772 17156
rect 45812 17116 45813 17156
rect 45771 17107 45813 17116
rect 51723 17156 51765 17165
rect 51723 17116 51724 17156
rect 51764 17116 51765 17156
rect 51723 17107 51765 17116
rect 4203 17072 4245 17081
rect 4203 17032 4204 17072
rect 4244 17032 4245 17072
rect 4203 17023 4245 17032
rect 4387 17072 4445 17073
rect 4387 17032 4396 17072
rect 4436 17032 4445 17072
rect 4387 17031 4445 17032
rect 23595 17072 23637 17081
rect 23595 17032 23596 17072
rect 23636 17032 23637 17072
rect 23595 17023 23637 17032
rect 23779 17072 23837 17073
rect 23779 17032 23788 17072
rect 23828 17032 23837 17072
rect 23779 17031 23837 17032
rect 27235 17072 27293 17073
rect 27235 17032 27244 17072
rect 27284 17032 27293 17072
rect 27235 17031 27293 17032
rect 27435 17072 27477 17081
rect 27435 17032 27436 17072
rect 27476 17032 27477 17072
rect 27435 17023 27477 17032
rect 30403 17072 30461 17073
rect 30403 17032 30412 17072
rect 30452 17032 30461 17072
rect 30403 17031 30461 17032
rect 30603 17072 30645 17081
rect 30603 17032 30604 17072
rect 30644 17032 30645 17072
rect 30603 17023 30645 17032
rect 33379 17072 33437 17073
rect 33379 17032 33388 17072
rect 33428 17032 33437 17072
rect 33379 17031 33437 17032
rect 33579 17072 33621 17081
rect 33579 17032 33580 17072
rect 33620 17032 33621 17072
rect 33579 17023 33621 17032
rect 33763 17072 33821 17073
rect 33763 17032 33772 17072
rect 33812 17032 33821 17072
rect 33763 17031 33821 17032
rect 33867 17072 33909 17081
rect 33867 17032 33868 17072
rect 33908 17032 33909 17072
rect 33867 17023 33909 17032
rect 34059 17072 34101 17081
rect 34059 17032 34060 17072
rect 34100 17032 34101 17072
rect 34059 17023 34101 17032
rect 34251 17072 34293 17081
rect 34251 17032 34252 17072
rect 34292 17032 34293 17072
rect 34251 17023 34293 17032
rect 34627 17072 34685 17073
rect 34627 17032 34636 17072
rect 34676 17032 34685 17072
rect 34627 17031 34685 17032
rect 35491 17072 35549 17073
rect 35491 17032 35500 17072
rect 35540 17032 35549 17072
rect 35491 17031 35549 17032
rect 36931 17072 36989 17073
rect 36931 17032 36940 17072
rect 36980 17032 36989 17072
rect 36931 17031 36989 17032
rect 37131 17072 37173 17081
rect 37131 17032 37132 17072
rect 37172 17032 37173 17072
rect 37131 17023 37173 17032
rect 37323 17072 37365 17081
rect 37323 17032 37324 17072
rect 37364 17032 37365 17072
rect 37323 17023 37365 17032
rect 37699 17072 37757 17073
rect 37699 17032 37708 17072
rect 37748 17032 37757 17072
rect 37699 17031 37757 17032
rect 38563 17072 38621 17073
rect 38563 17032 38572 17072
rect 38612 17032 38621 17072
rect 38563 17031 38621 17032
rect 41739 17072 41781 17081
rect 41739 17032 41740 17072
rect 41780 17032 41781 17072
rect 41739 17023 41781 17032
rect 41835 17072 41877 17081
rect 41835 17032 41836 17072
rect 41876 17032 41877 17072
rect 41835 17023 41877 17032
rect 41931 17072 41973 17081
rect 41931 17032 41932 17072
rect 41972 17032 41973 17072
rect 41931 17023 41973 17032
rect 42211 17072 42269 17073
rect 42211 17032 42220 17072
rect 42260 17032 42269 17072
rect 42211 17031 42269 17032
rect 42507 17072 42549 17081
rect 42507 17032 42508 17072
rect 42548 17032 42549 17072
rect 42507 17023 42549 17032
rect 43947 17072 43989 17081
rect 43947 17032 43948 17072
rect 43988 17032 43989 17072
rect 43947 17023 43989 17032
rect 44131 17072 44189 17073
rect 44131 17032 44140 17072
rect 44180 17032 44189 17072
rect 44131 17031 44189 17032
rect 45379 17072 45437 17073
rect 45379 17032 45388 17072
rect 45428 17032 45437 17072
rect 45379 17031 45437 17032
rect 45675 17072 45717 17081
rect 45675 17032 45676 17072
rect 45716 17032 45717 17072
rect 45675 17023 45717 17032
rect 46251 17072 46293 17081
rect 46251 17032 46252 17072
rect 46292 17032 46293 17072
rect 46251 17023 46293 17032
rect 46627 17072 46685 17073
rect 46627 17032 46636 17072
rect 46676 17032 46685 17072
rect 46627 17031 46685 17032
rect 47491 17072 47549 17073
rect 47491 17032 47500 17072
rect 47540 17032 47549 17072
rect 47491 17031 47549 17032
rect 49123 17072 49181 17073
rect 49123 17032 49132 17072
rect 49172 17032 49181 17072
rect 49123 17031 49181 17032
rect 49227 17072 49269 17081
rect 49227 17032 49228 17072
rect 49268 17032 49269 17072
rect 49227 17023 49269 17032
rect 49419 17072 49461 17081
rect 49419 17032 49420 17072
rect 49460 17032 49461 17072
rect 49419 17023 49461 17032
rect 49707 17072 49749 17081
rect 49707 17032 49708 17072
rect 49748 17032 49749 17072
rect 49707 17023 49749 17032
rect 49803 17072 49845 17081
rect 49803 17032 49804 17072
rect 49844 17032 49845 17072
rect 49803 17023 49845 17032
rect 49899 17072 49941 17081
rect 49899 17032 49900 17072
rect 49940 17032 49941 17072
rect 49899 17023 49941 17032
rect 49995 17072 50037 17081
rect 49995 17032 49996 17072
rect 50036 17032 50037 17072
rect 49995 17023 50037 17032
rect 50371 17072 50429 17073
rect 50371 17032 50380 17072
rect 50420 17032 50429 17072
rect 50371 17031 50429 17032
rect 50667 17072 50709 17081
rect 50667 17032 50668 17072
rect 50708 17032 50709 17072
rect 50667 17023 50709 17032
rect 50763 17072 50805 17081
rect 50763 17032 50764 17072
rect 50804 17032 50805 17072
rect 50763 17023 50805 17032
rect 51627 17072 51669 17081
rect 51627 17032 51628 17072
rect 51668 17032 51669 17072
rect 51627 17023 51669 17032
rect 51811 17072 51869 17073
rect 51811 17032 51820 17072
rect 51860 17032 51869 17072
rect 51811 17031 51869 17032
rect 52291 17072 52349 17073
rect 52291 17032 52300 17072
rect 52340 17032 52349 17072
rect 52291 17031 52349 17032
rect 52579 17072 52637 17073
rect 52579 17032 52588 17072
rect 52628 17032 52637 17072
rect 52579 17031 52637 17032
rect 2755 16988 2813 16989
rect 2755 16948 2764 16988
rect 2804 16948 2813 16988
rect 2755 16947 2813 16948
rect 3139 16988 3197 16989
rect 3139 16948 3148 16988
rect 3188 16948 3197 16988
rect 3139 16947 3197 16948
rect 4771 16988 4829 16989
rect 4771 16948 4780 16988
rect 4820 16948 4829 16988
rect 4771 16947 4829 16948
rect 23395 16988 23453 16989
rect 23395 16948 23404 16988
rect 23444 16948 23453 16988
rect 23395 16947 23453 16948
rect 40867 16988 40925 16989
rect 40867 16948 40876 16988
rect 40916 16948 40925 16988
rect 40867 16947 40925 16948
rect 41443 16988 41501 16989
rect 41443 16948 41452 16988
rect 41492 16948 41501 16988
rect 41443 16947 41501 16948
rect 43267 16988 43325 16989
rect 43267 16948 43276 16988
rect 43316 16948 43325 16988
rect 43267 16947 43325 16948
rect 44515 16988 44573 16989
rect 44515 16948 44524 16988
rect 44564 16948 44573 16988
rect 44515 16947 44573 16948
rect 44899 16988 44957 16989
rect 44899 16948 44908 16988
rect 44948 16948 44957 16988
rect 44899 16947 44957 16948
rect 48651 16988 48693 16997
rect 48651 16948 48652 16988
rect 48692 16948 48693 16988
rect 48651 16939 48693 16948
rect 51235 16988 51293 16989
rect 51235 16948 51244 16988
rect 51284 16948 51293 16988
rect 51235 16947 51293 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 2955 16904 2997 16913
rect 2955 16864 2956 16904
rect 2996 16864 2997 16904
rect 2955 16855 2997 16864
rect 3339 16904 3381 16913
rect 3339 16864 3340 16904
rect 3380 16864 3381 16904
rect 3339 16855 3381 16864
rect 4587 16904 4629 16913
rect 4587 16864 4588 16904
rect 4628 16864 4629 16904
rect 4587 16855 4629 16864
rect 23979 16904 24021 16913
rect 23979 16864 23980 16904
rect 24020 16864 24021 16904
rect 23979 16855 24021 16864
rect 27627 16904 27669 16913
rect 27627 16864 27628 16904
rect 27668 16864 27669 16904
rect 27627 16855 27669 16864
rect 30795 16904 30837 16913
rect 30795 16864 30796 16904
rect 30836 16864 30837 16904
rect 30795 16855 30837 16864
rect 31563 16904 31605 16913
rect 31563 16864 31564 16904
rect 31604 16864 31605 16904
rect 31563 16855 31605 16864
rect 33483 16904 33525 16913
rect 33483 16864 33484 16904
rect 33524 16864 33525 16904
rect 33483 16855 33525 16864
rect 34059 16904 34101 16913
rect 34059 16864 34060 16904
rect 34100 16864 34101 16904
rect 34059 16855 34101 16864
rect 39715 16904 39773 16905
rect 39715 16864 39724 16904
rect 39764 16864 39773 16904
rect 39715 16863 39773 16864
rect 41067 16904 41109 16913
rect 41067 16864 41068 16904
rect 41108 16864 41109 16904
rect 41067 16855 41109 16864
rect 42883 16904 42941 16905
rect 42883 16864 42892 16904
rect 42932 16864 42941 16904
rect 42883 16863 42941 16864
rect 43083 16904 43125 16913
rect 43083 16864 43084 16904
rect 43124 16864 43125 16904
rect 43083 16855 43125 16864
rect 43563 16904 43605 16913
rect 43563 16864 43564 16904
rect 43604 16864 43605 16904
rect 43563 16855 43605 16864
rect 44715 16904 44757 16913
rect 44715 16864 44716 16904
rect 44756 16864 44757 16904
rect 44715 16855 44757 16864
rect 51043 16904 51101 16905
rect 51043 16864 51052 16904
rect 51092 16864 51101 16904
rect 51043 16863 51101 16864
rect 4299 16820 4341 16829
rect 4299 16780 4300 16820
rect 4340 16780 4341 16820
rect 4299 16771 4341 16780
rect 36643 16820 36701 16821
rect 36643 16780 36652 16820
rect 36692 16780 36701 16820
rect 36643 16779 36701 16780
rect 37035 16820 37077 16829
rect 37035 16780 37036 16820
rect 37076 16780 37077 16820
rect 37035 16771 37077 16780
rect 41259 16820 41301 16829
rect 41259 16780 41260 16820
rect 41300 16780 41301 16820
rect 41259 16771 41301 16780
rect 45099 16820 45141 16829
rect 45099 16780 45100 16820
rect 45140 16780 45141 16820
rect 45099 16771 45141 16780
rect 46051 16820 46109 16821
rect 46051 16780 46060 16820
rect 46100 16780 46109 16820
rect 46051 16779 46109 16780
rect 49419 16820 49461 16829
rect 49419 16780 49420 16820
rect 49460 16780 49461 16820
rect 49419 16771 49461 16780
rect 51435 16820 51477 16829
rect 51435 16780 51436 16820
rect 51476 16780 51477 16820
rect 51435 16771 51477 16780
rect 52395 16820 52437 16829
rect 52395 16780 52396 16820
rect 52436 16780 52437 16820
rect 52395 16771 52437 16780
rect 576 16652 79584 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 79584 16652
rect 576 16588 79584 16612
rect 1995 16484 2037 16493
rect 1995 16444 1996 16484
rect 2036 16444 2037 16484
rect 1995 16435 2037 16444
rect 2571 16484 2613 16493
rect 2571 16444 2572 16484
rect 2612 16444 2613 16484
rect 2571 16435 2613 16444
rect 4011 16484 4053 16493
rect 4011 16444 4012 16484
rect 4052 16444 4053 16484
rect 4011 16435 4053 16444
rect 6979 16484 7037 16485
rect 6979 16444 6988 16484
rect 7028 16444 7037 16484
rect 6979 16443 7037 16444
rect 34731 16484 34773 16493
rect 34731 16444 34732 16484
rect 34772 16444 34773 16484
rect 34731 16435 34773 16444
rect 37995 16484 38037 16493
rect 37995 16444 37996 16484
rect 38036 16444 38037 16484
rect 37995 16435 38037 16444
rect 45763 16484 45821 16485
rect 45763 16444 45772 16484
rect 45812 16444 45821 16484
rect 45763 16443 45821 16444
rect 46251 16484 46293 16493
rect 46251 16444 46252 16484
rect 46292 16444 46293 16484
rect 46251 16435 46293 16444
rect 51043 16484 51101 16485
rect 51043 16444 51052 16484
rect 51092 16444 51101 16484
rect 51043 16443 51101 16444
rect 54795 16484 54837 16493
rect 54795 16444 54796 16484
rect 54836 16444 54837 16484
rect 54795 16435 54837 16444
rect 55083 16484 55125 16493
rect 55083 16444 55084 16484
rect 55124 16444 55125 16484
rect 55083 16435 55125 16444
rect 55371 16484 55413 16493
rect 55371 16444 55372 16484
rect 55412 16444 55413 16484
rect 55371 16435 55413 16444
rect 55755 16484 55797 16493
rect 55755 16444 55756 16484
rect 55796 16444 55797 16484
rect 55755 16435 55797 16444
rect 56619 16484 56661 16493
rect 56619 16444 56620 16484
rect 56660 16444 56661 16484
rect 56619 16435 56661 16444
rect 57387 16484 57429 16493
rect 57387 16444 57388 16484
rect 57428 16444 57429 16484
rect 57387 16435 57429 16444
rect 58059 16484 58101 16493
rect 58059 16444 58060 16484
rect 58100 16444 58101 16484
rect 58059 16435 58101 16444
rect 58347 16484 58389 16493
rect 58347 16444 58348 16484
rect 58388 16444 58389 16484
rect 58347 16435 58389 16444
rect 58635 16484 58677 16493
rect 58635 16444 58636 16484
rect 58676 16444 58677 16484
rect 58635 16435 58677 16444
rect 59019 16484 59061 16493
rect 59019 16444 59020 16484
rect 59060 16444 59061 16484
rect 59019 16435 59061 16444
rect 60171 16484 60213 16493
rect 60171 16444 60172 16484
rect 60212 16444 60213 16484
rect 60171 16435 60213 16444
rect 60555 16484 60597 16493
rect 60555 16444 60556 16484
rect 60596 16444 60597 16484
rect 60555 16435 60597 16444
rect 60843 16484 60885 16493
rect 60843 16444 60844 16484
rect 60884 16444 60885 16484
rect 60843 16435 60885 16444
rect 61515 16484 61557 16493
rect 61515 16444 61516 16484
rect 61556 16444 61557 16484
rect 61515 16435 61557 16444
rect 62187 16484 62229 16493
rect 62187 16444 62188 16484
rect 62228 16444 62229 16484
rect 62187 16435 62229 16444
rect 62475 16484 62517 16493
rect 62475 16444 62476 16484
rect 62516 16444 62517 16484
rect 62475 16435 62517 16444
rect 62763 16484 62805 16493
rect 62763 16444 62764 16484
rect 62804 16444 62805 16484
rect 62763 16435 62805 16444
rect 63051 16484 63093 16493
rect 63051 16444 63052 16484
rect 63092 16444 63093 16484
rect 63051 16435 63093 16444
rect 63435 16484 63477 16493
rect 63435 16444 63436 16484
rect 63476 16444 63477 16484
rect 63435 16435 63477 16444
rect 64587 16484 64629 16493
rect 64587 16444 64588 16484
rect 64628 16444 64629 16484
rect 64587 16435 64629 16444
rect 65067 16484 65109 16493
rect 65067 16444 65068 16484
rect 65108 16444 65109 16484
rect 65067 16435 65109 16444
rect 65451 16484 65493 16493
rect 65451 16444 65452 16484
rect 65492 16444 65493 16484
rect 65451 16435 65493 16444
rect 65835 16484 65877 16493
rect 65835 16444 65836 16484
rect 65876 16444 65877 16484
rect 65835 16435 65877 16444
rect 66603 16484 66645 16493
rect 66603 16444 66604 16484
rect 66644 16444 66645 16484
rect 66603 16435 66645 16444
rect 67083 16484 67125 16493
rect 67083 16444 67084 16484
rect 67124 16444 67125 16484
rect 67083 16435 67125 16444
rect 67467 16484 67509 16493
rect 67467 16444 67468 16484
rect 67508 16444 67509 16484
rect 67467 16435 67509 16444
rect 67851 16484 67893 16493
rect 67851 16444 67852 16484
rect 67892 16444 67893 16484
rect 67851 16435 67893 16444
rect 68235 16484 68277 16493
rect 68235 16444 68236 16484
rect 68276 16444 68277 16484
rect 68235 16435 68277 16444
rect 69003 16484 69045 16493
rect 69003 16444 69004 16484
rect 69044 16444 69045 16484
rect 69003 16435 69045 16444
rect 69483 16484 69525 16493
rect 69483 16444 69484 16484
rect 69524 16444 69525 16484
rect 69483 16435 69525 16444
rect 69867 16484 69909 16493
rect 69867 16444 69868 16484
rect 69908 16444 69909 16484
rect 69867 16435 69909 16444
rect 70251 16484 70293 16493
rect 70251 16444 70252 16484
rect 70292 16444 70293 16484
rect 70251 16435 70293 16444
rect 70635 16484 70677 16493
rect 70635 16444 70636 16484
rect 70676 16444 70677 16484
rect 70635 16435 70677 16444
rect 71019 16484 71061 16493
rect 71019 16444 71020 16484
rect 71060 16444 71061 16484
rect 71019 16435 71061 16444
rect 71403 16484 71445 16493
rect 71403 16444 71404 16484
rect 71444 16444 71445 16484
rect 71403 16435 71445 16444
rect 71883 16484 71925 16493
rect 71883 16444 71884 16484
rect 71924 16444 71925 16484
rect 71883 16435 71925 16444
rect 72267 16484 72309 16493
rect 72267 16444 72268 16484
rect 72308 16444 72309 16484
rect 72267 16435 72309 16444
rect 72651 16484 72693 16493
rect 72651 16444 72652 16484
rect 72692 16444 72693 16484
rect 72651 16435 72693 16444
rect 73035 16484 73077 16493
rect 73035 16444 73036 16484
rect 73076 16444 73077 16484
rect 73035 16435 73077 16444
rect 73419 16484 73461 16493
rect 73419 16444 73420 16484
rect 73460 16444 73461 16484
rect 73419 16435 73461 16444
rect 74283 16484 74325 16493
rect 74283 16444 74284 16484
rect 74324 16444 74325 16484
rect 74283 16435 74325 16444
rect 74667 16484 74709 16493
rect 74667 16444 74668 16484
rect 74708 16444 74709 16484
rect 74667 16435 74709 16444
rect 75051 16484 75093 16493
rect 75051 16444 75052 16484
rect 75092 16444 75093 16484
rect 75051 16435 75093 16444
rect 75435 16484 75477 16493
rect 75435 16444 75436 16484
rect 75476 16444 75477 16484
rect 75435 16435 75477 16444
rect 76491 16484 76533 16493
rect 76491 16444 76492 16484
rect 76532 16444 76533 16484
rect 76491 16435 76533 16444
rect 76875 16484 76917 16493
rect 76875 16444 76876 16484
rect 76916 16444 76917 16484
rect 76875 16435 76917 16444
rect 77259 16484 77301 16493
rect 77259 16444 77260 16484
rect 77300 16444 77301 16484
rect 77259 16435 77301 16444
rect 77643 16484 77685 16493
rect 77643 16444 77644 16484
rect 77684 16444 77685 16484
rect 77643 16435 77685 16444
rect 78027 16484 78069 16493
rect 78027 16444 78028 16484
rect 78068 16444 78069 16484
rect 78027 16435 78069 16444
rect 78315 16484 78357 16493
rect 78315 16444 78316 16484
rect 78356 16444 78357 16484
rect 78315 16435 78357 16444
rect 78699 16484 78741 16493
rect 78699 16444 78700 16484
rect 78740 16444 78741 16484
rect 78699 16435 78741 16444
rect 78987 16484 79029 16493
rect 78987 16444 78988 16484
rect 79028 16444 79029 16484
rect 78987 16435 79029 16444
rect 79275 16484 79317 16493
rect 79275 16444 79276 16484
rect 79316 16444 79317 16484
rect 79275 16435 79317 16444
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 1803 16400 1845 16409
rect 1803 16360 1804 16400
rect 1844 16360 1845 16400
rect 1803 16351 1845 16360
rect 4203 16400 4245 16409
rect 4203 16360 4204 16400
rect 4244 16360 4245 16400
rect 4203 16351 4245 16360
rect 34435 16400 34493 16401
rect 34435 16360 34444 16400
rect 34484 16360 34493 16400
rect 34435 16359 34493 16360
rect 37507 16400 37565 16401
rect 37507 16360 37516 16400
rect 37556 16360 37565 16400
rect 37507 16359 37565 16360
rect 43083 16400 43125 16409
rect 43083 16360 43084 16400
rect 43124 16360 43125 16400
rect 43083 16351 43125 16360
rect 46731 16400 46773 16409
rect 46731 16360 46732 16400
rect 46772 16360 46773 16400
rect 46731 16351 46773 16360
rect 52099 16400 52157 16401
rect 52099 16360 52108 16400
rect 52148 16360 52157 16400
rect 52099 16359 52157 16360
rect 53643 16400 53685 16409
rect 53643 16360 53644 16400
rect 53684 16360 53685 16400
rect 53643 16351 53685 16360
rect 53931 16400 53973 16409
rect 53931 16360 53932 16400
rect 53972 16360 53973 16400
rect 53931 16351 53973 16360
rect 54315 16400 54357 16409
rect 54315 16360 54316 16400
rect 54356 16360 54357 16400
rect 54315 16351 54357 16360
rect 57579 16400 57621 16409
rect 57579 16360 57580 16400
rect 57620 16360 57621 16400
rect 57579 16351 57621 16360
rect 61035 16400 61077 16409
rect 61035 16360 61036 16400
rect 61076 16360 61077 16400
rect 61035 16351 61077 16360
rect 2179 16316 2237 16317
rect 2179 16276 2188 16316
rect 2228 16276 2237 16316
rect 2179 16275 2237 16276
rect 2371 16316 2429 16317
rect 2371 16276 2380 16316
rect 2420 16276 2429 16316
rect 2371 16275 2429 16276
rect 3427 16316 3485 16317
rect 3427 16276 3436 16316
rect 3476 16276 3485 16316
rect 3427 16275 3485 16276
rect 3811 16316 3869 16317
rect 3811 16276 3820 16316
rect 3860 16276 3869 16316
rect 3811 16275 3869 16276
rect 4387 16316 4445 16317
rect 4387 16276 4396 16316
rect 4436 16276 4445 16316
rect 4387 16275 4445 16276
rect 61699 16316 61757 16317
rect 61699 16276 61708 16316
rect 61748 16276 61757 16316
rect 61699 16275 61757 16276
rect 36835 16249 36893 16250
rect 2763 16232 2805 16241
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 2955 16232 2997 16241
rect 2955 16192 2956 16232
rect 2996 16192 2997 16232
rect 2955 16183 2997 16192
rect 3043 16232 3101 16233
rect 3043 16192 3052 16232
rect 3092 16192 3101 16232
rect 3043 16191 3101 16192
rect 4963 16232 5021 16233
rect 4963 16192 4972 16232
rect 5012 16192 5021 16232
rect 4963 16191 5021 16192
rect 5827 16232 5885 16233
rect 5827 16192 5836 16232
rect 5876 16192 5885 16232
rect 5827 16191 5885 16192
rect 31459 16232 31517 16233
rect 31459 16192 31468 16232
rect 31508 16192 31517 16232
rect 31459 16191 31517 16192
rect 32323 16232 32381 16233
rect 32323 16192 32332 16232
rect 32372 16192 32381 16232
rect 32323 16191 32381 16192
rect 33763 16232 33821 16233
rect 33763 16192 33772 16232
rect 33812 16192 33821 16232
rect 33763 16191 33821 16192
rect 34059 16232 34101 16241
rect 34059 16192 34060 16232
rect 34100 16192 34101 16232
rect 34059 16183 34101 16192
rect 34635 16232 34677 16241
rect 34635 16192 34636 16232
rect 34676 16192 34677 16232
rect 34635 16183 34677 16192
rect 34819 16232 34877 16233
rect 34819 16192 34828 16232
rect 34868 16192 34877 16232
rect 36835 16209 36844 16249
rect 36884 16209 36893 16249
rect 43172 16247 43214 16256
rect 36835 16208 36893 16209
rect 37131 16232 37173 16241
rect 34819 16191 34877 16192
rect 37131 16192 37132 16232
rect 37172 16192 37173 16232
rect 37131 16183 37173 16192
rect 37699 16232 37757 16233
rect 37699 16192 37708 16232
rect 37748 16192 37757 16232
rect 37699 16191 37757 16192
rect 37803 16232 37845 16241
rect 37803 16192 37804 16232
rect 37844 16192 37845 16232
rect 37803 16183 37845 16192
rect 37995 16232 38037 16241
rect 37995 16192 37996 16232
rect 38036 16192 38037 16232
rect 37995 16183 38037 16192
rect 39819 16232 39861 16241
rect 39819 16192 39820 16232
rect 39860 16192 39861 16232
rect 39819 16183 39861 16192
rect 40003 16232 40061 16233
rect 40003 16192 40012 16232
rect 40052 16192 40061 16232
rect 40003 16191 40061 16192
rect 40579 16232 40637 16233
rect 40579 16192 40588 16232
rect 40628 16192 40637 16232
rect 40579 16191 40637 16192
rect 41443 16232 41501 16233
rect 41443 16192 41452 16232
rect 41492 16192 41501 16232
rect 41443 16191 41501 16192
rect 42979 16232 43037 16233
rect 42979 16192 42988 16232
rect 43028 16192 43037 16232
rect 43172 16207 43173 16247
rect 43213 16207 43214 16247
rect 43172 16198 43214 16207
rect 43747 16232 43805 16233
rect 42979 16191 43037 16192
rect 43747 16192 43756 16232
rect 43796 16192 43805 16232
rect 43747 16191 43805 16192
rect 44611 16232 44669 16233
rect 44611 16192 44620 16232
rect 44660 16192 44669 16232
rect 44611 16191 44669 16192
rect 45955 16232 46013 16233
rect 45955 16192 45964 16232
rect 46004 16192 46013 16232
rect 45955 16191 46013 16192
rect 46059 16232 46101 16241
rect 46059 16192 46060 16232
rect 46100 16192 46101 16232
rect 46059 16183 46101 16192
rect 46251 16232 46293 16241
rect 46251 16192 46252 16232
rect 46292 16192 46293 16232
rect 46251 16183 46293 16192
rect 47115 16232 47157 16241
rect 47115 16192 47116 16232
rect 47156 16192 47157 16232
rect 47115 16183 47157 16192
rect 47211 16232 47253 16241
rect 47211 16192 47212 16232
rect 47252 16192 47253 16232
rect 47211 16183 47253 16192
rect 47299 16232 47357 16233
rect 47299 16192 47308 16232
rect 47348 16192 47357 16232
rect 47299 16191 47357 16192
rect 48651 16232 48693 16241
rect 48651 16192 48652 16232
rect 48692 16192 48693 16232
rect 48651 16183 48693 16192
rect 49027 16232 49085 16233
rect 49027 16192 49036 16232
rect 49076 16192 49085 16232
rect 49027 16191 49085 16192
rect 49891 16232 49949 16233
rect 49891 16192 49900 16232
rect 49940 16192 49949 16232
rect 49891 16191 49949 16192
rect 51627 16232 51669 16241
rect 51627 16192 51628 16232
rect 51668 16192 51669 16232
rect 51627 16183 51669 16192
rect 51723 16232 51765 16241
rect 51723 16192 51724 16232
rect 51764 16192 51765 16232
rect 51723 16183 51765 16192
rect 51819 16232 51861 16241
rect 51819 16192 51820 16232
rect 51860 16192 51861 16232
rect 51819 16183 51861 16192
rect 52395 16232 52437 16241
rect 52395 16192 52396 16232
rect 52436 16192 52437 16232
rect 52395 16183 52437 16192
rect 52491 16232 52533 16241
rect 52491 16192 52492 16232
rect 52532 16192 52533 16232
rect 52491 16183 52533 16192
rect 52771 16232 52829 16233
rect 52771 16192 52780 16232
rect 52820 16192 52829 16232
rect 53347 16232 53405 16233
rect 52771 16191 52829 16192
rect 53067 16218 53109 16227
rect 53067 16178 53068 16218
rect 53108 16178 53109 16218
rect 53067 16169 53109 16178
rect 53259 16190 53301 16199
rect 53347 16192 53356 16232
rect 53396 16192 53405 16232
rect 53347 16191 53405 16192
rect 53539 16232 53597 16233
rect 53539 16192 53548 16232
rect 53588 16192 53597 16232
rect 53539 16191 53597 16192
rect 53739 16232 53781 16241
rect 53739 16192 53740 16232
rect 53780 16192 53781 16232
rect 4587 16148 4629 16157
rect 4587 16108 4588 16148
rect 4628 16108 4629 16148
rect 4587 16099 4629 16108
rect 31083 16148 31125 16157
rect 31083 16108 31084 16148
rect 31124 16108 31125 16148
rect 31083 16099 31125 16108
rect 34155 16148 34197 16157
rect 34155 16108 34156 16148
rect 34196 16108 34197 16148
rect 34155 16099 34197 16108
rect 37227 16148 37269 16157
rect 37227 16108 37228 16148
rect 37268 16108 37269 16148
rect 37227 16099 37269 16108
rect 39915 16148 39957 16157
rect 39915 16108 39916 16148
rect 39956 16108 39957 16148
rect 39915 16099 39957 16108
rect 40203 16148 40245 16157
rect 40203 16108 40204 16148
rect 40244 16108 40245 16148
rect 40203 16099 40245 16108
rect 43371 16148 43413 16157
rect 43371 16108 43372 16148
rect 43412 16108 43413 16148
rect 53259 16150 53260 16190
rect 53300 16150 53301 16190
rect 53739 16183 53781 16192
rect 54691 16232 54749 16233
rect 54691 16192 54700 16232
rect 54740 16192 54749 16232
rect 54691 16191 54749 16192
rect 54979 16232 55037 16233
rect 54979 16192 54988 16232
rect 55028 16192 55037 16232
rect 54979 16191 55037 16192
rect 55267 16232 55325 16233
rect 55267 16192 55276 16232
rect 55316 16192 55325 16232
rect 55267 16191 55325 16192
rect 55651 16232 55709 16233
rect 55651 16192 55660 16232
rect 55700 16192 55709 16232
rect 55651 16191 55709 16192
rect 56035 16232 56093 16233
rect 56035 16192 56044 16232
rect 56084 16192 56093 16232
rect 56035 16191 56093 16192
rect 56515 16232 56573 16233
rect 56515 16192 56524 16232
rect 56564 16192 56573 16232
rect 56515 16191 56573 16192
rect 56899 16232 56957 16233
rect 56899 16192 56908 16232
rect 56948 16192 56957 16232
rect 56899 16191 56957 16192
rect 57283 16232 57341 16233
rect 57283 16192 57292 16232
rect 57332 16192 57341 16232
rect 57283 16191 57341 16192
rect 57955 16232 58013 16233
rect 57955 16192 57964 16232
rect 58004 16192 58013 16232
rect 57955 16191 58013 16192
rect 58243 16232 58301 16233
rect 58243 16192 58252 16232
rect 58292 16192 58301 16232
rect 58243 16191 58301 16192
rect 58531 16232 58589 16233
rect 58531 16192 58540 16232
rect 58580 16192 58589 16232
rect 58531 16191 58589 16192
rect 58915 16232 58973 16233
rect 58915 16192 58924 16232
rect 58964 16192 58973 16232
rect 58915 16191 58973 16192
rect 59299 16232 59357 16233
rect 59299 16192 59308 16232
rect 59348 16192 59357 16232
rect 59299 16191 59357 16192
rect 59683 16232 59741 16233
rect 59683 16192 59692 16232
rect 59732 16192 59741 16232
rect 59683 16191 59741 16192
rect 60067 16232 60125 16233
rect 60067 16192 60076 16232
rect 60116 16192 60125 16232
rect 60067 16191 60125 16192
rect 60451 16232 60509 16233
rect 60451 16192 60460 16232
rect 60500 16192 60509 16232
rect 60451 16191 60509 16192
rect 60739 16232 60797 16233
rect 60739 16192 60748 16232
rect 60788 16192 60797 16232
rect 60739 16191 60797 16192
rect 61411 16232 61469 16233
rect 61411 16192 61420 16232
rect 61460 16192 61469 16232
rect 61411 16191 61469 16192
rect 62083 16232 62141 16233
rect 62083 16192 62092 16232
rect 62132 16192 62141 16232
rect 62083 16191 62141 16192
rect 62371 16232 62429 16233
rect 62371 16192 62380 16232
rect 62420 16192 62429 16232
rect 62371 16191 62429 16192
rect 62659 16232 62717 16233
rect 62659 16192 62668 16232
rect 62708 16192 62717 16232
rect 62659 16191 62717 16192
rect 62947 16232 63005 16233
rect 62947 16192 62956 16232
rect 62996 16192 63005 16232
rect 63715 16232 63773 16233
rect 62947 16191 63005 16192
rect 63326 16221 63368 16230
rect 63326 16181 63327 16221
rect 63367 16181 63368 16221
rect 63715 16192 63724 16232
rect 63764 16192 63773 16232
rect 63715 16191 63773 16192
rect 64099 16232 64157 16233
rect 64099 16192 64108 16232
rect 64148 16192 64157 16232
rect 64099 16191 64157 16192
rect 64483 16232 64541 16233
rect 64483 16192 64492 16232
rect 64532 16192 64541 16232
rect 64483 16191 64541 16192
rect 64963 16232 65021 16233
rect 64963 16192 64972 16232
rect 65012 16192 65021 16232
rect 64963 16191 65021 16192
rect 65347 16232 65405 16233
rect 65347 16192 65356 16232
rect 65396 16192 65405 16232
rect 65347 16191 65405 16192
rect 65731 16232 65789 16233
rect 65731 16192 65740 16232
rect 65780 16192 65789 16232
rect 65731 16191 65789 16192
rect 66115 16232 66173 16233
rect 66115 16192 66124 16232
rect 66164 16192 66173 16232
rect 66115 16191 66173 16192
rect 66499 16232 66557 16233
rect 66499 16192 66508 16232
rect 66548 16192 66557 16232
rect 66499 16191 66557 16192
rect 66979 16232 67037 16233
rect 66979 16192 66988 16232
rect 67028 16192 67037 16232
rect 66979 16191 67037 16192
rect 67363 16232 67421 16233
rect 67363 16192 67372 16232
rect 67412 16192 67421 16232
rect 67363 16191 67421 16192
rect 67747 16232 67805 16233
rect 67747 16192 67756 16232
rect 67796 16192 67805 16232
rect 67747 16191 67805 16192
rect 68131 16232 68189 16233
rect 68131 16192 68140 16232
rect 68180 16192 68189 16232
rect 68131 16191 68189 16192
rect 68515 16232 68573 16233
rect 68515 16192 68524 16232
rect 68564 16192 68573 16232
rect 68515 16191 68573 16192
rect 68899 16232 68957 16233
rect 68899 16192 68908 16232
rect 68948 16192 68957 16232
rect 68899 16191 68957 16192
rect 69379 16232 69437 16233
rect 69379 16192 69388 16232
rect 69428 16192 69437 16232
rect 69379 16191 69437 16192
rect 69763 16232 69821 16233
rect 69763 16192 69772 16232
rect 69812 16192 69821 16232
rect 69763 16191 69821 16192
rect 70147 16232 70205 16233
rect 70147 16192 70156 16232
rect 70196 16192 70205 16232
rect 70147 16191 70205 16192
rect 70531 16232 70589 16233
rect 70531 16192 70540 16232
rect 70580 16192 70589 16232
rect 70531 16191 70589 16192
rect 70915 16232 70973 16233
rect 70915 16192 70924 16232
rect 70964 16192 70973 16232
rect 70915 16191 70973 16192
rect 71299 16232 71357 16233
rect 71299 16192 71308 16232
rect 71348 16192 71357 16232
rect 71299 16191 71357 16192
rect 71779 16232 71837 16233
rect 71779 16192 71788 16232
rect 71828 16192 71837 16232
rect 71779 16191 71837 16192
rect 72163 16232 72221 16233
rect 72163 16192 72172 16232
rect 72212 16192 72221 16232
rect 72163 16191 72221 16192
rect 72547 16232 72605 16233
rect 72547 16192 72556 16232
rect 72596 16192 72605 16232
rect 72547 16191 72605 16192
rect 72931 16232 72989 16233
rect 72931 16192 72940 16232
rect 72980 16192 72989 16232
rect 72931 16191 72989 16192
rect 73315 16232 73373 16233
rect 73315 16192 73324 16232
rect 73364 16192 73373 16232
rect 73315 16191 73373 16192
rect 73699 16232 73757 16233
rect 73699 16192 73708 16232
rect 73748 16192 73757 16232
rect 73699 16191 73757 16192
rect 74179 16232 74237 16233
rect 74179 16192 74188 16232
rect 74228 16192 74237 16232
rect 74179 16191 74237 16192
rect 74563 16232 74621 16233
rect 74563 16192 74572 16232
rect 74612 16192 74621 16232
rect 74563 16191 74621 16192
rect 74947 16232 75005 16233
rect 74947 16192 74956 16232
rect 74996 16192 75005 16232
rect 74947 16191 75005 16192
rect 75331 16232 75389 16233
rect 75331 16192 75340 16232
rect 75380 16192 75389 16232
rect 75331 16191 75389 16192
rect 75715 16232 75773 16233
rect 75715 16192 75724 16232
rect 75764 16192 75773 16232
rect 75715 16191 75773 16192
rect 76579 16232 76637 16233
rect 76579 16192 76588 16232
rect 76628 16192 76637 16232
rect 76579 16191 76637 16192
rect 76963 16232 77021 16233
rect 76963 16192 76972 16232
rect 77012 16192 77021 16232
rect 76963 16191 77021 16192
rect 77155 16232 77213 16233
rect 77155 16192 77164 16232
rect 77204 16192 77213 16232
rect 77155 16191 77213 16192
rect 77539 16232 77597 16233
rect 77539 16192 77548 16232
rect 77588 16192 77597 16232
rect 77539 16191 77597 16192
rect 77923 16232 77981 16233
rect 77923 16192 77932 16232
rect 77972 16192 77981 16232
rect 77923 16191 77981 16192
rect 78211 16232 78269 16233
rect 78211 16192 78220 16232
rect 78260 16192 78269 16232
rect 78211 16191 78269 16192
rect 78595 16232 78653 16233
rect 78595 16192 78604 16232
rect 78644 16192 78653 16232
rect 78595 16191 78653 16192
rect 78883 16232 78941 16233
rect 78883 16192 78892 16232
rect 78932 16192 78941 16232
rect 78883 16191 78941 16192
rect 79171 16232 79229 16233
rect 79171 16192 79180 16232
rect 79220 16192 79229 16232
rect 79171 16191 79229 16192
rect 63326 16172 63368 16181
rect 53259 16141 53301 16150
rect 63819 16148 63861 16157
rect 43371 16099 43413 16108
rect 63819 16108 63820 16148
rect 63860 16108 63861 16148
rect 63819 16099 63861 16108
rect 1995 16064 2037 16073
rect 1995 16024 1996 16064
rect 2036 16024 2037 16064
rect 1995 16015 2037 16024
rect 2851 16064 2909 16065
rect 2851 16024 2860 16064
rect 2900 16024 2909 16064
rect 2851 16023 2909 16024
rect 3627 16064 3669 16073
rect 3627 16024 3628 16064
rect 3668 16024 3669 16064
rect 3627 16015 3669 16024
rect 33475 16064 33533 16065
rect 33475 16024 33484 16064
rect 33524 16024 33533 16064
rect 33475 16023 33533 16024
rect 42595 16064 42653 16065
rect 42595 16024 42604 16064
rect 42644 16024 42653 16064
rect 42595 16023 42653 16024
rect 45763 16064 45821 16065
rect 45763 16024 45772 16064
rect 45812 16024 45821 16064
rect 45763 16023 45821 16024
rect 51523 16064 51581 16065
rect 51523 16024 51532 16064
rect 51572 16024 51581 16064
rect 51523 16023 51581 16024
rect 53155 16064 53213 16065
rect 53155 16024 53164 16064
rect 53204 16024 53213 16064
rect 53155 16023 53213 16024
rect 56139 16064 56181 16073
rect 56139 16024 56140 16064
rect 56180 16024 56181 16064
rect 56139 16015 56181 16024
rect 57003 16064 57045 16073
rect 57003 16024 57004 16064
rect 57044 16024 57045 16064
rect 57003 16015 57045 16024
rect 59403 16064 59445 16073
rect 59403 16024 59404 16064
rect 59444 16024 59445 16064
rect 59403 16015 59445 16024
rect 59787 16064 59829 16073
rect 59787 16024 59788 16064
rect 59828 16024 59829 16064
rect 59787 16015 59829 16024
rect 61899 16064 61941 16073
rect 61899 16024 61900 16064
rect 61940 16024 61941 16064
rect 61899 16015 61941 16024
rect 64203 16064 64245 16073
rect 64203 16024 64204 16064
rect 64244 16024 64245 16064
rect 64203 16015 64245 16024
rect 66219 16064 66261 16073
rect 66219 16024 66220 16064
rect 66260 16024 66261 16064
rect 66219 16015 66261 16024
rect 68619 16064 68661 16073
rect 68619 16024 68620 16064
rect 68660 16024 68661 16064
rect 68619 16015 68661 16024
rect 73803 16064 73845 16073
rect 73803 16024 73804 16064
rect 73844 16024 73845 16064
rect 73803 16015 73845 16024
rect 75819 16064 75861 16073
rect 75819 16024 75820 16064
rect 75860 16024 75861 16064
rect 75819 16015 75861 16024
rect 576 15896 79584 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 79584 15896
rect 576 15832 79584 15856
rect 4483 15728 4541 15729
rect 4483 15688 4492 15728
rect 4532 15688 4541 15728
rect 4483 15687 4541 15688
rect 33955 15728 34013 15729
rect 33955 15688 33964 15728
rect 34004 15688 34013 15728
rect 33955 15687 34013 15688
rect 40483 15728 40541 15729
rect 40483 15688 40492 15728
rect 40532 15688 40541 15728
rect 40483 15687 40541 15688
rect 46051 15728 46109 15729
rect 46051 15688 46060 15728
rect 46100 15688 46109 15728
rect 46051 15687 46109 15688
rect 50187 15728 50229 15737
rect 50187 15688 50188 15728
rect 50228 15688 50229 15728
rect 50187 15679 50229 15688
rect 55459 15728 55517 15729
rect 55459 15688 55468 15728
rect 55508 15688 55517 15728
rect 55459 15687 55517 15688
rect 59491 15728 59549 15729
rect 59491 15688 59500 15728
rect 59540 15688 59549 15728
rect 59491 15687 59549 15688
rect 62947 15728 63005 15729
rect 62947 15688 62956 15728
rect 62996 15688 63005 15728
rect 62947 15687 63005 15688
rect 67843 15728 67901 15729
rect 67843 15688 67852 15728
rect 67892 15688 67901 15728
rect 67843 15687 67901 15688
rect 79467 15728 79509 15737
rect 79467 15688 79468 15728
rect 79508 15688 79509 15728
rect 79467 15679 79509 15688
rect 3531 15644 3573 15653
rect 3531 15604 3532 15644
rect 3572 15604 3573 15644
rect 3531 15595 3573 15604
rect 3819 15644 3861 15653
rect 3819 15604 3820 15644
rect 3860 15604 3861 15644
rect 3819 15595 3861 15604
rect 32139 15644 32181 15653
rect 32139 15604 32140 15644
rect 32180 15604 32181 15644
rect 32139 15595 32181 15604
rect 38379 15644 38421 15653
rect 38379 15604 38380 15644
rect 38420 15604 38421 15644
rect 38379 15595 38421 15604
rect 53067 15644 53109 15653
rect 53067 15604 53068 15644
rect 53108 15604 53109 15644
rect 53067 15595 53109 15604
rect 2275 15560 2333 15561
rect 2275 15520 2284 15560
rect 2324 15520 2333 15560
rect 2275 15519 2333 15520
rect 3139 15560 3197 15561
rect 3139 15520 3148 15560
rect 3188 15520 3197 15560
rect 3139 15519 3197 15520
rect 3723 15560 3765 15569
rect 3723 15520 3724 15560
rect 3764 15520 3765 15560
rect 3723 15511 3765 15520
rect 3907 15560 3965 15561
rect 3907 15520 3916 15560
rect 3956 15520 3965 15560
rect 3907 15519 3965 15520
rect 4291 15560 4349 15561
rect 4291 15520 4300 15560
rect 4340 15520 4349 15560
rect 4291 15519 4349 15520
rect 4395 15560 4437 15569
rect 4395 15520 4396 15560
rect 4436 15520 4437 15560
rect 4395 15511 4437 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 31563 15560 31605 15569
rect 31563 15520 31564 15560
rect 31604 15520 31605 15560
rect 31563 15511 31605 15520
rect 31755 15560 31797 15569
rect 31755 15520 31756 15560
rect 31796 15520 31797 15560
rect 31755 15511 31797 15520
rect 31843 15560 31901 15561
rect 31843 15520 31852 15560
rect 31892 15520 31901 15560
rect 31843 15519 31901 15520
rect 32035 15560 32093 15561
rect 32035 15520 32044 15560
rect 32084 15520 32093 15560
rect 32035 15519 32093 15520
rect 32235 15560 32277 15569
rect 32235 15520 32236 15560
rect 32276 15520 32277 15560
rect 32235 15511 32277 15520
rect 33387 15560 33429 15569
rect 33387 15520 33388 15560
rect 33428 15520 33429 15560
rect 33387 15511 33429 15520
rect 33483 15560 33525 15569
rect 33483 15520 33484 15560
rect 33524 15520 33525 15560
rect 33483 15511 33525 15520
rect 33579 15560 33621 15569
rect 33579 15520 33580 15560
rect 33620 15520 33621 15560
rect 33579 15511 33621 15520
rect 33675 15560 33717 15569
rect 33675 15520 33676 15560
rect 33716 15520 33717 15560
rect 33675 15511 33717 15520
rect 33867 15560 33909 15569
rect 33867 15520 33868 15560
rect 33908 15520 33909 15560
rect 33867 15511 33909 15520
rect 34059 15560 34101 15569
rect 34059 15520 34060 15560
rect 34100 15520 34101 15560
rect 34059 15511 34101 15520
rect 34147 15560 34205 15561
rect 34147 15520 34156 15560
rect 34196 15520 34205 15560
rect 34147 15519 34205 15520
rect 34923 15560 34965 15569
rect 34923 15520 34924 15560
rect 34964 15520 34965 15560
rect 34923 15511 34965 15520
rect 35115 15560 35157 15569
rect 35115 15520 35116 15560
rect 35156 15520 35157 15560
rect 35115 15511 35157 15520
rect 35203 15560 35261 15561
rect 35203 15520 35212 15560
rect 35252 15520 35261 15560
rect 35203 15519 35261 15520
rect 36267 15560 36309 15569
rect 36267 15520 36268 15560
rect 36308 15520 36309 15560
rect 36267 15511 36309 15520
rect 36363 15560 36405 15569
rect 36363 15520 36364 15560
rect 36404 15520 36405 15560
rect 36363 15511 36405 15520
rect 36459 15560 36501 15569
rect 36459 15520 36460 15560
rect 36500 15520 36501 15560
rect 36459 15511 36501 15520
rect 36555 15560 36597 15569
rect 36555 15520 36556 15560
rect 36596 15520 36597 15560
rect 36555 15511 36597 15520
rect 36747 15560 36789 15569
rect 36747 15520 36748 15560
rect 36788 15520 36789 15560
rect 36747 15511 36789 15520
rect 36939 15560 36981 15569
rect 36939 15520 36940 15560
rect 36980 15520 36981 15560
rect 36939 15511 36981 15520
rect 37027 15560 37085 15561
rect 37027 15520 37036 15560
rect 37076 15520 37085 15560
rect 37027 15519 37085 15520
rect 37515 15560 37557 15569
rect 37515 15520 37516 15560
rect 37556 15520 37557 15560
rect 37515 15511 37557 15520
rect 38275 15560 38333 15561
rect 38275 15520 38284 15560
rect 38324 15520 38333 15560
rect 38275 15519 38333 15520
rect 38475 15560 38517 15569
rect 38475 15520 38476 15560
rect 38516 15520 38517 15560
rect 38475 15511 38517 15520
rect 39051 15560 39093 15569
rect 39051 15520 39052 15560
rect 39092 15520 39093 15560
rect 39051 15511 39093 15520
rect 39147 15560 39189 15569
rect 39147 15520 39148 15560
rect 39188 15520 39189 15560
rect 39147 15511 39189 15520
rect 39235 15560 39293 15561
rect 39235 15520 39244 15560
rect 39284 15520 39293 15560
rect 39235 15519 39293 15520
rect 39723 15560 39765 15569
rect 39723 15520 39724 15560
rect 39764 15520 39765 15560
rect 39723 15511 39765 15520
rect 39819 15560 39861 15569
rect 39819 15520 39820 15560
rect 39860 15520 39861 15560
rect 39819 15511 39861 15520
rect 40099 15560 40157 15561
rect 40099 15520 40108 15560
rect 40148 15520 40157 15560
rect 40099 15519 40157 15520
rect 40395 15560 40437 15569
rect 40395 15520 40396 15560
rect 40436 15520 40437 15560
rect 40395 15511 40437 15520
rect 40587 15560 40629 15569
rect 40587 15520 40588 15560
rect 40628 15520 40629 15560
rect 40587 15511 40629 15520
rect 40675 15560 40733 15561
rect 40675 15520 40684 15560
rect 40724 15520 40733 15560
rect 40675 15519 40733 15520
rect 41835 15560 41877 15569
rect 41835 15520 41836 15560
rect 41876 15520 41877 15560
rect 41835 15511 41877 15520
rect 42027 15560 42069 15569
rect 42027 15520 42028 15560
rect 42068 15520 42069 15560
rect 42027 15511 42069 15520
rect 42115 15560 42173 15561
rect 42115 15520 42124 15560
rect 42164 15520 42173 15560
rect 42115 15519 42173 15520
rect 45483 15560 45525 15569
rect 45483 15520 45484 15560
rect 45524 15520 45525 15560
rect 45483 15511 45525 15520
rect 45579 15560 45621 15569
rect 45579 15520 45580 15560
rect 45620 15520 45621 15560
rect 45579 15511 45621 15520
rect 45675 15560 45717 15569
rect 45675 15520 45676 15560
rect 45716 15520 45717 15560
rect 45675 15511 45717 15520
rect 45771 15560 45813 15569
rect 45771 15520 45772 15560
rect 45812 15520 45813 15560
rect 45771 15511 45813 15520
rect 45963 15560 46005 15569
rect 45963 15520 45964 15560
rect 46004 15520 46005 15560
rect 45963 15511 46005 15520
rect 46155 15560 46197 15569
rect 46155 15520 46156 15560
rect 46196 15520 46197 15560
rect 46155 15511 46197 15520
rect 46243 15560 46301 15561
rect 46243 15520 46252 15560
rect 46292 15520 46301 15560
rect 46243 15519 46301 15520
rect 47491 15560 47549 15561
rect 47491 15520 47500 15560
rect 47540 15520 47549 15560
rect 47491 15519 47549 15520
rect 47691 15560 47733 15569
rect 47691 15520 47692 15560
rect 47732 15520 47733 15560
rect 47691 15511 47733 15520
rect 47875 15560 47933 15561
rect 47875 15520 47884 15560
rect 47924 15520 47933 15560
rect 47875 15519 47933 15520
rect 48075 15560 48117 15569
rect 48075 15520 48076 15560
rect 48116 15520 48117 15560
rect 48075 15511 48117 15520
rect 50755 15560 50813 15561
rect 50755 15520 50764 15560
rect 50804 15520 50813 15560
rect 50755 15519 50813 15520
rect 50859 15560 50901 15569
rect 50859 15520 50860 15560
rect 50900 15520 50901 15560
rect 50859 15511 50901 15520
rect 51051 15560 51093 15569
rect 51051 15520 51052 15560
rect 51092 15520 51093 15560
rect 51051 15511 51093 15520
rect 51235 15560 51293 15561
rect 51235 15520 51244 15560
rect 51284 15520 51293 15560
rect 51235 15519 51293 15520
rect 51715 15560 51773 15561
rect 51715 15520 51724 15560
rect 51764 15520 51773 15560
rect 51715 15519 51773 15520
rect 52675 15560 52733 15561
rect 52675 15520 52684 15560
rect 52724 15520 52733 15560
rect 52675 15519 52733 15520
rect 53443 15560 53501 15561
rect 53443 15520 53452 15560
rect 53492 15520 53501 15560
rect 53443 15519 53501 15520
rect 54307 15560 54365 15561
rect 54307 15520 54316 15560
rect 54356 15520 54365 15560
rect 54307 15519 54365 15520
rect 57099 15560 57141 15569
rect 57099 15520 57100 15560
rect 57140 15520 57141 15560
rect 57099 15511 57141 15520
rect 57475 15560 57533 15561
rect 57475 15520 57484 15560
rect 57524 15520 57533 15560
rect 57475 15519 57533 15520
rect 58339 15560 58397 15561
rect 58339 15520 58348 15560
rect 58388 15520 58397 15560
rect 58339 15519 58397 15520
rect 60555 15560 60597 15569
rect 60555 15520 60556 15560
rect 60596 15520 60597 15560
rect 60555 15511 60597 15520
rect 60931 15560 60989 15561
rect 60931 15520 60940 15560
rect 60980 15520 60989 15560
rect 60931 15519 60989 15520
rect 61795 15560 61853 15561
rect 61795 15520 61804 15560
rect 61844 15520 61853 15560
rect 61795 15519 61853 15520
rect 64875 15560 64917 15569
rect 64875 15520 64876 15560
rect 64916 15520 64917 15560
rect 64875 15511 64917 15520
rect 65059 15560 65117 15561
rect 65059 15520 65068 15560
rect 65108 15520 65117 15560
rect 65059 15519 65117 15520
rect 65451 15560 65493 15569
rect 65451 15520 65452 15560
rect 65492 15520 65493 15560
rect 65451 15511 65493 15520
rect 65827 15560 65885 15561
rect 65827 15520 65836 15560
rect 65876 15520 65885 15560
rect 65827 15519 65885 15520
rect 66691 15560 66749 15561
rect 66691 15520 66700 15560
rect 66740 15520 66749 15560
rect 66691 15519 66749 15520
rect 70051 15560 70109 15561
rect 70051 15520 70060 15560
rect 70100 15520 70109 15560
rect 70051 15519 70109 15520
rect 70155 15560 70197 15569
rect 70155 15520 70156 15560
rect 70196 15520 70197 15560
rect 70155 15511 70197 15520
rect 70347 15560 70389 15569
rect 70347 15520 70348 15560
rect 70388 15520 70389 15560
rect 70347 15511 70389 15520
rect 70915 15560 70973 15561
rect 70915 15520 70924 15560
rect 70964 15520 70973 15560
rect 70915 15519 70973 15520
rect 71019 15560 71061 15569
rect 71019 15520 71020 15560
rect 71060 15520 71061 15560
rect 71019 15511 71061 15520
rect 71115 15560 71157 15569
rect 71115 15520 71116 15560
rect 71156 15520 71157 15560
rect 71115 15511 71157 15520
rect 75139 15560 75197 15561
rect 75139 15520 75148 15560
rect 75188 15520 75197 15560
rect 75139 15519 75197 15520
rect 75339 15560 75381 15569
rect 75339 15520 75340 15560
rect 75380 15520 75381 15560
rect 75339 15511 75381 15520
rect 79363 15560 79421 15561
rect 79363 15520 79372 15560
rect 79412 15520 79421 15560
rect 79363 15519 79421 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 49987 15476 50045 15477
rect 49987 15436 49996 15476
rect 50036 15436 50045 15476
rect 49987 15435 50045 15436
rect 50371 15476 50429 15477
rect 50371 15436 50380 15476
rect 50420 15436 50429 15476
rect 50371 15435 50429 15436
rect 60355 15476 60413 15477
rect 60355 15436 60364 15476
rect 60404 15436 60413 15476
rect 60355 15435 60413 15436
rect 68707 15476 68765 15477
rect 68707 15436 68716 15476
rect 68756 15436 68765 15476
rect 68707 15435 68765 15436
rect 69859 15476 69917 15477
rect 69859 15436 69868 15476
rect 69908 15436 69917 15476
rect 69859 15435 69917 15436
rect 70723 15476 70781 15477
rect 70723 15436 70732 15476
rect 70772 15436 70781 15476
rect 70723 15435 70781 15436
rect 5067 15392 5109 15401
rect 5067 15352 5068 15392
rect 5108 15352 5109 15392
rect 5067 15343 5109 15352
rect 31563 15392 31605 15401
rect 31563 15352 31564 15392
rect 31604 15352 31605 15392
rect 31563 15343 31605 15352
rect 34923 15392 34965 15401
rect 34923 15352 34924 15392
rect 34964 15352 34965 15392
rect 34923 15343 34965 15352
rect 35691 15392 35733 15401
rect 35691 15352 35692 15392
rect 35732 15352 35733 15392
rect 35691 15343 35733 15352
rect 38091 15392 38133 15401
rect 38091 15352 38092 15392
rect 38132 15352 38133 15392
rect 38091 15343 38133 15352
rect 40875 15392 40917 15401
rect 40875 15352 40876 15392
rect 40916 15352 40917 15392
rect 40875 15343 40917 15352
rect 43851 15392 43893 15401
rect 43851 15352 43852 15392
rect 43892 15352 43893 15392
rect 43851 15343 43893 15352
rect 48459 15392 48501 15401
rect 48459 15352 48460 15392
rect 48500 15352 48501 15392
rect 48459 15343 48501 15352
rect 49131 15392 49173 15401
rect 49131 15352 49132 15392
rect 49172 15352 49173 15392
rect 49131 15343 49173 15352
rect 52011 15392 52053 15401
rect 52011 15352 52012 15392
rect 52052 15352 52053 15392
rect 52011 15343 52053 15352
rect 60171 15392 60213 15401
rect 60171 15352 60172 15392
rect 60212 15352 60213 15392
rect 60171 15343 60213 15352
rect 68043 15392 68085 15401
rect 68043 15352 68044 15392
rect 68084 15352 68085 15392
rect 68043 15343 68085 15352
rect 71307 15392 71349 15401
rect 71307 15352 71308 15392
rect 71348 15352 71349 15392
rect 71307 15343 71349 15352
rect 72651 15392 72693 15401
rect 72651 15352 72652 15392
rect 72692 15352 72693 15392
rect 72651 15343 72693 15352
rect 76683 15392 76725 15401
rect 76683 15352 76684 15392
rect 76724 15352 76725 15392
rect 76683 15343 76725 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 1123 15308 1181 15309
rect 1123 15268 1132 15308
rect 1172 15268 1181 15308
rect 1123 15267 1181 15268
rect 36747 15308 36789 15317
rect 36747 15268 36748 15308
rect 36788 15268 36789 15308
rect 36747 15259 36789 15268
rect 39427 15308 39485 15309
rect 39427 15268 39436 15308
rect 39476 15268 39485 15308
rect 39427 15267 39485 15268
rect 41835 15308 41877 15317
rect 41835 15268 41836 15308
rect 41876 15268 41877 15308
rect 41835 15259 41877 15268
rect 47595 15308 47637 15317
rect 47595 15268 47596 15308
rect 47636 15268 47637 15308
rect 47595 15259 47637 15268
rect 47979 15308 48021 15317
rect 47979 15268 47980 15308
rect 48020 15268 48021 15308
rect 47979 15259 48021 15268
rect 50187 15308 50229 15317
rect 50187 15268 50188 15308
rect 50228 15268 50229 15308
rect 50187 15259 50229 15268
rect 50571 15308 50613 15317
rect 50571 15268 50572 15308
rect 50612 15268 50613 15308
rect 50571 15259 50613 15268
rect 51051 15308 51093 15317
rect 51051 15268 51052 15308
rect 51092 15268 51093 15308
rect 51051 15259 51093 15268
rect 59491 15308 59549 15309
rect 59491 15268 59500 15308
rect 59540 15268 59549 15308
rect 59491 15267 59549 15268
rect 64971 15308 65013 15317
rect 64971 15268 64972 15308
rect 65012 15268 65013 15308
rect 64971 15259 65013 15268
rect 68907 15308 68949 15317
rect 68907 15268 68908 15308
rect 68948 15268 68949 15308
rect 68907 15259 68949 15268
rect 69675 15308 69717 15317
rect 69675 15268 69676 15308
rect 69716 15268 69717 15308
rect 69675 15259 69717 15268
rect 70347 15308 70389 15317
rect 70347 15268 70348 15308
rect 70388 15268 70389 15308
rect 70347 15259 70389 15268
rect 70539 15308 70581 15317
rect 70539 15268 70540 15308
rect 70580 15268 70581 15308
rect 70539 15259 70581 15268
rect 75243 15308 75285 15317
rect 75243 15268 75244 15308
rect 75284 15268 75285 15308
rect 75243 15259 75285 15268
rect 576 15140 79584 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79584 15140
rect 576 15076 79584 15100
rect 1515 14972 1557 14981
rect 1515 14932 1516 14972
rect 1556 14932 1557 14972
rect 1515 14923 1557 14932
rect 3619 14972 3677 14973
rect 3619 14932 3628 14972
rect 3668 14932 3677 14972
rect 3619 14931 3677 14932
rect 32907 14972 32949 14981
rect 32907 14932 32908 14972
rect 32948 14932 32949 14972
rect 32907 14923 32949 14932
rect 34819 14972 34877 14973
rect 34819 14932 34828 14972
rect 34868 14932 34877 14972
rect 34819 14931 34877 14932
rect 46347 14972 46389 14981
rect 46347 14932 46348 14972
rect 46388 14932 46389 14972
rect 46347 14923 46389 14932
rect 47683 14972 47741 14973
rect 47683 14932 47692 14972
rect 47732 14932 47741 14972
rect 47683 14931 47741 14932
rect 50371 14972 50429 14973
rect 50371 14932 50380 14972
rect 50420 14932 50429 14972
rect 50371 14931 50429 14932
rect 53155 14972 53213 14973
rect 53155 14932 53164 14972
rect 53204 14932 53213 14972
rect 53155 14931 53213 14932
rect 56907 14972 56949 14981
rect 56907 14932 56908 14972
rect 56948 14932 56949 14972
rect 56907 14923 56949 14932
rect 60555 14972 60597 14981
rect 60555 14932 60556 14972
rect 60596 14932 60597 14972
rect 60555 14923 60597 14932
rect 65451 14972 65493 14981
rect 65451 14932 65452 14972
rect 65492 14932 65493 14972
rect 65451 14923 65493 14932
rect 72739 14972 72797 14973
rect 72739 14932 72748 14972
rect 72788 14932 72797 14972
rect 72739 14931 72797 14932
rect 75331 14972 75389 14973
rect 75331 14932 75340 14972
rect 75380 14932 75389 14972
rect 75331 14931 75389 14932
rect 1995 14888 2037 14897
rect 1995 14848 1996 14888
rect 2036 14848 2037 14888
rect 1995 14839 2037 14848
rect 40011 14888 40053 14897
rect 40011 14848 40012 14888
rect 40052 14848 40053 14888
rect 40011 14839 40053 14848
rect 45099 14888 45141 14897
rect 45099 14848 45100 14888
rect 45140 14848 45141 14888
rect 45099 14839 45141 14848
rect 56707 14888 56765 14889
rect 56707 14848 56716 14888
rect 56756 14848 56765 14888
rect 56707 14847 56765 14848
rect 57483 14888 57525 14897
rect 57483 14848 57484 14888
rect 57524 14848 57525 14888
rect 57483 14839 57525 14848
rect 58635 14888 58677 14897
rect 58635 14848 58636 14888
rect 58676 14848 58677 14888
rect 58635 14839 58677 14848
rect 60171 14888 60213 14897
rect 60171 14848 60172 14888
rect 60212 14848 60213 14888
rect 60171 14839 60213 14848
rect 61795 14888 61853 14889
rect 61795 14848 61804 14888
rect 61844 14848 61853 14888
rect 61795 14847 61853 14848
rect 64195 14888 64253 14889
rect 64195 14848 64204 14888
rect 64244 14848 64253 14888
rect 64195 14847 64253 14848
rect 65931 14888 65973 14897
rect 65931 14848 65932 14888
rect 65972 14848 65973 14888
rect 65931 14839 65973 14848
rect 75531 14888 75573 14897
rect 75531 14848 75532 14888
rect 75572 14848 75573 14888
rect 75531 14839 75573 14848
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 1315 14804 1373 14805
rect 1315 14764 1324 14804
rect 1364 14764 1373 14804
rect 1315 14763 1373 14764
rect 1699 14804 1757 14805
rect 1699 14764 1708 14804
rect 1748 14764 1757 14804
rect 1699 14763 1757 14764
rect 2179 14804 2237 14805
rect 2179 14764 2188 14804
rect 2228 14764 2237 14804
rect 2179 14763 2237 14764
rect 60355 14804 60413 14805
rect 60355 14764 60364 14804
rect 60404 14764 60413 14804
rect 60355 14763 60413 14764
rect 62179 14804 62237 14805
rect 62179 14764 62188 14804
rect 62228 14764 62237 14804
rect 62179 14763 62237 14764
rect 62947 14804 63005 14805
rect 62947 14764 62956 14804
rect 62996 14764 63005 14804
rect 62947 14763 63005 14764
rect 63915 14804 63957 14813
rect 63915 14764 63916 14804
rect 63956 14764 63957 14804
rect 63915 14755 63957 14764
rect 67171 14804 67229 14805
rect 67171 14764 67180 14804
rect 67220 14764 67229 14804
rect 67171 14763 67229 14764
rect 2379 14720 2421 14729
rect 2379 14680 2380 14720
rect 2420 14680 2421 14720
rect 2379 14671 2421 14680
rect 2475 14720 2517 14729
rect 2475 14680 2476 14720
rect 2516 14680 2517 14720
rect 2475 14671 2517 14680
rect 2571 14720 2613 14729
rect 2571 14680 2572 14720
rect 2612 14680 2613 14720
rect 2571 14671 2613 14680
rect 2667 14720 2709 14729
rect 2667 14680 2668 14720
rect 2708 14680 2709 14720
rect 2667 14671 2709 14680
rect 2947 14720 3005 14721
rect 2947 14680 2956 14720
rect 2996 14680 3005 14720
rect 2947 14679 3005 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3339 14720 3381 14729
rect 3339 14680 3340 14720
rect 3380 14680 3381 14720
rect 3339 14671 3381 14680
rect 30219 14720 30261 14729
rect 30219 14680 30220 14720
rect 30260 14680 30261 14720
rect 30219 14671 30261 14680
rect 30595 14720 30653 14721
rect 30595 14680 30604 14720
rect 30644 14680 30653 14720
rect 30595 14679 30653 14680
rect 31459 14720 31517 14721
rect 31459 14680 31468 14720
rect 31508 14680 31517 14720
rect 31459 14679 31517 14680
rect 32803 14720 32861 14721
rect 32803 14680 32812 14720
rect 32852 14680 32861 14720
rect 32803 14679 32861 14680
rect 33003 14720 33045 14729
rect 33003 14680 33004 14720
rect 33044 14680 33045 14720
rect 33003 14671 33045 14680
rect 33195 14720 33237 14729
rect 33195 14680 33196 14720
rect 33236 14680 33237 14720
rect 33195 14671 33237 14680
rect 33387 14720 33429 14729
rect 33387 14680 33388 14720
rect 33428 14680 33429 14720
rect 33387 14671 33429 14680
rect 33475 14720 33533 14721
rect 33475 14680 33484 14720
rect 33524 14680 33533 14720
rect 33475 14679 33533 14680
rect 35971 14720 36029 14721
rect 35971 14680 35980 14720
rect 36020 14680 36029 14720
rect 35971 14679 36029 14680
rect 36835 14720 36893 14721
rect 36835 14680 36844 14720
rect 36884 14680 36893 14720
rect 36835 14679 36893 14680
rect 37227 14720 37269 14729
rect 37227 14680 37228 14720
rect 37268 14680 37269 14720
rect 37227 14671 37269 14680
rect 38563 14720 38621 14721
rect 38563 14680 38572 14720
rect 38612 14680 38621 14720
rect 38563 14679 38621 14680
rect 39427 14720 39485 14721
rect 39427 14680 39436 14720
rect 39476 14680 39485 14720
rect 39427 14679 39485 14680
rect 39819 14720 39861 14729
rect 39819 14680 39820 14720
rect 39860 14680 39861 14720
rect 39819 14671 39861 14680
rect 40011 14720 40053 14729
rect 40011 14680 40012 14720
rect 40052 14680 40053 14720
rect 40011 14671 40053 14680
rect 40203 14720 40245 14729
rect 40203 14680 40204 14720
rect 40244 14680 40245 14720
rect 40203 14671 40245 14680
rect 40291 14720 40349 14721
rect 40291 14680 40300 14720
rect 40340 14680 40349 14720
rect 40291 14679 40349 14680
rect 41163 14720 41205 14729
rect 41163 14680 41164 14720
rect 41204 14680 41205 14720
rect 41163 14671 41205 14680
rect 41259 14720 41301 14729
rect 41259 14680 41260 14720
rect 41300 14680 41301 14720
rect 41259 14671 41301 14680
rect 41355 14720 41397 14729
rect 41355 14680 41356 14720
rect 41396 14680 41397 14720
rect 41355 14671 41397 14680
rect 42699 14720 42741 14729
rect 42699 14680 42700 14720
rect 42740 14680 42741 14720
rect 42699 14671 42741 14680
rect 42891 14720 42933 14729
rect 42891 14680 42892 14720
rect 42932 14680 42933 14720
rect 42891 14671 42933 14680
rect 42979 14720 43037 14721
rect 42979 14680 42988 14720
rect 43028 14680 43037 14720
rect 42979 14679 43037 14680
rect 43171 14720 43229 14721
rect 43171 14680 43180 14720
rect 43220 14680 43229 14720
rect 43171 14679 43229 14680
rect 43275 14720 43317 14729
rect 43275 14680 43276 14720
rect 43316 14680 43317 14720
rect 43275 14671 43317 14680
rect 43371 14720 43413 14729
rect 43371 14680 43372 14720
rect 43412 14680 43413 14720
rect 43371 14671 43413 14680
rect 46051 14720 46109 14721
rect 46051 14680 46060 14720
rect 46100 14680 46109 14720
rect 46051 14679 46109 14680
rect 46155 14720 46197 14729
rect 46155 14680 46156 14720
rect 46196 14680 46197 14720
rect 46155 14671 46197 14680
rect 46347 14720 46389 14729
rect 46347 14680 46348 14720
rect 46388 14680 46389 14720
rect 46347 14671 46389 14680
rect 47011 14720 47069 14721
rect 47011 14680 47020 14720
rect 47060 14680 47069 14720
rect 47011 14679 47069 14680
rect 47307 14720 47349 14729
rect 47307 14680 47308 14720
rect 47348 14680 47349 14720
rect 47307 14671 47349 14680
rect 48355 14720 48413 14721
rect 48355 14680 48364 14720
rect 48404 14680 48413 14720
rect 48355 14679 48413 14680
rect 49219 14720 49277 14721
rect 49219 14680 49228 14720
rect 49268 14680 49277 14720
rect 49219 14679 49277 14680
rect 51139 14720 51197 14721
rect 51139 14680 51148 14720
rect 51188 14680 51197 14720
rect 51139 14679 51197 14680
rect 52003 14720 52061 14721
rect 52003 14680 52012 14720
rect 52052 14680 52061 14720
rect 52003 14679 52061 14680
rect 53443 14720 53501 14721
rect 53443 14680 53452 14720
rect 53492 14680 53501 14720
rect 53443 14679 53501 14680
rect 54891 14720 54933 14729
rect 54891 14680 54892 14720
rect 54932 14680 54933 14720
rect 54891 14671 54933 14680
rect 56035 14720 56093 14721
rect 56035 14680 56044 14720
rect 56084 14680 56093 14720
rect 56035 14679 56093 14680
rect 56331 14720 56373 14729
rect 56331 14680 56332 14720
rect 56372 14680 56373 14720
rect 56331 14671 56373 14680
rect 56907 14720 56949 14729
rect 56907 14680 56908 14720
rect 56948 14680 56949 14720
rect 56907 14671 56949 14680
rect 57099 14720 57141 14729
rect 57099 14680 57100 14720
rect 57140 14680 57141 14720
rect 57099 14671 57141 14680
rect 57187 14720 57245 14721
rect 57187 14680 57196 14720
rect 57236 14680 57245 14720
rect 57187 14679 57245 14680
rect 57379 14720 57437 14721
rect 57379 14680 57388 14720
rect 57428 14680 57437 14720
rect 57379 14679 57437 14680
rect 57579 14720 57621 14729
rect 57579 14680 57580 14720
rect 57620 14680 57621 14720
rect 57579 14671 57621 14680
rect 60555 14720 60597 14729
rect 60555 14680 60556 14720
rect 60596 14680 60597 14720
rect 60555 14671 60597 14680
rect 60747 14720 60789 14729
rect 60747 14680 60748 14720
rect 60788 14680 60789 14720
rect 60747 14671 60789 14680
rect 60835 14720 60893 14721
rect 60835 14680 60844 14720
rect 60884 14680 60893 14720
rect 60835 14679 60893 14680
rect 61123 14720 61181 14721
rect 61123 14680 61132 14720
rect 61172 14680 61181 14720
rect 61123 14679 61181 14680
rect 61419 14720 61461 14729
rect 61419 14680 61420 14720
rect 61460 14680 61461 14720
rect 61419 14671 61461 14680
rect 62371 14720 62429 14721
rect 62371 14680 62380 14720
rect 62420 14680 62429 14720
rect 62371 14679 62429 14680
rect 62475 14720 62517 14729
rect 62475 14680 62476 14720
rect 62516 14680 62517 14720
rect 62475 14671 62517 14680
rect 62571 14720 62613 14729
rect 62571 14680 62572 14720
rect 62612 14680 62613 14720
rect 62571 14671 62613 14680
rect 63811 14720 63869 14721
rect 63811 14680 63820 14720
rect 63860 14680 63869 14720
rect 63811 14679 63869 14680
rect 64011 14720 64053 14729
rect 64011 14680 64012 14720
rect 64052 14680 64053 14720
rect 64011 14671 64053 14680
rect 64587 14720 64629 14729
rect 64587 14680 64588 14720
rect 64628 14680 64629 14720
rect 64587 14671 64629 14680
rect 64867 14720 64925 14721
rect 64867 14680 64876 14720
rect 64916 14680 64925 14720
rect 64867 14679 64925 14680
rect 65155 14720 65213 14721
rect 65155 14680 65164 14720
rect 65204 14680 65213 14720
rect 65155 14679 65213 14680
rect 65259 14720 65301 14729
rect 65259 14680 65260 14720
rect 65300 14680 65301 14720
rect 65259 14671 65301 14680
rect 65451 14720 65493 14729
rect 65451 14680 65452 14720
rect 65492 14680 65493 14720
rect 65451 14671 65493 14680
rect 67939 14720 67997 14721
rect 67939 14680 67948 14720
rect 67988 14680 67997 14720
rect 67939 14679 67997 14680
rect 68803 14720 68861 14721
rect 68803 14680 68812 14720
rect 68852 14680 68861 14720
rect 68803 14679 68861 14680
rect 70347 14720 70389 14729
rect 70347 14680 70348 14720
rect 70388 14680 70389 14720
rect 70347 14671 70389 14680
rect 70723 14720 70781 14721
rect 70723 14680 70732 14720
rect 70772 14680 70781 14720
rect 70723 14679 70781 14680
rect 71587 14720 71645 14721
rect 71587 14680 71596 14720
rect 71636 14680 71645 14720
rect 71587 14679 71645 14680
rect 73611 14720 73653 14729
rect 73611 14680 73612 14720
rect 73652 14680 73653 14720
rect 73611 14671 73653 14680
rect 73803 14720 73845 14729
rect 73803 14680 73804 14720
rect 73844 14680 73845 14720
rect 73803 14671 73845 14680
rect 73891 14720 73949 14721
rect 73891 14680 73900 14720
rect 73940 14680 73949 14720
rect 73891 14679 73949 14680
rect 74091 14720 74133 14729
rect 74091 14680 74092 14720
rect 74132 14680 74133 14720
rect 74091 14671 74133 14680
rect 74187 14720 74229 14729
rect 74187 14680 74188 14720
rect 74228 14680 74229 14720
rect 74187 14671 74229 14680
rect 74283 14720 74325 14729
rect 74283 14680 74284 14720
rect 74324 14680 74325 14720
rect 74283 14671 74325 14680
rect 74379 14720 74421 14729
rect 74379 14680 74380 14720
rect 74420 14680 74421 14720
rect 74379 14671 74421 14680
rect 74659 14720 74717 14721
rect 74659 14680 74668 14720
rect 74708 14680 74717 14720
rect 74659 14679 74717 14680
rect 74955 14720 74997 14729
rect 74955 14680 74956 14720
rect 74996 14680 74997 14720
rect 75723 14720 75765 14729
rect 74955 14671 74997 14680
rect 75531 14678 75573 14687
rect 47403 14636 47445 14645
rect 47403 14596 47404 14636
rect 47444 14596 47445 14636
rect 47403 14587 47445 14596
rect 47979 14636 48021 14645
rect 47979 14596 47980 14636
rect 48020 14596 48021 14636
rect 47979 14587 48021 14596
rect 50763 14636 50805 14645
rect 50763 14596 50764 14636
rect 50804 14596 50805 14636
rect 50763 14587 50805 14596
rect 56427 14636 56469 14645
rect 56427 14596 56428 14636
rect 56468 14596 56469 14636
rect 56427 14587 56469 14596
rect 61515 14636 61557 14645
rect 61515 14596 61516 14636
rect 61556 14596 61557 14636
rect 61515 14587 61557 14596
rect 64491 14636 64533 14645
rect 64491 14596 64492 14636
rect 64532 14596 64533 14636
rect 64491 14587 64533 14596
rect 67563 14636 67605 14645
rect 67563 14596 67564 14636
rect 67604 14596 67605 14636
rect 67563 14587 67605 14596
rect 75051 14636 75093 14645
rect 75051 14596 75052 14636
rect 75092 14596 75093 14636
rect 75531 14638 75532 14678
rect 75572 14638 75573 14678
rect 75723 14680 75724 14720
rect 75764 14680 75765 14720
rect 75723 14671 75765 14680
rect 75811 14720 75869 14721
rect 75811 14680 75820 14720
rect 75860 14680 75869 14720
rect 75811 14679 75869 14680
rect 76203 14720 76245 14729
rect 76203 14680 76204 14720
rect 76244 14680 76245 14720
rect 76203 14671 76245 14680
rect 76579 14720 76637 14721
rect 76579 14680 76588 14720
rect 76628 14680 76637 14720
rect 76579 14679 76637 14680
rect 77443 14720 77501 14721
rect 77443 14680 77452 14720
rect 77492 14680 77501 14720
rect 77443 14679 77501 14680
rect 75531 14629 75573 14638
rect 75051 14587 75093 14596
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 1131 14552 1173 14561
rect 1131 14512 1132 14552
rect 1172 14512 1173 14552
rect 1131 14503 1173 14512
rect 32611 14552 32669 14553
rect 32611 14512 32620 14552
rect 32660 14512 32669 14552
rect 32611 14511 32669 14512
rect 33283 14552 33341 14553
rect 33283 14512 33292 14552
rect 33332 14512 33341 14552
rect 33283 14511 33341 14512
rect 37411 14552 37469 14553
rect 37411 14512 37420 14552
rect 37460 14512 37469 14552
rect 37411 14511 37469 14512
rect 41443 14552 41501 14553
rect 41443 14512 41452 14552
rect 41492 14512 41501 14552
rect 41443 14511 41501 14512
rect 42787 14552 42845 14553
rect 42787 14512 42796 14552
rect 42836 14512 42845 14552
rect 42787 14511 42845 14512
rect 53155 14552 53213 14553
rect 53155 14512 53164 14552
rect 53204 14512 53213 14552
rect 53155 14511 53213 14512
rect 61995 14552 62037 14561
rect 61995 14512 61996 14552
rect 62036 14512 62037 14552
rect 61995 14503 62037 14512
rect 62763 14552 62805 14561
rect 62763 14512 62764 14552
rect 62804 14512 62805 14552
rect 62763 14503 62805 14512
rect 67371 14552 67413 14561
rect 67371 14512 67372 14552
rect 67412 14512 67413 14552
rect 67371 14503 67413 14512
rect 69955 14552 70013 14553
rect 69955 14512 69964 14552
rect 70004 14512 70013 14552
rect 69955 14511 70013 14512
rect 73699 14552 73757 14553
rect 73699 14512 73708 14552
rect 73748 14512 73757 14552
rect 73699 14511 73757 14512
rect 78595 14552 78653 14553
rect 78595 14512 78604 14552
rect 78644 14512 78653 14552
rect 78595 14511 78653 14512
rect 576 14384 79584 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79584 14384
rect 576 14320 79584 14344
rect 1323 14216 1365 14225
rect 1323 14176 1324 14216
rect 1364 14176 1365 14216
rect 1323 14167 1365 14176
rect 2851 14216 2909 14217
rect 2851 14176 2860 14216
rect 2900 14176 2909 14216
rect 2851 14175 2909 14176
rect 7267 14216 7325 14217
rect 7267 14176 7276 14216
rect 7316 14176 7325 14216
rect 7267 14175 7325 14176
rect 38563 14216 38621 14217
rect 38563 14176 38572 14216
rect 38612 14176 38621 14216
rect 38563 14175 38621 14176
rect 39427 14216 39485 14217
rect 39427 14176 39436 14216
rect 39476 14176 39485 14216
rect 39427 14175 39485 14176
rect 40003 14216 40061 14217
rect 40003 14176 40012 14216
rect 40052 14176 40061 14216
rect 40003 14175 40061 14176
rect 42691 14216 42749 14217
rect 42691 14176 42700 14216
rect 42740 14176 42749 14216
rect 42691 14175 42749 14176
rect 47011 14216 47069 14217
rect 47011 14176 47020 14216
rect 47060 14176 47069 14216
rect 47011 14175 47069 14176
rect 56131 14216 56189 14217
rect 56131 14176 56140 14216
rect 56180 14176 56189 14216
rect 56131 14175 56189 14176
rect 60547 14216 60605 14217
rect 60547 14176 60556 14216
rect 60596 14176 60605 14216
rect 60547 14175 60605 14176
rect 61035 14216 61077 14225
rect 61035 14176 61036 14216
rect 61076 14176 61077 14216
rect 61035 14167 61077 14176
rect 66979 14216 67037 14217
rect 66979 14176 66988 14216
rect 67028 14176 67037 14216
rect 66979 14175 67037 14176
rect 69003 14216 69045 14225
rect 69003 14176 69004 14216
rect 69044 14176 69045 14216
rect 69003 14167 69045 14176
rect 70731 14216 70773 14225
rect 70731 14176 70732 14216
rect 70772 14176 70773 14216
rect 70731 14167 70773 14176
rect 71115 14216 71157 14225
rect 71115 14176 71116 14216
rect 71156 14176 71157 14216
rect 71115 14167 71157 14176
rect 79363 14216 79421 14217
rect 79363 14176 79372 14216
rect 79412 14176 79421 14216
rect 79363 14175 79421 14176
rect 43179 14132 43221 14141
rect 43179 14092 43180 14132
rect 43220 14092 43221 14132
rect 43179 14083 43221 14092
rect 47691 14132 47733 14141
rect 47691 14092 47692 14132
rect 47732 14092 47733 14132
rect 47691 14083 47733 14092
rect 52587 14132 52629 14141
rect 52587 14092 52588 14132
rect 52628 14092 52629 14132
rect 52587 14083 52629 14092
rect 67467 14132 67509 14141
rect 67467 14092 67468 14132
rect 67508 14092 67509 14132
rect 67467 14083 67509 14092
rect 70059 14132 70101 14141
rect 70059 14092 70060 14132
rect 70100 14092 70101 14132
rect 70059 14083 70101 14092
rect 72171 14132 72213 14141
rect 72171 14092 72172 14132
rect 72212 14092 72213 14132
rect 72171 14083 72213 14092
rect 75915 14132 75957 14141
rect 75915 14092 75916 14132
rect 75956 14092 75957 14132
rect 75915 14083 75957 14092
rect 57763 14069 57821 14070
rect 53241 14063 53299 14064
rect 2091 14048 2133 14057
rect 2091 14008 2092 14048
rect 2132 14008 2133 14048
rect 2091 13999 2133 14008
rect 2187 14048 2229 14057
rect 2187 14008 2188 14048
rect 2228 14008 2229 14048
rect 2187 13999 2229 14008
rect 2283 14048 2325 14057
rect 2283 14008 2284 14048
rect 2324 14008 2325 14048
rect 2283 13999 2325 14008
rect 2379 14048 2421 14057
rect 2379 14008 2380 14048
rect 2420 14008 2421 14048
rect 2379 13999 2421 14008
rect 2659 14048 2717 14049
rect 2659 14008 2668 14048
rect 2708 14008 2717 14048
rect 2659 14007 2717 14008
rect 2763 14048 2805 14057
rect 2763 14008 2764 14048
rect 2804 14008 2805 14048
rect 2763 13999 2805 14008
rect 2955 14048 2997 14057
rect 2955 14008 2956 14048
rect 2996 14008 2997 14048
rect 2955 13999 2997 14008
rect 3235 14048 3293 14049
rect 3235 14008 3244 14048
rect 3284 14008 3293 14048
rect 3235 14007 3293 14008
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 3531 13999 3573 14008
rect 3627 14048 3669 14057
rect 3627 14008 3628 14048
rect 3668 14008 3669 14048
rect 3627 13999 3669 14008
rect 4387 14048 4445 14049
rect 4387 14008 4396 14048
rect 4436 14008 4445 14048
rect 4387 14007 4445 14008
rect 4491 14048 4533 14057
rect 4491 14008 4492 14048
rect 4532 14008 4533 14048
rect 4491 13999 4533 14008
rect 4683 14048 4725 14057
rect 4683 14008 4684 14048
rect 4724 14008 4725 14048
rect 4683 13999 4725 14008
rect 4875 14048 4917 14057
rect 4875 14008 4876 14048
rect 4916 14008 4917 14048
rect 4875 13999 4917 14008
rect 5251 14048 5309 14049
rect 5251 14008 5260 14048
rect 5300 14008 5309 14048
rect 5251 14007 5309 14008
rect 6115 14048 6173 14049
rect 6115 14008 6124 14048
rect 6164 14008 6173 14048
rect 6115 14007 6173 14008
rect 31659 14048 31701 14057
rect 31659 14008 31660 14048
rect 31700 14008 31701 14048
rect 31659 13999 31701 14008
rect 31755 14048 31797 14057
rect 31755 14008 31756 14048
rect 31796 14008 31797 14048
rect 31755 13999 31797 14008
rect 31851 14048 31893 14057
rect 31851 14008 31852 14048
rect 31892 14008 31893 14048
rect 31851 13999 31893 14008
rect 31947 14048 31989 14057
rect 31947 14008 31948 14048
rect 31988 14008 31989 14048
rect 31947 13999 31989 14008
rect 32227 14048 32285 14049
rect 32227 14008 32236 14048
rect 32276 14008 32285 14048
rect 32227 14007 32285 14008
rect 32523 14048 32565 14057
rect 32523 14008 32524 14048
rect 32564 14008 32565 14048
rect 32523 13999 32565 14008
rect 32619 14048 32661 14057
rect 32619 14008 32620 14048
rect 32660 14008 32661 14048
rect 33475 14048 33533 14049
rect 32619 13999 32661 14008
rect 33099 14006 33141 14015
rect 33475 14008 33484 14048
rect 33524 14008 33533 14048
rect 33475 14007 33533 14008
rect 34339 14048 34397 14049
rect 34339 14008 34348 14048
rect 34388 14008 34397 14048
rect 34339 14007 34397 14008
rect 37315 14048 37373 14049
rect 37315 14008 37324 14048
rect 37364 14008 37373 14048
rect 37315 14007 37373 14008
rect 38275 14048 38333 14049
rect 38275 14008 38284 14048
rect 38324 14008 38333 14048
rect 38275 14007 38333 14008
rect 38475 14048 38517 14057
rect 38475 14008 38476 14048
rect 38516 14008 38517 14048
rect 33099 13966 33100 14006
rect 33140 13966 33141 14006
rect 38475 13999 38517 14008
rect 38667 14048 38709 14057
rect 38667 14008 38668 14048
rect 38708 14008 38709 14048
rect 38667 13999 38709 14008
rect 38755 14048 38813 14049
rect 38755 14008 38764 14048
rect 38804 14008 38813 14048
rect 38755 14007 38813 14008
rect 39147 14048 39189 14057
rect 39147 14008 39148 14048
rect 39188 14008 39189 14048
rect 39147 13999 39189 14008
rect 39243 14048 39285 14057
rect 39243 14008 39244 14048
rect 39284 14008 39285 14048
rect 39243 13999 39285 14008
rect 39339 14048 39381 14057
rect 39339 14008 39340 14048
rect 39380 14008 39381 14048
rect 39339 13999 39381 14008
rect 39811 14048 39869 14049
rect 39811 14008 39820 14048
rect 39860 14008 39869 14048
rect 39811 14007 39869 14008
rect 39915 14048 39957 14057
rect 39915 14008 39916 14048
rect 39956 14008 39957 14048
rect 39915 13999 39957 14008
rect 40107 14048 40149 14057
rect 40107 14008 40108 14048
rect 40148 14008 40149 14048
rect 40107 13999 40149 14008
rect 40299 14048 40341 14057
rect 40299 14008 40300 14048
rect 40340 14008 40341 14048
rect 40299 13999 40341 14008
rect 40675 14048 40733 14049
rect 40675 14008 40684 14048
rect 40724 14008 40733 14048
rect 40675 14007 40733 14008
rect 41539 14048 41597 14049
rect 41539 14008 41548 14048
rect 41588 14008 41597 14048
rect 41539 14007 41597 14008
rect 43275 14048 43317 14057
rect 43275 14008 43276 14048
rect 43316 14008 43317 14048
rect 43275 13999 43317 14008
rect 43555 14048 43613 14049
rect 43555 14008 43564 14048
rect 43604 14008 43613 14048
rect 43555 14007 43613 14008
rect 44619 14048 44661 14057
rect 44619 14008 44620 14048
rect 44660 14008 44661 14048
rect 44619 13999 44661 14008
rect 44995 14048 45053 14049
rect 44995 14008 45004 14048
rect 45044 14008 45053 14048
rect 44995 14007 45053 14008
rect 45859 14048 45917 14049
rect 45859 14008 45868 14048
rect 45908 14008 45917 14048
rect 45859 14007 45917 14008
rect 47203 14048 47261 14049
rect 47203 14008 47212 14048
rect 47252 14008 47261 14048
rect 47203 14007 47261 14008
rect 47595 14048 47637 14057
rect 47595 14008 47596 14048
rect 47636 14008 47637 14048
rect 47595 13999 47637 14008
rect 47787 14048 47829 14057
rect 47787 14008 47788 14048
rect 47828 14008 47829 14048
rect 47787 13999 47829 14008
rect 47875 14048 47933 14049
rect 47875 14008 47884 14048
rect 47924 14008 47933 14048
rect 47875 14007 47933 14008
rect 51139 14048 51197 14049
rect 51139 14008 51148 14048
rect 51188 14008 51197 14048
rect 51139 14007 51197 14008
rect 51243 14048 51285 14057
rect 51243 14008 51244 14048
rect 51284 14008 51285 14048
rect 51243 13999 51285 14008
rect 51435 14048 51477 14057
rect 51435 14008 51436 14048
rect 51476 14008 51477 14048
rect 51435 13999 51477 14008
rect 52491 14048 52533 14057
rect 52491 14008 52492 14048
rect 52532 14008 52533 14048
rect 52491 13999 52533 14008
rect 52675 14048 52733 14049
rect 52675 14008 52684 14048
rect 52724 14008 52733 14048
rect 53241 14023 53250 14063
rect 53290 14023 53299 14063
rect 53241 14022 53299 14023
rect 53355 14048 53397 14057
rect 52675 14007 52733 14008
rect 53355 14008 53356 14048
rect 53396 14008 53397 14048
rect 53355 13999 53397 14008
rect 53547 14048 53589 14057
rect 53547 14008 53548 14048
rect 53588 14008 53589 14048
rect 53547 13999 53589 14008
rect 53739 14048 53781 14057
rect 53739 14008 53740 14048
rect 53780 14008 53781 14048
rect 53739 13999 53781 14008
rect 54115 14048 54173 14049
rect 54115 14008 54124 14048
rect 54164 14008 54173 14048
rect 54115 14007 54173 14008
rect 54979 14048 55037 14049
rect 54979 14008 54988 14048
rect 55028 14008 55037 14048
rect 54979 14007 55037 14008
rect 56419 14048 56477 14049
rect 56419 14008 56428 14048
rect 56468 14008 56477 14048
rect 56419 14007 56477 14008
rect 56619 14048 56661 14057
rect 56619 14008 56620 14048
rect 56660 14008 56661 14048
rect 57763 14029 57772 14069
rect 57812 14029 57821 14069
rect 57763 14028 57821 14029
rect 57963 14048 58005 14057
rect 56619 13999 56661 14008
rect 57963 14008 57964 14048
rect 58004 14008 58005 14048
rect 57963 13999 58005 14008
rect 58155 14048 58197 14057
rect 58155 14008 58156 14048
rect 58196 14008 58197 14048
rect 58155 13999 58197 14008
rect 58531 14048 58589 14049
rect 58531 14008 58540 14048
rect 58580 14008 58589 14048
rect 58531 14007 58589 14008
rect 59395 14048 59453 14049
rect 59395 14008 59404 14048
rect 59444 14008 59453 14048
rect 59395 14007 59453 14008
rect 61227 14048 61269 14057
rect 61227 14008 61228 14048
rect 61268 14008 61269 14048
rect 61227 13999 61269 14008
rect 61603 14048 61661 14049
rect 61603 14008 61612 14048
rect 61652 14008 61661 14048
rect 61603 14007 61661 14008
rect 62467 14048 62525 14049
rect 62467 14008 62476 14048
rect 62516 14008 62525 14048
rect 62467 14007 62525 14008
rect 63811 14048 63869 14049
rect 63811 14008 63820 14048
rect 63860 14008 63869 14048
rect 63811 14007 63869 14008
rect 63915 14048 63957 14057
rect 63915 14008 63916 14048
rect 63956 14008 63957 14048
rect 63915 13999 63957 14008
rect 64107 14048 64149 14057
rect 64107 14008 64108 14048
rect 64148 14008 64149 14048
rect 64107 13999 64149 14008
rect 64587 14048 64629 14057
rect 64587 14008 64588 14048
rect 64628 14008 64629 14048
rect 64587 13999 64629 14008
rect 64963 14048 65021 14049
rect 64963 14008 64972 14048
rect 65012 14008 65021 14048
rect 64963 14007 65021 14008
rect 65827 14048 65885 14049
rect 65827 14008 65836 14048
rect 65876 14008 65885 14048
rect 65827 14007 65885 14008
rect 67267 14048 67325 14049
rect 67267 14008 67276 14048
rect 67316 14008 67325 14048
rect 67267 14007 67325 14008
rect 67371 14048 67413 14057
rect 67371 14008 67372 14048
rect 67412 14008 67413 14048
rect 67371 13999 67413 14008
rect 67563 14048 67605 14057
rect 67563 14008 67564 14048
rect 67604 14008 67605 14048
rect 67563 13999 67605 14008
rect 68035 14048 68093 14049
rect 68035 14008 68044 14048
rect 68084 14008 68093 14048
rect 68035 14007 68093 14008
rect 68139 14048 68181 14057
rect 68139 14008 68140 14048
rect 68180 14008 68181 14048
rect 68139 13999 68181 14008
rect 68331 14048 68373 14057
rect 68331 14008 68332 14048
rect 68372 14008 68373 14048
rect 68331 13999 68373 14008
rect 68523 14048 68565 14057
rect 68523 14008 68524 14048
rect 68564 14008 68565 14048
rect 68523 13999 68565 14008
rect 68619 14048 68661 14057
rect 68619 14008 68620 14048
rect 68660 14008 68661 14048
rect 68619 13999 68661 14008
rect 68715 14048 68757 14057
rect 68715 14008 68716 14048
rect 68756 14008 68757 14048
rect 68715 13999 68757 14008
rect 68811 14048 68853 14057
rect 68811 14008 68812 14048
rect 68852 14008 68853 14048
rect 68811 13999 68853 14008
rect 69667 14048 69725 14049
rect 69667 14008 69676 14048
rect 69716 14008 69725 14048
rect 69667 14007 69725 14008
rect 69963 14048 70005 14057
rect 69963 14008 69964 14048
rect 70004 14008 70005 14048
rect 69963 13999 70005 14008
rect 72547 14048 72605 14049
rect 72547 14008 72556 14048
rect 72596 14008 72605 14048
rect 72547 14007 72605 14008
rect 73436 14048 73494 14049
rect 73436 14008 73445 14048
rect 73485 14008 73494 14048
rect 73436 14007 73494 14008
rect 74763 14048 74805 14057
rect 74763 14008 74764 14048
rect 74804 14008 74805 14048
rect 74763 13999 74805 14008
rect 74955 14048 74997 14057
rect 74955 14008 74956 14048
rect 74996 14008 74997 14048
rect 74955 13999 74997 14008
rect 75043 14048 75101 14049
rect 75043 14008 75052 14048
rect 75092 14008 75101 14048
rect 75043 14007 75101 14008
rect 75811 14048 75869 14049
rect 75811 14008 75820 14048
rect 75860 14008 75869 14048
rect 75811 14007 75869 14008
rect 76011 14048 76053 14057
rect 76011 14008 76012 14048
rect 76052 14008 76053 14048
rect 76011 13999 76053 14008
rect 76971 14048 77013 14057
rect 76971 14008 76972 14048
rect 77012 14008 77013 14048
rect 76971 13999 77013 14008
rect 77347 14048 77405 14049
rect 77347 14008 77356 14048
rect 77396 14008 77405 14048
rect 77347 14007 77405 14008
rect 78211 14048 78269 14049
rect 78211 14008 78220 14048
rect 78260 14008 78269 14048
rect 78211 14007 78269 14008
rect 1507 13964 1565 13965
rect 1507 13924 1516 13964
rect 1556 13924 1565 13964
rect 33099 13957 33141 13966
rect 60835 13964 60893 13965
rect 1507 13923 1565 13924
rect 60835 13924 60844 13964
rect 60884 13924 60893 13964
rect 60835 13923 60893 13924
rect 63627 13964 63669 13973
rect 63627 13924 63628 13964
rect 63668 13924 63669 13964
rect 63627 13915 63669 13924
rect 69187 13964 69245 13965
rect 69187 13924 69196 13964
rect 69236 13924 69245 13964
rect 69187 13923 69245 13924
rect 70531 13964 70589 13965
rect 70531 13924 70540 13964
rect 70580 13924 70589 13964
rect 70531 13923 70589 13924
rect 70915 13964 70973 13965
rect 70915 13924 70924 13964
rect 70964 13924 70973 13964
rect 70915 13923 70973 13924
rect 1899 13880 1941 13889
rect 1899 13840 1900 13880
rect 1940 13840 1941 13880
rect 1899 13831 1941 13840
rect 4683 13880 4725 13889
rect 4683 13840 4684 13880
rect 4724 13840 4725 13880
rect 4683 13831 4725 13840
rect 30699 13880 30741 13889
rect 30699 13840 30700 13880
rect 30740 13840 30741 13880
rect 30699 13831 30741 13840
rect 32899 13880 32957 13881
rect 32899 13840 32908 13880
rect 32948 13840 32957 13880
rect 32899 13839 32957 13840
rect 43851 13880 43893 13889
rect 43851 13840 43852 13880
rect 43892 13840 43893 13880
rect 43851 13831 43893 13840
rect 51627 13880 51669 13889
rect 51627 13840 51628 13880
rect 51668 13840 51669 13880
rect 51627 13831 51669 13840
rect 74763 13880 74805 13889
rect 74763 13840 74764 13880
rect 74804 13840 74805 13880
rect 74763 13831 74805 13840
rect 3907 13796 3965 13797
rect 3907 13756 3916 13796
rect 3956 13756 3965 13796
rect 3907 13755 3965 13756
rect 35491 13796 35549 13797
rect 35491 13756 35500 13796
rect 35540 13756 35549 13796
rect 35491 13755 35549 13756
rect 42883 13796 42941 13797
rect 42883 13756 42892 13796
rect 42932 13756 42941 13796
rect 42883 13755 42941 13756
rect 51435 13796 51477 13805
rect 51435 13756 51436 13796
rect 51476 13756 51477 13796
rect 51435 13747 51477 13756
rect 53547 13796 53589 13805
rect 53547 13756 53548 13796
rect 53588 13756 53589 13796
rect 53547 13747 53589 13756
rect 56131 13796 56189 13797
rect 56131 13756 56140 13796
rect 56180 13756 56189 13796
rect 56131 13755 56189 13756
rect 56523 13796 56565 13805
rect 56523 13756 56524 13796
rect 56564 13756 56565 13796
rect 56523 13747 56565 13756
rect 57867 13796 57909 13805
rect 57867 13756 57868 13796
rect 57908 13756 57909 13796
rect 57867 13747 57909 13756
rect 61035 13796 61077 13805
rect 61035 13756 61036 13796
rect 61076 13756 61077 13796
rect 61035 13747 61077 13756
rect 64107 13796 64149 13805
rect 64107 13756 64108 13796
rect 64148 13756 64149 13796
rect 64107 13747 64149 13756
rect 68331 13796 68373 13805
rect 68331 13756 68332 13796
rect 68372 13756 68373 13796
rect 68331 13747 68373 13756
rect 70339 13796 70397 13797
rect 70339 13756 70348 13796
rect 70388 13756 70397 13796
rect 70339 13755 70397 13756
rect 70731 13796 70773 13805
rect 70731 13756 70732 13796
rect 70772 13756 70773 13796
rect 70731 13747 70773 13756
rect 71115 13796 71157 13805
rect 71115 13756 71116 13796
rect 71156 13756 71157 13796
rect 71115 13747 71157 13756
rect 74563 13796 74621 13797
rect 74563 13756 74572 13796
rect 74612 13756 74621 13796
rect 74563 13755 74621 13756
rect 576 13628 79584 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79584 13628
rect 576 13564 79584 13588
rect 3811 13460 3869 13461
rect 3811 13420 3820 13460
rect 3860 13420 3869 13460
rect 3811 13419 3869 13420
rect 4299 13460 4341 13469
rect 4299 13420 4300 13460
rect 4340 13420 4341 13460
rect 4299 13411 4341 13420
rect 32811 13460 32853 13469
rect 32811 13420 32812 13460
rect 32852 13420 32853 13460
rect 32811 13411 32853 13420
rect 42795 13460 42837 13469
rect 42795 13420 42796 13460
rect 42836 13420 42837 13460
rect 42795 13411 42837 13420
rect 45475 13460 45533 13461
rect 45475 13420 45484 13460
rect 45524 13420 45533 13460
rect 45475 13419 45533 13420
rect 46155 13460 46197 13469
rect 46155 13420 46156 13460
rect 46196 13420 46197 13460
rect 46155 13411 46197 13420
rect 47211 13460 47253 13469
rect 47211 13420 47212 13460
rect 47252 13420 47253 13460
rect 47211 13411 47253 13420
rect 51619 13460 51677 13461
rect 51619 13420 51628 13460
rect 51668 13420 51677 13460
rect 51619 13419 51677 13420
rect 58923 13460 58965 13469
rect 58923 13420 58924 13460
rect 58964 13420 58965 13460
rect 58923 13411 58965 13420
rect 61131 13460 61173 13469
rect 61131 13420 61132 13460
rect 61172 13420 61173 13460
rect 61131 13411 61173 13420
rect 61899 13460 61941 13469
rect 61899 13420 61900 13460
rect 61940 13420 61941 13460
rect 64491 13460 64533 13469
rect 61899 13411 61941 13420
rect 62187 13418 62229 13427
rect 1035 13376 1077 13385
rect 1035 13336 1036 13376
rect 1076 13336 1077 13376
rect 1035 13327 1077 13336
rect 5547 13376 5589 13385
rect 5547 13336 5548 13376
rect 5588 13336 5589 13376
rect 5547 13327 5589 13336
rect 33579 13376 33621 13385
rect 33579 13336 33580 13376
rect 33620 13336 33621 13376
rect 33579 13327 33621 13336
rect 39331 13376 39389 13377
rect 39331 13336 39340 13376
rect 39380 13336 39389 13376
rect 39331 13335 39389 13336
rect 40779 13376 40821 13385
rect 40779 13336 40780 13376
rect 40820 13336 40821 13376
rect 40779 13327 40821 13336
rect 47403 13376 47445 13385
rect 47403 13336 47404 13376
rect 47444 13336 47445 13376
rect 47403 13327 47445 13336
rect 52491 13376 52533 13385
rect 52491 13336 52492 13376
rect 52532 13336 52533 13376
rect 52491 13327 52533 13336
rect 56331 13376 56373 13385
rect 62187 13378 62188 13418
rect 62228 13378 62229 13418
rect 64491 13420 64492 13460
rect 64532 13420 64533 13460
rect 64491 13411 64533 13420
rect 70155 13460 70197 13469
rect 70155 13420 70156 13460
rect 70196 13420 70197 13460
rect 70155 13411 70197 13420
rect 76491 13460 76533 13469
rect 76491 13420 76492 13460
rect 76532 13420 76533 13460
rect 76491 13411 76533 13420
rect 56331 13336 56332 13376
rect 56372 13336 56373 13376
rect 56331 13327 56373 13336
rect 58435 13376 58493 13377
rect 58435 13336 58444 13376
rect 58484 13336 58493 13376
rect 62187 13369 62229 13378
rect 65163 13376 65205 13385
rect 58435 13335 58493 13336
rect 65163 13336 65164 13376
rect 65204 13336 65205 13376
rect 65163 13327 65205 13336
rect 70923 13376 70965 13385
rect 70923 13336 70924 13376
rect 70964 13336 70965 13376
rect 70923 13327 70965 13336
rect 72075 13376 72117 13385
rect 72075 13336 72076 13376
rect 72116 13336 72117 13376
rect 72075 13327 72117 13336
rect 76099 13376 76157 13377
rect 76099 13336 76108 13376
rect 76148 13336 76157 13376
rect 76099 13335 76157 13336
rect 77067 13376 77109 13385
rect 77067 13336 77068 13376
rect 77108 13336 77109 13376
rect 77067 13327 77109 13336
rect 77451 13376 77493 13385
rect 77451 13336 77452 13376
rect 77492 13336 77493 13376
rect 77451 13327 77493 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1219 13292 1277 13293
rect 1219 13252 1228 13292
rect 1268 13252 1277 13292
rect 74667 13292 74709 13301
rect 1219 13251 1277 13252
rect 61515 13245 61557 13254
rect 33117 13219 33159 13228
rect 1795 13208 1853 13209
rect 1795 13168 1804 13208
rect 1844 13168 1853 13208
rect 1795 13167 1853 13168
rect 2659 13208 2717 13209
rect 2659 13168 2668 13208
rect 2708 13168 2717 13208
rect 2659 13167 2717 13168
rect 4203 13208 4245 13217
rect 4203 13168 4204 13208
rect 4244 13168 4245 13208
rect 4203 13159 4245 13168
rect 4387 13208 4445 13209
rect 4387 13168 4396 13208
rect 4436 13168 4445 13208
rect 4387 13167 4445 13168
rect 4971 13208 5013 13217
rect 4971 13168 4972 13208
rect 5012 13168 5013 13208
rect 4971 13159 5013 13168
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 33003 13208 33045 13217
rect 33003 13168 33004 13208
rect 33044 13168 33045 13208
rect 33117 13179 33118 13219
rect 33158 13179 33159 13219
rect 33117 13170 33159 13179
rect 34915 13208 34973 13209
rect 33003 13159 33045 13168
rect 34915 13168 34924 13208
rect 34964 13168 34973 13208
rect 34915 13167 34973 13168
rect 35019 13208 35061 13217
rect 35019 13168 35020 13208
rect 35060 13168 35061 13208
rect 35019 13159 35061 13168
rect 35211 13208 35253 13217
rect 35211 13168 35212 13208
rect 35252 13168 35253 13208
rect 35211 13159 35253 13168
rect 36547 13208 36605 13209
rect 36547 13168 36556 13208
rect 36596 13168 36605 13208
rect 36547 13167 36605 13168
rect 36747 13208 36789 13217
rect 36747 13168 36748 13208
rect 36788 13168 36789 13208
rect 36747 13159 36789 13168
rect 37315 13208 37373 13209
rect 37315 13168 37324 13208
rect 37364 13168 37373 13208
rect 37315 13167 37373 13168
rect 38179 13208 38237 13209
rect 38179 13168 38188 13208
rect 38228 13168 38237 13208
rect 38179 13167 38237 13168
rect 41451 13208 41493 13217
rect 41451 13168 41452 13208
rect 41492 13168 41493 13208
rect 41451 13159 41493 13168
rect 41643 13208 41685 13217
rect 41643 13168 41644 13208
rect 41684 13168 41685 13208
rect 41643 13159 41685 13168
rect 41731 13208 41789 13209
rect 41731 13168 41740 13208
rect 41780 13168 41789 13208
rect 41731 13167 41789 13168
rect 42691 13208 42749 13209
rect 42691 13168 42700 13208
rect 42740 13168 42749 13208
rect 42691 13167 42749 13168
rect 42891 13208 42933 13217
rect 42891 13168 42892 13208
rect 42932 13168 42933 13208
rect 42891 13159 42933 13168
rect 43083 13208 43125 13217
rect 43083 13168 43084 13208
rect 43124 13168 43125 13208
rect 43083 13159 43125 13168
rect 43459 13208 43517 13209
rect 43459 13168 43468 13208
rect 43508 13168 43517 13208
rect 43459 13167 43517 13168
rect 44323 13208 44381 13209
rect 44323 13168 44332 13208
rect 44372 13168 44381 13208
rect 44323 13167 44381 13168
rect 45675 13208 45717 13217
rect 45675 13168 45676 13208
rect 45716 13168 45717 13208
rect 45675 13159 45717 13168
rect 45771 13208 45813 13217
rect 45771 13168 45772 13208
rect 45812 13168 45813 13208
rect 45771 13159 45813 13168
rect 45867 13208 45909 13217
rect 45867 13168 45868 13208
rect 45908 13168 45909 13208
rect 45867 13159 45909 13168
rect 45963 13208 46005 13217
rect 45963 13168 45964 13208
rect 46004 13168 46005 13208
rect 45963 13159 46005 13168
rect 46155 13208 46197 13217
rect 46155 13168 46156 13208
rect 46196 13168 46197 13208
rect 46155 13159 46197 13168
rect 46347 13208 46389 13217
rect 46347 13168 46348 13208
rect 46388 13168 46389 13208
rect 46347 13159 46389 13168
rect 46435 13208 46493 13209
rect 46435 13168 46444 13208
rect 46484 13168 46493 13208
rect 46435 13167 46493 13168
rect 46827 13208 46869 13217
rect 46827 13168 46828 13208
rect 46868 13168 46869 13208
rect 46827 13159 46869 13168
rect 47883 13208 47925 13217
rect 47883 13168 47884 13208
rect 47924 13168 47925 13208
rect 47883 13159 47925 13168
rect 48075 13208 48117 13217
rect 48075 13168 48076 13208
rect 48116 13168 48117 13208
rect 48075 13159 48117 13168
rect 48163 13208 48221 13209
rect 48163 13168 48172 13208
rect 48212 13168 48221 13208
rect 48163 13167 48221 13168
rect 48547 13208 48605 13209
rect 48547 13168 48556 13208
rect 48596 13168 48605 13208
rect 48547 13167 48605 13168
rect 48747 13208 48789 13217
rect 48747 13168 48748 13208
rect 48788 13168 48789 13208
rect 48747 13159 48789 13168
rect 49603 13208 49661 13209
rect 49603 13168 49612 13208
rect 49652 13168 49661 13208
rect 49603 13167 49661 13168
rect 50467 13208 50525 13209
rect 50467 13168 50476 13208
rect 50516 13168 50525 13208
rect 50467 13167 50525 13168
rect 51915 13208 51957 13217
rect 51915 13168 51916 13208
rect 51956 13168 51957 13208
rect 51915 13159 51957 13168
rect 52099 13208 52157 13209
rect 52099 13168 52108 13208
rect 52148 13168 52157 13208
rect 52099 13167 52157 13168
rect 54403 13208 54461 13209
rect 54403 13168 54412 13208
rect 54452 13168 54461 13208
rect 54403 13167 54461 13168
rect 54507 13208 54549 13217
rect 54507 13168 54508 13208
rect 54548 13168 54549 13208
rect 54507 13159 54549 13168
rect 54699 13208 54741 13217
rect 54699 13168 54700 13208
rect 54740 13168 54741 13208
rect 54699 13159 54741 13168
rect 55083 13208 55125 13217
rect 55083 13168 55084 13208
rect 55124 13168 55125 13208
rect 55083 13159 55125 13168
rect 55179 13208 55221 13217
rect 55179 13168 55180 13208
rect 55220 13168 55221 13208
rect 55179 13159 55221 13168
rect 55275 13208 55317 13217
rect 55275 13168 55276 13208
rect 55316 13168 55317 13208
rect 55275 13159 55317 13168
rect 55371 13208 55413 13217
rect 55371 13168 55372 13208
rect 55412 13168 55413 13208
rect 55371 13159 55413 13168
rect 56035 13208 56093 13209
rect 56035 13168 56044 13208
rect 56084 13168 56093 13208
rect 56035 13167 56093 13168
rect 56139 13208 56181 13217
rect 56139 13168 56140 13208
rect 56180 13168 56181 13208
rect 56139 13159 56181 13168
rect 56331 13208 56373 13217
rect 56331 13168 56332 13208
rect 56372 13168 56373 13208
rect 56331 13159 56373 13168
rect 56523 13208 56565 13217
rect 56523 13168 56524 13208
rect 56564 13168 56565 13208
rect 56803 13208 56861 13209
rect 56523 13159 56565 13168
rect 56715 13194 56757 13203
rect 56715 13154 56716 13194
rect 56756 13154 56757 13194
rect 56803 13168 56812 13208
rect 56852 13168 56861 13208
rect 56803 13167 56861 13168
rect 57763 13208 57821 13209
rect 57763 13168 57772 13208
rect 57812 13168 57821 13208
rect 57763 13167 57821 13168
rect 58059 13208 58101 13217
rect 58059 13168 58060 13208
rect 58100 13168 58101 13208
rect 58059 13159 58101 13168
rect 58627 13208 58685 13209
rect 58627 13168 58636 13208
rect 58676 13168 58685 13208
rect 58627 13167 58685 13168
rect 58731 13208 58773 13217
rect 58731 13168 58732 13208
rect 58772 13168 58773 13208
rect 58731 13159 58773 13168
rect 58923 13208 58965 13217
rect 58923 13168 58924 13208
rect 58964 13168 58965 13208
rect 58923 13159 58965 13168
rect 60835 13208 60893 13209
rect 60835 13168 60844 13208
rect 60884 13168 60893 13208
rect 60835 13167 60893 13168
rect 60939 13208 60981 13217
rect 60939 13168 60940 13208
rect 60980 13168 60981 13208
rect 60939 13159 60981 13168
rect 61131 13208 61173 13217
rect 61131 13168 61132 13208
rect 61172 13168 61173 13208
rect 61131 13159 61173 13168
rect 61323 13208 61365 13217
rect 61323 13168 61324 13208
rect 61364 13168 61365 13208
rect 61323 13159 61365 13168
rect 61419 13208 61461 13217
rect 61419 13168 61420 13208
rect 61460 13168 61461 13208
rect 61515 13205 61516 13245
rect 61556 13205 61557 13245
rect 74667 13252 74668 13292
rect 74708 13252 74709 13292
rect 74667 13243 74709 13252
rect 61515 13196 61557 13205
rect 61611 13208 61653 13217
rect 61419 13159 61461 13168
rect 61611 13168 61612 13208
rect 61652 13168 61653 13208
rect 61611 13159 61653 13168
rect 61803 13208 61845 13217
rect 61803 13168 61804 13208
rect 61844 13168 61845 13208
rect 61803 13159 61845 13168
rect 61987 13208 62045 13209
rect 61987 13168 61996 13208
rect 62036 13168 62045 13208
rect 61987 13167 62045 13168
rect 64195 13208 64253 13209
rect 64195 13168 64204 13208
rect 64244 13168 64253 13208
rect 64195 13167 64253 13168
rect 64299 13208 64341 13217
rect 64299 13168 64300 13208
rect 64340 13168 64341 13208
rect 64299 13159 64341 13168
rect 64491 13208 64533 13217
rect 64491 13168 64492 13208
rect 64532 13168 64533 13208
rect 64491 13159 64533 13168
rect 64683 13208 64725 13217
rect 64683 13168 64684 13208
rect 64724 13168 64725 13208
rect 64683 13159 64725 13168
rect 64779 13208 64821 13217
rect 64779 13168 64780 13208
rect 64820 13168 64821 13208
rect 64779 13159 64821 13168
rect 64875 13208 64917 13217
rect 64875 13168 64876 13208
rect 64916 13168 64917 13208
rect 64875 13159 64917 13168
rect 64971 13208 65013 13217
rect 64971 13168 64972 13208
rect 65012 13168 65013 13208
rect 64971 13159 65013 13168
rect 68619 13208 68661 13217
rect 68619 13168 68620 13208
rect 68660 13168 68661 13208
rect 68619 13159 68661 13168
rect 68715 13208 68757 13217
rect 68715 13168 68716 13208
rect 68756 13168 68757 13208
rect 68715 13159 68757 13168
rect 68811 13208 68853 13217
rect 68811 13168 68812 13208
rect 68852 13168 68853 13208
rect 68811 13159 68853 13168
rect 68995 13208 69053 13209
rect 68995 13168 69004 13208
rect 69044 13168 69053 13208
rect 68995 13167 69053 13168
rect 69099 13208 69141 13217
rect 69099 13168 69100 13208
rect 69140 13168 69141 13208
rect 69099 13159 69141 13168
rect 69291 13208 69333 13217
rect 69291 13168 69292 13208
rect 69332 13168 69333 13208
rect 69291 13159 69333 13168
rect 69667 13208 69725 13209
rect 69667 13168 69676 13208
rect 69716 13168 69725 13208
rect 69667 13167 69725 13168
rect 69867 13208 69909 13217
rect 69867 13168 69868 13208
rect 69908 13168 69909 13208
rect 69867 13159 69909 13168
rect 70051 13208 70109 13209
rect 70051 13168 70060 13208
rect 70100 13168 70109 13208
rect 70051 13167 70109 13168
rect 70251 13208 70293 13217
rect 70251 13168 70252 13208
rect 70292 13168 70293 13208
rect 70251 13159 70293 13168
rect 72643 13208 72701 13209
rect 72643 13168 72652 13208
rect 72692 13168 72701 13208
rect 72643 13167 72701 13168
rect 73507 13208 73565 13209
rect 73507 13168 73516 13208
rect 73556 13168 73565 13208
rect 73507 13167 73565 13168
rect 74955 13208 74997 13217
rect 74955 13168 74956 13208
rect 74996 13168 74997 13208
rect 74955 13159 74997 13168
rect 75051 13208 75093 13217
rect 75051 13168 75052 13208
rect 75092 13168 75093 13208
rect 75051 13159 75093 13168
rect 75147 13208 75189 13217
rect 75147 13168 75148 13208
rect 75188 13168 75189 13208
rect 75147 13159 75189 13168
rect 75427 13208 75485 13209
rect 75427 13168 75436 13208
rect 75476 13168 75485 13208
rect 75427 13167 75485 13168
rect 75723 13208 75765 13217
rect 75723 13168 75724 13208
rect 75764 13168 75765 13208
rect 75723 13159 75765 13168
rect 75819 13208 75861 13217
rect 75819 13168 75820 13208
rect 75860 13168 75861 13208
rect 75819 13159 75861 13168
rect 76491 13208 76533 13217
rect 76491 13168 76492 13208
rect 76532 13168 76533 13208
rect 76491 13159 76533 13168
rect 76683 13208 76725 13217
rect 76683 13168 76684 13208
rect 76724 13168 76725 13208
rect 76683 13159 76725 13168
rect 76771 13208 76829 13209
rect 76771 13168 76780 13208
rect 76820 13168 76829 13208
rect 76771 13167 76829 13168
rect 76963 13208 77021 13209
rect 76963 13168 76972 13208
rect 77012 13168 77021 13208
rect 76963 13167 77021 13168
rect 77163 13208 77205 13217
rect 77163 13168 77164 13208
rect 77204 13168 77205 13208
rect 77163 13159 77205 13168
rect 56715 13145 56757 13154
rect 1419 13124 1461 13133
rect 1419 13084 1420 13124
rect 1460 13084 1461 13124
rect 1419 13075 1461 13084
rect 36651 13124 36693 13133
rect 36651 13084 36652 13124
rect 36692 13084 36693 13124
rect 36651 13075 36693 13084
rect 36939 13124 36981 13133
rect 36939 13084 36940 13124
rect 36980 13084 36981 13124
rect 36939 13075 36981 13084
rect 41547 13124 41589 13133
rect 41547 13084 41548 13124
rect 41588 13084 41589 13124
rect 41547 13075 41589 13084
rect 47979 13124 48021 13133
rect 47979 13084 47980 13124
rect 48020 13084 48021 13124
rect 47979 13075 48021 13084
rect 48651 13124 48693 13133
rect 48651 13084 48652 13124
rect 48692 13084 48693 13124
rect 48651 13075 48693 13084
rect 49227 13124 49269 13133
rect 49227 13084 49228 13124
rect 49268 13084 49269 13124
rect 49227 13075 49269 13084
rect 52011 13124 52053 13133
rect 52011 13084 52012 13124
rect 52052 13084 52053 13124
rect 52011 13075 52053 13084
rect 54603 13124 54645 13133
rect 54603 13084 54604 13124
rect 54644 13084 54645 13124
rect 54603 13075 54645 13084
rect 58155 13124 58197 13133
rect 58155 13084 58156 13124
rect 58196 13084 58197 13124
rect 58155 13075 58197 13084
rect 69771 13124 69813 13133
rect 69771 13084 69772 13124
rect 69812 13084 69813 13124
rect 69771 13075 69813 13084
rect 72267 13124 72309 13133
rect 72267 13084 72268 13124
rect 72308 13084 72309 13124
rect 72267 13075 72309 13084
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 35107 13040 35165 13041
rect 35107 13000 35116 13040
rect 35156 13000 35165 13040
rect 35107 12999 35165 13000
rect 51619 13040 51677 13041
rect 51619 13000 51628 13040
rect 51668 13000 51677 13040
rect 51619 12999 51677 13000
rect 56611 13040 56669 13041
rect 56611 13000 56620 13040
rect 56660 13000 56669 13040
rect 56611 12999 56669 13000
rect 68515 13040 68573 13041
rect 68515 13000 68524 13040
rect 68564 13000 68573 13040
rect 68515 12999 68573 13000
rect 69187 13040 69245 13041
rect 69187 13000 69196 13040
rect 69236 13000 69245 13040
rect 69187 12999 69245 13000
rect 74851 13040 74909 13041
rect 74851 13000 74860 13040
rect 74900 13000 74909 13040
rect 74851 12999 74909 13000
rect 576 12872 79584 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79584 12872
rect 576 12808 79584 12832
rect 2371 12704 2429 12705
rect 2371 12664 2380 12704
rect 2420 12664 2429 12704
rect 2371 12663 2429 12664
rect 47683 12704 47741 12705
rect 47683 12664 47692 12704
rect 47732 12664 47741 12704
rect 47683 12663 47741 12664
rect 48931 12704 48989 12705
rect 48931 12664 48940 12704
rect 48980 12664 48989 12704
rect 48931 12663 48989 12664
rect 54403 12704 54461 12705
rect 54403 12664 54412 12704
rect 54452 12664 54461 12704
rect 54403 12663 54461 12664
rect 57187 12704 57245 12705
rect 57187 12664 57196 12704
rect 57236 12664 57245 12704
rect 57187 12663 57245 12664
rect 57963 12704 58005 12713
rect 57963 12664 57964 12704
rect 58004 12664 58005 12704
rect 57963 12655 58005 12664
rect 62083 12704 62141 12705
rect 62083 12664 62092 12704
rect 62132 12664 62141 12704
rect 62083 12663 62141 12664
rect 67171 12704 67229 12705
rect 67171 12664 67180 12704
rect 67220 12664 67229 12704
rect 67171 12663 67229 12664
rect 72835 12704 72893 12705
rect 72835 12664 72844 12704
rect 72884 12664 72893 12704
rect 72835 12663 72893 12664
rect 74371 12704 74429 12705
rect 74371 12664 74380 12704
rect 74420 12664 74429 12704
rect 74371 12663 74429 12664
rect 4107 12620 4149 12629
rect 4107 12580 4108 12620
rect 4148 12580 4149 12620
rect 4107 12571 4149 12580
rect 48363 12620 48405 12629
rect 48363 12580 48364 12620
rect 48404 12580 48405 12620
rect 48363 12571 48405 12580
rect 54795 12620 54837 12629
rect 54795 12580 54796 12620
rect 54836 12580 54837 12620
rect 76107 12620 76149 12629
rect 54795 12571 54837 12580
rect 70251 12578 70293 12587
rect 59508 12549 59550 12558
rect 2283 12536 2325 12545
rect 2283 12496 2284 12536
rect 2324 12496 2325 12536
rect 2283 12487 2325 12496
rect 2475 12536 2517 12545
rect 2475 12496 2476 12536
rect 2516 12496 2517 12536
rect 2475 12487 2517 12496
rect 2563 12536 2621 12537
rect 2563 12496 2572 12536
rect 2612 12496 2621 12536
rect 2563 12495 2621 12496
rect 2763 12536 2805 12545
rect 2763 12496 2764 12536
rect 2804 12496 2805 12536
rect 2763 12487 2805 12496
rect 2955 12536 2997 12545
rect 2955 12496 2956 12536
rect 2996 12496 2997 12536
rect 2955 12487 2997 12496
rect 3043 12536 3101 12537
rect 3043 12496 3052 12536
rect 3092 12496 3101 12536
rect 3043 12495 3101 12496
rect 4011 12536 4053 12545
rect 4011 12496 4012 12536
rect 4052 12496 4053 12536
rect 4011 12487 4053 12496
rect 4195 12536 4253 12537
rect 4195 12496 4204 12536
rect 4244 12496 4253 12536
rect 4195 12495 4253 12496
rect 4779 12536 4821 12545
rect 4779 12496 4780 12536
rect 4820 12496 4821 12536
rect 4779 12487 4821 12496
rect 5635 12536 5693 12537
rect 5635 12496 5644 12536
rect 5684 12496 5693 12536
rect 5635 12495 5693 12496
rect 29931 12536 29973 12545
rect 29931 12496 29932 12536
rect 29972 12496 29973 12536
rect 29931 12487 29973 12496
rect 31363 12536 31421 12537
rect 31363 12496 31372 12536
rect 31412 12496 31421 12536
rect 31363 12495 31421 12496
rect 33867 12536 33909 12545
rect 33867 12496 33868 12536
rect 33908 12496 33909 12536
rect 33867 12487 33909 12496
rect 34243 12536 34301 12537
rect 34243 12496 34252 12536
rect 34292 12496 34301 12536
rect 34243 12495 34301 12496
rect 35107 12536 35165 12537
rect 35107 12496 35116 12536
rect 35156 12496 35165 12536
rect 35107 12495 35165 12496
rect 36747 12536 36789 12545
rect 36747 12496 36748 12536
rect 36788 12496 36789 12536
rect 36747 12487 36789 12496
rect 36843 12536 36885 12545
rect 36843 12496 36844 12536
rect 36884 12496 36885 12536
rect 36843 12487 36885 12496
rect 37123 12536 37181 12537
rect 37123 12496 37132 12536
rect 37172 12496 37181 12536
rect 37123 12495 37181 12496
rect 39147 12536 39189 12545
rect 39147 12496 39148 12536
rect 39188 12496 39189 12536
rect 39147 12487 39189 12496
rect 39523 12536 39581 12537
rect 39523 12496 39532 12536
rect 39572 12496 39581 12536
rect 39523 12495 39581 12496
rect 40387 12536 40445 12537
rect 40387 12496 40396 12536
rect 40436 12496 40445 12536
rect 40387 12495 40445 12496
rect 41923 12536 41981 12537
rect 41923 12496 41932 12536
rect 41972 12496 41981 12536
rect 41923 12495 41981 12496
rect 42027 12536 42069 12545
rect 42027 12496 42028 12536
rect 42068 12496 42069 12536
rect 42027 12487 42069 12496
rect 42219 12536 42261 12545
rect 42219 12496 42220 12536
rect 42260 12496 42261 12536
rect 42219 12487 42261 12496
rect 42403 12536 42461 12537
rect 42403 12496 42412 12536
rect 42452 12496 42461 12536
rect 42403 12495 42461 12496
rect 42507 12536 42549 12545
rect 42507 12496 42508 12536
rect 42548 12496 42549 12536
rect 42507 12487 42549 12496
rect 42603 12536 42645 12545
rect 42603 12496 42604 12536
rect 42644 12496 42645 12536
rect 42603 12487 42645 12496
rect 45291 12536 45333 12545
rect 45291 12496 45292 12536
rect 45332 12496 45333 12536
rect 45291 12487 45333 12496
rect 45667 12536 45725 12537
rect 45667 12496 45676 12536
rect 45716 12496 45725 12536
rect 45667 12495 45725 12496
rect 46531 12536 46589 12537
rect 46531 12496 46540 12536
rect 46580 12496 46589 12536
rect 46531 12495 46589 12496
rect 47971 12536 48029 12537
rect 47971 12496 47980 12536
rect 48020 12496 48029 12536
rect 47971 12495 48029 12496
rect 48267 12536 48309 12545
rect 48267 12496 48268 12536
rect 48308 12496 48309 12536
rect 48267 12487 48309 12496
rect 48843 12536 48885 12545
rect 48843 12496 48844 12536
rect 48884 12496 48885 12536
rect 48843 12487 48885 12496
rect 49035 12536 49077 12545
rect 49035 12496 49036 12536
rect 49076 12496 49077 12536
rect 49035 12487 49077 12496
rect 49123 12536 49181 12537
rect 49123 12496 49132 12536
rect 49172 12496 49181 12536
rect 49123 12495 49181 12496
rect 49315 12536 49373 12537
rect 49315 12496 49324 12536
rect 49364 12496 49373 12536
rect 49315 12495 49373 12496
rect 49515 12536 49557 12545
rect 49515 12496 49516 12536
rect 49556 12496 49557 12536
rect 49515 12487 49557 12496
rect 52011 12536 52053 12545
rect 52011 12496 52012 12536
rect 52052 12496 52053 12536
rect 52011 12487 52053 12496
rect 52387 12536 52445 12537
rect 52387 12496 52396 12536
rect 52436 12496 52445 12536
rect 52387 12495 52445 12496
rect 53292 12536 53334 12545
rect 53292 12496 53293 12536
rect 53333 12496 53334 12536
rect 53292 12487 53334 12496
rect 55171 12536 55229 12537
rect 55171 12496 55180 12536
rect 55220 12496 55229 12536
rect 55171 12495 55229 12496
rect 56035 12536 56093 12537
rect 56035 12496 56044 12536
rect 56084 12496 56093 12536
rect 56035 12495 56093 12496
rect 58147 12536 58205 12537
rect 58147 12496 58156 12536
rect 58196 12496 58205 12536
rect 58147 12495 58205 12496
rect 58347 12536 58389 12545
rect 58347 12496 58348 12536
rect 58388 12496 58389 12536
rect 58347 12487 58389 12496
rect 59299 12536 59357 12537
rect 59299 12496 59308 12536
rect 59348 12496 59357 12536
rect 59508 12509 59509 12549
rect 59549 12509 59550 12549
rect 59508 12500 59550 12509
rect 61995 12536 62037 12545
rect 59299 12495 59357 12496
rect 61995 12496 61996 12536
rect 62036 12496 62037 12536
rect 61995 12487 62037 12496
rect 62187 12536 62229 12545
rect 62187 12496 62188 12536
rect 62228 12496 62229 12536
rect 62187 12487 62229 12496
rect 62275 12536 62333 12537
rect 62275 12496 62284 12536
rect 62324 12496 62333 12536
rect 62275 12495 62333 12496
rect 63295 12536 63337 12545
rect 63295 12496 63296 12536
rect 63336 12496 63337 12536
rect 63295 12487 63337 12496
rect 63627 12536 63669 12545
rect 63627 12496 63628 12536
rect 63668 12496 63669 12536
rect 63627 12487 63669 12496
rect 63723 12536 63765 12545
rect 63723 12496 63724 12536
rect 63764 12496 63765 12536
rect 63723 12487 63765 12496
rect 64395 12536 64437 12545
rect 64395 12496 64396 12536
rect 64436 12496 64437 12536
rect 64395 12487 64437 12496
rect 64579 12536 64637 12537
rect 64579 12496 64588 12536
rect 64628 12496 64637 12536
rect 64579 12495 64637 12496
rect 64779 12536 64821 12545
rect 64779 12496 64780 12536
rect 64820 12496 64821 12536
rect 64779 12487 64821 12496
rect 65155 12536 65213 12537
rect 65155 12496 65164 12536
rect 65204 12496 65213 12536
rect 65155 12495 65213 12496
rect 66019 12536 66077 12537
rect 66019 12496 66028 12536
rect 66068 12496 66077 12536
rect 66019 12495 66077 12496
rect 67371 12536 67413 12545
rect 67371 12496 67372 12536
rect 67412 12496 67413 12536
rect 67371 12487 67413 12496
rect 67747 12536 67805 12537
rect 67747 12496 67756 12536
rect 67796 12496 67805 12536
rect 67747 12495 67805 12496
rect 68611 12536 68669 12537
rect 68611 12496 68620 12536
rect 68660 12496 68669 12536
rect 68611 12495 68669 12496
rect 69955 12536 70013 12537
rect 69955 12496 69964 12536
rect 70004 12496 70013 12536
rect 69955 12495 70013 12496
rect 70059 12536 70101 12545
rect 70059 12496 70060 12536
rect 70100 12496 70101 12536
rect 70251 12538 70252 12578
rect 70292 12538 70293 12578
rect 76107 12580 76108 12620
rect 76148 12580 76149 12620
rect 76107 12571 76149 12580
rect 70251 12529 70293 12538
rect 70443 12536 70485 12545
rect 70059 12487 70101 12496
rect 70443 12496 70444 12536
rect 70484 12496 70485 12536
rect 70443 12487 70485 12496
rect 70819 12536 70877 12537
rect 70819 12496 70828 12536
rect 70868 12496 70877 12536
rect 70819 12495 70877 12496
rect 71683 12536 71741 12537
rect 71683 12496 71692 12536
rect 71732 12496 71741 12536
rect 71683 12495 71741 12496
rect 74283 12536 74325 12545
rect 74283 12496 74284 12536
rect 74324 12496 74325 12536
rect 74283 12487 74325 12496
rect 74475 12536 74517 12545
rect 74475 12496 74476 12536
rect 74516 12496 74517 12536
rect 74475 12487 74517 12496
rect 74563 12536 74621 12537
rect 74563 12496 74572 12536
rect 74612 12496 74621 12536
rect 74563 12495 74621 12496
rect 74763 12536 74805 12545
rect 74763 12496 74764 12536
rect 74804 12496 74805 12536
rect 74763 12487 74805 12496
rect 74955 12536 74997 12545
rect 74955 12496 74956 12536
rect 74996 12496 74997 12536
rect 74955 12487 74997 12496
rect 75043 12536 75101 12537
rect 75043 12496 75052 12536
rect 75092 12496 75101 12536
rect 75043 12495 75101 12496
rect 76003 12536 76061 12537
rect 76003 12496 76012 12536
rect 76052 12496 76061 12536
rect 76003 12495 76061 12496
rect 76203 12536 76245 12545
rect 76203 12496 76204 12536
rect 76244 12496 76245 12536
rect 76203 12487 76245 12496
rect 76875 12536 76917 12545
rect 76875 12496 76876 12536
rect 76916 12496 76917 12536
rect 76875 12487 76917 12496
rect 77251 12536 77309 12537
rect 77251 12496 77260 12536
rect 77300 12496 77309 12536
rect 77251 12495 77309 12496
rect 78115 12536 78173 12537
rect 78115 12496 78124 12536
rect 78164 12496 78173 12536
rect 78115 12495 78173 12496
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1315 12452 1373 12453
rect 1315 12412 1324 12452
rect 1364 12412 1373 12452
rect 1315 12411 1373 12412
rect 1699 12452 1757 12453
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 1699 12411 1757 12412
rect 49419 12452 49461 12461
rect 49419 12412 49420 12452
rect 49460 12412 49461 12452
rect 49419 12403 49461 12412
rect 50275 12452 50333 12453
rect 50275 12412 50284 12452
rect 50324 12412 50333 12452
rect 50275 12411 50333 12412
rect 51139 12452 51197 12453
rect 51139 12412 51148 12452
rect 51188 12412 51197 12452
rect 51139 12411 51197 12412
rect 51619 12452 51677 12453
rect 51619 12412 51628 12452
rect 51668 12412 51677 12452
rect 51619 12411 51677 12412
rect 57763 12452 57821 12453
rect 57763 12412 57772 12452
rect 57812 12412 57821 12452
rect 57763 12411 57821 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 1131 12368 1173 12377
rect 1131 12328 1132 12368
rect 1172 12328 1173 12368
rect 1131 12319 1173 12328
rect 1899 12368 1941 12377
rect 1899 12328 1900 12368
rect 1940 12328 1941 12368
rect 1899 12319 1941 12328
rect 2763 12368 2805 12377
rect 2763 12328 2764 12368
rect 2804 12328 2805 12368
rect 2763 12319 2805 12328
rect 4971 12368 5013 12377
rect 4971 12328 4972 12368
rect 5012 12328 5013 12368
rect 4971 12319 5013 12328
rect 5835 12368 5877 12377
rect 5835 12328 5836 12368
rect 5876 12328 5877 12368
rect 5835 12319 5877 12328
rect 36259 12368 36317 12369
rect 36259 12328 36268 12368
rect 36308 12328 36317 12368
rect 36259 12327 36317 12328
rect 37419 12368 37461 12377
rect 37419 12328 37420 12368
rect 37460 12328 37461 12368
rect 37419 12319 37461 12328
rect 41539 12368 41597 12369
rect 41539 12328 41548 12368
rect 41588 12328 41597 12368
rect 41539 12327 41597 12328
rect 42891 12368 42933 12377
rect 42891 12328 42892 12368
rect 42932 12328 42933 12368
rect 42891 12319 42933 12328
rect 48643 12368 48701 12369
rect 48643 12328 48652 12368
rect 48692 12328 48701 12368
rect 48643 12327 48701 12328
rect 49707 12368 49749 12377
rect 49707 12328 49708 12368
rect 49748 12328 49749 12368
rect 49707 12319 49749 12328
rect 58251 12368 58293 12377
rect 58251 12328 58252 12368
rect 58292 12328 58293 12368
rect 58251 12319 58293 12328
rect 59787 12368 59829 12377
rect 59787 12328 59788 12368
rect 59828 12328 59829 12368
rect 59787 12319 59829 12328
rect 70251 12368 70293 12377
rect 70251 12328 70252 12368
rect 70292 12328 70293 12368
rect 70251 12319 70293 12328
rect 74763 12368 74805 12377
rect 74763 12328 74764 12368
rect 74804 12328 74805 12368
rect 74763 12319 74805 12328
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 36451 12284 36509 12285
rect 36451 12244 36460 12284
rect 36500 12244 36509 12284
rect 36451 12243 36509 12244
rect 42219 12284 42261 12293
rect 42219 12244 42220 12284
rect 42260 12244 42261 12284
rect 42219 12235 42261 12244
rect 47683 12284 47741 12285
rect 47683 12244 47692 12284
rect 47732 12244 47741 12284
rect 47683 12243 47741 12244
rect 50091 12284 50133 12293
rect 50091 12244 50092 12284
rect 50132 12244 50133 12284
rect 50091 12235 50133 12244
rect 50955 12284 50997 12293
rect 50955 12244 50956 12284
rect 50996 12244 50997 12284
rect 50955 12235 50997 12244
rect 51819 12284 51861 12293
rect 51819 12244 51820 12284
rect 51860 12244 51861 12284
rect 51819 12235 51861 12244
rect 57963 12284 58005 12293
rect 57963 12244 57964 12284
rect 58004 12244 58005 12284
rect 57963 12235 58005 12244
rect 59403 12284 59445 12293
rect 59403 12244 59404 12284
rect 59444 12244 59445 12284
rect 59403 12235 59445 12244
rect 64003 12284 64061 12285
rect 64003 12244 64012 12284
rect 64052 12244 64061 12284
rect 64003 12243 64061 12244
rect 64491 12284 64533 12293
rect 64491 12244 64492 12284
rect 64532 12244 64533 12284
rect 64491 12235 64533 12244
rect 69763 12284 69821 12285
rect 69763 12244 69772 12284
rect 69812 12244 69821 12284
rect 69763 12243 69821 12244
rect 79267 12284 79325 12285
rect 79267 12244 79276 12284
rect 79316 12244 79325 12284
rect 79267 12243 79325 12244
rect 576 12116 79584 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79584 12116
rect 576 12052 79584 12076
rect 7363 11948 7421 11949
rect 7363 11908 7372 11948
rect 7412 11908 7421 11948
rect 7363 11907 7421 11908
rect 34827 11948 34869 11957
rect 34827 11908 34828 11948
rect 34868 11908 34869 11948
rect 34827 11899 34869 11908
rect 36843 11948 36885 11957
rect 36843 11908 36844 11948
rect 36884 11908 36885 11948
rect 36843 11899 36885 11908
rect 38859 11948 38901 11957
rect 38859 11908 38860 11948
rect 38900 11908 38901 11948
rect 38859 11899 38901 11908
rect 44803 11948 44861 11949
rect 44803 11908 44812 11948
rect 44852 11908 44861 11948
rect 44803 11907 44861 11908
rect 48267 11948 48309 11957
rect 48267 11908 48268 11948
rect 48308 11908 48309 11948
rect 48267 11899 48309 11908
rect 51723 11948 51765 11957
rect 51723 11908 51724 11948
rect 51764 11908 51765 11948
rect 51723 11899 51765 11908
rect 61699 11948 61757 11949
rect 61699 11908 61708 11948
rect 61748 11908 61757 11948
rect 61699 11907 61757 11908
rect 64203 11948 64245 11957
rect 64203 11908 64204 11948
rect 64244 11908 64245 11948
rect 64203 11899 64245 11908
rect 68907 11948 68949 11957
rect 68907 11908 68908 11948
rect 68948 11908 68949 11948
rect 68907 11899 68949 11908
rect 70147 11948 70205 11949
rect 70147 11908 70156 11948
rect 70196 11908 70205 11948
rect 70147 11907 70205 11908
rect 70539 11948 70581 11957
rect 70539 11908 70540 11948
rect 70580 11908 70581 11948
rect 70539 11899 70581 11908
rect 74947 11948 75005 11949
rect 74947 11908 74956 11948
rect 74996 11908 75005 11948
rect 74947 11907 75005 11908
rect 76491 11948 76533 11957
rect 76491 11908 76492 11948
rect 76532 11908 76533 11948
rect 76491 11899 76533 11908
rect 34347 11864 34389 11873
rect 34347 11824 34348 11864
rect 34388 11824 34389 11864
rect 34347 11815 34389 11824
rect 36267 11864 36309 11873
rect 36267 11824 36268 11864
rect 36308 11824 36309 11864
rect 36267 11815 36309 11824
rect 37035 11864 37077 11873
rect 37035 11824 37036 11864
rect 37076 11824 37077 11864
rect 37035 11815 37077 11824
rect 39435 11864 39477 11873
rect 39435 11824 39436 11864
rect 39476 11824 39477 11864
rect 39435 11815 39477 11824
rect 39723 11864 39765 11873
rect 39723 11824 39724 11864
rect 39764 11824 39765 11864
rect 39723 11815 39765 11824
rect 42211 11864 42269 11865
rect 42211 11824 42220 11864
rect 42260 11824 42269 11864
rect 42211 11823 42269 11824
rect 45003 11864 45045 11873
rect 45003 11824 45004 11864
rect 45044 11824 45045 11864
rect 45003 11815 45045 11824
rect 45771 11864 45813 11873
rect 45771 11824 45772 11864
rect 45812 11824 45813 11864
rect 45771 11815 45813 11824
rect 48939 11864 48981 11873
rect 48939 11824 48940 11864
rect 48980 11824 48981 11864
rect 48939 11815 48981 11824
rect 49227 11864 49269 11873
rect 49227 11824 49228 11864
rect 49268 11824 49269 11864
rect 49227 11815 49269 11824
rect 51523 11864 51581 11865
rect 51523 11824 51532 11864
rect 51572 11824 51581 11864
rect 51523 11823 51581 11824
rect 55275 11864 55317 11873
rect 55275 11824 55276 11864
rect 55316 11824 55317 11864
rect 55275 11815 55317 11824
rect 56331 11864 56373 11873
rect 56331 11824 56332 11864
rect 56372 11824 56373 11864
rect 56331 11815 56373 11824
rect 57291 11864 57333 11873
rect 57291 11824 57292 11864
rect 57332 11824 57333 11864
rect 57291 11815 57333 11824
rect 62091 11864 62133 11873
rect 62091 11824 62092 11864
rect 62132 11824 62133 11864
rect 62091 11815 62133 11824
rect 65259 11864 65301 11873
rect 65259 11824 65260 11864
rect 65300 11824 65301 11864
rect 65259 11815 65301 11824
rect 67467 11864 67509 11873
rect 67467 11824 67468 11864
rect 67508 11824 67509 11864
rect 67467 11815 67509 11824
rect 76003 11864 76061 11865
rect 76003 11824 76012 11864
rect 76052 11824 76061 11864
rect 76003 11823 76061 11824
rect 77355 11864 77397 11873
rect 77355 11824 77356 11864
rect 77396 11824 77397 11864
rect 77355 11815 77397 11824
rect 1123 11780 1181 11781
rect 1123 11740 1132 11780
rect 1172 11740 1181 11780
rect 1123 11739 1181 11740
rect 57475 11780 57533 11781
rect 57475 11740 57484 11780
rect 57524 11740 57533 11780
rect 57475 11739 57533 11740
rect 1699 11696 1757 11697
rect 1699 11656 1708 11696
rect 1748 11656 1757 11696
rect 1699 11655 1757 11656
rect 2563 11696 2621 11697
rect 2563 11656 2572 11696
rect 2612 11656 2621 11696
rect 2563 11655 2621 11656
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 4099 11696 4157 11697
rect 4099 11656 4108 11696
rect 4148 11656 4157 11696
rect 4099 11655 4157 11656
rect 4491 11696 4533 11705
rect 4491 11656 4492 11696
rect 4532 11656 4533 11696
rect 4491 11647 4533 11656
rect 4683 11696 4725 11705
rect 4683 11656 4684 11696
rect 4724 11656 4725 11696
rect 4683 11647 4725 11656
rect 4771 11696 4829 11697
rect 4771 11656 4780 11696
rect 4820 11656 4829 11696
rect 4771 11655 4829 11656
rect 4971 11696 5013 11705
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 5347 11696 5405 11697
rect 5347 11656 5356 11696
rect 5396 11656 5405 11696
rect 5347 11655 5405 11656
rect 6211 11696 6269 11697
rect 6211 11656 6220 11696
rect 6260 11656 6269 11696
rect 6211 11655 6269 11656
rect 34827 11696 34869 11705
rect 34827 11656 34828 11696
rect 34868 11656 34869 11696
rect 34827 11647 34869 11656
rect 35019 11696 35061 11705
rect 35019 11656 35020 11696
rect 35060 11656 35061 11696
rect 35019 11647 35061 11656
rect 35107 11696 35165 11697
rect 35107 11656 35116 11696
rect 35156 11656 35165 11696
rect 35107 11655 35165 11656
rect 35307 11696 35349 11705
rect 35307 11656 35308 11696
rect 35348 11656 35349 11696
rect 35307 11647 35349 11656
rect 35403 11696 35445 11705
rect 35403 11656 35404 11696
rect 35444 11656 35445 11696
rect 35403 11647 35445 11656
rect 35499 11696 35541 11705
rect 35499 11656 35500 11696
rect 35540 11656 35541 11696
rect 35499 11647 35541 11656
rect 35595 11696 35637 11705
rect 35595 11656 35596 11696
rect 35636 11656 35637 11696
rect 35595 11647 35637 11656
rect 36163 11696 36221 11697
rect 36163 11656 36172 11696
rect 36212 11656 36221 11696
rect 36163 11655 36221 11656
rect 36363 11696 36405 11705
rect 36363 11656 36364 11696
rect 36404 11656 36405 11696
rect 36363 11647 36405 11656
rect 36547 11696 36605 11697
rect 36547 11656 36556 11696
rect 36596 11656 36605 11696
rect 36547 11655 36605 11656
rect 36651 11696 36693 11705
rect 36651 11656 36652 11696
rect 36692 11656 36693 11696
rect 36651 11647 36693 11656
rect 36843 11696 36885 11705
rect 36843 11656 36844 11696
rect 36884 11656 36885 11696
rect 36843 11647 36885 11656
rect 38859 11696 38901 11705
rect 38859 11656 38860 11696
rect 38900 11656 38901 11696
rect 38859 11647 38901 11656
rect 39051 11696 39093 11705
rect 39051 11656 39052 11696
rect 39092 11656 39093 11696
rect 39051 11647 39093 11656
rect 39139 11696 39197 11697
rect 39139 11656 39148 11696
rect 39188 11656 39197 11696
rect 39139 11655 39197 11656
rect 39331 11696 39389 11697
rect 39331 11656 39340 11696
rect 39380 11656 39389 11696
rect 39331 11655 39389 11656
rect 39531 11696 39573 11705
rect 39531 11656 39532 11696
rect 39572 11656 39573 11696
rect 39531 11647 39573 11656
rect 41539 11696 41597 11697
rect 41539 11656 41548 11696
rect 41588 11656 41597 11696
rect 41539 11655 41597 11656
rect 41835 11696 41877 11705
rect 41835 11656 41836 11696
rect 41876 11656 41877 11696
rect 41835 11647 41877 11656
rect 42411 11696 42453 11705
rect 42411 11656 42412 11696
rect 42452 11656 42453 11696
rect 42411 11647 42453 11656
rect 42787 11696 42845 11697
rect 42787 11656 42796 11696
rect 42836 11656 42845 11696
rect 42787 11655 42845 11656
rect 43651 11696 43709 11697
rect 43651 11656 43660 11696
rect 43700 11656 43709 11696
rect 43651 11655 43709 11656
rect 47787 11696 47829 11705
rect 47787 11656 47788 11696
rect 47828 11656 47829 11696
rect 47787 11647 47829 11656
rect 47883 11696 47925 11705
rect 47883 11656 47884 11696
rect 47924 11656 47925 11696
rect 47883 11647 47925 11656
rect 47979 11696 48021 11705
rect 47979 11656 47980 11696
rect 48020 11656 48021 11696
rect 47979 11647 48021 11656
rect 48075 11696 48117 11705
rect 48075 11656 48076 11696
rect 48116 11656 48117 11696
rect 48075 11647 48117 11656
rect 48267 11696 48309 11705
rect 48267 11656 48268 11696
rect 48308 11656 48309 11696
rect 48267 11647 48309 11656
rect 48459 11696 48501 11705
rect 48459 11656 48460 11696
rect 48500 11656 48501 11696
rect 48459 11647 48501 11656
rect 48547 11696 48605 11697
rect 48547 11656 48556 11696
rect 48596 11656 48605 11696
rect 48547 11655 48605 11656
rect 49227 11696 49269 11705
rect 49227 11656 49228 11696
rect 49268 11656 49269 11696
rect 49227 11647 49269 11656
rect 49419 11696 49461 11705
rect 49419 11656 49420 11696
rect 49460 11656 49461 11696
rect 49419 11647 49461 11656
rect 49507 11696 49565 11697
rect 49507 11656 49516 11696
rect 49556 11656 49565 11696
rect 49507 11655 49565 11656
rect 50851 11696 50909 11697
rect 50851 11656 50860 11696
rect 50900 11656 50909 11696
rect 50851 11655 50909 11656
rect 51147 11696 51189 11705
rect 51147 11656 51148 11696
rect 51188 11656 51189 11696
rect 51147 11647 51189 11656
rect 51723 11696 51765 11705
rect 51723 11656 51724 11696
rect 51764 11656 51765 11696
rect 51723 11647 51765 11656
rect 51915 11696 51957 11705
rect 51915 11656 51916 11696
rect 51956 11656 51957 11696
rect 51915 11647 51957 11656
rect 52003 11696 52061 11697
rect 52003 11656 52012 11696
rect 52052 11656 52061 11696
rect 52003 11655 52061 11656
rect 52203 11696 52245 11705
rect 52203 11656 52204 11696
rect 52244 11656 52245 11696
rect 52203 11647 52245 11656
rect 52387 11696 52445 11697
rect 52387 11656 52396 11696
rect 52436 11656 52445 11696
rect 52387 11655 52445 11656
rect 56523 11696 56565 11705
rect 56523 11656 56524 11696
rect 56564 11656 56565 11696
rect 56523 11647 56565 11656
rect 56619 11696 56661 11705
rect 56619 11656 56620 11696
rect 56660 11656 56661 11696
rect 56619 11647 56661 11656
rect 56715 11696 56757 11705
rect 56715 11656 56716 11696
rect 56756 11656 56757 11696
rect 56715 11647 56757 11656
rect 56811 11696 56853 11705
rect 56811 11656 56812 11696
rect 56852 11656 56853 11696
rect 56811 11647 56853 11656
rect 57675 11696 57717 11705
rect 57675 11656 57676 11696
rect 57716 11656 57717 11696
rect 57675 11647 57717 11656
rect 57867 11696 57909 11705
rect 57867 11656 57868 11696
rect 57908 11656 57909 11696
rect 57867 11647 57909 11656
rect 57955 11696 58013 11697
rect 57955 11656 57964 11696
rect 58004 11656 58013 11696
rect 57955 11655 58013 11656
rect 58251 11696 58293 11705
rect 58251 11656 58252 11696
rect 58292 11656 58293 11696
rect 58251 11647 58293 11656
rect 58347 11696 58389 11705
rect 58347 11656 58348 11696
rect 58388 11656 58389 11696
rect 58347 11647 58389 11656
rect 58443 11696 58485 11705
rect 58443 11656 58444 11696
rect 58484 11656 58485 11696
rect 58443 11647 58485 11656
rect 58827 11696 58869 11705
rect 58827 11656 58828 11696
rect 58868 11656 58869 11696
rect 58827 11647 58869 11656
rect 59019 11696 59061 11705
rect 59019 11656 59020 11696
rect 59060 11656 59061 11696
rect 59019 11647 59061 11656
rect 59107 11696 59165 11697
rect 59107 11656 59116 11696
rect 59156 11656 59165 11696
rect 59107 11655 59165 11656
rect 59683 11696 59741 11697
rect 59683 11656 59692 11696
rect 59732 11656 59741 11696
rect 59683 11655 59741 11656
rect 60547 11696 60605 11697
rect 60547 11656 60556 11696
rect 60596 11656 60605 11696
rect 60547 11655 60605 11656
rect 62763 11696 62805 11705
rect 62763 11656 62764 11696
rect 62804 11656 62805 11696
rect 62763 11647 62805 11656
rect 62859 11696 62901 11705
rect 62859 11656 62860 11696
rect 62900 11656 62901 11696
rect 62859 11647 62901 11656
rect 62955 11696 62997 11705
rect 62955 11656 62956 11696
rect 62996 11656 62997 11696
rect 62955 11647 62997 11656
rect 63051 11696 63093 11705
rect 63051 11656 63052 11696
rect 63092 11656 63093 11696
rect 63051 11647 63093 11656
rect 63243 11696 63285 11705
rect 63243 11656 63244 11696
rect 63284 11656 63285 11696
rect 63243 11647 63285 11656
rect 63435 11696 63477 11705
rect 63435 11656 63436 11696
rect 63476 11656 63477 11696
rect 63435 11647 63477 11656
rect 63523 11696 63581 11697
rect 63523 11656 63532 11696
rect 63572 11656 63581 11696
rect 63523 11655 63581 11656
rect 63811 11696 63869 11697
rect 63811 11656 63820 11696
rect 63860 11656 63869 11696
rect 63811 11655 63869 11656
rect 63915 11696 63957 11705
rect 63915 11656 63916 11696
rect 63956 11656 63957 11696
rect 63915 11647 63957 11656
rect 64011 11696 64053 11705
rect 64011 11656 64012 11696
rect 64052 11656 64053 11696
rect 64011 11647 64053 11656
rect 64203 11696 64245 11705
rect 64203 11656 64204 11696
rect 64244 11656 64245 11696
rect 64203 11647 64245 11656
rect 64395 11696 64437 11705
rect 64395 11656 64396 11696
rect 64436 11656 64437 11696
rect 64395 11647 64437 11656
rect 64483 11696 64541 11697
rect 64483 11656 64492 11696
rect 64532 11656 64541 11696
rect 64483 11655 64541 11656
rect 68907 11696 68949 11705
rect 68907 11656 68908 11696
rect 68948 11656 68949 11696
rect 68907 11647 68949 11656
rect 69099 11696 69141 11705
rect 69099 11656 69100 11696
rect 69140 11656 69141 11696
rect 69099 11647 69141 11656
rect 69187 11696 69245 11697
rect 69187 11656 69196 11696
rect 69236 11656 69245 11696
rect 69187 11655 69245 11656
rect 69475 11696 69533 11697
rect 69475 11656 69484 11696
rect 69524 11656 69533 11696
rect 69475 11655 69533 11656
rect 69771 11696 69813 11705
rect 69771 11656 69772 11696
rect 69812 11656 69813 11696
rect 69771 11647 69813 11656
rect 70435 11696 70493 11697
rect 70435 11656 70444 11696
rect 70484 11656 70493 11696
rect 70435 11655 70493 11656
rect 70635 11696 70677 11705
rect 70635 11656 70636 11696
rect 70676 11656 70677 11696
rect 70635 11647 70677 11656
rect 72931 11696 72989 11697
rect 72931 11656 72940 11696
rect 72980 11656 72989 11696
rect 72931 11655 72989 11656
rect 73795 11696 73853 11697
rect 73795 11656 73804 11696
rect 73844 11656 73853 11696
rect 73795 11655 73853 11656
rect 75331 11696 75389 11697
rect 75331 11656 75340 11696
rect 75380 11656 75389 11696
rect 75331 11655 75389 11656
rect 75627 11696 75669 11705
rect 75627 11656 75628 11696
rect 75668 11656 75669 11696
rect 75627 11647 75669 11656
rect 75723 11696 75765 11705
rect 75723 11656 75724 11696
rect 75764 11656 75765 11696
rect 75723 11647 75765 11656
rect 76491 11696 76533 11705
rect 76491 11656 76492 11696
rect 76532 11656 76533 11696
rect 76491 11647 76533 11656
rect 76683 11696 76725 11705
rect 76683 11656 76684 11696
rect 76724 11656 76725 11696
rect 76683 11647 76725 11656
rect 76771 11696 76829 11697
rect 76771 11656 76780 11696
rect 76820 11656 76829 11696
rect 76771 11655 76829 11656
rect 76963 11696 77021 11697
rect 76963 11656 76972 11696
rect 77012 11656 77021 11696
rect 76963 11655 77021 11656
rect 77163 11696 77205 11705
rect 77163 11656 77164 11696
rect 77204 11656 77205 11696
rect 77163 11647 77205 11656
rect 1323 11612 1365 11621
rect 1323 11572 1324 11612
rect 1364 11572 1365 11612
rect 1323 11563 1365 11572
rect 4011 11612 4053 11621
rect 4011 11572 4012 11612
rect 4052 11572 4053 11612
rect 4011 11563 4053 11572
rect 4587 11612 4629 11621
rect 4587 11572 4588 11612
rect 4628 11572 4629 11612
rect 4587 11563 4629 11572
rect 41931 11612 41973 11621
rect 41931 11572 41932 11612
rect 41972 11572 41973 11612
rect 41931 11563 41973 11572
rect 51243 11612 51285 11621
rect 51243 11572 51244 11612
rect 51284 11572 51285 11612
rect 51243 11563 51285 11572
rect 52299 11612 52341 11621
rect 52299 11572 52300 11612
rect 52340 11572 52341 11612
rect 52299 11563 52341 11572
rect 58923 11612 58965 11621
rect 58923 11572 58924 11612
rect 58964 11572 58965 11612
rect 58923 11563 58965 11572
rect 59307 11612 59349 11621
rect 59307 11572 59308 11612
rect 59348 11572 59349 11612
rect 59307 11563 59349 11572
rect 69867 11612 69909 11621
rect 69867 11572 69868 11612
rect 69908 11572 69909 11612
rect 69867 11563 69909 11572
rect 72555 11612 72597 11621
rect 72555 11572 72556 11612
rect 72596 11572 72597 11612
rect 72555 11563 72597 11572
rect 77067 11612 77109 11621
rect 77067 11572 77068 11612
rect 77108 11572 77109 11612
rect 77067 11563 77109 11572
rect 939 11528 981 11537
rect 939 11488 940 11528
rect 980 11488 981 11528
rect 939 11479 981 11488
rect 3715 11528 3773 11529
rect 3715 11488 3724 11528
rect 3764 11488 3773 11528
rect 3715 11487 3773 11488
rect 7363 11528 7421 11529
rect 7363 11488 7372 11528
rect 7412 11488 7421 11528
rect 7363 11487 7421 11488
rect 57763 11528 57821 11529
rect 57763 11488 57772 11528
rect 57812 11488 57821 11528
rect 57763 11487 57821 11488
rect 58147 11528 58205 11529
rect 58147 11488 58156 11528
rect 58196 11488 58205 11528
rect 58147 11487 58205 11488
rect 63331 11528 63389 11529
rect 63331 11488 63340 11528
rect 63380 11488 63389 11528
rect 63331 11487 63389 11488
rect 74947 11528 75005 11529
rect 74947 11488 74956 11528
rect 74996 11488 75005 11528
rect 74947 11487 75005 11488
rect 576 11360 79584 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79584 11360
rect 576 11296 79584 11320
rect 651 11192 693 11201
rect 651 11152 652 11192
rect 692 11152 693 11192
rect 651 11143 693 11152
rect 42603 11192 42645 11201
rect 42603 11152 42604 11192
rect 42644 11152 42645 11192
rect 42603 11143 42645 11152
rect 46723 11192 46781 11193
rect 46723 11152 46732 11192
rect 46772 11152 46781 11192
rect 46723 11151 46781 11152
rect 48163 11192 48221 11193
rect 48163 11152 48172 11192
rect 48212 11152 48221 11192
rect 48163 11151 48221 11152
rect 56323 11192 56381 11193
rect 56323 11152 56332 11192
rect 56372 11152 56381 11192
rect 56323 11151 56381 11152
rect 58915 11192 58973 11193
rect 58915 11152 58924 11192
rect 58964 11152 58973 11192
rect 58915 11151 58973 11152
rect 60931 11192 60989 11193
rect 60931 11152 60940 11192
rect 60980 11152 60989 11192
rect 60931 11151 60989 11152
rect 75235 11192 75293 11193
rect 75235 11152 75244 11192
rect 75284 11152 75293 11192
rect 75235 11151 75293 11152
rect 3531 11108 3573 11117
rect 3531 11068 3532 11108
rect 3572 11068 3573 11108
rect 3531 11059 3573 11068
rect 4971 11108 5013 11117
rect 4971 11068 4972 11108
rect 5012 11068 5013 11108
rect 4971 11059 5013 11068
rect 59403 11108 59445 11117
rect 59403 11068 59404 11108
rect 59444 11068 59445 11108
rect 59403 11059 59445 11068
rect 63339 11108 63381 11117
rect 63339 11068 63340 11108
rect 63380 11068 63381 11108
rect 63339 11059 63381 11068
rect 76203 11108 76245 11117
rect 76203 11068 76204 11108
rect 76244 11068 76245 11108
rect 76203 11059 76245 11068
rect 1803 11024 1845 11033
rect 1803 10984 1804 11024
rect 1844 10984 1845 11024
rect 1803 10975 1845 10984
rect 1899 11024 1941 11033
rect 1899 10984 1900 11024
rect 1940 10984 1941 11024
rect 1899 10975 1941 10984
rect 1995 11024 2037 11033
rect 1995 10984 1996 11024
rect 2036 10984 2037 11024
rect 1995 10975 2037 10984
rect 2091 11024 2133 11033
rect 2091 10984 2092 11024
rect 2132 10984 2133 11024
rect 2091 10975 2133 10984
rect 2283 11024 2325 11033
rect 2283 10984 2284 11024
rect 2324 10984 2325 11024
rect 2283 10975 2325 10984
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2563 11024 2621 11025
rect 2563 10984 2572 11024
rect 2612 10984 2621 11024
rect 2563 10983 2621 10984
rect 3139 11024 3197 11025
rect 3139 10984 3148 11024
rect 3188 10984 3197 11024
rect 3139 10983 3197 10984
rect 3435 11024 3477 11033
rect 3435 10984 3436 11024
rect 3476 10984 3477 11024
rect 3435 10975 3477 10984
rect 4867 11024 4925 11025
rect 4867 10984 4876 11024
rect 4916 10984 4925 11024
rect 4867 10983 4925 10984
rect 5067 11024 5109 11033
rect 5067 10984 5068 11024
rect 5108 10984 5109 11024
rect 5067 10975 5109 10984
rect 36451 11024 36509 11025
rect 36451 10984 36460 11024
rect 36500 10984 36509 11024
rect 36451 10983 36509 10984
rect 36555 11024 36597 11033
rect 36555 10984 36556 11024
rect 36596 10984 36597 11024
rect 36555 10975 36597 10984
rect 36747 11024 36789 11033
rect 36747 10984 36748 11024
rect 36788 10984 36789 11024
rect 36747 10975 36789 10984
rect 36931 11024 36989 11025
rect 36931 10984 36940 11024
rect 36980 10984 36989 11024
rect 36931 10983 36989 10984
rect 37035 11024 37077 11033
rect 37035 10984 37036 11024
rect 37076 10984 37077 11024
rect 37035 10975 37077 10984
rect 37227 11024 37269 11033
rect 37227 10984 37228 11024
rect 37268 10984 37269 11024
rect 37227 10975 37269 10984
rect 37419 11024 37461 11033
rect 37419 10984 37420 11024
rect 37460 10984 37461 11024
rect 37419 10975 37461 10984
rect 37515 11024 37557 11033
rect 37515 10984 37516 11024
rect 37556 10984 37557 11024
rect 37515 10975 37557 10984
rect 37611 11024 37653 11033
rect 37611 10984 37612 11024
rect 37652 10984 37653 11024
rect 37611 10975 37653 10984
rect 37707 11024 37749 11033
rect 37707 10984 37708 11024
rect 37748 10984 37749 11024
rect 37707 10975 37749 10984
rect 38563 11024 38621 11025
rect 38563 10984 38572 11024
rect 38612 10984 38621 11024
rect 38563 10983 38621 10984
rect 38859 11024 38901 11033
rect 38859 10984 38860 11024
rect 38900 10984 38901 11024
rect 38859 10975 38901 10984
rect 38955 11024 38997 11033
rect 38955 10984 38956 11024
rect 38996 10984 38997 11024
rect 38955 10975 38997 10984
rect 39427 11024 39485 11025
rect 39427 10984 39436 11024
rect 39476 10984 39485 11024
rect 39427 10983 39485 10984
rect 39627 11024 39669 11033
rect 39627 10984 39628 11024
rect 39668 10984 39669 11024
rect 39627 10975 39669 10984
rect 40675 11024 40733 11025
rect 40675 10984 40684 11024
rect 40724 10984 40733 11024
rect 40675 10983 40733 10984
rect 42891 11024 42933 11033
rect 42891 10984 42892 11024
rect 42932 10984 42933 11024
rect 42891 10975 42933 10984
rect 43075 11024 43133 11025
rect 43075 10984 43084 11024
rect 43124 10984 43133 11024
rect 43075 10983 43133 10984
rect 43947 11024 43989 11033
rect 43947 10984 43948 11024
rect 43988 10984 43989 11024
rect 43947 10975 43989 10984
rect 44131 11024 44189 11025
rect 44131 10984 44140 11024
rect 44180 10984 44189 11024
rect 44131 10983 44189 10984
rect 44331 11024 44373 11033
rect 44331 10984 44332 11024
rect 44372 10984 44373 11024
rect 44331 10975 44373 10984
rect 44707 11024 44765 11025
rect 44707 10984 44716 11024
rect 44756 10984 44765 11024
rect 44707 10983 44765 10984
rect 45571 11024 45629 11025
rect 45571 10984 45580 11024
rect 45620 10984 45629 11024
rect 45571 10983 45629 10984
rect 46915 11024 46973 11025
rect 46915 10984 46924 11024
rect 46964 10984 46973 11024
rect 46915 10983 46973 10984
rect 47115 11024 47157 11033
rect 47115 10984 47116 11024
rect 47156 10984 47157 11024
rect 47115 10975 47157 10984
rect 49315 11024 49373 11025
rect 49315 10984 49324 11024
rect 49364 10984 49373 11024
rect 49315 10983 49373 10984
rect 50179 11024 50237 11025
rect 50179 10984 50188 11024
rect 50228 10984 50237 11024
rect 50179 10983 50237 10984
rect 50571 11024 50613 11033
rect 50571 10984 50572 11024
rect 50612 10984 50613 11024
rect 50571 10975 50613 10984
rect 50763 11024 50805 11033
rect 50763 10984 50764 11024
rect 50804 10984 50805 11024
rect 50763 10975 50805 10984
rect 50859 11024 50901 11033
rect 50859 10984 50860 11024
rect 50900 10984 50901 11024
rect 50859 10975 50901 10984
rect 50955 11024 50997 11033
rect 50955 10984 50956 11024
rect 50996 10984 50997 11024
rect 50955 10975 50997 10984
rect 51051 11024 51093 11033
rect 51051 10984 51052 11024
rect 51092 10984 51093 11024
rect 51051 10975 51093 10984
rect 51243 11024 51285 11033
rect 51243 10984 51244 11024
rect 51284 10984 51285 11024
rect 51243 10975 51285 10984
rect 51435 11024 51477 11033
rect 51435 10984 51436 11024
rect 51476 10984 51477 11024
rect 51435 10975 51477 10984
rect 51523 11024 51581 11025
rect 51523 10984 51532 11024
rect 51572 10984 51581 11024
rect 51523 10983 51581 10984
rect 52491 11024 52533 11033
rect 52491 10984 52492 11024
rect 52532 10984 52533 11024
rect 52491 10975 52533 10984
rect 52683 11024 52725 11033
rect 52683 10984 52684 11024
rect 52724 10984 52725 11024
rect 52683 10975 52725 10984
rect 52771 11024 52829 11025
rect 52771 10984 52780 11024
rect 52820 10984 52829 11024
rect 52771 10983 52829 10984
rect 53067 11024 53109 11033
rect 53067 10984 53068 11024
rect 53108 10984 53109 11024
rect 53067 10975 53109 10984
rect 53163 11024 53205 11033
rect 53163 10984 53164 11024
rect 53204 10984 53205 11024
rect 53443 11024 53501 11025
rect 53163 10975 53205 10984
rect 53251 11001 53309 11002
rect 53251 10961 53260 11001
rect 53300 10961 53309 11001
rect 53443 10984 53452 11024
rect 53492 10984 53501 11024
rect 53443 10983 53501 10984
rect 53547 11024 53589 11033
rect 53547 10984 53548 11024
rect 53588 10984 53589 11024
rect 53547 10975 53589 10984
rect 53739 11024 53781 11033
rect 53739 10984 53740 11024
rect 53780 10984 53781 11024
rect 53739 10975 53781 10984
rect 53931 11024 53973 11033
rect 53931 10984 53932 11024
rect 53972 10984 53973 11024
rect 53931 10975 53973 10984
rect 54307 11024 54365 11025
rect 54307 10984 54316 11024
rect 54356 10984 54365 11024
rect 54307 10983 54365 10984
rect 55171 11024 55229 11025
rect 55171 10984 55180 11024
rect 55220 10984 55229 11024
rect 55171 10983 55229 10984
rect 56523 11024 56565 11033
rect 56523 10984 56524 11024
rect 56564 10984 56565 11024
rect 56523 10975 56565 10984
rect 56899 11024 56957 11025
rect 56899 10984 56908 11024
rect 56948 10984 56957 11024
rect 56899 10983 56957 10984
rect 57763 11024 57821 11025
rect 57763 10984 57772 11024
rect 57812 10984 57821 11024
rect 57763 10983 57821 10984
rect 59499 11024 59541 11033
rect 59499 10984 59500 11024
rect 59540 10984 59541 11024
rect 59499 10975 59541 10984
rect 59779 11024 59837 11025
rect 59779 10984 59788 11024
rect 59828 10984 59837 11024
rect 59779 10983 59837 10984
rect 62083 11024 62141 11025
rect 62083 10984 62092 11024
rect 62132 10984 62141 11024
rect 62083 10983 62141 10984
rect 62947 11024 63005 11025
rect 62947 10984 62956 11024
rect 62996 10984 63005 11024
rect 62947 10983 63005 10984
rect 64491 11024 64533 11033
rect 64491 10984 64492 11024
rect 64532 10984 64533 11024
rect 64491 10975 64533 10984
rect 64675 11024 64733 11025
rect 64675 10984 64684 11024
rect 64724 10984 64733 11024
rect 64675 10983 64733 10984
rect 64875 11024 64917 11033
rect 64875 10984 64876 11024
rect 64916 10984 64917 11024
rect 64875 10975 64917 10984
rect 65067 11024 65109 11033
rect 65067 10984 65068 11024
rect 65108 10984 65109 11024
rect 65067 10975 65109 10984
rect 65155 11024 65213 11025
rect 65155 10984 65164 11024
rect 65204 10984 65213 11024
rect 65155 10983 65213 10984
rect 68907 11024 68949 11033
rect 68907 10984 68908 11024
rect 68948 10984 68949 11024
rect 68907 10975 68949 10984
rect 69099 11024 69141 11033
rect 69099 10984 69100 11024
rect 69140 10984 69141 11024
rect 69099 10975 69141 10984
rect 69187 11024 69245 11025
rect 69187 10984 69196 11024
rect 69236 10984 69245 11024
rect 69187 10983 69245 10984
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 74763 11024 74805 11033
rect 74763 10984 74764 11024
rect 74804 10984 74805 11024
rect 74763 10975 74805 10984
rect 74859 11024 74901 11033
rect 74859 10984 74860 11024
rect 74900 10984 74901 11024
rect 74859 10975 74901 10984
rect 74955 11024 74997 11033
rect 74955 10984 74956 11024
rect 74996 10984 74997 11024
rect 74955 10975 74997 10984
rect 75147 11024 75189 11033
rect 75147 10984 75148 11024
rect 75188 10984 75189 11024
rect 75147 10975 75189 10984
rect 75339 11024 75381 11033
rect 75339 10984 75340 11024
rect 75380 10984 75381 11024
rect 75339 10975 75381 10984
rect 75427 11024 75485 11025
rect 75427 10984 75436 11024
rect 75476 10984 75485 11024
rect 75427 10983 75485 10984
rect 75627 11024 75669 11033
rect 75627 10984 75628 11024
rect 75668 10984 75669 11024
rect 75627 10975 75669 10984
rect 75819 11024 75861 11033
rect 75819 10984 75820 11024
rect 75860 10984 75861 11024
rect 75819 10975 75861 10984
rect 75907 11024 75965 11025
rect 75907 10984 75916 11024
rect 75956 10984 75965 11024
rect 75907 10983 75965 10984
rect 76107 11024 76149 11033
rect 76107 10984 76108 11024
rect 76148 10984 76149 11024
rect 76107 10975 76149 10984
rect 76310 11023 76352 11032
rect 76310 10983 76311 11023
rect 76351 10983 76352 11023
rect 76310 10974 76352 10983
rect 77067 11024 77109 11033
rect 77067 10984 77068 11024
rect 77108 10984 77109 11024
rect 77067 10975 77109 10984
rect 77251 11024 77309 11025
rect 77251 10984 77260 11024
rect 77300 10984 77309 11024
rect 77251 10983 77309 10984
rect 53251 10960 53309 10961
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 1219 10940 1277 10941
rect 1219 10900 1228 10940
rect 1268 10900 1277 10940
rect 1219 10899 1277 10900
rect 1603 10940 1661 10941
rect 1603 10900 1612 10940
rect 1652 10900 1661 10940
rect 1603 10899 1661 10900
rect 39531 10940 39573 10949
rect 39531 10900 39532 10940
rect 39572 10900 39573 10940
rect 39531 10891 39573 10900
rect 51907 10940 51965 10941
rect 51907 10900 51916 10940
rect 51956 10900 51965 10940
rect 51907 10899 51965 10900
rect 64587 10940 64629 10949
rect 64587 10900 64588 10940
rect 64628 10900 64629 10940
rect 64587 10891 64629 10900
rect 69571 10940 69629 10941
rect 69571 10900 69580 10940
rect 69620 10900 69629 10940
rect 69571 10899 69629 10900
rect 69955 10940 70013 10941
rect 69955 10900 69964 10940
rect 70004 10900 70013 10940
rect 69955 10899 70013 10900
rect 70339 10940 70397 10941
rect 70339 10900 70348 10940
rect 70388 10900 70397 10940
rect 70339 10899 70397 10900
rect 70531 10940 70589 10941
rect 70531 10900 70540 10940
rect 70580 10900 70589 10940
rect 70531 10899 70589 10900
rect 71107 10940 71165 10941
rect 71107 10900 71116 10940
rect 71156 10900 71165 10940
rect 71107 10899 71165 10900
rect 76483 10929 76541 10930
rect 76483 10889 76492 10929
rect 76532 10889 76541 10929
rect 76483 10888 76541 10889
rect 1419 10856 1461 10865
rect 1419 10816 1420 10856
rect 1460 10816 1461 10856
rect 1419 10807 1461 10816
rect 2283 10856 2325 10865
rect 2283 10816 2284 10856
rect 2324 10816 2325 10856
rect 2283 10807 2325 10816
rect 3811 10856 3869 10857
rect 3811 10816 3820 10856
rect 3860 10816 3869 10856
rect 3811 10815 3869 10816
rect 36747 10856 36789 10865
rect 36747 10816 36748 10856
rect 36788 10816 36789 10856
rect 36747 10807 36789 10816
rect 39235 10856 39293 10857
rect 39235 10816 39244 10856
rect 39284 10816 39293 10856
rect 39235 10815 39293 10816
rect 40011 10856 40053 10865
rect 40011 10816 40012 10856
rect 40052 10816 40053 10856
rect 40011 10807 40053 10816
rect 51243 10856 51285 10865
rect 51243 10816 51244 10856
rect 51284 10816 51285 10856
rect 51243 10807 51285 10816
rect 53739 10856 53781 10865
rect 53739 10816 53740 10856
rect 53780 10816 53781 10856
rect 53739 10807 53781 10816
rect 65739 10856 65781 10865
rect 65739 10816 65740 10856
rect 65780 10816 65781 10856
rect 65739 10807 65781 10816
rect 71307 10856 71349 10865
rect 71307 10816 71308 10856
rect 71348 10816 71349 10856
rect 71307 10807 71349 10816
rect 73035 10856 73077 10865
rect 73035 10816 73036 10856
rect 73076 10816 73077 10856
rect 73035 10807 73077 10816
rect 75627 10856 75669 10865
rect 75627 10816 75628 10856
rect 75668 10816 75669 10856
rect 75627 10807 75669 10816
rect 77643 10856 77685 10865
rect 77643 10816 77644 10856
rect 77684 10816 77685 10856
rect 77643 10807 77685 10816
rect 1035 10772 1077 10781
rect 1035 10732 1036 10772
rect 1076 10732 1077 10772
rect 1035 10723 1077 10732
rect 37227 10772 37269 10781
rect 37227 10732 37228 10772
rect 37268 10732 37269 10772
rect 37227 10723 37269 10732
rect 42987 10772 43029 10781
rect 42987 10732 42988 10772
rect 43028 10732 43029 10772
rect 42987 10723 43029 10732
rect 44043 10772 44085 10781
rect 44043 10732 44044 10772
rect 44084 10732 44085 10772
rect 44043 10723 44085 10732
rect 47019 10772 47061 10781
rect 47019 10732 47020 10772
rect 47060 10732 47061 10772
rect 47019 10723 47061 10732
rect 51723 10772 51765 10781
rect 51723 10732 51724 10772
rect 51764 10732 51765 10772
rect 51723 10723 51765 10732
rect 52491 10772 52533 10781
rect 52491 10732 52492 10772
rect 52532 10732 52533 10772
rect 52491 10723 52533 10732
rect 59107 10772 59165 10773
rect 59107 10732 59116 10772
rect 59156 10732 59165 10772
rect 59107 10731 59165 10732
rect 64875 10772 64917 10781
rect 64875 10732 64876 10772
rect 64916 10732 64917 10772
rect 64875 10723 64917 10732
rect 68907 10772 68949 10781
rect 68907 10732 68908 10772
rect 68948 10732 68949 10772
rect 68907 10723 68949 10732
rect 69387 10772 69429 10781
rect 69387 10732 69388 10772
rect 69428 10732 69429 10772
rect 69387 10723 69429 10732
rect 69771 10772 69813 10781
rect 69771 10732 69772 10772
rect 69812 10732 69813 10772
rect 69771 10723 69813 10732
rect 70155 10772 70197 10781
rect 70155 10732 70156 10772
rect 70196 10732 70197 10772
rect 70155 10723 70197 10732
rect 70731 10772 70773 10781
rect 70731 10732 70732 10772
rect 70772 10732 70773 10772
rect 70731 10723 70773 10732
rect 70923 10772 70965 10781
rect 70923 10732 70924 10772
rect 70964 10732 70965 10772
rect 70923 10723 70965 10732
rect 76683 10772 76725 10781
rect 76683 10732 76684 10772
rect 76724 10732 76725 10772
rect 76683 10723 76725 10732
rect 77163 10772 77205 10781
rect 77163 10732 77164 10772
rect 77204 10732 77205 10772
rect 77163 10723 77205 10732
rect 576 10604 79584 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79584 10604
rect 576 10540 79584 10564
rect 2571 10436 2613 10445
rect 2571 10396 2572 10436
rect 2612 10396 2613 10436
rect 2571 10387 2613 10396
rect 38851 10436 38909 10437
rect 38851 10396 38860 10436
rect 38900 10396 38909 10436
rect 38851 10395 38909 10396
rect 41827 10436 41885 10437
rect 41827 10396 41836 10436
rect 41876 10396 41885 10436
rect 41827 10395 41885 10396
rect 42315 10436 42357 10445
rect 42315 10396 42316 10436
rect 42356 10396 42357 10436
rect 42315 10387 42357 10396
rect 44811 10436 44853 10445
rect 44811 10396 44812 10436
rect 44852 10396 44853 10436
rect 44811 10387 44853 10396
rect 49219 10436 49277 10437
rect 49219 10396 49228 10436
rect 49268 10396 49277 10436
rect 49219 10395 49277 10396
rect 53739 10436 53781 10445
rect 53739 10396 53740 10436
rect 53780 10396 53781 10436
rect 53739 10387 53781 10396
rect 58059 10436 58101 10445
rect 58059 10396 58060 10436
rect 58100 10396 58101 10436
rect 58059 10387 58101 10396
rect 63435 10436 63477 10445
rect 63435 10396 63436 10436
rect 63476 10396 63477 10436
rect 63435 10387 63477 10396
rect 64195 10436 64253 10437
rect 64195 10396 64204 10436
rect 64244 10396 64253 10436
rect 64195 10395 64253 10396
rect 67651 10436 67709 10437
rect 67651 10396 67660 10436
rect 67700 10396 67709 10436
rect 67651 10395 67709 10396
rect 72931 10436 72989 10437
rect 72931 10396 72940 10436
rect 72980 10396 72989 10436
rect 72931 10395 72989 10396
rect 75907 10436 75965 10437
rect 75907 10396 75916 10436
rect 75956 10396 75965 10436
rect 75907 10395 75965 10396
rect 76867 10436 76925 10437
rect 76867 10396 76876 10436
rect 76916 10396 76925 10436
rect 76867 10395 76925 10396
rect 1515 10352 1557 10361
rect 1515 10312 1516 10352
rect 1556 10312 1557 10352
rect 1515 10303 1557 10312
rect 3051 10352 3093 10361
rect 3051 10312 3052 10352
rect 3092 10312 3093 10352
rect 3051 10303 3093 10312
rect 43555 10352 43613 10353
rect 43555 10312 43564 10352
rect 43604 10312 43613 10352
rect 43555 10311 43613 10312
rect 53443 10352 53501 10353
rect 53443 10312 53452 10352
rect 53492 10312 53501 10352
rect 53443 10311 53501 10312
rect 54411 10352 54453 10361
rect 54411 10312 54412 10352
rect 54452 10312 54453 10352
rect 54411 10303 54453 10312
rect 57579 10352 57621 10361
rect 57579 10312 57580 10352
rect 57620 10312 57621 10352
rect 57579 10303 57621 10312
rect 58731 10352 58773 10361
rect 58731 10312 58732 10352
rect 58772 10312 58773 10352
rect 58731 10303 58773 10312
rect 62379 10352 62421 10361
rect 62379 10312 62380 10352
rect 62420 10312 62421 10352
rect 62379 10303 62421 10312
rect 67851 10352 67893 10361
rect 67851 10312 67852 10352
rect 67892 10312 67893 10352
rect 67851 10303 67893 10312
rect 69955 10352 70013 10353
rect 69955 10312 69964 10352
rect 70004 10312 70013 10352
rect 69955 10311 70013 10312
rect 70347 10352 70389 10361
rect 70347 10312 70348 10352
rect 70388 10312 70389 10352
rect 70347 10303 70389 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 1699 10268 1757 10269
rect 1699 10228 1708 10268
rect 1748 10228 1757 10268
rect 1699 10227 1757 10228
rect 3235 10268 3293 10269
rect 3235 10228 3244 10268
rect 3284 10228 3293 10268
rect 3235 10227 3293 10228
rect 7179 10268 7221 10277
rect 7179 10228 7180 10268
rect 7220 10228 7221 10268
rect 7179 10219 7221 10228
rect 42115 10268 42173 10269
rect 42115 10228 42124 10268
rect 42164 10228 42173 10268
rect 42115 10227 42173 10228
rect 57379 10268 57437 10269
rect 57379 10228 57388 10268
rect 57428 10228 57437 10268
rect 57379 10227 57437 10228
rect 58915 10268 58973 10269
rect 58915 10228 58924 10268
rect 58964 10228 58973 10268
rect 58915 10227 58973 10228
rect 70147 10268 70205 10269
rect 70147 10228 70156 10268
rect 70196 10228 70205 10268
rect 70147 10227 70205 10228
rect 79467 10268 79509 10277
rect 79467 10228 79468 10268
rect 79508 10228 79509 10268
rect 79467 10219 79509 10228
rect 2571 10184 2613 10193
rect 2571 10144 2572 10184
rect 2612 10144 2613 10184
rect 2571 10135 2613 10144
rect 2763 10184 2805 10193
rect 2763 10144 2764 10184
rect 2804 10144 2805 10184
rect 5155 10184 5213 10185
rect 2763 10135 2805 10144
rect 2861 10169 2919 10170
rect 2861 10129 2870 10169
rect 2910 10129 2919 10169
rect 5155 10144 5164 10184
rect 5204 10144 5213 10184
rect 5155 10143 5213 10144
rect 6019 10184 6077 10185
rect 6019 10144 6028 10184
rect 6068 10144 6077 10184
rect 6019 10143 6077 10144
rect 36459 10184 36501 10193
rect 36459 10144 36460 10184
rect 36500 10144 36501 10184
rect 36459 10135 36501 10144
rect 36835 10184 36893 10185
rect 36835 10144 36844 10184
rect 36884 10144 36893 10184
rect 36835 10143 36893 10144
rect 37699 10184 37757 10185
rect 37699 10144 37708 10184
rect 37748 10144 37757 10184
rect 37699 10143 37757 10144
rect 39811 10184 39869 10185
rect 39811 10144 39820 10184
rect 39860 10144 39869 10184
rect 39811 10143 39869 10144
rect 40675 10184 40733 10185
rect 40675 10144 40684 10184
rect 40724 10144 40733 10184
rect 40675 10143 40733 10144
rect 43947 10184 43989 10193
rect 43947 10144 43948 10184
rect 43988 10144 43989 10184
rect 43947 10135 43989 10144
rect 44227 10184 44285 10185
rect 44227 10144 44236 10184
rect 44276 10144 44285 10184
rect 44227 10143 44285 10144
rect 44515 10184 44573 10185
rect 44515 10144 44524 10184
rect 44564 10144 44573 10184
rect 44515 10143 44573 10144
rect 44619 10184 44661 10193
rect 44619 10144 44620 10184
rect 44660 10144 44661 10184
rect 44619 10135 44661 10144
rect 44811 10184 44853 10193
rect 44811 10144 44812 10184
rect 44852 10144 44853 10184
rect 44811 10135 44853 10144
rect 46347 10184 46389 10193
rect 46347 10144 46348 10184
rect 46388 10144 46389 10184
rect 46347 10135 46389 10144
rect 46539 10184 46581 10193
rect 46539 10144 46540 10184
rect 46580 10144 46581 10184
rect 46539 10135 46581 10144
rect 46627 10184 46685 10185
rect 46627 10144 46636 10184
rect 46676 10144 46685 10184
rect 46627 10143 46685 10144
rect 46827 10184 46869 10193
rect 46827 10144 46828 10184
rect 46868 10144 46869 10184
rect 46827 10135 46869 10144
rect 47203 10184 47261 10185
rect 47203 10144 47212 10184
rect 47252 10144 47261 10184
rect 47203 10143 47261 10144
rect 48067 10184 48125 10185
rect 48067 10144 48076 10184
rect 48116 10144 48125 10184
rect 48067 10143 48125 10144
rect 49803 10184 49845 10193
rect 49803 10144 49804 10184
rect 49844 10144 49845 10184
rect 49803 10135 49845 10144
rect 50179 10184 50237 10185
rect 50179 10144 50188 10184
rect 50228 10144 50237 10184
rect 50179 10143 50237 10144
rect 51043 10184 51101 10185
rect 51043 10144 51052 10184
rect 51092 10144 51101 10184
rect 51043 10143 51101 10144
rect 52771 10184 52829 10185
rect 52771 10144 52780 10184
rect 52820 10144 52829 10184
rect 52771 10143 52829 10144
rect 53067 10184 53109 10193
rect 53067 10144 53068 10184
rect 53108 10144 53109 10184
rect 53067 10135 53109 10144
rect 53643 10184 53685 10193
rect 53643 10144 53644 10184
rect 53684 10144 53685 10184
rect 53643 10135 53685 10144
rect 53827 10184 53885 10185
rect 53827 10144 53836 10184
rect 53876 10144 53885 10184
rect 53827 10143 53885 10144
rect 57763 10184 57821 10185
rect 57763 10144 57772 10184
rect 57812 10144 57821 10184
rect 57763 10143 57821 10144
rect 57867 10184 57909 10193
rect 57867 10144 57868 10184
rect 57908 10144 57909 10184
rect 57867 10135 57909 10144
rect 58059 10184 58101 10193
rect 58059 10144 58060 10184
rect 58100 10144 58101 10184
rect 58059 10135 58101 10144
rect 58251 10184 58293 10193
rect 58251 10144 58252 10184
rect 58292 10144 58293 10184
rect 58251 10135 58293 10144
rect 58443 10184 58485 10193
rect 58443 10144 58444 10184
rect 58484 10144 58485 10184
rect 58443 10135 58485 10144
rect 58531 10184 58589 10185
rect 58531 10144 58540 10184
rect 58580 10144 58589 10184
rect 58531 10143 58589 10144
rect 59115 10184 59157 10193
rect 59115 10144 59116 10184
rect 59156 10144 59157 10184
rect 59115 10135 59157 10144
rect 59299 10184 59357 10185
rect 59299 10144 59308 10184
rect 59348 10144 59357 10184
rect 59299 10143 59357 10144
rect 59491 10184 59549 10185
rect 59491 10144 59500 10184
rect 59540 10144 59549 10184
rect 59491 10143 59549 10144
rect 59691 10184 59733 10193
rect 59691 10144 59692 10184
rect 59732 10144 59733 10184
rect 59691 10135 59733 10144
rect 63435 10184 63477 10193
rect 63435 10144 63436 10184
rect 63476 10144 63477 10184
rect 63435 10135 63477 10144
rect 63627 10184 63669 10193
rect 63627 10144 63628 10184
rect 63668 10144 63669 10184
rect 63627 10135 63669 10144
rect 63715 10184 63773 10185
rect 63715 10144 63724 10184
rect 63764 10144 63773 10184
rect 63715 10143 63773 10144
rect 64587 10184 64629 10193
rect 64587 10144 64588 10184
rect 64628 10144 64629 10184
rect 64587 10135 64629 10144
rect 64867 10184 64925 10185
rect 64867 10144 64876 10184
rect 64916 10144 64925 10184
rect 64867 10143 64925 10144
rect 65259 10184 65301 10193
rect 65259 10144 65260 10184
rect 65300 10144 65301 10184
rect 65259 10135 65301 10144
rect 65635 10184 65693 10185
rect 65635 10144 65644 10184
rect 65684 10144 65693 10184
rect 65635 10143 65693 10144
rect 66499 10184 66557 10185
rect 66499 10144 66508 10184
rect 66548 10144 66557 10184
rect 66499 10143 66557 10144
rect 68331 10184 68373 10193
rect 68331 10144 68332 10184
rect 68372 10144 68373 10184
rect 68331 10135 68373 10144
rect 68427 10184 68469 10193
rect 68427 10144 68428 10184
rect 68468 10144 68469 10184
rect 68427 10135 68469 10144
rect 68523 10184 68565 10193
rect 68523 10144 68524 10184
rect 68564 10144 68565 10184
rect 68523 10135 68565 10144
rect 68715 10184 68757 10193
rect 68715 10144 68716 10184
rect 68756 10144 68757 10184
rect 68715 10135 68757 10144
rect 68907 10184 68949 10193
rect 68907 10144 68908 10184
rect 68948 10144 68949 10184
rect 68907 10135 68949 10144
rect 68995 10184 69053 10185
rect 68995 10144 69004 10184
rect 69044 10144 69053 10184
rect 68995 10143 69053 10144
rect 69283 10184 69341 10185
rect 69283 10144 69292 10184
rect 69332 10144 69341 10184
rect 69283 10143 69341 10144
rect 69579 10184 69621 10193
rect 69579 10144 69580 10184
rect 69620 10144 69621 10184
rect 69579 10135 69621 10144
rect 69675 10184 69717 10193
rect 69675 10144 69676 10184
rect 69716 10144 69717 10184
rect 69675 10135 69717 10144
rect 70915 10184 70973 10185
rect 70915 10144 70924 10184
rect 70964 10144 70973 10184
rect 70915 10143 70973 10144
rect 71779 10184 71837 10185
rect 71779 10144 71788 10184
rect 71828 10144 71837 10184
rect 71779 10143 71837 10144
rect 73891 10184 73949 10185
rect 73891 10144 73900 10184
rect 73940 10144 73949 10184
rect 73891 10143 73949 10144
rect 74755 10184 74813 10185
rect 74755 10144 74764 10184
rect 74804 10144 74813 10184
rect 74755 10143 74813 10144
rect 76195 10184 76253 10185
rect 76195 10144 76204 10184
rect 76244 10144 76253 10184
rect 76195 10143 76253 10144
rect 76491 10184 76533 10193
rect 76491 10144 76492 10184
rect 76532 10144 76533 10184
rect 76491 10135 76533 10144
rect 76587 10184 76629 10193
rect 76587 10144 76588 10184
rect 76628 10144 76629 10184
rect 76587 10135 76629 10144
rect 77443 10184 77501 10185
rect 77443 10144 77452 10184
rect 77492 10144 77501 10184
rect 77443 10143 77501 10144
rect 78307 10184 78365 10185
rect 78307 10144 78316 10184
rect 78356 10144 78365 10184
rect 78307 10143 78365 10144
rect 2861 10128 2919 10129
rect 4779 10100 4821 10109
rect 4779 10060 4780 10100
rect 4820 10060 4821 10100
rect 4779 10051 4821 10060
rect 39435 10100 39477 10109
rect 39435 10060 39436 10100
rect 39476 10060 39477 10100
rect 39435 10051 39477 10060
rect 43851 10100 43893 10109
rect 43851 10060 43852 10100
rect 43892 10060 43893 10100
rect 43851 10051 43893 10060
rect 46443 10100 46485 10109
rect 46443 10060 46444 10100
rect 46484 10060 46485 10100
rect 46443 10051 46485 10060
rect 53163 10100 53205 10109
rect 53163 10060 53164 10100
rect 53204 10060 53205 10100
rect 53163 10051 53205 10060
rect 59211 10100 59253 10109
rect 59211 10060 59212 10100
rect 59252 10060 59253 10100
rect 59211 10051 59253 10060
rect 59595 10100 59637 10109
rect 59595 10060 59596 10100
rect 59636 10060 59637 10100
rect 59595 10051 59637 10060
rect 64491 10100 64533 10109
rect 64491 10060 64492 10100
rect 64532 10060 64533 10100
rect 64491 10051 64533 10060
rect 68235 10100 68277 10109
rect 68235 10060 68236 10100
rect 68276 10060 68277 10100
rect 68235 10051 68277 10060
rect 68811 10100 68853 10109
rect 68811 10060 68812 10100
rect 68852 10060 68853 10100
rect 68811 10051 68853 10060
rect 70539 10100 70581 10109
rect 70539 10060 70540 10100
rect 70580 10060 70581 10100
rect 70539 10051 70581 10060
rect 73515 10100 73557 10109
rect 73515 10060 73516 10100
rect 73556 10060 73557 10100
rect 73515 10051 73557 10060
rect 77067 10100 77109 10109
rect 77067 10060 77068 10100
rect 77108 10060 77109 10100
rect 77067 10051 77109 10060
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 52195 10016 52253 10017
rect 52195 9976 52204 10016
rect 52244 9976 52253 10016
rect 52195 9975 52253 9976
rect 58339 10016 58397 10017
rect 58339 9976 58348 10016
rect 58388 9976 58397 10016
rect 58339 9975 58397 9976
rect 75907 10016 75965 10017
rect 75907 9976 75916 10016
rect 75956 9976 75965 10016
rect 75907 9975 75965 9976
rect 576 9848 79584 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79584 9848
rect 576 9784 79584 9808
rect 651 9680 693 9689
rect 651 9640 652 9680
rect 692 9640 693 9680
rect 651 9631 693 9640
rect 3427 9680 3485 9681
rect 3427 9640 3436 9680
rect 3476 9640 3485 9680
rect 3427 9639 3485 9640
rect 4483 9680 4541 9681
rect 4483 9640 4492 9680
rect 4532 9640 4541 9680
rect 4483 9639 4541 9640
rect 40195 9680 40253 9681
rect 40195 9640 40204 9680
rect 40244 9640 40253 9680
rect 40195 9639 40253 9640
rect 42787 9680 42845 9681
rect 42787 9640 42796 9680
rect 42836 9640 42845 9680
rect 42787 9639 42845 9640
rect 51523 9680 51581 9681
rect 51523 9640 51532 9680
rect 51572 9640 51581 9680
rect 51523 9639 51581 9640
rect 52483 9680 52541 9681
rect 52483 9640 52492 9680
rect 52532 9640 52541 9680
rect 52483 9639 52541 9640
rect 52771 9680 52829 9681
rect 52771 9640 52780 9680
rect 52820 9640 52829 9680
rect 52771 9639 52829 9640
rect 61987 9680 62045 9681
rect 61987 9640 61996 9680
rect 62036 9640 62045 9680
rect 61987 9639 62045 9640
rect 64579 9680 64637 9681
rect 64579 9640 64588 9680
rect 64628 9640 64637 9680
rect 64579 9639 64637 9640
rect 69283 9680 69341 9681
rect 69283 9640 69292 9680
rect 69332 9640 69341 9680
rect 69283 9639 69341 9640
rect 70635 9680 70677 9689
rect 70635 9640 70636 9680
rect 70676 9640 70677 9680
rect 70635 9631 70677 9640
rect 75523 9680 75581 9681
rect 75523 9640 75532 9680
rect 75572 9640 75581 9680
rect 75523 9639 75581 9640
rect 77155 9680 77213 9681
rect 77155 9640 77164 9680
rect 77204 9640 77213 9680
rect 77155 9639 77213 9640
rect 62187 9596 62229 9605
rect 62187 9556 62188 9596
rect 62228 9556 62229 9596
rect 62187 9547 62229 9556
rect 64875 9596 64917 9605
rect 64875 9556 64876 9596
rect 64916 9556 64917 9596
rect 64875 9547 64917 9556
rect 65355 9596 65397 9605
rect 65355 9556 65356 9596
rect 65396 9556 65397 9596
rect 65355 9547 65397 9556
rect 66891 9596 66933 9605
rect 66891 9556 66892 9596
rect 66932 9556 66933 9596
rect 66891 9547 66933 9556
rect 1035 9512 1077 9521
rect 1035 9472 1036 9512
rect 1076 9472 1077 9512
rect 1035 9463 1077 9472
rect 1411 9512 1469 9513
rect 1411 9472 1420 9512
rect 1460 9472 1469 9512
rect 1411 9471 1469 9472
rect 2275 9512 2333 9513
rect 2275 9472 2284 9512
rect 2324 9472 2333 9512
rect 2275 9471 2333 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3811 9512 3869 9513
rect 3811 9472 3820 9512
rect 3860 9472 3869 9512
rect 3811 9471 3869 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 4867 9512 4925 9513
rect 4867 9472 4876 9512
rect 4916 9472 4925 9512
rect 4867 9471 4925 9472
rect 5067 9512 5109 9521
rect 5067 9472 5068 9512
rect 5108 9472 5109 9512
rect 5067 9463 5109 9472
rect 39235 9512 39293 9513
rect 39235 9472 39244 9512
rect 39284 9472 39293 9512
rect 39235 9471 39293 9472
rect 39339 9512 39381 9521
rect 39339 9472 39340 9512
rect 39380 9472 39381 9512
rect 39339 9463 39381 9472
rect 39531 9512 39573 9521
rect 39531 9472 39532 9512
rect 39572 9472 39573 9512
rect 39531 9463 39573 9472
rect 40003 9512 40061 9513
rect 40003 9472 40012 9512
rect 40052 9472 40061 9512
rect 40003 9471 40061 9472
rect 40107 9512 40149 9521
rect 40107 9472 40108 9512
rect 40148 9472 40149 9512
rect 40107 9463 40149 9472
rect 40299 9512 40341 9521
rect 40299 9472 40300 9512
rect 40340 9472 40341 9512
rect 40299 9463 40341 9472
rect 40683 9512 40725 9521
rect 40683 9472 40684 9512
rect 40724 9472 40725 9512
rect 40683 9463 40725 9472
rect 40779 9512 40821 9521
rect 40779 9472 40780 9512
rect 40820 9472 40821 9512
rect 40779 9463 40821 9472
rect 40875 9512 40917 9521
rect 40875 9472 40876 9512
rect 40916 9472 40917 9512
rect 40875 9463 40917 9472
rect 40971 9512 41013 9521
rect 40971 9472 40972 9512
rect 41012 9472 41013 9512
rect 40971 9463 41013 9472
rect 41731 9512 41789 9513
rect 41731 9472 41740 9512
rect 41780 9472 41789 9512
rect 41731 9471 41789 9472
rect 41835 9512 41877 9521
rect 41835 9472 41836 9512
rect 41876 9472 41877 9512
rect 41835 9463 41877 9472
rect 42027 9512 42069 9521
rect 42027 9472 42028 9512
rect 42068 9472 42069 9512
rect 42027 9463 42069 9472
rect 42211 9512 42269 9513
rect 42211 9472 42220 9512
rect 42260 9472 42269 9512
rect 42211 9471 42269 9472
rect 42315 9512 42357 9521
rect 42315 9472 42316 9512
rect 42356 9472 42357 9512
rect 42315 9463 42357 9472
rect 42507 9512 42549 9521
rect 42507 9472 42508 9512
rect 42548 9472 42549 9512
rect 42507 9463 42549 9472
rect 42891 9512 42933 9521
rect 42891 9472 42892 9512
rect 42932 9472 42933 9512
rect 42891 9463 42933 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43083 9512 43125 9521
rect 43083 9472 43084 9512
rect 43124 9472 43125 9512
rect 43083 9463 43125 9472
rect 43947 9512 43989 9521
rect 43947 9472 43948 9512
rect 43988 9472 43989 9512
rect 43947 9463 43989 9472
rect 44131 9512 44189 9513
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44131 9471 44189 9472
rect 46635 9512 46677 9521
rect 46635 9472 46636 9512
rect 46676 9472 46677 9512
rect 46635 9463 46677 9472
rect 46731 9512 46773 9521
rect 46731 9472 46732 9512
rect 46772 9472 46773 9512
rect 46731 9463 46773 9472
rect 47011 9512 47069 9513
rect 47011 9472 47020 9512
rect 47060 9472 47069 9512
rect 47011 9471 47069 9472
rect 51435 9512 51477 9521
rect 51435 9472 51436 9512
rect 51476 9472 51477 9512
rect 51435 9463 51477 9472
rect 51627 9512 51669 9521
rect 51627 9472 51628 9512
rect 51668 9472 51669 9512
rect 51627 9463 51669 9472
rect 51715 9512 51773 9513
rect 51715 9472 51724 9512
rect 51764 9472 51773 9512
rect 51715 9471 51773 9472
rect 52203 9512 52245 9521
rect 52203 9472 52204 9512
rect 52244 9472 52245 9512
rect 52203 9463 52245 9472
rect 52299 9512 52341 9521
rect 52299 9472 52300 9512
rect 52340 9472 52341 9512
rect 52299 9463 52341 9472
rect 52395 9512 52437 9521
rect 52395 9472 52396 9512
rect 52436 9472 52437 9512
rect 52395 9463 52437 9472
rect 52683 9512 52725 9521
rect 52683 9472 52684 9512
rect 52724 9472 52725 9512
rect 52683 9463 52725 9472
rect 52875 9512 52917 9521
rect 52875 9472 52876 9512
rect 52916 9472 52917 9512
rect 52875 9463 52917 9472
rect 52963 9512 53021 9513
rect 52963 9472 52972 9512
rect 53012 9472 53021 9512
rect 52963 9471 53021 9472
rect 53635 9512 53693 9513
rect 53635 9472 53644 9512
rect 53684 9472 53693 9512
rect 53635 9471 53693 9472
rect 53835 9512 53877 9521
rect 53835 9472 53836 9512
rect 53876 9472 53877 9512
rect 53835 9463 53877 9472
rect 54123 9512 54165 9521
rect 54123 9472 54124 9512
rect 54164 9472 54165 9512
rect 54123 9463 54165 9472
rect 54307 9512 54365 9513
rect 54307 9472 54316 9512
rect 54356 9472 54365 9512
rect 54307 9471 54365 9472
rect 57771 9512 57813 9521
rect 57771 9472 57772 9512
rect 57812 9472 57813 9512
rect 57771 9463 57813 9472
rect 57963 9512 58005 9521
rect 57963 9472 57964 9512
rect 58004 9472 58005 9512
rect 57963 9463 58005 9472
rect 58051 9512 58109 9513
rect 58051 9472 58060 9512
rect 58100 9472 58109 9512
rect 58051 9471 58109 9472
rect 58339 9512 58397 9513
rect 58339 9472 58348 9512
rect 58388 9472 58397 9512
rect 58339 9471 58397 9472
rect 58635 9512 58677 9521
rect 58635 9472 58636 9512
rect 58676 9472 58677 9512
rect 58635 9463 58677 9472
rect 58731 9512 58773 9521
rect 58731 9472 58732 9512
rect 58772 9472 58773 9512
rect 58731 9463 58773 9472
rect 59595 9512 59637 9521
rect 59595 9472 59596 9512
rect 59636 9472 59637 9512
rect 59595 9463 59637 9472
rect 59971 9512 60029 9513
rect 59971 9472 59980 9512
rect 60020 9472 60029 9512
rect 59971 9471 60029 9472
rect 60835 9512 60893 9513
rect 60835 9472 60844 9512
rect 60884 9472 60893 9512
rect 60835 9471 60893 9472
rect 62563 9512 62621 9513
rect 62563 9472 62572 9512
rect 62612 9472 62621 9512
rect 62563 9471 62621 9472
rect 63427 9512 63485 9513
rect 63427 9472 63436 9512
rect 63476 9472 63485 9512
rect 63427 9471 63485 9472
rect 64779 9512 64821 9521
rect 64779 9472 64780 9512
rect 64820 9472 64821 9512
rect 64779 9463 64821 9472
rect 64971 9512 65013 9521
rect 64971 9472 64972 9512
rect 65012 9472 65013 9512
rect 64971 9463 65013 9472
rect 65059 9512 65117 9513
rect 65059 9472 65068 9512
rect 65108 9472 65117 9512
rect 65059 9471 65117 9472
rect 65251 9512 65309 9513
rect 65251 9472 65260 9512
rect 65300 9472 65309 9512
rect 65251 9471 65309 9472
rect 65451 9512 65493 9521
rect 65451 9472 65452 9512
rect 65492 9472 65493 9512
rect 65451 9463 65493 9472
rect 67267 9512 67325 9513
rect 67267 9472 67276 9512
rect 67316 9472 67325 9512
rect 67267 9471 67325 9472
rect 68131 9512 68189 9513
rect 68131 9472 68140 9512
rect 68180 9472 68189 9512
rect 68131 9471 68189 9472
rect 69475 9512 69533 9513
rect 69475 9472 69484 9512
rect 69524 9472 69533 9512
rect 69475 9471 69533 9472
rect 69579 9512 69621 9521
rect 69579 9472 69580 9512
rect 69620 9472 69621 9512
rect 69579 9463 69621 9472
rect 69771 9512 69813 9521
rect 69771 9472 69772 9512
rect 69812 9472 69813 9512
rect 69771 9463 69813 9472
rect 69963 9512 70005 9521
rect 69963 9472 69964 9512
rect 70004 9472 70005 9512
rect 69963 9463 70005 9472
rect 70155 9512 70197 9521
rect 70155 9472 70156 9512
rect 70196 9472 70197 9512
rect 70155 9463 70197 9472
rect 70243 9512 70301 9513
rect 70243 9472 70252 9512
rect 70292 9472 70301 9512
rect 70243 9471 70301 9472
rect 70819 9512 70877 9513
rect 70819 9472 70828 9512
rect 70868 9472 70877 9512
rect 70819 9471 70877 9472
rect 70923 9512 70965 9521
rect 70923 9472 70924 9512
rect 70964 9472 70965 9512
rect 70923 9463 70965 9472
rect 71019 9512 71061 9521
rect 71019 9472 71020 9512
rect 71060 9472 71061 9512
rect 71019 9463 71061 9472
rect 71299 9512 71357 9513
rect 71299 9472 71308 9512
rect 71348 9472 71357 9512
rect 71299 9471 71357 9472
rect 71499 9512 71541 9521
rect 71499 9472 71500 9512
rect 71540 9472 71541 9512
rect 71499 9463 71541 9472
rect 71683 9512 71741 9513
rect 71683 9472 71692 9512
rect 71732 9472 71741 9512
rect 71683 9471 71741 9472
rect 71883 9512 71925 9521
rect 71883 9472 71884 9512
rect 71924 9472 71925 9512
rect 71883 9463 71925 9472
rect 75627 9512 75669 9521
rect 75627 9472 75628 9512
rect 75668 9472 75669 9512
rect 75627 9463 75669 9472
rect 75723 9512 75765 9521
rect 75723 9472 75724 9512
rect 75764 9472 75765 9512
rect 75723 9463 75765 9472
rect 75819 9512 75861 9521
rect 75819 9472 75820 9512
rect 75860 9472 75861 9512
rect 75819 9463 75861 9472
rect 76011 9512 76053 9521
rect 76011 9472 76012 9512
rect 76052 9472 76053 9512
rect 76291 9512 76349 9513
rect 76011 9463 76053 9472
rect 76195 9498 76253 9499
rect 76195 9458 76204 9498
rect 76244 9458 76253 9498
rect 76291 9472 76300 9512
rect 76340 9472 76349 9512
rect 76291 9471 76349 9472
rect 77067 9512 77109 9521
rect 77067 9472 77068 9512
rect 77108 9472 77109 9512
rect 77067 9463 77109 9472
rect 77259 9512 77301 9521
rect 77259 9472 77260 9512
rect 77300 9472 77301 9512
rect 77259 9463 77301 9472
rect 77347 9512 77405 9513
rect 77347 9472 77356 9512
rect 77396 9472 77405 9512
rect 77347 9471 77405 9472
rect 77539 9512 77597 9513
rect 77539 9472 77548 9512
rect 77588 9472 77597 9512
rect 77539 9471 77597 9472
rect 77643 9512 77685 9521
rect 77643 9472 77644 9512
rect 77684 9472 77685 9512
rect 77643 9463 77685 9472
rect 77739 9512 77781 9521
rect 77739 9472 77740 9512
rect 77780 9472 77781 9512
rect 77739 9463 77781 9472
rect 76195 9457 76253 9458
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 57379 9428 57437 9429
rect 57379 9388 57388 9428
rect 57428 9388 57437 9428
rect 57379 9387 57437 9388
rect 59395 9428 59453 9429
rect 59395 9388 59404 9428
rect 59444 9388 59453 9428
rect 59395 9387 59453 9388
rect 70435 9428 70493 9429
rect 70435 9388 70444 9428
rect 70484 9388 70493 9428
rect 70435 9387 70493 9388
rect 76483 9428 76541 9429
rect 76483 9388 76492 9428
rect 76532 9388 76541 9428
rect 76483 9387 76541 9388
rect 4971 9344 5013 9353
rect 4971 9304 4972 9344
rect 5012 9304 5013 9344
rect 4971 9295 5013 9304
rect 5259 9344 5301 9353
rect 5259 9304 5260 9344
rect 5300 9304 5301 9344
rect 5259 9295 5301 9304
rect 39531 9344 39573 9353
rect 39531 9304 39532 9344
rect 39572 9304 39573 9344
rect 39531 9295 39573 9304
rect 41547 9344 41589 9353
rect 41547 9304 41548 9344
rect 41588 9304 41589 9344
rect 41547 9295 41589 9304
rect 42027 9344 42069 9353
rect 42027 9304 42028 9344
rect 42068 9304 42069 9344
rect 42027 9295 42069 9304
rect 44619 9344 44661 9353
rect 44619 9304 44620 9344
rect 44660 9304 44661 9344
rect 44619 9295 44661 9304
rect 47307 9344 47349 9353
rect 47307 9304 47308 9344
rect 47348 9304 47349 9344
rect 47307 9295 47349 9304
rect 50379 9344 50421 9353
rect 50379 9304 50380 9344
rect 50420 9304 50421 9344
rect 50379 9295 50421 9304
rect 54795 9344 54837 9353
rect 54795 9304 54796 9344
rect 54836 9304 54837 9344
rect 54795 9295 54837 9304
rect 56427 9344 56469 9353
rect 56427 9304 56428 9344
rect 56468 9304 56469 9344
rect 56427 9295 56469 9304
rect 69963 9344 70005 9353
rect 69963 9304 69964 9344
rect 70004 9304 70005 9344
rect 69963 9295 70005 9304
rect 72171 9344 72213 9353
rect 72171 9304 72172 9344
rect 72212 9304 72213 9344
rect 72171 9295 72213 9304
rect 73995 9344 74037 9353
rect 73995 9304 73996 9344
rect 74036 9304 74037 9344
rect 73995 9295 74037 9304
rect 76683 9344 76725 9353
rect 76683 9304 76684 9344
rect 76724 9304 76725 9344
rect 76683 9295 76725 9304
rect 3723 9260 3765 9269
rect 3723 9220 3724 9260
rect 3764 9220 3765 9260
rect 3723 9211 3765 9220
rect 42507 9260 42549 9269
rect 42507 9220 42508 9260
rect 42548 9220 42549 9260
rect 42507 9211 42549 9220
rect 44043 9260 44085 9269
rect 44043 9220 44044 9260
rect 44084 9220 44085 9260
rect 44043 9211 44085 9220
rect 46339 9260 46397 9261
rect 46339 9220 46348 9260
rect 46388 9220 46397 9260
rect 46339 9219 46397 9220
rect 53739 9260 53781 9269
rect 53739 9220 53740 9260
rect 53780 9220 53781 9260
rect 53739 9211 53781 9220
rect 54219 9260 54261 9269
rect 54219 9220 54220 9260
rect 54260 9220 54261 9260
rect 54219 9211 54261 9220
rect 57579 9260 57621 9269
rect 57579 9220 57580 9260
rect 57620 9220 57621 9260
rect 57579 9211 57621 9220
rect 57771 9260 57813 9269
rect 57771 9220 57772 9260
rect 57812 9220 57813 9260
rect 57771 9211 57813 9220
rect 59011 9260 59069 9261
rect 59011 9220 59020 9260
rect 59060 9220 59069 9260
rect 59011 9219 59069 9220
rect 59211 9260 59253 9269
rect 59211 9220 59212 9260
rect 59252 9220 59253 9260
rect 59211 9211 59253 9220
rect 64579 9260 64637 9261
rect 64579 9220 64588 9260
rect 64628 9220 64637 9260
rect 64579 9219 64637 9220
rect 69771 9260 69813 9269
rect 69771 9220 69772 9260
rect 69812 9220 69813 9260
rect 69771 9211 69813 9220
rect 70635 9260 70677 9269
rect 70635 9220 70636 9260
rect 70676 9220 70677 9260
rect 70635 9211 70677 9220
rect 71403 9260 71445 9269
rect 71403 9220 71404 9260
rect 71444 9220 71445 9260
rect 71403 9211 71445 9220
rect 71787 9260 71829 9269
rect 71787 9220 71788 9260
rect 71828 9220 71829 9260
rect 71787 9211 71829 9220
rect 76011 9260 76053 9269
rect 76011 9220 76012 9260
rect 76052 9220 76053 9260
rect 76011 9211 76053 9220
rect 576 9092 79584 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79584 9092
rect 576 9028 79584 9052
rect 651 8924 693 8933
rect 651 8884 652 8924
rect 692 8884 693 8924
rect 651 8875 693 8884
rect 3427 8924 3485 8925
rect 3427 8884 3436 8924
rect 3476 8884 3485 8924
rect 3427 8883 3485 8884
rect 43939 8924 43997 8925
rect 43939 8884 43948 8924
rect 43988 8884 43997 8924
rect 43939 8883 43997 8884
rect 46531 8924 46589 8925
rect 46531 8884 46540 8924
rect 46580 8884 46589 8924
rect 46531 8883 46589 8884
rect 53827 8924 53885 8925
rect 53827 8884 53836 8924
rect 53876 8884 53885 8924
rect 53827 8883 53885 8884
rect 56707 8924 56765 8925
rect 56707 8884 56716 8924
rect 56756 8884 56765 8924
rect 56707 8883 56765 8884
rect 59499 8924 59541 8933
rect 59499 8884 59500 8924
rect 59540 8884 59541 8924
rect 59499 8875 59541 8884
rect 68419 8924 68477 8925
rect 68419 8884 68428 8924
rect 68468 8884 68477 8924
rect 68419 8883 68477 8884
rect 69867 8924 69909 8933
rect 69867 8884 69868 8924
rect 69908 8884 69909 8924
rect 69867 8875 69909 8884
rect 71491 8924 71549 8925
rect 71491 8884 71500 8924
rect 71540 8884 71549 8924
rect 71491 8883 71549 8884
rect 74083 8924 74141 8925
rect 74083 8884 74092 8924
rect 74132 8884 74141 8924
rect 74083 8883 74141 8884
rect 75915 8924 75957 8933
rect 75915 8884 75916 8924
rect 75956 8884 75957 8924
rect 75915 8875 75957 8884
rect 79459 8924 79517 8925
rect 79459 8884 79468 8924
rect 79508 8884 79517 8924
rect 79459 8883 79517 8884
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 5259 8840 5301 8849
rect 5259 8800 5260 8840
rect 5300 8800 5301 8840
rect 5259 8791 5301 8800
rect 49323 8840 49365 8849
rect 49323 8800 49324 8840
rect 49364 8800 49365 8840
rect 49323 8791 49365 8800
rect 50955 8840 50997 8849
rect 50955 8800 50956 8840
rect 50996 8800 50997 8840
rect 50955 8791 50997 8800
rect 60075 8840 60117 8849
rect 60075 8800 60076 8840
rect 60116 8800 60117 8840
rect 60075 8791 60117 8800
rect 64971 8840 65013 8849
rect 64971 8800 64972 8840
rect 65012 8800 65013 8840
rect 64971 8791 65013 8800
rect 70155 8840 70197 8849
rect 70155 8800 70156 8840
rect 70196 8800 70197 8840
rect 70155 8791 70197 8800
rect 74283 8840 74325 8849
rect 74283 8800 74284 8840
rect 74324 8800 74325 8840
rect 74283 8791 74325 8800
rect 76867 8840 76925 8841
rect 76867 8800 76876 8840
rect 76916 8800 76925 8840
rect 76867 8799 76925 8800
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 58243 8756 58301 8757
rect 58243 8716 58252 8756
rect 58292 8716 58301 8756
rect 58243 8715 58301 8716
rect 58731 8756 58773 8765
rect 58731 8716 58732 8756
rect 58772 8716 58773 8756
rect 58731 8707 58773 8716
rect 59683 8756 59741 8757
rect 59683 8716 59692 8756
rect 59732 8716 59741 8756
rect 59683 8715 59741 8716
rect 64771 8756 64829 8757
rect 64771 8716 64780 8756
rect 64820 8716 64829 8756
rect 64771 8715 64829 8716
rect 68899 8756 68957 8757
rect 68899 8716 68908 8756
rect 68948 8716 68957 8756
rect 68899 8715 68957 8716
rect 1707 8672 1749 8681
rect 1707 8632 1708 8672
rect 1748 8632 1749 8672
rect 1707 8623 1749 8632
rect 1803 8672 1845 8681
rect 1803 8632 1804 8672
rect 1844 8632 1845 8672
rect 1803 8623 1845 8632
rect 1899 8672 1941 8681
rect 1899 8632 1900 8672
rect 1940 8632 1941 8672
rect 1899 8623 1941 8632
rect 2187 8672 2229 8681
rect 2187 8632 2188 8672
rect 2228 8632 2229 8672
rect 2187 8623 2229 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2467 8672 2525 8673
rect 2467 8632 2476 8672
rect 2516 8632 2525 8672
rect 2467 8631 2525 8632
rect 2755 8672 2813 8673
rect 2755 8632 2764 8672
rect 2804 8632 2813 8672
rect 2755 8631 2813 8632
rect 3051 8672 3093 8681
rect 3051 8632 3052 8672
rect 3092 8632 3093 8672
rect 3051 8623 3093 8632
rect 3147 8672 3189 8681
rect 3147 8632 3148 8672
rect 3188 8632 3189 8672
rect 3147 8623 3189 8632
rect 41923 8672 41981 8673
rect 41923 8632 41932 8672
rect 41972 8632 41981 8672
rect 41923 8631 41981 8632
rect 42787 8672 42845 8673
rect 42787 8632 42796 8672
rect 42836 8632 42845 8672
rect 42787 8631 42845 8632
rect 44515 8672 44573 8673
rect 44515 8632 44524 8672
rect 44564 8632 44573 8672
rect 44515 8631 44573 8632
rect 45379 8672 45437 8673
rect 45379 8632 45388 8672
rect 45428 8632 45437 8672
rect 45379 8631 45437 8632
rect 46731 8672 46773 8681
rect 46731 8632 46732 8672
rect 46772 8632 46773 8672
rect 46731 8623 46773 8632
rect 46915 8672 46973 8673
rect 46915 8632 46924 8672
rect 46964 8632 46973 8672
rect 46915 8631 46973 8632
rect 48451 8672 48509 8673
rect 48451 8632 48460 8672
rect 48500 8632 48509 8672
rect 48451 8631 48509 8632
rect 48651 8672 48693 8681
rect 48651 8632 48652 8672
rect 48692 8632 48693 8672
rect 48651 8623 48693 8632
rect 48843 8672 48885 8681
rect 48843 8632 48844 8672
rect 48884 8632 48885 8672
rect 48843 8623 48885 8632
rect 49035 8672 49077 8681
rect 49035 8632 49036 8672
rect 49076 8632 49077 8672
rect 49035 8623 49077 8632
rect 49123 8672 49181 8673
rect 49123 8632 49132 8672
rect 49172 8632 49181 8672
rect 49123 8631 49181 8632
rect 53155 8672 53213 8673
rect 53155 8632 53164 8672
rect 53204 8632 53213 8672
rect 53155 8631 53213 8632
rect 53451 8672 53493 8681
rect 53451 8632 53452 8672
rect 53492 8632 53493 8672
rect 53451 8623 53493 8632
rect 54691 8672 54749 8673
rect 54691 8632 54700 8672
rect 54740 8632 54749 8672
rect 54691 8631 54749 8632
rect 55555 8672 55613 8673
rect 55555 8632 55564 8672
rect 55604 8632 55613 8672
rect 55555 8631 55613 8632
rect 57771 8672 57813 8681
rect 57771 8632 57772 8672
rect 57812 8632 57813 8672
rect 57771 8623 57813 8632
rect 57867 8672 57909 8681
rect 57867 8632 57868 8672
rect 57908 8632 57909 8672
rect 57867 8623 57909 8632
rect 57963 8672 58005 8681
rect 57963 8632 57964 8672
rect 58004 8632 58005 8672
rect 57963 8623 58005 8632
rect 58059 8672 58101 8681
rect 58059 8632 58060 8672
rect 58100 8632 58101 8672
rect 58059 8623 58101 8632
rect 58627 8672 58685 8673
rect 58627 8632 58636 8672
rect 58676 8632 58685 8672
rect 58627 8631 58685 8632
rect 58827 8672 58869 8681
rect 58827 8632 58828 8672
rect 58868 8632 58869 8672
rect 58827 8623 58869 8632
rect 59019 8672 59061 8681
rect 59019 8632 59020 8672
rect 59060 8632 59061 8672
rect 59019 8623 59061 8632
rect 59211 8672 59253 8681
rect 59211 8632 59212 8672
rect 59252 8632 59253 8672
rect 59211 8623 59253 8632
rect 59299 8672 59357 8673
rect 59299 8632 59308 8672
rect 59348 8632 59357 8672
rect 59299 8631 59357 8632
rect 60451 8672 60509 8673
rect 60451 8632 60460 8672
rect 60500 8632 60509 8672
rect 60451 8631 60509 8632
rect 60651 8672 60693 8681
rect 60651 8632 60652 8672
rect 60692 8632 60693 8672
rect 60651 8623 60693 8632
rect 63819 8672 63861 8681
rect 63819 8632 63820 8672
rect 63860 8632 63861 8672
rect 63819 8623 63861 8632
rect 63915 8672 63957 8681
rect 63915 8632 63916 8672
rect 63956 8632 63957 8672
rect 63915 8623 63957 8632
rect 64011 8672 64053 8681
rect 64011 8632 64012 8672
rect 64052 8632 64053 8672
rect 64011 8623 64053 8632
rect 64107 8672 64149 8681
rect 64107 8632 64108 8672
rect 64148 8632 64149 8672
rect 64107 8623 64149 8632
rect 64299 8672 64341 8681
rect 64299 8632 64300 8672
rect 64340 8632 64341 8672
rect 64299 8623 64341 8632
rect 64491 8672 64533 8681
rect 64491 8632 64492 8672
rect 64532 8632 64533 8672
rect 64491 8623 64533 8632
rect 64579 8672 64637 8673
rect 64579 8632 64588 8672
rect 64628 8632 64637 8672
rect 64579 8631 64637 8632
rect 66403 8672 66461 8673
rect 66403 8632 66412 8672
rect 66452 8632 66461 8672
rect 66403 8631 66461 8632
rect 67267 8672 67325 8673
rect 67267 8632 67276 8672
rect 67316 8632 67325 8672
rect 67267 8631 67325 8632
rect 69291 8672 69333 8681
rect 69291 8632 69292 8672
rect 69332 8632 69333 8672
rect 69291 8623 69333 8632
rect 69483 8672 69525 8681
rect 69483 8632 69484 8672
rect 69524 8632 69525 8672
rect 69483 8623 69525 8632
rect 69571 8672 69629 8673
rect 69571 8632 69580 8672
rect 69620 8632 69629 8672
rect 69571 8631 69629 8632
rect 69763 8672 69821 8673
rect 69763 8632 69772 8672
rect 69812 8632 69821 8672
rect 69763 8631 69821 8632
rect 69963 8672 70005 8681
rect 69963 8632 69964 8672
rect 70004 8632 70005 8672
rect 69963 8623 70005 8632
rect 70819 8672 70877 8673
rect 70819 8632 70828 8672
rect 70868 8632 70877 8672
rect 70819 8631 70877 8632
rect 71115 8672 71157 8681
rect 71115 8632 71116 8672
rect 71156 8632 71157 8672
rect 71115 8623 71157 8632
rect 72067 8672 72125 8673
rect 72067 8632 72076 8672
rect 72116 8632 72125 8672
rect 72067 8631 72125 8632
rect 72931 8672 72989 8673
rect 72931 8632 72940 8672
rect 72980 8632 72989 8672
rect 72931 8631 72989 8632
rect 75619 8672 75677 8673
rect 75619 8632 75628 8672
rect 75668 8632 75677 8672
rect 75619 8631 75677 8632
rect 75723 8672 75765 8681
rect 75723 8632 75724 8672
rect 75764 8632 75765 8672
rect 75723 8623 75765 8632
rect 75915 8672 75957 8681
rect 75915 8632 75916 8672
rect 75956 8632 75957 8672
rect 75915 8623 75957 8632
rect 76195 8672 76253 8673
rect 76195 8632 76204 8672
rect 76244 8632 76253 8672
rect 76195 8631 76253 8632
rect 76491 8672 76533 8681
rect 76491 8632 76492 8672
rect 76532 8632 76533 8672
rect 76491 8623 76533 8632
rect 77443 8672 77501 8673
rect 77443 8632 77452 8672
rect 77492 8632 77501 8672
rect 77443 8631 77501 8632
rect 78307 8672 78365 8673
rect 78307 8632 78316 8672
rect 78356 8632 78365 8672
rect 78307 8631 78365 8632
rect 1995 8588 2037 8597
rect 1995 8548 1996 8588
rect 2036 8548 2037 8588
rect 1995 8539 2037 8548
rect 2283 8588 2325 8597
rect 2283 8548 2284 8588
rect 2324 8548 2325 8588
rect 2283 8539 2325 8548
rect 41547 8588 41589 8597
rect 41547 8548 41548 8588
rect 41588 8548 41589 8588
rect 41547 8539 41589 8548
rect 44139 8588 44181 8597
rect 44139 8548 44140 8588
rect 44180 8548 44181 8588
rect 44139 8539 44181 8548
rect 46827 8588 46869 8597
rect 46827 8548 46828 8588
rect 46868 8548 46869 8588
rect 46827 8539 46869 8548
rect 48555 8588 48597 8597
rect 48555 8548 48556 8588
rect 48596 8548 48597 8588
rect 48555 8539 48597 8548
rect 53547 8588 53589 8597
rect 53547 8548 53548 8588
rect 53588 8548 53589 8588
rect 53547 8539 53589 8548
rect 54315 8588 54357 8597
rect 54315 8548 54316 8588
rect 54356 8548 54357 8588
rect 54315 8539 54357 8548
rect 60555 8588 60597 8597
rect 60555 8548 60556 8588
rect 60596 8548 60597 8588
rect 60555 8539 60597 8548
rect 64395 8588 64437 8597
rect 64395 8548 64396 8588
rect 64436 8548 64437 8588
rect 64395 8539 64437 8548
rect 66027 8588 66069 8597
rect 66027 8548 66028 8588
rect 66068 8548 66069 8588
rect 66027 8539 66069 8548
rect 71211 8588 71253 8597
rect 71211 8548 71212 8588
rect 71252 8548 71253 8588
rect 71211 8539 71253 8548
rect 71691 8588 71733 8597
rect 71691 8548 71692 8588
rect 71732 8548 71733 8588
rect 71691 8539 71733 8548
rect 76587 8588 76629 8597
rect 76587 8548 76588 8588
rect 76628 8548 76629 8588
rect 76587 8539 76629 8548
rect 77067 8588 77109 8597
rect 77067 8548 77068 8588
rect 77108 8548 77109 8588
rect 77067 8539 77109 8548
rect 43939 8504 43997 8505
rect 43939 8464 43948 8504
rect 43988 8464 43997 8504
rect 43939 8463 43997 8464
rect 46531 8504 46589 8505
rect 46531 8464 46540 8504
rect 46580 8464 46589 8504
rect 46531 8463 46589 8464
rect 48931 8504 48989 8505
rect 48931 8464 48940 8504
rect 48980 8464 48989 8504
rect 48931 8463 48989 8464
rect 58443 8504 58485 8513
rect 58443 8464 58444 8504
rect 58484 8464 58485 8504
rect 58443 8455 58485 8464
rect 59107 8504 59165 8505
rect 59107 8464 59116 8504
rect 59156 8464 59165 8504
rect 59107 8463 59165 8464
rect 68419 8504 68477 8505
rect 68419 8464 68428 8504
rect 68468 8464 68477 8504
rect 68419 8463 68477 8464
rect 69099 8504 69141 8513
rect 69099 8464 69100 8504
rect 69140 8464 69141 8504
rect 69099 8455 69141 8464
rect 69379 8504 69437 8505
rect 69379 8464 69388 8504
rect 69428 8464 69437 8504
rect 69379 8463 69437 8464
rect 576 8336 79584 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79584 8336
rect 576 8272 79584 8296
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 4387 8168 4445 8169
rect 4387 8128 4396 8168
rect 4436 8128 4445 8168
rect 4387 8127 4445 8128
rect 7171 8168 7229 8169
rect 7171 8128 7180 8168
rect 7220 8128 7229 8168
rect 7171 8127 7229 8128
rect 44899 8168 44957 8169
rect 44899 8128 44908 8168
rect 44948 8128 44957 8168
rect 44899 8127 44957 8128
rect 52867 8168 52925 8169
rect 52867 8128 52876 8168
rect 52916 8128 52925 8168
rect 52867 8127 52925 8128
rect 62851 8168 62909 8169
rect 62851 8128 62860 8168
rect 62900 8128 62909 8168
rect 62851 8127 62909 8128
rect 64099 8168 64157 8169
rect 64099 8128 64108 8168
rect 64148 8128 64157 8168
rect 64099 8127 64157 8128
rect 65635 8168 65693 8169
rect 65635 8128 65644 8168
rect 65684 8128 65693 8168
rect 65635 8127 65693 8128
rect 70723 8168 70781 8169
rect 70723 8128 70732 8168
rect 70772 8128 70781 8168
rect 70723 8127 70781 8128
rect 71491 8168 71549 8169
rect 71491 8128 71500 8168
rect 71540 8128 71549 8168
rect 71491 8127 71549 8128
rect 77059 8168 77117 8169
rect 77059 8128 77068 8168
rect 77108 8128 77117 8168
rect 77059 8127 77117 8128
rect 4779 8084 4821 8093
rect 4779 8044 4780 8084
rect 4820 8044 4821 8084
rect 4779 8035 4821 8044
rect 54027 8084 54069 8093
rect 54027 8044 54028 8084
rect 54068 8044 54069 8084
rect 54027 8035 54069 8044
rect 55947 8084 55989 8093
rect 55947 8044 55948 8084
rect 55988 8044 55989 8084
rect 55947 8035 55989 8044
rect 68331 8084 68373 8093
rect 68331 8044 68332 8084
rect 68372 8044 68373 8084
rect 68331 8035 68373 8044
rect 73611 8084 73653 8093
rect 73611 8044 73612 8084
rect 73652 8044 73653 8084
rect 73611 8035 73653 8044
rect 76299 8084 76341 8093
rect 76299 8044 76300 8084
rect 76340 8044 76341 8084
rect 76299 8035 76341 8044
rect 48843 8013 48885 8022
rect 1995 8000 2037 8009
rect 1995 7960 1996 8000
rect 2036 7960 2037 8000
rect 1995 7951 2037 7960
rect 2091 8000 2133 8009
rect 2091 7960 2092 8000
rect 2132 7960 2133 8000
rect 2091 7951 2133 7960
rect 2187 8000 2229 8009
rect 2187 7960 2188 8000
rect 2228 7960 2229 8000
rect 2187 7951 2229 7960
rect 2283 8000 2325 8009
rect 2283 7960 2284 8000
rect 2324 7960 2325 8000
rect 2283 7951 2325 7960
rect 2571 8000 2613 8009
rect 2571 7960 2572 8000
rect 2612 7960 2613 8000
rect 2571 7951 2613 7960
rect 2763 8000 2805 8009
rect 2763 7960 2764 8000
rect 2804 7960 2805 8000
rect 2763 7951 2805 7960
rect 2877 8000 2919 8009
rect 2877 7960 2878 8000
rect 2918 7960 2919 8000
rect 2877 7951 2919 7960
rect 3331 8000 3389 8001
rect 3331 7960 3340 8000
rect 3380 7960 3389 8000
rect 3331 7959 3389 7960
rect 3627 8000 3669 8009
rect 3627 7960 3628 8000
rect 3668 7960 3669 8000
rect 3627 7951 3669 7960
rect 3723 8000 3765 8009
rect 3723 7960 3724 8000
rect 3764 7960 3765 8000
rect 3723 7951 3765 7960
rect 4299 8000 4341 8009
rect 4299 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4579 8000 4637 8001
rect 4579 7960 4588 8000
rect 4628 7960 4637 8000
rect 4579 7959 4637 7960
rect 5155 8000 5213 8001
rect 5155 7960 5164 8000
rect 5204 7960 5213 8000
rect 5155 7959 5213 7960
rect 6019 8000 6077 8001
rect 6019 7960 6028 8000
rect 6068 7960 6077 8000
rect 6019 7959 6077 7960
rect 44131 8000 44189 8001
rect 44131 7960 44140 8000
rect 44180 7960 44189 8000
rect 44131 7959 44189 7960
rect 44235 8000 44277 8009
rect 44235 7960 44236 8000
rect 44276 7960 44277 8000
rect 44235 7951 44277 7960
rect 44427 8000 44469 8009
rect 44427 7960 44428 8000
rect 44468 7960 44469 8000
rect 44427 7951 44469 7960
rect 44707 8000 44765 8001
rect 44707 7960 44716 8000
rect 44756 7960 44765 8000
rect 44707 7959 44765 7960
rect 44811 8000 44853 8009
rect 44811 7960 44812 8000
rect 44852 7960 44853 8000
rect 44811 7951 44853 7960
rect 45003 8000 45045 8009
rect 45003 7960 45004 8000
rect 45044 7960 45045 8000
rect 45003 7951 45045 7960
rect 45387 8000 45429 8009
rect 45387 7960 45388 8000
rect 45428 7960 45429 8000
rect 45387 7951 45429 7960
rect 45483 8000 45525 8009
rect 45483 7960 45484 8000
rect 45524 7960 45525 8000
rect 45483 7951 45525 7960
rect 45579 8000 45621 8009
rect 45579 7960 45580 8000
rect 45620 7960 45621 8000
rect 45579 7951 45621 7960
rect 45675 8000 45717 8009
rect 45675 7960 45676 8000
rect 45716 7960 45717 8000
rect 45675 7951 45717 7960
rect 46723 8000 46781 8001
rect 46723 7960 46732 8000
rect 46772 7960 46781 8000
rect 46723 7959 46781 7960
rect 46827 8000 46869 8009
rect 46827 7960 46828 8000
rect 46868 7960 46869 8000
rect 46827 7951 46869 7960
rect 47019 8000 47061 8009
rect 47019 7960 47020 8000
rect 47060 7960 47061 8000
rect 47019 7951 47061 7960
rect 47203 8000 47261 8001
rect 47203 7960 47212 8000
rect 47252 7960 47261 8000
rect 47203 7959 47261 7960
rect 47307 8000 47349 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 47499 8000 47541 8009
rect 47499 7960 47500 8000
rect 47540 7960 47541 8000
rect 47499 7951 47541 7960
rect 47971 8000 48029 8001
rect 47971 7960 47980 8000
rect 48020 7960 48029 8000
rect 47971 7959 48029 7960
rect 48267 8000 48309 8009
rect 48267 7960 48268 8000
rect 48308 7960 48309 8000
rect 48267 7951 48309 7960
rect 48363 8000 48405 8009
rect 48363 7960 48364 8000
rect 48404 7960 48405 8000
rect 48843 7973 48844 8013
rect 48884 7973 48885 8013
rect 53259 8021 53301 8030
rect 48843 7964 48885 7973
rect 49027 8000 49085 8001
rect 48363 7951 48405 7960
rect 49027 7960 49036 8000
rect 49076 7960 49085 8000
rect 49027 7959 49085 7960
rect 49419 8000 49461 8009
rect 49419 7960 49420 8000
rect 49460 7960 49461 8000
rect 49419 7951 49461 7960
rect 50475 8000 50517 8009
rect 50475 7960 50476 8000
rect 50516 7960 50517 8000
rect 50475 7951 50517 7960
rect 50851 8000 50909 8001
rect 50851 7960 50860 8000
rect 50900 7960 50909 8000
rect 50851 7959 50909 7960
rect 51715 8000 51773 8001
rect 51715 7960 51724 8000
rect 51764 7960 51773 8000
rect 51715 7959 51773 7960
rect 53067 8000 53109 8009
rect 53067 7960 53068 8000
rect 53108 7960 53109 8000
rect 53067 7951 53109 7960
rect 53163 8000 53205 8009
rect 53163 7960 53164 8000
rect 53204 7960 53205 8000
rect 53259 7981 53260 8021
rect 53300 7981 53301 8021
rect 53259 7972 53301 7981
rect 53355 8000 53397 8009
rect 53163 7951 53205 7960
rect 53355 7960 53356 8000
rect 53396 7960 53397 8000
rect 53355 7951 53397 7960
rect 53931 8000 53973 8009
rect 53931 7960 53932 8000
rect 53972 7960 53973 8000
rect 53931 7951 53973 7960
rect 54123 8000 54165 8009
rect 54123 7960 54124 8000
rect 54164 7960 54165 8000
rect 54123 7951 54165 7960
rect 54211 8000 54269 8001
rect 54211 7960 54220 8000
rect 54260 7960 54269 8000
rect 54211 7959 54269 7960
rect 56323 8000 56381 8001
rect 56323 7960 56332 8000
rect 56372 7960 56381 8000
rect 56323 7959 56381 7960
rect 57187 8000 57245 8001
rect 57187 7960 57196 8000
rect 57236 7960 57245 8000
rect 57187 7959 57245 7960
rect 58531 8000 58589 8001
rect 58531 7960 58540 8000
rect 58580 7960 58589 8000
rect 58531 7959 58589 7960
rect 58635 8000 58677 8009
rect 58635 7960 58636 8000
rect 58676 7960 58677 8000
rect 58635 7951 58677 7960
rect 58827 8000 58869 8009
rect 58827 7960 58828 8000
rect 58868 7960 58869 8000
rect 58827 7951 58869 7960
rect 60459 8000 60501 8009
rect 60459 7960 60460 8000
rect 60500 7960 60501 8000
rect 60459 7951 60501 7960
rect 60835 8000 60893 8001
rect 60835 7960 60844 8000
rect 60884 7960 60893 8000
rect 60835 7959 60893 7960
rect 61699 8000 61757 8001
rect 61699 7960 61708 8000
rect 61748 7960 61757 8000
rect 61699 7959 61757 7960
rect 63627 8000 63669 8009
rect 63627 7960 63628 8000
rect 63668 7960 63669 8000
rect 63627 7951 63669 7960
rect 63819 8000 63861 8009
rect 63819 7960 63820 8000
rect 63860 7960 63861 8000
rect 63819 7951 63861 7960
rect 63907 8000 63965 8001
rect 63907 7960 63916 8000
rect 63956 7960 63965 8000
rect 63907 7959 63965 7960
rect 64203 8000 64245 8009
rect 64203 7960 64204 8000
rect 64244 7960 64245 8000
rect 64203 7951 64245 7960
rect 64299 8000 64341 8009
rect 64299 7960 64300 8000
rect 64340 7960 64341 8000
rect 64299 7951 64341 7960
rect 64395 8000 64437 8009
rect 64395 7960 64396 8000
rect 64436 7960 64437 8000
rect 64395 7951 64437 7960
rect 64675 8000 64733 8001
rect 64675 7960 64684 8000
rect 64724 7960 64733 8000
rect 64675 7959 64733 7960
rect 64971 8000 65013 8009
rect 64971 7960 64972 8000
rect 65012 7960 65013 8000
rect 64971 7951 65013 7960
rect 65067 8000 65109 8009
rect 65067 7960 65068 8000
rect 65108 7960 65109 8000
rect 65067 7951 65109 7960
rect 65547 8000 65589 8009
rect 65547 7960 65548 8000
rect 65588 7960 65589 8000
rect 65547 7951 65589 7960
rect 65739 8000 65781 8009
rect 65739 7960 65740 8000
rect 65780 7960 65781 8000
rect 65739 7951 65781 7960
rect 65827 8000 65885 8001
rect 65827 7960 65836 8000
rect 65876 7960 65885 8000
rect 65827 7959 65885 7960
rect 66019 8000 66077 8001
rect 66019 7960 66028 8000
rect 66068 7960 66077 8000
rect 66019 7959 66077 7960
rect 66219 8000 66261 8009
rect 66219 7960 66220 8000
rect 66260 7960 66261 8000
rect 66219 7951 66261 7960
rect 68707 8000 68765 8001
rect 68707 7960 68716 8000
rect 68756 7960 68765 8000
rect 68707 7959 68765 7960
rect 69571 8000 69629 8001
rect 69571 7960 69580 8000
rect 69620 7960 69629 8000
rect 69571 7959 69629 7960
rect 71403 8000 71445 8009
rect 71403 7960 71404 8000
rect 71444 7960 71445 8000
rect 71403 7951 71445 7960
rect 71595 8000 71637 8009
rect 71595 7960 71596 8000
rect 71636 7960 71637 8000
rect 71595 7951 71637 7960
rect 71683 8000 71741 8001
rect 71683 7960 71692 8000
rect 71732 7960 71741 8000
rect 71683 7959 71741 7960
rect 73987 8000 74045 8001
rect 73987 7960 73996 8000
rect 74036 7960 74045 8000
rect 73987 7959 74045 7960
rect 74851 8000 74909 8001
rect 74851 7960 74860 8000
rect 74900 7960 74909 8000
rect 74851 7959 74909 7960
rect 76203 8000 76245 8009
rect 76203 7960 76204 8000
rect 76244 7960 76245 8000
rect 76203 7951 76245 7960
rect 76395 8000 76437 8009
rect 76395 7960 76396 8000
rect 76436 7960 76437 8000
rect 76395 7951 76437 7960
rect 76483 8000 76541 8001
rect 76483 7960 76492 8000
rect 76532 7960 76541 8000
rect 76483 7959 76541 7960
rect 76971 8000 77013 8009
rect 76971 7960 76972 8000
rect 77012 7960 77013 8000
rect 76971 7951 77013 7960
rect 77163 8000 77205 8009
rect 77163 7960 77164 8000
rect 77204 7960 77205 8000
rect 77163 7951 77205 7960
rect 77251 8000 77309 8001
rect 77251 7960 77260 8000
rect 77300 7960 77309 8000
rect 77251 7959 77309 7960
rect 77443 8000 77501 8001
rect 77443 7960 77452 8000
rect 77492 7960 77501 8000
rect 77443 7959 77501 7960
rect 77547 8000 77589 8009
rect 77547 7960 77548 8000
rect 77588 7960 77589 8000
rect 77547 7951 77589 7960
rect 77643 8000 77685 8009
rect 77643 7960 77644 8000
rect 77684 7960 77685 8000
rect 77643 7951 77685 7960
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 1699 7916 1757 7917
rect 1699 7876 1708 7916
rect 1748 7876 1757 7916
rect 1699 7875 1757 7876
rect 58347 7916 58389 7925
rect 58347 7876 58348 7916
rect 58388 7876 58389 7916
rect 58347 7867 58389 7876
rect 59875 7916 59933 7917
rect 59875 7876 59884 7916
rect 59924 7876 59933 7916
rect 59875 7875 59933 7876
rect 60259 7916 60317 7917
rect 60259 7876 60268 7916
rect 60308 7876 60317 7916
rect 60259 7875 60317 7876
rect 1323 7832 1365 7841
rect 1323 7792 1324 7832
rect 1364 7792 1365 7832
rect 1323 7783 1365 7792
rect 44427 7832 44469 7841
rect 44427 7792 44428 7832
rect 44468 7792 44469 7832
rect 44427 7783 44469 7792
rect 45963 7832 46005 7841
rect 45963 7792 45964 7832
rect 46004 7792 46005 7832
rect 45963 7783 46005 7792
rect 47019 7832 47061 7841
rect 47019 7792 47020 7832
rect 47060 7792 47061 7832
rect 47019 7783 47061 7792
rect 48643 7832 48701 7833
rect 48643 7792 48652 7832
rect 48692 7792 48701 7832
rect 48643 7791 48701 7792
rect 48939 7832 48981 7841
rect 48939 7792 48940 7832
rect 48980 7792 48981 7832
rect 48939 7783 48981 7792
rect 63051 7832 63093 7841
rect 63051 7792 63052 7832
rect 63092 7792 63093 7832
rect 63051 7783 63093 7792
rect 66123 7832 66165 7841
rect 66123 7792 66124 7832
rect 66164 7792 66165 7832
rect 66123 7783 66165 7792
rect 66507 7832 66549 7841
rect 66507 7792 66508 7832
rect 66548 7792 66549 7832
rect 66507 7783 66549 7792
rect 77835 7832 77877 7841
rect 77835 7792 77836 7832
rect 77876 7792 77877 7832
rect 77835 7783 77877 7792
rect 1515 7748 1557 7757
rect 1515 7708 1516 7748
rect 1556 7708 1557 7748
rect 1515 7699 1557 7708
rect 2571 7748 2613 7757
rect 2571 7708 2572 7748
rect 2612 7708 2613 7748
rect 2571 7699 2613 7708
rect 4003 7748 4061 7749
rect 4003 7708 4012 7748
rect 4052 7708 4061 7748
rect 4003 7707 4061 7708
rect 7171 7748 7229 7749
rect 7171 7708 7180 7748
rect 7220 7708 7229 7748
rect 7171 7707 7229 7708
rect 47499 7748 47541 7757
rect 47499 7708 47500 7748
rect 47540 7708 47541 7748
rect 47499 7699 47541 7708
rect 49611 7748 49653 7757
rect 49611 7708 49612 7748
rect 49652 7708 49653 7748
rect 49611 7699 49653 7708
rect 58827 7748 58869 7757
rect 58827 7708 58828 7748
rect 58868 7708 58869 7748
rect 58827 7699 58869 7708
rect 59691 7748 59733 7757
rect 59691 7708 59692 7748
rect 59732 7708 59733 7748
rect 59691 7699 59733 7708
rect 60075 7748 60117 7757
rect 60075 7708 60076 7748
rect 60116 7708 60117 7748
rect 60075 7699 60117 7708
rect 63627 7748 63669 7757
rect 63627 7708 63628 7748
rect 63668 7708 63669 7748
rect 63627 7699 63669 7708
rect 65347 7748 65405 7749
rect 65347 7708 65356 7748
rect 65396 7708 65405 7748
rect 65347 7707 65405 7708
rect 70723 7748 70781 7749
rect 70723 7708 70732 7748
rect 70772 7708 70781 7748
rect 70723 7707 70781 7708
rect 76003 7748 76061 7749
rect 76003 7708 76012 7748
rect 76052 7708 76061 7748
rect 76003 7707 76061 7708
rect 576 7580 79584 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79584 7580
rect 576 7516 79584 7540
rect 3715 7412 3773 7413
rect 3715 7372 3724 7412
rect 3764 7372 3773 7412
rect 3715 7371 3773 7372
rect 4875 7412 4917 7421
rect 4875 7372 4876 7412
rect 4916 7372 4917 7412
rect 4875 7363 4917 7372
rect 47779 7412 47837 7413
rect 47779 7372 47788 7412
rect 47828 7372 47837 7412
rect 47779 7371 47837 7372
rect 51139 7412 51197 7413
rect 51139 7372 51148 7412
rect 51188 7372 51197 7412
rect 51139 7371 51197 7372
rect 64579 7412 64637 7413
rect 64579 7372 64588 7412
rect 64628 7372 64637 7412
rect 64579 7371 64637 7372
rect 65355 7412 65397 7421
rect 65355 7372 65356 7412
rect 65396 7372 65397 7412
rect 65355 7363 65397 7372
rect 77451 7412 77493 7421
rect 77451 7372 77452 7412
rect 77492 7372 77493 7412
rect 77451 7363 77493 7372
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 51915 7328 51957 7337
rect 51915 7288 51916 7328
rect 51956 7288 51957 7328
rect 51915 7279 51957 7288
rect 55275 7328 55317 7337
rect 55275 7288 55276 7328
rect 55316 7288 55317 7328
rect 55275 7279 55317 7288
rect 61035 7328 61077 7337
rect 61035 7288 61036 7328
rect 61076 7288 61077 7328
rect 61035 7279 61077 7288
rect 69387 7328 69429 7337
rect 69387 7288 69388 7328
rect 69428 7288 69429 7328
rect 69387 7279 69429 7288
rect 72363 7328 72405 7337
rect 72363 7288 72364 7328
rect 72404 7288 72405 7328
rect 72363 7279 72405 7288
rect 77835 7328 77877 7337
rect 77835 7288 77836 7328
rect 77876 7288 77877 7328
rect 77835 7279 77877 7288
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 54883 7244 54941 7245
rect 54883 7204 54892 7244
rect 54932 7204 54941 7244
rect 54883 7203 54941 7204
rect 70339 7179 70397 7180
rect 1699 7160 1757 7161
rect 1699 7120 1708 7160
rect 1748 7120 1757 7160
rect 1699 7119 1757 7120
rect 2563 7160 2621 7161
rect 2563 7120 2572 7160
rect 2612 7120 2621 7160
rect 2563 7119 2621 7120
rect 4011 7160 4053 7169
rect 4011 7120 4012 7160
rect 4052 7120 4053 7160
rect 4011 7111 4053 7120
rect 4195 7160 4253 7161
rect 4195 7120 4204 7160
rect 4244 7120 4253 7160
rect 4195 7119 4253 7120
rect 4771 7160 4829 7161
rect 4771 7120 4780 7160
rect 4820 7120 4829 7160
rect 4771 7119 4829 7120
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4971 7111 5013 7120
rect 45387 7160 45429 7169
rect 45387 7120 45388 7160
rect 45428 7120 45429 7160
rect 45387 7111 45429 7120
rect 45763 7160 45821 7161
rect 45763 7120 45772 7160
rect 45812 7120 45821 7160
rect 45763 7119 45821 7120
rect 46627 7160 46685 7161
rect 46627 7120 46636 7160
rect 46676 7120 46685 7160
rect 46627 7119 46685 7120
rect 48355 7160 48413 7161
rect 48355 7120 48364 7160
rect 48404 7120 48413 7160
rect 48355 7119 48413 7120
rect 48747 7160 48789 7169
rect 48747 7120 48748 7160
rect 48788 7120 48789 7160
rect 48747 7111 48789 7120
rect 49123 7160 49181 7161
rect 49123 7120 49132 7160
rect 49172 7120 49181 7160
rect 49123 7119 49181 7120
rect 49987 7160 50045 7161
rect 49987 7120 49996 7160
rect 50036 7120 50045 7160
rect 49987 7119 50045 7120
rect 52779 7160 52821 7169
rect 52779 7120 52780 7160
rect 52820 7120 52821 7160
rect 52779 7111 52821 7120
rect 52971 7160 53013 7169
rect 52971 7120 52972 7160
rect 53012 7120 53013 7160
rect 52971 7111 53013 7120
rect 53059 7160 53117 7161
rect 53059 7120 53068 7160
rect 53108 7120 53117 7160
rect 53451 7160 53493 7169
rect 53059 7119 53117 7120
rect 53259 7118 53301 7127
rect 1323 7076 1365 7085
rect 1323 7036 1324 7076
rect 1364 7036 1365 7076
rect 1323 7027 1365 7036
rect 4107 7076 4149 7085
rect 4107 7036 4108 7076
rect 4148 7036 4149 7076
rect 4107 7027 4149 7036
rect 52875 7076 52917 7085
rect 52875 7036 52876 7076
rect 52916 7036 52917 7076
rect 53259 7078 53260 7118
rect 53300 7078 53301 7118
rect 53451 7120 53452 7160
rect 53492 7120 53493 7160
rect 53451 7111 53493 7120
rect 53539 7160 53597 7161
rect 53539 7120 53548 7160
rect 53588 7120 53597 7160
rect 53539 7119 53597 7120
rect 54211 7160 54269 7161
rect 54211 7120 54220 7160
rect 54260 7120 54269 7160
rect 54211 7119 54269 7120
rect 54411 7160 54453 7169
rect 54411 7120 54412 7160
rect 54452 7120 54453 7160
rect 54411 7111 54453 7120
rect 57283 7160 57341 7161
rect 57283 7120 57292 7160
rect 57332 7120 57341 7160
rect 57283 7119 57341 7120
rect 58147 7160 58205 7161
rect 58147 7120 58156 7160
rect 58196 7120 58205 7160
rect 58147 7119 58205 7120
rect 59683 7160 59741 7161
rect 59683 7120 59692 7160
rect 59732 7120 59741 7160
rect 59683 7119 59741 7120
rect 59979 7160 60021 7169
rect 59979 7120 59980 7160
rect 60020 7120 60021 7160
rect 59979 7111 60021 7120
rect 60547 7160 60605 7161
rect 60547 7120 60556 7160
rect 60596 7120 60605 7160
rect 60547 7119 60605 7120
rect 60651 7160 60693 7169
rect 60651 7120 60652 7160
rect 60692 7120 60693 7160
rect 60651 7111 60693 7120
rect 60843 7160 60885 7169
rect 60843 7120 60844 7160
rect 60884 7120 60885 7160
rect 60843 7111 60885 7120
rect 62187 7160 62229 7169
rect 62187 7120 62188 7160
rect 62228 7120 62229 7160
rect 62187 7111 62229 7120
rect 62563 7160 62621 7161
rect 62563 7120 62572 7160
rect 62612 7120 62621 7160
rect 62563 7119 62621 7120
rect 63427 7160 63485 7161
rect 63427 7120 63436 7160
rect 63476 7120 63485 7160
rect 63427 7119 63485 7120
rect 64779 7160 64821 7169
rect 64779 7120 64780 7160
rect 64820 7120 64821 7160
rect 64779 7111 64821 7120
rect 64971 7160 65013 7169
rect 64971 7120 64972 7160
rect 65012 7120 65013 7160
rect 64971 7111 65013 7120
rect 65059 7160 65117 7161
rect 65059 7120 65068 7160
rect 65108 7120 65117 7160
rect 65059 7119 65117 7120
rect 65251 7160 65309 7161
rect 65251 7120 65260 7160
rect 65300 7120 65309 7160
rect 65251 7119 65309 7120
rect 65451 7160 65493 7169
rect 65451 7120 65452 7160
rect 65492 7120 65493 7160
rect 65451 7111 65493 7120
rect 66211 7160 66269 7161
rect 66211 7120 66220 7160
rect 66260 7120 66269 7160
rect 66211 7119 66269 7120
rect 66411 7160 66453 7169
rect 66411 7120 66412 7160
rect 66452 7120 66453 7160
rect 66411 7111 66453 7120
rect 66691 7160 66749 7161
rect 66691 7120 66700 7160
rect 66740 7120 66749 7160
rect 66691 7119 66749 7120
rect 66891 7160 66933 7169
rect 66891 7120 66892 7160
rect 66932 7120 66933 7160
rect 66891 7111 66933 7120
rect 69675 7160 69717 7169
rect 69675 7120 69676 7160
rect 69716 7120 69717 7160
rect 69675 7111 69717 7120
rect 69771 7160 69813 7169
rect 69771 7120 69772 7160
rect 69812 7120 69813 7160
rect 69771 7111 69813 7120
rect 69867 7160 69909 7169
rect 69867 7120 69868 7160
rect 69908 7120 69909 7160
rect 69867 7111 69909 7120
rect 70059 7160 70101 7169
rect 70059 7120 70060 7160
rect 70100 7120 70101 7160
rect 70059 7111 70101 7120
rect 70251 7160 70293 7169
rect 70251 7120 70252 7160
rect 70292 7120 70293 7160
rect 70339 7139 70348 7179
rect 70388 7139 70397 7179
rect 70339 7138 70397 7139
rect 71211 7160 71253 7169
rect 70251 7111 70293 7120
rect 71211 7120 71212 7160
rect 71252 7120 71253 7160
rect 71211 7111 71253 7120
rect 71395 7160 71453 7161
rect 71395 7120 71404 7160
rect 71444 7120 71453 7160
rect 71395 7119 71453 7120
rect 71595 7160 71637 7169
rect 71595 7120 71596 7160
rect 71636 7120 71637 7160
rect 71595 7111 71637 7120
rect 71787 7160 71829 7169
rect 71787 7120 71788 7160
rect 71828 7120 71829 7160
rect 71787 7111 71829 7120
rect 71875 7160 71933 7161
rect 71875 7120 71884 7160
rect 71924 7120 71933 7160
rect 71875 7119 71933 7120
rect 75435 7160 75477 7169
rect 75435 7120 75436 7160
rect 75476 7120 75477 7160
rect 75435 7111 75477 7120
rect 75531 7160 75573 7169
rect 75531 7120 75532 7160
rect 75572 7120 75573 7160
rect 75531 7111 75573 7120
rect 75627 7160 75669 7169
rect 75627 7120 75628 7160
rect 75668 7120 75669 7160
rect 75627 7111 75669 7120
rect 75723 7160 75765 7169
rect 75723 7120 75724 7160
rect 75764 7120 75765 7160
rect 75723 7111 75765 7120
rect 75915 7160 75957 7169
rect 75915 7120 75916 7160
rect 75956 7120 75957 7160
rect 75915 7111 75957 7120
rect 76107 7160 76149 7169
rect 76107 7120 76108 7160
rect 76148 7120 76149 7160
rect 76107 7111 76149 7120
rect 76195 7160 76253 7161
rect 76195 7120 76204 7160
rect 76244 7120 76253 7160
rect 76195 7119 76253 7120
rect 76875 7160 76917 7169
rect 76875 7120 76876 7160
rect 76916 7120 76917 7160
rect 76875 7111 76917 7120
rect 77059 7160 77117 7161
rect 77059 7120 77068 7160
rect 77108 7120 77117 7160
rect 77059 7119 77117 7120
rect 77347 7160 77405 7161
rect 77347 7120 77356 7160
rect 77396 7120 77405 7160
rect 77347 7119 77405 7120
rect 77547 7160 77589 7169
rect 77547 7120 77548 7160
rect 77588 7120 77589 7160
rect 77547 7111 77589 7120
rect 53259 7069 53301 7078
rect 53355 7076 53397 7085
rect 52875 7027 52917 7036
rect 53355 7036 53356 7076
rect 53396 7036 53397 7076
rect 53355 7027 53397 7036
rect 54315 7076 54357 7085
rect 54315 7036 54316 7076
rect 54356 7036 54357 7076
rect 54315 7027 54357 7036
rect 56907 7076 56949 7085
rect 56907 7036 56908 7076
rect 56948 7036 56949 7076
rect 56907 7027 56949 7036
rect 60075 7076 60117 7085
rect 60075 7036 60076 7076
rect 60116 7036 60117 7076
rect 60075 7027 60117 7036
rect 64875 7076 64917 7085
rect 64875 7036 64876 7076
rect 64916 7036 64917 7076
rect 64875 7027 64917 7036
rect 66315 7076 66357 7085
rect 66315 7036 66316 7076
rect 66356 7036 66357 7076
rect 66315 7027 66357 7036
rect 66795 7076 66837 7085
rect 66795 7036 66796 7076
rect 66836 7036 66837 7076
rect 66795 7027 66837 7036
rect 71307 7076 71349 7085
rect 71307 7036 71308 7076
rect 71348 7036 71349 7076
rect 71307 7027 71349 7036
rect 76011 7076 76053 7085
rect 76011 7036 76012 7076
rect 76052 7036 76053 7076
rect 76011 7027 76053 7036
rect 76971 7076 77013 7085
rect 76971 7036 76972 7076
rect 77012 7036 77013 7076
rect 76971 7027 77013 7036
rect 55083 6992 55125 7001
rect 55083 6952 55084 6992
rect 55124 6952 55125 6992
rect 55083 6943 55125 6952
rect 59299 6992 59357 6993
rect 59299 6952 59308 6992
rect 59348 6952 59357 6992
rect 60739 6992 60797 6993
rect 59299 6951 59357 6952
rect 60363 6950 60405 6959
rect 60739 6952 60748 6992
rect 60788 6952 60797 6992
rect 60739 6951 60797 6952
rect 69571 6992 69629 6993
rect 69571 6952 69580 6992
rect 69620 6952 69629 6992
rect 69571 6951 69629 6952
rect 70147 6992 70205 6993
rect 70147 6952 70156 6992
rect 70196 6952 70205 6992
rect 70147 6951 70205 6952
rect 71683 6992 71741 6993
rect 71683 6952 71692 6992
rect 71732 6952 71741 6992
rect 71683 6951 71741 6952
rect 60363 6910 60364 6950
rect 60404 6910 60405 6950
rect 60363 6901 60405 6910
rect 576 6824 79584 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79584 6824
rect 576 6760 79584 6784
rect 47203 6656 47261 6657
rect 47203 6616 47212 6656
rect 47252 6616 47261 6656
rect 47203 6615 47261 6616
rect 56995 6656 57053 6657
rect 56995 6616 57004 6656
rect 57044 6616 57053 6656
rect 56995 6615 57053 6616
rect 69091 6656 69149 6657
rect 69091 6616 69100 6656
rect 69140 6616 69149 6656
rect 69091 6615 69149 6616
rect 74275 6656 74333 6657
rect 74275 6616 74284 6656
rect 74324 6616 74333 6656
rect 74275 6615 74333 6616
rect 54219 6572 54261 6581
rect 2859 6530 2901 6539
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2467 6488 2525 6489
rect 2467 6448 2476 6488
rect 2516 6448 2525 6488
rect 2467 6447 2525 6448
rect 2667 6488 2709 6497
rect 2667 6448 2668 6488
rect 2708 6448 2709 6488
rect 2859 6490 2860 6530
rect 2900 6490 2901 6530
rect 54219 6532 54220 6572
rect 54260 6532 54261 6572
rect 54219 6523 54261 6532
rect 54603 6572 54645 6581
rect 54603 6532 54604 6572
rect 54644 6532 54645 6572
rect 54603 6523 54645 6532
rect 58539 6572 58581 6581
rect 58539 6532 58540 6572
rect 58580 6532 58581 6572
rect 58539 6523 58581 6532
rect 66123 6572 66165 6581
rect 66123 6532 66124 6572
rect 66164 6532 66165 6572
rect 66123 6523 66165 6532
rect 71883 6572 71925 6581
rect 71883 6532 71884 6572
rect 71924 6532 71925 6572
rect 71883 6523 71925 6532
rect 2859 6481 2901 6490
rect 2947 6488 3005 6489
rect 2667 6439 2709 6448
rect 2947 6448 2956 6488
rect 2996 6448 3005 6488
rect 2947 6447 3005 6448
rect 4107 6488 4149 6497
rect 4107 6448 4108 6488
rect 4148 6448 4149 6488
rect 4107 6439 4149 6448
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 4483 6488 4541 6489
rect 4483 6448 4492 6488
rect 4532 6448 4541 6488
rect 4483 6447 4541 6448
rect 4867 6488 4925 6489
rect 4867 6448 4876 6488
rect 4916 6448 4925 6488
rect 4867 6447 4925 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 47307 6488 47349 6497
rect 47307 6448 47308 6488
rect 47348 6448 47349 6488
rect 47307 6439 47349 6448
rect 47403 6488 47445 6497
rect 47403 6448 47404 6488
rect 47444 6448 47445 6488
rect 47403 6439 47445 6448
rect 47499 6488 47541 6497
rect 47499 6448 47500 6488
rect 47540 6448 47541 6488
rect 47499 6439 47541 6448
rect 47691 6488 47733 6497
rect 47691 6448 47692 6488
rect 47732 6448 47733 6488
rect 47691 6439 47733 6448
rect 47883 6488 47925 6497
rect 47883 6448 47884 6488
rect 47924 6448 47925 6488
rect 47883 6439 47925 6448
rect 47971 6488 48029 6489
rect 47971 6448 47980 6488
rect 48020 6448 48029 6488
rect 47971 6447 48029 6448
rect 48843 6488 48885 6497
rect 48843 6448 48844 6488
rect 48884 6448 48885 6488
rect 48843 6439 48885 6448
rect 49219 6488 49277 6489
rect 49219 6448 49228 6488
rect 49268 6448 49277 6488
rect 49219 6447 49277 6448
rect 50083 6488 50141 6489
rect 50083 6448 50092 6488
rect 50132 6448 50141 6488
rect 50083 6447 50141 6448
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51811 6488 51869 6489
rect 51811 6448 51820 6488
rect 51860 6448 51869 6488
rect 51811 6447 51869 6448
rect 52675 6488 52733 6489
rect 52675 6448 52684 6488
rect 52724 6448 52733 6488
rect 52675 6447 52733 6448
rect 54123 6488 54165 6497
rect 54123 6448 54124 6488
rect 54164 6448 54165 6488
rect 54123 6439 54165 6448
rect 54315 6488 54357 6497
rect 54315 6448 54316 6488
rect 54356 6448 54357 6488
rect 54315 6439 54357 6448
rect 54403 6488 54461 6489
rect 54403 6448 54412 6488
rect 54452 6448 54461 6488
rect 54403 6447 54461 6448
rect 54979 6488 55037 6489
rect 54979 6448 54988 6488
rect 55028 6448 55037 6488
rect 54979 6447 55037 6448
rect 55843 6488 55901 6489
rect 55843 6448 55852 6488
rect 55892 6448 55901 6488
rect 55843 6447 55901 6448
rect 58059 6488 58101 6497
rect 58059 6448 58060 6488
rect 58100 6448 58101 6488
rect 58059 6439 58101 6448
rect 58251 6488 58293 6497
rect 58251 6448 58252 6488
rect 58292 6448 58293 6488
rect 58251 6439 58293 6448
rect 58339 6488 58397 6489
rect 58339 6448 58348 6488
rect 58388 6448 58397 6488
rect 58339 6447 58397 6448
rect 58635 6488 58677 6497
rect 58635 6448 58636 6488
rect 58676 6448 58677 6488
rect 58635 6439 58677 6448
rect 58731 6488 58773 6497
rect 58731 6448 58732 6488
rect 58772 6448 58773 6488
rect 58731 6439 58773 6448
rect 58827 6488 58869 6497
rect 58827 6448 58828 6488
rect 58868 6448 58869 6488
rect 58827 6439 58869 6448
rect 59203 6488 59261 6489
rect 59203 6448 59212 6488
rect 59252 6448 59261 6488
rect 59203 6447 59261 6448
rect 59307 6488 59349 6497
rect 59307 6448 59308 6488
rect 59348 6448 59349 6488
rect 59307 6439 59349 6448
rect 59499 6488 59541 6497
rect 59499 6448 59500 6488
rect 59540 6448 59541 6488
rect 59499 6439 59541 6448
rect 60163 6488 60221 6489
rect 60163 6448 60172 6488
rect 60212 6448 60221 6488
rect 60163 6447 60221 6448
rect 60363 6488 60405 6497
rect 60363 6448 60364 6488
rect 60404 6448 60405 6488
rect 60363 6439 60405 6448
rect 61411 6488 61469 6489
rect 61411 6448 61420 6488
rect 61460 6448 61469 6488
rect 61411 6447 61469 6448
rect 61611 6488 61653 6497
rect 61611 6448 61612 6488
rect 61652 6448 61653 6488
rect 61611 6439 61653 6448
rect 65731 6488 65789 6489
rect 65731 6448 65740 6488
rect 65780 6448 65789 6488
rect 65731 6447 65789 6448
rect 66027 6488 66069 6497
rect 66027 6448 66028 6488
rect 66068 6448 66069 6488
rect 66027 6439 66069 6448
rect 66699 6488 66741 6497
rect 66699 6448 66700 6488
rect 66740 6448 66741 6488
rect 66699 6439 66741 6448
rect 67075 6488 67133 6489
rect 67075 6448 67084 6488
rect 67124 6448 67133 6488
rect 67075 6447 67133 6448
rect 67939 6488 67997 6489
rect 67939 6448 67948 6488
rect 67988 6448 67997 6488
rect 67939 6447 67997 6448
rect 69291 6488 69333 6497
rect 69291 6448 69292 6488
rect 69332 6448 69333 6488
rect 69291 6439 69333 6448
rect 69667 6488 69725 6489
rect 69667 6448 69676 6488
rect 69716 6448 69725 6488
rect 69667 6447 69725 6448
rect 70531 6488 70589 6489
rect 70531 6448 70540 6488
rect 70580 6448 70589 6488
rect 70531 6447 70589 6448
rect 72259 6488 72317 6489
rect 72259 6448 72268 6488
rect 72308 6448 72317 6488
rect 72259 6447 72317 6448
rect 73123 6488 73181 6489
rect 73123 6448 73132 6488
rect 73172 6448 73181 6488
rect 73123 6447 73181 6448
rect 75627 6488 75669 6497
rect 75627 6448 75628 6488
rect 75668 6448 75669 6488
rect 75627 6439 75669 6448
rect 75723 6488 75765 6497
rect 75723 6448 75724 6488
rect 75764 6448 75765 6488
rect 75723 6439 75765 6448
rect 75819 6488 75861 6497
rect 75819 6448 75820 6488
rect 75860 6448 75861 6488
rect 76195 6488 76253 6489
rect 75819 6439 75861 6448
rect 75915 6451 75957 6460
rect 75915 6411 75916 6451
rect 75956 6411 75957 6451
rect 76195 6448 76204 6488
rect 76244 6448 76253 6488
rect 76195 6447 76253 6448
rect 76491 6488 76533 6497
rect 76491 6448 76492 6488
rect 76532 6448 76533 6488
rect 76491 6439 76533 6448
rect 76587 6488 76629 6497
rect 76587 6448 76588 6488
rect 76628 6448 76629 6488
rect 76587 6439 76629 6448
rect 77067 6488 77109 6497
rect 77067 6448 77068 6488
rect 77108 6448 77109 6488
rect 77067 6439 77109 6448
rect 77443 6488 77501 6489
rect 77443 6448 77452 6488
rect 77492 6448 77501 6488
rect 77443 6447 77501 6448
rect 78307 6488 78365 6489
rect 78307 6448 78316 6488
rect 78356 6448 78365 6488
rect 78307 6447 78365 6448
rect 835 6404 893 6405
rect 835 6364 844 6404
rect 884 6364 893 6404
rect 75915 6402 75957 6411
rect 835 6363 893 6364
rect 651 6320 693 6329
rect 651 6280 652 6320
rect 692 6280 693 6320
rect 651 6271 693 6280
rect 1707 6320 1749 6329
rect 1707 6280 1708 6320
rect 1748 6280 1749 6320
rect 1707 6271 1749 6280
rect 2187 6320 2229 6329
rect 2187 6280 2188 6320
rect 2228 6280 2229 6320
rect 2187 6271 2229 6280
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 5451 6320 5493 6329
rect 5451 6280 5452 6320
rect 5492 6280 5493 6320
rect 5451 6271 5493 6280
rect 57387 6320 57429 6329
rect 57387 6280 57388 6320
rect 57428 6280 57429 6320
rect 57387 6271 57429 6280
rect 58059 6320 58101 6329
rect 58059 6280 58060 6320
rect 58100 6280 58101 6320
rect 58059 6271 58101 6280
rect 60267 6320 60309 6329
rect 60267 6280 60268 6320
rect 60308 6280 60309 6320
rect 60267 6271 60309 6280
rect 63627 6320 63669 6329
rect 63627 6280 63628 6320
rect 63668 6280 63669 6320
rect 63627 6271 63669 6280
rect 66403 6320 66461 6321
rect 66403 6280 66412 6320
rect 66452 6280 66461 6320
rect 66403 6279 66461 6280
rect 74475 6320 74517 6329
rect 74475 6280 74476 6320
rect 74516 6280 74517 6320
rect 74475 6271 74517 6280
rect 76867 6320 76925 6321
rect 76867 6280 76876 6320
rect 76916 6280 76925 6320
rect 76867 6279 76925 6280
rect 3811 6236 3869 6237
rect 3811 6196 3820 6236
rect 3860 6196 3869 6236
rect 3811 6195 3869 6196
rect 4971 6236 5013 6245
rect 4971 6196 4972 6236
rect 5012 6196 5013 6236
rect 4971 6187 5013 6196
rect 47691 6236 47733 6245
rect 47691 6196 47692 6236
rect 47732 6196 47733 6236
rect 47691 6187 47733 6196
rect 51235 6236 51293 6237
rect 51235 6196 51244 6236
rect 51284 6196 51293 6236
rect 51235 6195 51293 6196
rect 53827 6236 53885 6237
rect 53827 6196 53836 6236
rect 53876 6196 53885 6236
rect 53827 6195 53885 6196
rect 56995 6236 57053 6237
rect 56995 6196 57004 6236
rect 57044 6196 57053 6236
rect 56995 6195 57053 6196
rect 59499 6236 59541 6245
rect 59499 6196 59500 6236
rect 59540 6196 59541 6236
rect 59499 6187 59541 6196
rect 61515 6236 61557 6245
rect 61515 6196 61516 6236
rect 61556 6196 61557 6236
rect 61515 6187 61557 6196
rect 71683 6236 71741 6237
rect 71683 6196 71692 6236
rect 71732 6196 71741 6236
rect 71683 6195 71741 6196
rect 74275 6236 74333 6237
rect 74275 6196 74284 6236
rect 74324 6196 74333 6236
rect 74275 6195 74333 6196
rect 79459 6236 79517 6237
rect 79459 6196 79468 6236
rect 79508 6196 79517 6236
rect 79459 6195 79517 6196
rect 576 6068 79584 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79584 6068
rect 576 6004 79584 6028
rect 7363 5900 7421 5901
rect 7363 5860 7372 5900
rect 7412 5860 7421 5900
rect 7363 5859 7421 5860
rect 49035 5900 49077 5909
rect 49035 5860 49036 5900
rect 49076 5860 49077 5900
rect 49035 5851 49077 5860
rect 54499 5900 54557 5901
rect 54499 5860 54508 5900
rect 54548 5860 54557 5900
rect 54499 5859 54557 5860
rect 66411 5900 66453 5909
rect 66411 5860 66412 5900
rect 66452 5860 66453 5900
rect 66411 5851 66453 5860
rect 69771 5900 69813 5909
rect 69771 5860 69772 5900
rect 69812 5860 69813 5900
rect 69771 5851 69813 5860
rect 71107 5900 71165 5901
rect 71107 5860 71116 5900
rect 71156 5860 71165 5900
rect 71107 5859 71165 5860
rect 76003 5900 76061 5901
rect 76003 5860 76012 5900
rect 76052 5860 76061 5900
rect 76003 5859 76061 5860
rect 77067 5900 77109 5909
rect 77067 5860 77068 5900
rect 77108 5860 77109 5900
rect 77067 5851 77109 5860
rect 46347 5816 46389 5825
rect 46347 5776 46348 5816
rect 46388 5776 46389 5816
rect 46347 5767 46389 5776
rect 48835 5816 48893 5817
rect 48835 5776 48844 5816
rect 48884 5776 48893 5816
rect 48835 5775 48893 5776
rect 49515 5816 49557 5825
rect 49515 5776 49516 5816
rect 49556 5776 49557 5816
rect 49515 5767 49557 5776
rect 56619 5816 56661 5825
rect 56619 5776 56620 5816
rect 56660 5776 56661 5816
rect 56619 5767 56661 5776
rect 59691 5816 59733 5825
rect 59691 5776 59692 5816
rect 59732 5776 59733 5816
rect 59691 5767 59733 5776
rect 67179 5816 67221 5825
rect 67179 5776 67180 5816
rect 67220 5776 67221 5816
rect 67179 5767 67221 5776
rect 1027 5732 1085 5733
rect 1027 5692 1036 5732
rect 1076 5692 1085 5732
rect 1027 5691 1085 5692
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 54795 5732 54837 5741
rect 54795 5692 54796 5732
rect 54836 5692 54837 5732
rect 54795 5683 54837 5692
rect 63723 5732 63765 5741
rect 63723 5692 63724 5732
rect 63764 5692 63765 5732
rect 63723 5683 63765 5692
rect 72171 5732 72213 5741
rect 72171 5692 72172 5732
rect 72212 5692 72213 5732
rect 72171 5683 72213 5692
rect 1603 5648 1661 5649
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1603 5607 1661 5608
rect 2467 5648 2525 5649
rect 2467 5608 2476 5648
rect 2516 5608 2525 5648
rect 2467 5607 2525 5608
rect 4099 5648 4157 5649
rect 4099 5608 4108 5648
rect 4148 5608 4157 5648
rect 4099 5607 4157 5608
rect 5347 5648 5405 5649
rect 5347 5608 5356 5648
rect 5396 5608 5405 5648
rect 5347 5607 5405 5608
rect 6211 5648 6269 5649
rect 6211 5608 6220 5648
rect 6260 5608 6269 5648
rect 6211 5607 6269 5608
rect 47211 5648 47253 5657
rect 47211 5608 47212 5648
rect 47252 5608 47253 5648
rect 47211 5599 47253 5608
rect 47403 5648 47445 5657
rect 47403 5608 47404 5648
rect 47444 5608 47445 5648
rect 47403 5599 47445 5608
rect 47491 5648 47549 5649
rect 47491 5608 47500 5648
rect 47540 5608 47549 5648
rect 47491 5607 47549 5608
rect 48163 5648 48221 5649
rect 48163 5608 48172 5648
rect 48212 5608 48221 5648
rect 48163 5607 48221 5608
rect 48459 5648 48501 5657
rect 48459 5608 48460 5648
rect 48500 5608 48501 5648
rect 48459 5599 48501 5608
rect 49035 5648 49077 5657
rect 49035 5608 49036 5648
rect 49076 5608 49077 5648
rect 49035 5599 49077 5608
rect 49227 5648 49269 5657
rect 49227 5608 49228 5648
rect 49268 5608 49269 5648
rect 49227 5599 49269 5608
rect 49315 5648 49373 5649
rect 49315 5608 49324 5648
rect 49364 5608 49373 5648
rect 49315 5607 49373 5608
rect 49891 5648 49949 5649
rect 49891 5608 49900 5648
rect 49940 5608 49949 5648
rect 49891 5607 49949 5608
rect 50091 5648 50133 5657
rect 50091 5608 50092 5648
rect 50132 5608 50133 5648
rect 50091 5599 50133 5608
rect 52291 5648 52349 5649
rect 52291 5608 52300 5648
rect 52340 5608 52349 5648
rect 52291 5607 52349 5608
rect 52395 5648 52437 5657
rect 52395 5608 52396 5648
rect 52436 5608 52437 5648
rect 52395 5599 52437 5608
rect 52587 5648 52629 5657
rect 52587 5608 52588 5648
rect 52628 5608 52629 5648
rect 52587 5599 52629 5608
rect 52779 5648 52821 5657
rect 52779 5608 52780 5648
rect 52820 5608 52821 5648
rect 52779 5599 52821 5608
rect 52875 5648 52917 5657
rect 52875 5608 52876 5648
rect 52916 5608 52917 5648
rect 52875 5599 52917 5608
rect 52971 5648 53013 5657
rect 52971 5608 52972 5648
rect 53012 5608 53013 5648
rect 52971 5599 53013 5608
rect 53067 5648 53109 5657
rect 53067 5608 53068 5648
rect 53108 5608 53109 5648
rect 53067 5599 53109 5608
rect 53827 5648 53885 5649
rect 53827 5608 53836 5648
rect 53876 5608 53885 5648
rect 53827 5607 53885 5608
rect 54123 5648 54165 5657
rect 54123 5608 54124 5648
rect 54164 5608 54165 5648
rect 54123 5599 54165 5608
rect 54219 5648 54261 5657
rect 54219 5608 54220 5648
rect 54260 5608 54261 5648
rect 54219 5599 54261 5608
rect 54699 5648 54741 5657
rect 54699 5608 54700 5648
rect 54740 5608 54741 5648
rect 54699 5599 54741 5608
rect 54883 5648 54941 5649
rect 54883 5608 54892 5648
rect 54932 5608 54941 5648
rect 54883 5607 54941 5608
rect 56227 5648 56285 5649
rect 56227 5608 56236 5648
rect 56276 5608 56285 5648
rect 56227 5607 56285 5608
rect 56427 5648 56469 5657
rect 56427 5608 56428 5648
rect 56468 5608 56469 5648
rect 56427 5599 56469 5608
rect 59211 5648 59253 5657
rect 59211 5608 59212 5648
rect 59252 5608 59253 5648
rect 59211 5599 59253 5608
rect 59403 5648 59445 5657
rect 59403 5608 59404 5648
rect 59444 5608 59445 5648
rect 59403 5599 59445 5608
rect 59491 5648 59549 5649
rect 59491 5608 59500 5648
rect 59540 5608 59549 5648
rect 59491 5607 59549 5608
rect 60843 5648 60885 5657
rect 60843 5608 60844 5648
rect 60884 5608 60885 5648
rect 60843 5599 60885 5608
rect 61035 5648 61077 5657
rect 61035 5608 61036 5648
rect 61076 5608 61077 5648
rect 61035 5599 61077 5608
rect 61123 5648 61181 5649
rect 61123 5608 61132 5648
rect 61172 5608 61181 5648
rect 61123 5607 61181 5608
rect 61699 5648 61757 5649
rect 61699 5608 61708 5648
rect 61748 5608 61757 5648
rect 61699 5607 61757 5608
rect 62563 5648 62621 5649
rect 62563 5608 62572 5648
rect 62612 5608 62621 5648
rect 62563 5607 62621 5608
rect 64587 5648 64629 5657
rect 64587 5608 64588 5648
rect 64628 5608 64629 5648
rect 64587 5599 64629 5608
rect 64779 5648 64821 5657
rect 64779 5608 64780 5648
rect 64820 5608 64821 5648
rect 64779 5599 64821 5608
rect 64867 5648 64925 5649
rect 64867 5608 64876 5648
rect 64916 5608 64925 5648
rect 64867 5607 64925 5608
rect 65067 5648 65109 5657
rect 65067 5608 65068 5648
rect 65108 5608 65109 5648
rect 65067 5599 65109 5608
rect 65163 5648 65205 5657
rect 65163 5608 65164 5648
rect 65204 5608 65205 5648
rect 65163 5599 65205 5608
rect 65259 5648 65301 5657
rect 65259 5608 65260 5648
rect 65300 5608 65301 5648
rect 65259 5599 65301 5608
rect 65355 5648 65397 5657
rect 65355 5608 65356 5648
rect 65396 5608 65397 5648
rect 65355 5599 65397 5608
rect 66411 5648 66453 5657
rect 66411 5608 66412 5648
rect 66452 5608 66453 5648
rect 66411 5599 66453 5608
rect 66603 5648 66645 5657
rect 66603 5608 66604 5648
rect 66644 5608 66645 5648
rect 66603 5599 66645 5608
rect 66691 5648 66749 5649
rect 66691 5608 66700 5648
rect 66740 5608 66749 5648
rect 66691 5607 66749 5608
rect 69291 5648 69333 5657
rect 69291 5608 69292 5648
rect 69332 5608 69333 5648
rect 69291 5599 69333 5608
rect 69387 5648 69429 5657
rect 69387 5608 69388 5648
rect 69428 5608 69429 5648
rect 69387 5599 69429 5608
rect 69483 5648 69525 5657
rect 69483 5608 69484 5648
rect 69524 5608 69525 5648
rect 69483 5599 69525 5608
rect 69579 5648 69621 5657
rect 69579 5608 69580 5648
rect 69620 5608 69621 5648
rect 69579 5599 69621 5608
rect 69771 5648 69813 5657
rect 69771 5608 69772 5648
rect 69812 5608 69813 5648
rect 69771 5599 69813 5608
rect 69963 5648 70005 5657
rect 69963 5608 69964 5648
rect 70004 5608 70005 5648
rect 69963 5599 70005 5608
rect 70051 5648 70109 5649
rect 70051 5608 70060 5648
rect 70100 5608 70109 5648
rect 70051 5607 70109 5608
rect 71403 5648 71445 5657
rect 71403 5608 71404 5648
rect 71444 5608 71445 5648
rect 71403 5599 71445 5608
rect 71499 5648 71541 5657
rect 71499 5608 71500 5648
rect 71540 5608 71541 5648
rect 71499 5599 71541 5608
rect 71779 5648 71837 5649
rect 71779 5608 71788 5648
rect 71828 5608 71837 5648
rect 71779 5607 71837 5608
rect 72067 5648 72125 5649
rect 72067 5608 72076 5648
rect 72116 5608 72125 5648
rect 72067 5607 72125 5608
rect 72267 5648 72309 5657
rect 72267 5608 72268 5648
rect 72308 5608 72309 5648
rect 72267 5599 72309 5608
rect 73987 5648 74045 5649
rect 73987 5608 73996 5648
rect 74036 5608 74045 5648
rect 73987 5607 74045 5608
rect 74851 5648 74909 5649
rect 74851 5608 74860 5648
rect 74900 5608 74909 5648
rect 74851 5607 74909 5608
rect 76203 5648 76245 5657
rect 76203 5608 76204 5648
rect 76244 5608 76245 5648
rect 76203 5599 76245 5608
rect 76395 5648 76437 5657
rect 76395 5608 76396 5648
rect 76436 5608 76437 5648
rect 76395 5599 76437 5608
rect 76483 5648 76541 5649
rect 76483 5608 76492 5648
rect 76532 5608 76541 5648
rect 76483 5607 76541 5608
rect 77067 5648 77109 5657
rect 77067 5608 77068 5648
rect 77108 5608 77109 5648
rect 77067 5599 77109 5608
rect 77259 5648 77301 5657
rect 77259 5608 77260 5648
rect 77300 5608 77301 5648
rect 77259 5599 77301 5608
rect 77347 5648 77405 5649
rect 77347 5608 77356 5648
rect 77396 5608 77405 5648
rect 77347 5607 77405 5608
rect 77539 5648 77597 5649
rect 77539 5608 77548 5648
rect 77588 5608 77597 5648
rect 77539 5607 77597 5608
rect 77739 5648 77781 5657
rect 77739 5608 77740 5648
rect 77780 5608 77781 5648
rect 77739 5599 77781 5608
rect 1227 5564 1269 5573
rect 1227 5524 1228 5564
rect 1268 5524 1269 5564
rect 1227 5515 1269 5524
rect 4971 5564 5013 5573
rect 4971 5524 4972 5564
rect 5012 5524 5013 5564
rect 4971 5515 5013 5524
rect 48555 5564 48597 5573
rect 48555 5524 48556 5564
rect 48596 5524 48597 5564
rect 48555 5515 48597 5524
rect 49995 5564 50037 5573
rect 49995 5524 49996 5564
rect 50036 5524 50037 5564
rect 49995 5515 50037 5524
rect 52491 5564 52533 5573
rect 52491 5524 52492 5564
rect 52532 5524 52533 5564
rect 52491 5515 52533 5524
rect 56331 5564 56373 5573
rect 56331 5524 56332 5564
rect 56372 5524 56373 5564
rect 56331 5515 56373 5524
rect 61323 5564 61365 5573
rect 61323 5524 61324 5564
rect 61364 5524 61365 5564
rect 61323 5515 61365 5524
rect 73611 5564 73653 5573
rect 73611 5524 73612 5564
rect 73652 5524 73653 5564
rect 73611 5515 73653 5524
rect 76299 5564 76341 5573
rect 76299 5524 76300 5564
rect 76340 5524 76341 5564
rect 76299 5515 76341 5524
rect 77643 5564 77685 5573
rect 77643 5524 77644 5564
rect 77684 5524 77685 5564
rect 77643 5515 77685 5524
rect 843 5480 885 5489
rect 843 5440 844 5480
rect 884 5440 885 5480
rect 843 5431 885 5440
rect 7363 5480 7421 5481
rect 7363 5440 7372 5480
rect 7412 5440 7421 5480
rect 7363 5439 7421 5440
rect 47299 5480 47357 5481
rect 47299 5440 47308 5480
rect 47348 5440 47357 5480
rect 47299 5439 47357 5440
rect 59299 5480 59357 5481
rect 59299 5440 59308 5480
rect 59348 5440 59357 5480
rect 59299 5439 59357 5440
rect 60931 5480 60989 5481
rect 60931 5440 60940 5480
rect 60980 5440 60989 5480
rect 60931 5439 60989 5440
rect 64675 5480 64733 5481
rect 64675 5440 64684 5480
rect 64724 5440 64733 5480
rect 64675 5439 64733 5440
rect 576 5312 79584 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79584 5312
rect 576 5248 79584 5272
rect 651 5144 693 5153
rect 651 5104 652 5144
rect 692 5104 693 5144
rect 651 5095 693 5104
rect 2275 5144 2333 5145
rect 2275 5104 2284 5144
rect 2324 5104 2333 5144
rect 2275 5103 2333 5104
rect 52195 5144 52253 5145
rect 52195 5104 52204 5144
rect 52244 5104 52253 5144
rect 52195 5103 52253 5104
rect 55747 5144 55805 5145
rect 55747 5104 55756 5144
rect 55796 5104 55805 5144
rect 55747 5103 55805 5104
rect 65539 5144 65597 5145
rect 65539 5104 65548 5144
rect 65588 5104 65597 5144
rect 65539 5103 65597 5104
rect 65827 5144 65885 5145
rect 65827 5104 65836 5144
rect 65876 5104 65885 5144
rect 65827 5103 65885 5104
rect 71683 5144 71741 5145
rect 71683 5104 71692 5144
rect 71732 5104 71741 5144
rect 71683 5103 71741 5104
rect 76099 5144 76157 5145
rect 76099 5104 76108 5144
rect 76148 5104 76157 5144
rect 76099 5103 76157 5104
rect 1995 5060 2037 5069
rect 1995 5020 1996 5060
rect 2036 5020 2037 5060
rect 45867 5060 45909 5069
rect 1995 5011 2037 5020
rect 2187 5018 2229 5027
rect 1707 4976 1749 4985
rect 1707 4936 1708 4976
rect 1748 4936 1749 4976
rect 1707 4927 1749 4936
rect 1803 4976 1845 4985
rect 1803 4936 1804 4976
rect 1844 4936 1845 4976
rect 1803 4927 1845 4936
rect 1899 4976 1941 4985
rect 1899 4936 1900 4976
rect 1940 4936 1941 4976
rect 2187 4978 2188 5018
rect 2228 4978 2229 5018
rect 45867 5020 45868 5060
rect 45908 5020 45909 5060
rect 45867 5011 45909 5020
rect 56139 5060 56181 5069
rect 56139 5020 56140 5060
rect 56180 5020 56181 5060
rect 56139 5011 56181 5020
rect 58923 5060 58965 5069
rect 58923 5020 58924 5060
rect 58964 5020 58965 5060
rect 58923 5011 58965 5020
rect 62283 5060 62325 5069
rect 62283 5020 62284 5060
rect 62324 5020 62325 5060
rect 62283 5011 62325 5020
rect 63147 5060 63189 5069
rect 63147 5020 63148 5060
rect 63188 5020 63189 5060
rect 63147 5011 63189 5020
rect 66315 5060 66357 5069
rect 66315 5020 66316 5060
rect 66356 5020 66357 5060
rect 66315 5011 66357 5020
rect 76962 4989 77004 4998
rect 2187 4969 2229 4978
rect 2379 4976 2421 4985
rect 1899 4927 1941 4936
rect 2379 4936 2380 4976
rect 2420 4936 2421 4976
rect 2379 4927 2421 4936
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 3723 4976 3765 4985
rect 3723 4936 3724 4976
rect 3764 4936 3765 4976
rect 3723 4927 3765 4936
rect 3907 4976 3965 4977
rect 3907 4936 3916 4976
rect 3956 4936 3965 4976
rect 3907 4935 3965 4936
rect 4099 4976 4157 4977
rect 4099 4936 4108 4976
rect 4148 4936 4157 4976
rect 4099 4935 4157 4936
rect 5059 4976 5117 4977
rect 5059 4936 5068 4976
rect 5108 4936 5117 4976
rect 5059 4935 5117 4936
rect 46243 4976 46301 4977
rect 46243 4936 46252 4976
rect 46292 4936 46301 4976
rect 46243 4935 46301 4936
rect 47107 4976 47165 4977
rect 47107 4936 47116 4976
rect 47156 4936 47165 4976
rect 47107 4935 47165 4936
rect 48451 4976 48509 4977
rect 48451 4936 48460 4976
rect 48500 4936 48509 4976
rect 48451 4935 48509 4936
rect 48651 4976 48693 4985
rect 48651 4936 48652 4976
rect 48692 4936 48693 4976
rect 48651 4927 48693 4936
rect 48835 4976 48893 4977
rect 48835 4936 48844 4976
rect 48884 4936 48893 4976
rect 48835 4935 48893 4936
rect 48939 4976 48981 4985
rect 48939 4936 48940 4976
rect 48980 4936 48981 4976
rect 48939 4927 48981 4936
rect 49131 4976 49173 4985
rect 49131 4936 49132 4976
rect 49172 4936 49173 4976
rect 49131 4927 49173 4936
rect 51523 4976 51581 4977
rect 51523 4936 51532 4976
rect 51572 4936 51581 4976
rect 51523 4935 51581 4936
rect 51627 4976 51669 4985
rect 51627 4936 51628 4976
rect 51668 4936 51669 4976
rect 51627 4927 51669 4936
rect 51819 4976 51861 4985
rect 51819 4936 51820 4976
rect 51860 4936 51861 4976
rect 51819 4927 51861 4936
rect 52003 4976 52061 4977
rect 52003 4936 52012 4976
rect 52052 4936 52061 4976
rect 52003 4935 52061 4936
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 52299 4976 52341 4985
rect 52299 4936 52300 4976
rect 52340 4936 52341 4976
rect 52299 4927 52341 4936
rect 52491 4976 52533 4985
rect 52491 4936 52492 4976
rect 52532 4936 52533 4976
rect 52491 4927 52533 4936
rect 52675 4976 52733 4977
rect 52675 4936 52684 4976
rect 52724 4936 52733 4976
rect 52675 4935 52733 4936
rect 55659 4976 55701 4985
rect 55659 4936 55660 4976
rect 55700 4936 55701 4976
rect 55659 4927 55701 4936
rect 55851 4976 55893 4985
rect 55851 4936 55852 4976
rect 55892 4936 55893 4976
rect 55851 4927 55893 4936
rect 55939 4976 55997 4977
rect 55939 4936 55948 4976
rect 55988 4936 55997 4976
rect 55939 4935 55997 4936
rect 56515 4976 56573 4977
rect 56515 4936 56524 4976
rect 56564 4936 56573 4976
rect 56515 4935 56573 4936
rect 57379 4976 57437 4977
rect 57379 4936 57388 4976
rect 57428 4936 57437 4976
rect 57379 4935 57437 4936
rect 59299 4976 59357 4977
rect 59299 4936 59308 4976
rect 59348 4936 59357 4976
rect 59299 4935 59357 4936
rect 60163 4976 60221 4977
rect 60163 4936 60172 4976
rect 60212 4936 60221 4976
rect 60163 4935 60221 4936
rect 62187 4976 62229 4985
rect 62187 4936 62188 4976
rect 62228 4936 62229 4976
rect 62187 4927 62229 4936
rect 62371 4976 62429 4977
rect 62371 4936 62380 4976
rect 62420 4936 62429 4976
rect 62371 4935 62429 4936
rect 63523 4976 63581 4977
rect 63523 4936 63532 4976
rect 63572 4936 63581 4976
rect 63523 4935 63581 4936
rect 64387 4976 64445 4977
rect 64387 4936 64396 4976
rect 64436 4936 64445 4976
rect 64387 4935 64445 4936
rect 65739 4976 65781 4985
rect 65739 4936 65740 4976
rect 65780 4936 65781 4976
rect 65739 4927 65781 4936
rect 65931 4976 65973 4985
rect 65931 4936 65932 4976
rect 65972 4936 65973 4976
rect 65931 4927 65973 4936
rect 66019 4976 66077 4977
rect 66019 4936 66028 4976
rect 66068 4936 66077 4976
rect 66019 4935 66077 4936
rect 66211 4976 66269 4977
rect 66211 4936 66220 4976
rect 66260 4936 66269 4976
rect 66211 4935 66269 4936
rect 66411 4976 66453 4985
rect 66411 4936 66412 4976
rect 66452 4936 66453 4976
rect 66411 4927 66453 4936
rect 68907 4976 68949 4985
rect 68907 4936 68908 4976
rect 68948 4936 68949 4976
rect 68907 4927 68949 4936
rect 69099 4976 69141 4985
rect 69099 4936 69100 4976
rect 69140 4936 69141 4976
rect 69099 4927 69141 4936
rect 69187 4976 69245 4977
rect 69187 4936 69196 4976
rect 69236 4936 69245 4976
rect 69187 4935 69245 4936
rect 71595 4976 71637 4985
rect 71595 4936 71596 4976
rect 71636 4936 71637 4976
rect 71595 4927 71637 4936
rect 71787 4976 71829 4985
rect 71787 4936 71788 4976
rect 71828 4936 71829 4976
rect 71787 4927 71829 4936
rect 71875 4976 71933 4977
rect 71875 4936 71884 4976
rect 71924 4936 71933 4976
rect 71875 4935 71933 4936
rect 72067 4976 72125 4977
rect 72067 4936 72076 4976
rect 72116 4936 72125 4976
rect 72067 4935 72125 4936
rect 72171 4976 72213 4985
rect 72171 4936 72172 4976
rect 72212 4936 72213 4976
rect 72171 4927 72213 4936
rect 72267 4976 72309 4985
rect 72267 4936 72268 4976
rect 72308 4936 72309 4976
rect 72267 4927 72309 4936
rect 75907 4976 75965 4977
rect 75907 4936 75916 4976
rect 75956 4936 75965 4976
rect 75907 4935 75965 4936
rect 76011 4976 76053 4985
rect 76011 4936 76012 4976
rect 76052 4936 76053 4976
rect 76011 4927 76053 4936
rect 76203 4976 76245 4985
rect 76203 4936 76204 4976
rect 76244 4936 76245 4976
rect 76962 4949 76963 4989
rect 77003 4949 77004 4989
rect 77643 4989 77685 4998
rect 76962 4940 77004 4949
rect 77155 4976 77213 4977
rect 76203 4927 76245 4936
rect 77155 4936 77164 4976
rect 77204 4936 77213 4976
rect 77155 4935 77213 4936
rect 77443 4976 77501 4977
rect 77443 4936 77452 4976
rect 77492 4936 77501 4976
rect 77643 4949 77644 4989
rect 77684 4949 77685 4989
rect 77643 4940 77685 4949
rect 77443 4935 77501 4936
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 1507 4892 1565 4893
rect 1507 4852 1516 4892
rect 1556 4852 1565 4892
rect 1507 4851 1565 4852
rect 3819 4808 3861 4817
rect 3819 4768 3820 4808
rect 3860 4768 3861 4808
rect 3819 4759 3861 4768
rect 5547 4808 5589 4817
rect 5547 4768 5548 4808
rect 5588 4768 5589 4808
rect 5547 4759 5589 4768
rect 48555 4808 48597 4817
rect 48555 4768 48556 4808
rect 48596 4768 48597 4808
rect 48555 4759 48597 4768
rect 50187 4808 50229 4817
rect 50187 4768 50188 4808
rect 50228 4768 50229 4808
rect 50187 4759 50229 4768
rect 52875 4808 52917 4817
rect 52875 4768 52876 4808
rect 52916 4768 52917 4808
rect 52875 4759 52917 4768
rect 58531 4808 58589 4809
rect 58531 4768 58540 4808
rect 58580 4768 58589 4808
rect 58531 4767 58589 4768
rect 61803 4808 61845 4817
rect 61803 4768 61804 4808
rect 61844 4768 61845 4808
rect 61803 4759 61845 4768
rect 66891 4808 66933 4817
rect 66891 4768 66892 4808
rect 66932 4768 66933 4808
rect 66891 4759 66933 4768
rect 69387 4808 69429 4817
rect 69387 4768 69388 4808
rect 69428 4768 69429 4808
rect 69387 4759 69429 4768
rect 72459 4808 72501 4817
rect 72459 4768 72460 4808
rect 72500 4768 72501 4808
rect 72459 4759 72501 4768
rect 74283 4808 74325 4817
rect 74283 4768 74284 4808
rect 74324 4768 74325 4808
rect 74283 4759 74325 4768
rect 77835 4808 77877 4817
rect 77835 4768 77836 4808
rect 77876 4768 77877 4808
rect 77835 4759 77877 4768
rect 1323 4724 1365 4733
rect 1323 4684 1324 4724
rect 1364 4684 1365 4724
rect 1323 4675 1365 4684
rect 48259 4724 48317 4725
rect 48259 4684 48268 4724
rect 48308 4684 48317 4724
rect 48259 4683 48317 4684
rect 49131 4724 49173 4733
rect 49131 4684 49132 4724
rect 49172 4684 49173 4724
rect 49131 4675 49173 4684
rect 51819 4724 51861 4733
rect 51819 4684 51820 4724
rect 51860 4684 51861 4724
rect 51819 4675 51861 4684
rect 52587 4724 52629 4733
rect 52587 4684 52588 4724
rect 52628 4684 52629 4724
rect 52587 4675 52629 4684
rect 61315 4724 61373 4725
rect 61315 4684 61324 4724
rect 61364 4684 61373 4724
rect 61315 4683 61373 4684
rect 68907 4724 68949 4733
rect 68907 4684 68908 4724
rect 68948 4684 68949 4724
rect 68907 4675 68949 4684
rect 77067 4724 77109 4733
rect 77067 4684 77068 4724
rect 77108 4684 77109 4724
rect 77067 4675 77109 4684
rect 77547 4724 77589 4733
rect 77547 4684 77548 4724
rect 77588 4684 77589 4724
rect 77547 4675 77589 4684
rect 576 4556 79584 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79584 4556
rect 576 4492 79584 4516
rect 2571 4388 2613 4397
rect 2571 4348 2572 4388
rect 2612 4348 2613 4388
rect 2571 4339 2613 4348
rect 52003 4388 52061 4389
rect 52003 4348 52012 4388
rect 52052 4348 52061 4388
rect 52003 4347 52061 4348
rect 61507 4388 61565 4389
rect 61507 4348 61516 4388
rect 61556 4348 61565 4388
rect 61507 4347 61565 4348
rect 66211 4388 66269 4389
rect 66211 4348 66220 4388
rect 66260 4348 66269 4388
rect 66211 4347 66269 4348
rect 76867 4388 76925 4389
rect 76867 4348 76876 4388
rect 76916 4348 76925 4388
rect 76867 4347 76925 4348
rect 651 4304 693 4313
rect 651 4264 652 4304
rect 692 4264 693 4304
rect 651 4255 693 4264
rect 1899 4304 1941 4313
rect 1899 4264 1900 4304
rect 1940 4264 1941 4304
rect 1899 4255 1941 4264
rect 4195 4304 4253 4305
rect 4195 4264 4204 4304
rect 4244 4264 4253 4304
rect 4195 4263 4253 4264
rect 7459 4304 7517 4305
rect 7459 4264 7468 4304
rect 7508 4264 7517 4304
rect 7459 4263 7517 4264
rect 55179 4304 55221 4313
rect 55179 4264 55180 4304
rect 55220 4264 55221 4304
rect 55179 4255 55221 4264
rect 56899 4304 56957 4305
rect 56899 4264 56908 4304
rect 56948 4264 56957 4304
rect 56899 4263 56957 4264
rect 57963 4304 58005 4313
rect 57963 4264 57964 4304
rect 58004 4264 58005 4304
rect 57963 4255 58005 4264
rect 60171 4304 60213 4313
rect 60171 4264 60172 4304
rect 60212 4264 60213 4304
rect 60171 4255 60213 4264
rect 68803 4304 68861 4305
rect 68803 4264 68812 4304
rect 68852 4264 68861 4304
rect 68803 4263 68861 4264
rect 74371 4304 74429 4305
rect 74371 4264 74380 4304
rect 74420 4264 74429 4304
rect 74371 4263 74429 4264
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 1219 4220 1277 4221
rect 1219 4180 1228 4220
rect 1268 4180 1277 4220
rect 1219 4179 1277 4180
rect 79467 4220 79509 4229
rect 79467 4180 79468 4220
rect 79508 4180 79509 4220
rect 79467 4171 79509 4180
rect 2091 4136 2133 4145
rect 2091 4096 2092 4136
rect 2132 4096 2133 4136
rect 2091 4087 2133 4096
rect 2187 4136 2229 4145
rect 2187 4096 2188 4136
rect 2228 4096 2229 4136
rect 2187 4087 2229 4096
rect 2283 4136 2325 4145
rect 2283 4096 2284 4136
rect 2324 4096 2325 4136
rect 2283 4087 2325 4096
rect 2571 4136 2613 4145
rect 2571 4096 2572 4136
rect 2612 4096 2613 4136
rect 2571 4087 2613 4096
rect 2763 4136 2805 4145
rect 2763 4096 2764 4136
rect 2804 4096 2805 4136
rect 2763 4087 2805 4096
rect 2877 4136 2919 4145
rect 2877 4096 2878 4136
rect 2918 4096 2919 4136
rect 2877 4087 2919 4096
rect 3523 4136 3581 4137
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 3523 4095 3581 4096
rect 3819 4136 3861 4145
rect 3819 4096 3820 4136
rect 3860 4096 3861 4136
rect 3819 4087 3861 4096
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4779 4136 4821 4145
rect 4779 4096 4780 4136
rect 4820 4096 4821 4136
rect 4779 4087 4821 4096
rect 4867 4136 4925 4137
rect 4867 4096 4876 4136
rect 4916 4096 4925 4136
rect 4867 4095 4925 4096
rect 5443 4136 5501 4137
rect 5443 4096 5452 4136
rect 5492 4096 5501 4136
rect 5443 4095 5501 4096
rect 6307 4136 6365 4137
rect 6307 4096 6316 4136
rect 6356 4096 6365 4136
rect 6307 4095 6365 4096
rect 47403 4136 47445 4145
rect 47403 4096 47404 4136
rect 47444 4096 47445 4136
rect 47403 4087 47445 4096
rect 47499 4136 47541 4145
rect 47499 4096 47500 4136
rect 47540 4096 47541 4136
rect 47499 4087 47541 4096
rect 47595 4136 47637 4145
rect 47595 4096 47596 4136
rect 47636 4096 47637 4136
rect 47595 4087 47637 4096
rect 47691 4136 47733 4145
rect 47691 4096 47692 4136
rect 47732 4096 47733 4136
rect 47691 4087 47733 4096
rect 49987 4136 50045 4137
rect 49987 4096 49996 4136
rect 50036 4096 50045 4136
rect 49987 4095 50045 4096
rect 50851 4136 50909 4137
rect 50851 4096 50860 4136
rect 50900 4096 50909 4136
rect 50851 4095 50909 4096
rect 52395 4136 52437 4145
rect 52395 4096 52396 4136
rect 52436 4096 52437 4136
rect 52395 4087 52437 4096
rect 52771 4136 52829 4137
rect 52771 4096 52780 4136
rect 52820 4096 52829 4136
rect 52771 4095 52829 4096
rect 53635 4136 53693 4137
rect 53635 4096 53644 4136
rect 53684 4096 53693 4136
rect 53635 4095 53693 4096
rect 55659 4136 55701 4145
rect 55659 4096 55660 4136
rect 55700 4096 55701 4136
rect 55659 4087 55701 4096
rect 55755 4136 55797 4145
rect 55755 4096 55756 4136
rect 55796 4096 55797 4136
rect 55755 4087 55797 4096
rect 55851 4136 55893 4145
rect 55851 4096 55852 4136
rect 55892 4096 55893 4136
rect 55851 4087 55893 4096
rect 55947 4136 55989 4145
rect 55947 4096 55948 4136
rect 55988 4096 55989 4136
rect 55947 4087 55989 4096
rect 56227 4136 56285 4137
rect 56227 4096 56236 4136
rect 56276 4096 56285 4136
rect 56227 4095 56285 4096
rect 56523 4136 56565 4145
rect 56523 4096 56524 4136
rect 56564 4096 56565 4136
rect 56523 4087 56565 4096
rect 57099 4136 57141 4145
rect 57099 4096 57100 4136
rect 57140 4096 57141 4136
rect 57099 4087 57141 4096
rect 57291 4136 57333 4145
rect 57291 4096 57292 4136
rect 57332 4096 57333 4136
rect 57291 4087 57333 4096
rect 57379 4136 57437 4137
rect 57379 4096 57388 4136
rect 57428 4096 57437 4136
rect 57379 4095 57437 4096
rect 57963 4136 58005 4145
rect 57963 4096 57964 4136
rect 58004 4096 58005 4136
rect 57963 4087 58005 4096
rect 58155 4136 58197 4145
rect 58155 4096 58156 4136
rect 58196 4096 58197 4136
rect 58155 4087 58197 4096
rect 58243 4136 58301 4137
rect 58243 4096 58252 4136
rect 58292 4096 58301 4136
rect 58243 4095 58301 4096
rect 59019 4136 59061 4145
rect 59019 4096 59020 4136
rect 59060 4096 59061 4136
rect 59019 4087 59061 4096
rect 59115 4136 59157 4145
rect 59115 4096 59116 4136
rect 59156 4096 59157 4136
rect 59115 4087 59157 4096
rect 59211 4136 59253 4145
rect 59211 4096 59212 4136
rect 59252 4096 59253 4136
rect 59211 4087 59253 4096
rect 59307 4136 59349 4145
rect 59307 4096 59308 4136
rect 59348 4096 59349 4136
rect 59307 4087 59349 4096
rect 60835 4136 60893 4137
rect 60835 4096 60844 4136
rect 60884 4096 60893 4136
rect 60835 4095 60893 4096
rect 61131 4136 61173 4145
rect 61131 4096 61132 4136
rect 61172 4096 61173 4136
rect 61131 4087 61173 4096
rect 61227 4136 61269 4145
rect 61227 4096 61228 4136
rect 61268 4096 61269 4136
rect 61227 4087 61269 4096
rect 63235 4136 63293 4137
rect 63235 4096 63244 4136
rect 63284 4096 63293 4136
rect 63235 4095 63293 4096
rect 64099 4136 64157 4137
rect 64099 4096 64108 4136
rect 64148 4096 64157 4136
rect 64099 4095 64157 4096
rect 65539 4136 65597 4137
rect 65539 4096 65548 4136
rect 65588 4096 65597 4136
rect 65539 4095 65597 4096
rect 65835 4136 65877 4145
rect 65835 4096 65836 4136
rect 65876 4096 65877 4136
rect 65835 4087 65877 4096
rect 66787 4136 66845 4137
rect 66787 4096 66796 4136
rect 66836 4096 66845 4136
rect 66787 4095 66845 4096
rect 67651 4136 67709 4137
rect 67651 4096 67660 4136
rect 67700 4096 67709 4136
rect 67651 4095 67709 4096
rect 69379 4136 69437 4137
rect 69379 4096 69388 4136
rect 69428 4096 69437 4136
rect 69379 4095 69437 4096
rect 70243 4136 70301 4137
rect 70243 4096 70252 4136
rect 70292 4096 70301 4136
rect 70243 4095 70301 4096
rect 71587 4136 71645 4137
rect 71587 4096 71596 4136
rect 71636 4096 71645 4136
rect 71587 4095 71645 4096
rect 71787 4136 71829 4145
rect 71787 4096 71788 4136
rect 71828 4096 71829 4136
rect 71787 4087 71829 4096
rect 71979 4136 72021 4145
rect 71979 4096 71980 4136
rect 72020 4096 72021 4136
rect 71979 4087 72021 4096
rect 72355 4136 72413 4137
rect 72355 4096 72364 4136
rect 72404 4096 72413 4136
rect 72355 4095 72413 4096
rect 73219 4136 73277 4137
rect 73219 4096 73228 4136
rect 73268 4096 73277 4136
rect 73219 4095 73277 4096
rect 75147 4136 75189 4145
rect 75147 4096 75148 4136
rect 75188 4096 75189 4136
rect 75147 4087 75189 4096
rect 75339 4136 75381 4145
rect 75339 4096 75340 4136
rect 75380 4096 75381 4136
rect 75339 4087 75381 4096
rect 75427 4136 75485 4137
rect 75427 4096 75436 4136
rect 75476 4096 75485 4136
rect 75427 4095 75485 4096
rect 75627 4136 75669 4145
rect 75627 4096 75628 4136
rect 75668 4096 75669 4136
rect 75627 4087 75669 4096
rect 75723 4136 75765 4145
rect 75723 4096 75724 4136
rect 75764 4096 75765 4136
rect 75723 4087 75765 4096
rect 75819 4136 75861 4145
rect 75819 4096 75820 4136
rect 75860 4096 75861 4136
rect 75819 4087 75861 4096
rect 75915 4136 75957 4145
rect 75915 4096 75916 4136
rect 75956 4096 75957 4136
rect 75915 4087 75957 4096
rect 76195 4136 76253 4137
rect 76195 4096 76204 4136
rect 76244 4096 76253 4136
rect 76195 4095 76253 4096
rect 76491 4136 76533 4145
rect 76491 4096 76492 4136
rect 76532 4096 76533 4136
rect 76491 4087 76533 4096
rect 76587 4136 76629 4145
rect 76587 4096 76588 4136
rect 76628 4096 76629 4136
rect 76587 4087 76629 4096
rect 77443 4136 77501 4137
rect 77443 4096 77452 4136
rect 77492 4096 77501 4136
rect 77443 4095 77501 4096
rect 78307 4136 78365 4137
rect 78307 4096 78316 4136
rect 78356 4096 78365 4136
rect 78307 4095 78365 4096
rect 3915 4052 3957 4061
rect 3915 4012 3916 4052
rect 3956 4012 3957 4052
rect 3915 4003 3957 4012
rect 5067 4052 5109 4061
rect 5067 4012 5068 4052
rect 5108 4012 5109 4052
rect 5067 4003 5109 4012
rect 49611 4052 49653 4061
rect 49611 4012 49612 4052
rect 49652 4012 49653 4052
rect 49611 4003 49653 4012
rect 56619 4052 56661 4061
rect 56619 4012 56620 4052
rect 56660 4012 56661 4052
rect 56619 4003 56661 4012
rect 62859 4052 62901 4061
rect 62859 4012 62860 4052
rect 62900 4012 62901 4052
rect 62859 4003 62901 4012
rect 65931 4052 65973 4061
rect 65931 4012 65932 4052
rect 65972 4012 65973 4052
rect 65931 4003 65973 4012
rect 66411 4052 66453 4061
rect 66411 4012 66412 4052
rect 66452 4012 66453 4052
rect 66411 4003 66453 4012
rect 69003 4052 69045 4061
rect 69003 4012 69004 4052
rect 69044 4012 69045 4052
rect 69003 4003 69045 4012
rect 71691 4052 71733 4061
rect 71691 4012 71692 4052
rect 71732 4012 71733 4052
rect 71691 4003 71733 4012
rect 77067 4052 77109 4061
rect 77067 4012 77068 4052
rect 77108 4012 77109 4052
rect 77067 4003 77109 4012
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 2371 3968 2429 3969
rect 2371 3928 2380 3968
rect 2420 3928 2429 3968
rect 2371 3927 2429 3928
rect 4675 3968 4733 3969
rect 4675 3928 4684 3968
rect 4724 3928 4733 3968
rect 4675 3927 4733 3928
rect 52003 3968 52061 3969
rect 52003 3928 52012 3968
rect 52052 3928 52061 3968
rect 52003 3927 52061 3928
rect 54787 3968 54845 3969
rect 54787 3928 54796 3968
rect 54836 3928 54845 3968
rect 54787 3927 54845 3928
rect 57187 3968 57245 3969
rect 57187 3928 57196 3968
rect 57236 3928 57245 3968
rect 57187 3927 57245 3928
rect 65251 3968 65309 3969
rect 65251 3928 65260 3968
rect 65300 3928 65309 3968
rect 65251 3927 65309 3928
rect 71395 3968 71453 3969
rect 71395 3928 71404 3968
rect 71444 3928 71453 3968
rect 71395 3927 71453 3928
rect 75235 3968 75293 3969
rect 75235 3928 75244 3968
rect 75284 3928 75293 3968
rect 75235 3927 75293 3928
rect 576 3800 79584 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79584 3800
rect 576 3736 79584 3760
rect 3811 3632 3869 3633
rect 3811 3592 3820 3632
rect 3860 3592 3869 3632
rect 3811 3591 3869 3592
rect 4675 3632 4733 3633
rect 4675 3592 4684 3632
rect 4724 3592 4733 3632
rect 4675 3591 4733 3592
rect 50275 3632 50333 3633
rect 50275 3592 50284 3632
rect 50324 3592 50333 3632
rect 50275 3591 50333 3592
rect 53923 3632 53981 3633
rect 53923 3592 53932 3632
rect 53972 3592 53981 3632
rect 53923 3591 53981 3592
rect 62083 3632 62141 3633
rect 62083 3592 62092 3632
rect 62132 3592 62141 3632
rect 62083 3591 62141 3592
rect 64003 3632 64061 3633
rect 64003 3592 64012 3632
rect 64052 3592 64061 3632
rect 64003 3591 64061 3592
rect 66211 3632 66269 3633
rect 66211 3592 66220 3632
rect 66260 3592 66269 3632
rect 66211 3591 66269 3592
rect 69379 3632 69437 3633
rect 69379 3592 69388 3632
rect 69428 3592 69437 3632
rect 69379 3591 69437 3592
rect 76195 3632 76253 3633
rect 76195 3592 76204 3632
rect 76244 3592 76253 3632
rect 76195 3591 76253 3592
rect 76483 3632 76541 3633
rect 76483 3592 76492 3632
rect 76532 3592 76541 3632
rect 76483 3591 76541 3592
rect 77251 3632 77309 3633
rect 77251 3592 77260 3632
rect 77300 3592 77309 3632
rect 77251 3591 77309 3592
rect 52107 3548 52149 3557
rect 52107 3508 52108 3548
rect 52148 3508 52149 3548
rect 52107 3499 52149 3508
rect 52683 3548 52725 3557
rect 52683 3508 52684 3548
rect 52724 3508 52725 3548
rect 52683 3499 52725 3508
rect 56331 3548 56373 3557
rect 56331 3508 56332 3548
rect 56372 3508 56373 3548
rect 56331 3499 56373 3508
rect 56811 3548 56853 3557
rect 56811 3508 56812 3548
rect 56852 3508 56853 3548
rect 56811 3499 56853 3508
rect 73803 3548 73845 3557
rect 73803 3508 73804 3548
rect 73844 3508 73845 3548
rect 73803 3499 73845 3508
rect 1419 3464 1461 3473
rect 1419 3424 1420 3464
rect 1460 3424 1461 3464
rect 1419 3415 1461 3424
rect 1795 3464 1853 3465
rect 1795 3424 1804 3464
rect 1844 3424 1853 3464
rect 1795 3423 1853 3424
rect 2659 3464 2717 3465
rect 2659 3424 2668 3464
rect 2708 3424 2717 3464
rect 2659 3423 2717 3424
rect 4203 3464 4245 3473
rect 4203 3424 4204 3464
rect 4244 3424 4245 3464
rect 4203 3415 4245 3424
rect 4387 3464 4445 3465
rect 4387 3424 4396 3464
rect 4436 3424 4445 3464
rect 4779 3464 4821 3473
rect 4387 3423 4445 3424
rect 4587 3453 4629 3462
rect 4587 3413 4588 3453
rect 4628 3413 4629 3453
rect 4779 3424 4780 3464
rect 4820 3424 4821 3464
rect 4779 3415 4821 3424
rect 4867 3464 4925 3465
rect 4867 3424 4876 3464
rect 4916 3424 4925 3464
rect 4867 3423 4925 3424
rect 5059 3464 5117 3465
rect 5059 3424 5068 3464
rect 5108 3424 5117 3464
rect 5059 3423 5117 3424
rect 5259 3464 5301 3473
rect 5259 3424 5260 3464
rect 5300 3424 5301 3464
rect 5259 3415 5301 3424
rect 50083 3464 50141 3465
rect 50083 3424 50092 3464
rect 50132 3424 50141 3464
rect 50083 3423 50141 3424
rect 50187 3464 50229 3473
rect 50187 3424 50188 3464
rect 50228 3424 50229 3464
rect 50187 3415 50229 3424
rect 50379 3464 50421 3473
rect 50379 3424 50380 3464
rect 50420 3424 50421 3464
rect 50379 3415 50421 3424
rect 50667 3464 50709 3473
rect 50667 3424 50668 3464
rect 50708 3424 50709 3464
rect 50667 3415 50709 3424
rect 50763 3464 50805 3473
rect 50763 3424 50764 3464
rect 50804 3424 50805 3464
rect 50763 3415 50805 3424
rect 50859 3464 50901 3473
rect 50859 3424 50860 3464
rect 50900 3424 50901 3464
rect 50859 3415 50901 3424
rect 50955 3464 50997 3473
rect 50955 3424 50956 3464
rect 50996 3424 50997 3464
rect 50955 3415 50997 3424
rect 51715 3464 51773 3465
rect 51715 3424 51724 3464
rect 51764 3424 51773 3464
rect 51715 3423 51773 3424
rect 52011 3464 52053 3473
rect 52011 3424 52012 3464
rect 52052 3424 52053 3464
rect 52011 3415 52053 3424
rect 52579 3464 52637 3465
rect 52579 3424 52588 3464
rect 52628 3424 52637 3464
rect 52579 3423 52637 3424
rect 52779 3464 52821 3473
rect 52779 3424 52780 3464
rect 52820 3424 52821 3464
rect 52779 3415 52821 3424
rect 55075 3464 55133 3465
rect 55075 3424 55084 3464
rect 55124 3424 55133 3464
rect 55075 3423 55133 3424
rect 55939 3464 55997 3465
rect 55939 3424 55948 3464
rect 55988 3424 55997 3464
rect 55939 3423 55997 3424
rect 56707 3464 56765 3465
rect 56707 3424 56716 3464
rect 56756 3424 56765 3464
rect 56707 3423 56765 3424
rect 56907 3464 56949 3473
rect 56907 3424 56908 3464
rect 56948 3424 56949 3464
rect 56907 3415 56949 3424
rect 59299 3464 59357 3465
rect 59299 3424 59308 3464
rect 59348 3424 59357 3464
rect 59299 3423 59357 3424
rect 59499 3464 59541 3473
rect 59499 3424 59500 3464
rect 59540 3424 59541 3464
rect 59499 3415 59541 3424
rect 59691 3464 59733 3473
rect 59691 3424 59692 3464
rect 59732 3424 59733 3464
rect 59691 3415 59733 3424
rect 60067 3464 60125 3465
rect 60067 3424 60076 3464
rect 60116 3424 60125 3464
rect 60067 3423 60125 3424
rect 60931 3464 60989 3465
rect 60931 3424 60940 3464
rect 60980 3424 60989 3464
rect 60931 3423 60989 3424
rect 63811 3464 63869 3465
rect 63811 3424 63820 3464
rect 63860 3424 63869 3464
rect 63811 3423 63869 3424
rect 63915 3464 63957 3473
rect 63915 3424 63916 3464
rect 63956 3424 63957 3464
rect 63915 3415 63957 3424
rect 64107 3464 64149 3473
rect 64107 3424 64108 3464
rect 64148 3424 64149 3464
rect 64107 3415 64149 3424
rect 64299 3464 64341 3473
rect 64299 3424 64300 3464
rect 64340 3424 64341 3464
rect 64299 3415 64341 3424
rect 64395 3464 64437 3473
rect 64395 3424 64396 3464
rect 64436 3424 64437 3464
rect 64395 3415 64437 3424
rect 64491 3464 64533 3473
rect 64491 3424 64492 3464
rect 64532 3424 64533 3464
rect 64491 3415 64533 3424
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 66123 3464 66165 3473
rect 66123 3424 66124 3464
rect 66164 3424 66165 3464
rect 66123 3415 66165 3424
rect 66315 3464 66357 3473
rect 66315 3424 66316 3464
rect 66356 3424 66357 3464
rect 66315 3415 66357 3424
rect 66403 3464 66461 3465
rect 66403 3424 66412 3464
rect 66452 3424 66461 3464
rect 66403 3423 66461 3424
rect 66595 3464 66653 3465
rect 66595 3424 66604 3464
rect 66644 3424 66653 3464
rect 66595 3423 66653 3424
rect 66795 3464 66837 3473
rect 66795 3424 66796 3464
rect 66836 3424 66837 3464
rect 66795 3415 66837 3424
rect 68611 3464 68669 3465
rect 68611 3424 68620 3464
rect 68660 3424 68669 3464
rect 68611 3423 68669 3424
rect 68715 3464 68757 3473
rect 68715 3424 68716 3464
rect 68756 3424 68757 3464
rect 68715 3415 68757 3424
rect 68907 3464 68949 3473
rect 68907 3424 68908 3464
rect 68948 3424 68949 3464
rect 68907 3415 68949 3424
rect 69187 3464 69245 3465
rect 69187 3424 69196 3464
rect 69236 3424 69245 3464
rect 69187 3423 69245 3424
rect 69291 3464 69333 3473
rect 69291 3424 69292 3464
rect 69332 3424 69333 3464
rect 69291 3415 69333 3424
rect 69483 3464 69525 3473
rect 69483 3424 69484 3464
rect 69524 3424 69525 3464
rect 69483 3415 69525 3424
rect 69771 3464 69813 3473
rect 69771 3424 69772 3464
rect 69812 3424 69813 3464
rect 69771 3415 69813 3424
rect 69867 3464 69909 3473
rect 69867 3424 69868 3464
rect 69908 3424 69909 3464
rect 69867 3415 69909 3424
rect 69963 3464 70005 3473
rect 69963 3424 69964 3464
rect 70004 3424 70005 3464
rect 69963 3415 70005 3424
rect 70059 3464 70101 3473
rect 70059 3424 70060 3464
rect 70100 3424 70101 3464
rect 70059 3415 70101 3424
rect 71203 3464 71261 3465
rect 71203 3424 71212 3464
rect 71252 3424 71261 3464
rect 71203 3423 71261 3424
rect 71499 3464 71541 3473
rect 71499 3424 71500 3464
rect 71540 3424 71541 3464
rect 71499 3415 71541 3424
rect 71595 3464 71637 3473
rect 71595 3424 71596 3464
rect 71636 3424 71637 3464
rect 71595 3415 71637 3424
rect 72067 3464 72125 3465
rect 72067 3424 72076 3464
rect 72116 3424 72125 3464
rect 72067 3423 72125 3424
rect 72171 3464 72213 3473
rect 72171 3424 72172 3464
rect 72212 3424 72213 3464
rect 72171 3415 72213 3424
rect 72363 3464 72405 3473
rect 72363 3424 72364 3464
rect 72404 3424 72405 3464
rect 72363 3415 72405 3424
rect 74179 3464 74237 3465
rect 74179 3424 74188 3464
rect 74228 3424 74237 3464
rect 74179 3423 74237 3424
rect 75043 3464 75101 3465
rect 75043 3424 75052 3464
rect 75092 3424 75101 3464
rect 75043 3423 75101 3424
rect 76395 3464 76437 3473
rect 76395 3424 76396 3464
rect 76436 3424 76437 3464
rect 76395 3415 76437 3424
rect 76587 3464 76629 3473
rect 76587 3424 76588 3464
rect 76628 3424 76629 3464
rect 76587 3415 76629 3424
rect 76675 3464 76733 3465
rect 76675 3424 76684 3464
rect 76724 3424 76733 3464
rect 76675 3423 76733 3424
rect 77163 3464 77205 3473
rect 77163 3424 77164 3464
rect 77204 3424 77205 3464
rect 77163 3415 77205 3424
rect 77355 3464 77397 3473
rect 77355 3424 77356 3464
rect 77396 3424 77397 3464
rect 77355 3415 77397 3424
rect 77443 3464 77501 3465
rect 77443 3424 77452 3464
rect 77492 3424 77501 3464
rect 77443 3423 77501 3424
rect 4587 3404 4629 3413
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 1219 3380 1277 3381
rect 1219 3340 1228 3380
rect 1268 3340 1277 3380
rect 1219 3339 1277 3340
rect 63339 3338 63381 3347
rect 1035 3296 1077 3305
rect 1035 3256 1036 3296
rect 1076 3256 1077 3296
rect 1035 3247 1077 3256
rect 5163 3296 5205 3305
rect 63339 3298 63340 3338
rect 63380 3298 63381 3338
rect 5163 3256 5164 3296
rect 5204 3256 5205 3296
rect 5163 3247 5205 3256
rect 52387 3296 52445 3297
rect 52387 3256 52396 3296
rect 52436 3256 52445 3296
rect 63339 3289 63381 3298
rect 66699 3296 66741 3305
rect 52387 3255 52445 3256
rect 66699 3256 66700 3296
rect 66740 3256 66741 3296
rect 66699 3247 66741 3256
rect 68907 3296 68949 3305
rect 68907 3256 68908 3296
rect 68948 3256 68949 3296
rect 68907 3247 68949 3256
rect 71875 3296 71933 3297
rect 71875 3256 71884 3296
rect 71924 3256 71933 3296
rect 71875 3255 71933 3256
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 4299 3212 4341 3221
rect 4299 3172 4300 3212
rect 4340 3172 4341 3212
rect 4299 3163 4341 3172
rect 59403 3212 59445 3221
rect 59403 3172 59404 3212
rect 59444 3172 59445 3212
rect 59403 3163 59445 3172
rect 72363 3212 72405 3221
rect 72363 3172 72364 3212
rect 72404 3172 72405 3212
rect 72363 3163 72405 3172
rect 576 3044 79584 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79584 3044
rect 576 2980 79584 3004
rect 59115 2876 59157 2885
rect 59115 2836 59116 2876
rect 59156 2836 59157 2876
rect 59115 2827 59157 2836
rect 64011 2876 64053 2885
rect 64011 2836 64012 2876
rect 64052 2836 64053 2876
rect 64011 2827 64053 2836
rect 73515 2876 73557 2885
rect 73515 2836 73516 2876
rect 73556 2836 73557 2876
rect 73515 2827 73557 2836
rect 1515 2792 1557 2801
rect 1515 2752 1516 2792
rect 1556 2752 1557 2792
rect 1515 2743 1557 2752
rect 54027 2792 54069 2801
rect 54027 2752 54028 2792
rect 54068 2752 54069 2792
rect 54027 2743 54069 2752
rect 56811 2792 56853 2801
rect 56811 2752 56812 2792
rect 56852 2752 56853 2792
rect 56811 2743 56853 2752
rect 57099 2792 57141 2801
rect 57099 2752 57100 2792
rect 57140 2752 57141 2792
rect 57099 2743 57141 2752
rect 60067 2792 60125 2793
rect 60067 2752 60076 2792
rect 60116 2752 60125 2792
rect 60067 2751 60125 2752
rect 62187 2792 62229 2801
rect 62187 2752 62188 2792
rect 62228 2752 62229 2792
rect 62187 2743 62229 2752
rect 66507 2792 66549 2801
rect 66507 2752 66508 2792
rect 66548 2752 66549 2792
rect 66507 2743 66549 2752
rect 68715 2792 68757 2801
rect 68715 2752 68716 2792
rect 68756 2752 68757 2792
rect 68715 2743 68757 2752
rect 71499 2792 71541 2801
rect 71499 2752 71500 2792
rect 71540 2752 71541 2792
rect 71499 2743 71541 2752
rect 72931 2792 72989 2793
rect 72931 2752 72940 2792
rect 72980 2752 72989 2792
rect 72931 2751 72989 2752
rect 74955 2792 74997 2801
rect 74955 2752 74956 2792
rect 74996 2752 74997 2792
rect 74955 2743 74997 2752
rect 76107 2792 76149 2801
rect 76107 2752 76108 2792
rect 76148 2752 76149 2792
rect 76107 2743 76149 2752
rect 77443 2792 77501 2793
rect 77443 2752 77452 2792
rect 77492 2752 77501 2792
rect 77443 2751 77501 2752
rect 78219 2792 78261 2801
rect 78219 2752 78220 2792
rect 78260 2752 78261 2792
rect 78219 2743 78261 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 1699 2708 1757 2709
rect 1699 2668 1708 2708
rect 1748 2668 1757 2708
rect 1699 2667 1757 2668
rect 64779 2708 64821 2717
rect 64779 2668 64780 2708
rect 64820 2668 64821 2708
rect 64779 2659 64821 2668
rect 2379 2624 2421 2633
rect 2379 2584 2380 2624
rect 2420 2584 2421 2624
rect 2379 2575 2421 2584
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2659 2624 2717 2625
rect 2659 2584 2668 2624
rect 2708 2584 2717 2624
rect 2659 2583 2717 2584
rect 2859 2624 2901 2633
rect 2859 2584 2860 2624
rect 2900 2584 2901 2624
rect 2859 2575 2901 2584
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 3051 2575 3093 2584
rect 3139 2624 3197 2625
rect 3139 2584 3148 2624
rect 3188 2584 3197 2624
rect 3139 2583 3197 2584
rect 55371 2624 55413 2633
rect 55371 2584 55372 2624
rect 55412 2584 55413 2624
rect 55371 2575 55413 2584
rect 55467 2624 55509 2633
rect 55467 2584 55468 2624
rect 55508 2584 55509 2624
rect 55467 2575 55509 2584
rect 55563 2624 55605 2633
rect 55563 2584 55564 2624
rect 55604 2584 55605 2624
rect 55563 2575 55605 2584
rect 55755 2624 55797 2633
rect 55755 2584 55756 2624
rect 55796 2584 55797 2624
rect 55755 2575 55797 2584
rect 55947 2624 55989 2633
rect 55947 2584 55948 2624
rect 55988 2584 55989 2624
rect 55947 2575 55989 2584
rect 56035 2624 56093 2625
rect 56035 2584 56044 2624
rect 56084 2584 56093 2624
rect 56035 2583 56093 2584
rect 56235 2624 56277 2633
rect 56235 2584 56236 2624
rect 56276 2584 56277 2624
rect 56235 2575 56277 2584
rect 56427 2624 56469 2633
rect 56427 2584 56428 2624
rect 56468 2584 56469 2624
rect 56427 2575 56469 2584
rect 56515 2624 56573 2625
rect 56515 2584 56524 2624
rect 56564 2584 56573 2624
rect 56515 2583 56573 2584
rect 56707 2624 56765 2625
rect 56707 2584 56716 2624
rect 56756 2584 56765 2624
rect 56707 2583 56765 2584
rect 56907 2624 56949 2633
rect 56907 2584 56908 2624
rect 56948 2584 56949 2624
rect 56907 2575 56949 2584
rect 58819 2624 58877 2625
rect 58819 2584 58828 2624
rect 58868 2584 58877 2624
rect 58819 2583 58877 2584
rect 58923 2624 58965 2633
rect 58923 2584 58924 2624
rect 58964 2584 58965 2624
rect 58923 2575 58965 2584
rect 59115 2624 59157 2633
rect 59115 2584 59116 2624
rect 59156 2584 59157 2624
rect 59115 2575 59157 2584
rect 59395 2624 59453 2625
rect 59395 2584 59404 2624
rect 59444 2584 59453 2624
rect 59395 2583 59453 2584
rect 59691 2624 59733 2633
rect 59691 2584 59692 2624
rect 59732 2584 59733 2624
rect 59691 2575 59733 2584
rect 60267 2624 60309 2633
rect 60267 2584 60268 2624
rect 60308 2584 60309 2624
rect 60267 2575 60309 2584
rect 60363 2624 60405 2633
rect 60363 2584 60364 2624
rect 60404 2584 60405 2624
rect 60363 2575 60405 2584
rect 60451 2624 60509 2625
rect 60451 2584 60460 2624
rect 60500 2584 60509 2624
rect 60451 2583 60509 2584
rect 63715 2624 63773 2625
rect 63715 2584 63724 2624
rect 63764 2584 63773 2624
rect 63715 2583 63773 2584
rect 63819 2624 63861 2633
rect 63819 2584 63820 2624
rect 63860 2584 63861 2624
rect 63819 2575 63861 2584
rect 64011 2624 64053 2633
rect 64011 2584 64012 2624
rect 64052 2584 64053 2624
rect 64011 2575 64053 2584
rect 64203 2624 64245 2633
rect 64203 2584 64204 2624
rect 64244 2584 64245 2624
rect 64203 2575 64245 2584
rect 64395 2624 64437 2633
rect 64395 2584 64396 2624
rect 64436 2584 64437 2624
rect 64395 2575 64437 2584
rect 64483 2624 64541 2625
rect 64483 2584 64492 2624
rect 64532 2584 64541 2624
rect 64483 2583 64541 2584
rect 64675 2624 64733 2625
rect 64675 2584 64684 2624
rect 64724 2584 64733 2624
rect 64675 2583 64733 2584
rect 64875 2624 64917 2633
rect 64875 2584 64876 2624
rect 64916 2584 64917 2624
rect 64875 2575 64917 2584
rect 68235 2624 68277 2633
rect 68235 2584 68236 2624
rect 68276 2584 68277 2624
rect 68235 2575 68277 2584
rect 68331 2624 68373 2633
rect 68331 2584 68332 2624
rect 68372 2584 68373 2624
rect 68331 2575 68373 2584
rect 68427 2624 68469 2633
rect 68427 2584 68428 2624
rect 68468 2584 68469 2624
rect 68427 2575 68469 2584
rect 68619 2624 68661 2633
rect 68619 2584 68620 2624
rect 68660 2584 68661 2624
rect 68619 2575 68661 2584
rect 68803 2624 68861 2625
rect 68803 2584 68812 2624
rect 68852 2584 68861 2624
rect 68803 2583 68861 2584
rect 68995 2624 69053 2625
rect 68995 2584 69004 2624
rect 69044 2584 69053 2624
rect 68995 2583 69053 2584
rect 69195 2624 69237 2633
rect 69195 2584 69196 2624
rect 69236 2584 69237 2624
rect 69195 2575 69237 2584
rect 71787 2624 71829 2633
rect 71787 2584 71788 2624
rect 71828 2584 71829 2624
rect 71787 2575 71829 2584
rect 71883 2624 71925 2633
rect 71883 2584 71884 2624
rect 71924 2584 71925 2624
rect 71883 2575 71925 2584
rect 71979 2624 72021 2633
rect 71979 2584 71980 2624
rect 72020 2584 72021 2624
rect 71979 2575 72021 2584
rect 72259 2624 72317 2625
rect 72259 2584 72268 2624
rect 72308 2584 72317 2624
rect 72259 2583 72317 2584
rect 72555 2624 72597 2633
rect 72555 2584 72556 2624
rect 72596 2584 72597 2624
rect 72555 2575 72597 2584
rect 72651 2624 72693 2633
rect 72651 2584 72652 2624
rect 72692 2584 72693 2624
rect 72651 2575 72693 2584
rect 73219 2624 73277 2625
rect 73219 2584 73228 2624
rect 73268 2584 73277 2624
rect 73219 2583 73277 2584
rect 74179 2624 74237 2625
rect 74179 2584 74188 2624
rect 74228 2584 74237 2624
rect 74179 2583 74237 2584
rect 74379 2624 74421 2633
rect 74379 2584 74380 2624
rect 74420 2584 74421 2624
rect 74379 2575 74421 2584
rect 74563 2624 74621 2625
rect 74563 2584 74572 2624
rect 74612 2584 74621 2624
rect 74563 2583 74621 2584
rect 75147 2624 75189 2633
rect 75147 2584 75148 2624
rect 75188 2584 75189 2624
rect 75147 2575 75189 2584
rect 75331 2624 75389 2625
rect 75331 2584 75340 2624
rect 75380 2584 75389 2624
rect 75331 2583 75389 2584
rect 76771 2624 76829 2625
rect 76771 2584 76780 2624
rect 76820 2584 76829 2624
rect 76771 2583 76829 2584
rect 77067 2624 77109 2633
rect 77067 2584 77068 2624
rect 77108 2584 77109 2624
rect 77067 2575 77109 2584
rect 77643 2624 77685 2633
rect 77643 2584 77644 2624
rect 77684 2584 77685 2624
rect 77643 2575 77685 2584
rect 77827 2624 77885 2625
rect 77827 2584 77836 2624
rect 77876 2584 77885 2624
rect 77827 2583 77885 2584
rect 2475 2540 2517 2549
rect 2475 2500 2476 2540
rect 2516 2500 2517 2540
rect 2475 2491 2517 2500
rect 59787 2540 59829 2549
rect 59787 2500 59788 2540
rect 59828 2500 59829 2540
rect 59787 2491 59829 2500
rect 69099 2540 69141 2549
rect 69099 2500 69100 2540
rect 69140 2500 69141 2540
rect 69099 2491 69141 2500
rect 74475 2540 74517 2549
rect 74475 2500 74476 2540
rect 74516 2500 74517 2540
rect 74475 2491 74517 2500
rect 75243 2540 75285 2549
rect 75243 2500 75244 2540
rect 75284 2500 75285 2540
rect 75243 2491 75285 2500
rect 77163 2540 77205 2549
rect 77163 2500 77164 2540
rect 77204 2500 77205 2540
rect 77163 2491 77205 2500
rect 77739 2540 77781 2549
rect 77739 2500 77740 2540
rect 77780 2500 77781 2540
rect 77739 2491 77781 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 2947 2456 3005 2457
rect 2947 2416 2956 2456
rect 2996 2416 3005 2456
rect 2947 2415 3005 2416
rect 55267 2456 55325 2457
rect 55267 2416 55276 2456
rect 55316 2416 55325 2456
rect 55267 2415 55325 2416
rect 55843 2456 55901 2457
rect 55843 2416 55852 2456
rect 55892 2416 55901 2456
rect 55843 2415 55901 2416
rect 56323 2456 56381 2457
rect 56323 2416 56332 2456
rect 56372 2416 56381 2456
rect 56323 2415 56381 2416
rect 64291 2456 64349 2457
rect 64291 2416 64300 2456
rect 64340 2416 64349 2456
rect 64291 2415 64349 2416
rect 68131 2456 68189 2457
rect 68131 2416 68140 2456
rect 68180 2416 68189 2456
rect 68131 2415 68189 2416
rect 71683 2456 71741 2457
rect 71683 2416 71692 2456
rect 71732 2416 71741 2456
rect 71683 2415 71741 2416
rect 576 2288 79584 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79584 2288
rect 576 2224 79584 2248
rect 55939 2120 55997 2121
rect 55939 2080 55948 2120
rect 55988 2080 55997 2120
rect 55939 2079 55997 2080
rect 58915 2120 58973 2121
rect 58915 2080 58924 2120
rect 58964 2080 58973 2120
rect 58915 2079 58973 2080
rect 61507 2120 61565 2121
rect 61507 2080 61516 2120
rect 61556 2080 61565 2120
rect 61507 2079 61565 2080
rect 64099 2120 64157 2121
rect 64099 2080 64108 2120
rect 64148 2080 64157 2120
rect 64099 2079 64157 2080
rect 66883 2120 66941 2121
rect 66883 2080 66892 2120
rect 66932 2080 66941 2120
rect 66883 2079 66941 2080
rect 71203 2120 71261 2121
rect 71203 2080 71212 2120
rect 71252 2080 71261 2120
rect 71203 2079 71261 2080
rect 73795 2120 73853 2121
rect 73795 2080 73804 2120
rect 73844 2080 73853 2120
rect 73795 2079 73853 2080
rect 78019 2120 78077 2121
rect 78019 2080 78028 2120
rect 78068 2080 78077 2120
rect 78019 2079 78077 2080
rect 56523 2036 56565 2045
rect 56523 1996 56524 2036
rect 56564 1996 56565 2036
rect 56523 1987 56565 1996
rect 53547 1952 53589 1961
rect 53547 1912 53548 1952
rect 53588 1912 53589 1952
rect 53547 1903 53589 1912
rect 53923 1952 53981 1953
rect 53923 1912 53932 1952
rect 53972 1912 53981 1952
rect 53923 1911 53981 1912
rect 54787 1952 54845 1953
rect 54787 1912 54796 1952
rect 54836 1912 54845 1952
rect 54787 1911 54845 1912
rect 56139 1952 56181 1961
rect 56139 1912 56140 1952
rect 56180 1912 56181 1952
rect 56139 1903 56181 1912
rect 56323 1952 56381 1953
rect 56323 1912 56332 1952
rect 56372 1912 56381 1952
rect 56323 1911 56381 1912
rect 56899 1952 56957 1953
rect 56899 1912 56908 1952
rect 56948 1912 56957 1952
rect 56899 1911 56957 1912
rect 57763 1952 57821 1953
rect 57763 1912 57772 1952
rect 57812 1912 57821 1952
rect 57763 1911 57821 1912
rect 59115 1952 59157 1961
rect 59115 1912 59116 1952
rect 59156 1912 59157 1952
rect 59115 1903 59157 1912
rect 59491 1952 59549 1953
rect 59491 1912 59500 1952
rect 59540 1912 59549 1952
rect 59491 1911 59549 1912
rect 60355 1952 60413 1953
rect 60355 1912 60364 1952
rect 60404 1912 60413 1952
rect 60355 1911 60413 1912
rect 61707 1952 61749 1961
rect 61707 1912 61708 1952
rect 61748 1912 61749 1952
rect 61707 1903 61749 1912
rect 62083 1952 62141 1953
rect 62083 1912 62092 1952
rect 62132 1912 62141 1952
rect 62083 1911 62141 1912
rect 62947 1952 63005 1953
rect 62947 1912 62956 1952
rect 62996 1912 63005 1952
rect 62947 1911 63005 1912
rect 64491 1952 64533 1961
rect 64491 1912 64492 1952
rect 64532 1912 64533 1952
rect 64491 1903 64533 1912
rect 64867 1952 64925 1953
rect 64867 1912 64876 1952
rect 64916 1912 64925 1952
rect 64867 1911 64925 1912
rect 65731 1952 65789 1953
rect 65731 1912 65740 1952
rect 65780 1912 65789 1952
rect 65731 1911 65789 1912
rect 67371 1952 67413 1961
rect 67371 1912 67372 1952
rect 67412 1912 67413 1952
rect 67371 1903 67413 1912
rect 67563 1952 67605 1961
rect 67563 1912 67564 1952
rect 67604 1912 67605 1952
rect 67563 1903 67605 1912
rect 67651 1952 67709 1953
rect 67651 1912 67660 1952
rect 67700 1912 67709 1952
rect 67651 1911 67709 1912
rect 67939 1952 67997 1953
rect 67939 1912 67948 1952
rect 67988 1912 67997 1952
rect 67939 1911 67997 1912
rect 68235 1952 68277 1961
rect 68235 1912 68236 1952
rect 68276 1912 68277 1952
rect 68235 1903 68277 1912
rect 68331 1952 68373 1961
rect 68331 1912 68332 1952
rect 68372 1912 68373 1952
rect 68331 1903 68373 1912
rect 68811 1952 68853 1961
rect 68811 1912 68812 1952
rect 68852 1912 68853 1952
rect 68811 1903 68853 1912
rect 69187 1952 69245 1953
rect 69187 1912 69196 1952
rect 69236 1912 69245 1952
rect 69187 1911 69245 1912
rect 70051 1952 70109 1953
rect 70051 1912 70060 1952
rect 70100 1912 70109 1952
rect 70051 1911 70109 1912
rect 71403 1952 71445 1961
rect 71403 1912 71404 1952
rect 71444 1912 71445 1952
rect 71403 1903 71445 1912
rect 71779 1952 71837 1953
rect 71779 1912 71788 1952
rect 71828 1912 71837 1952
rect 71779 1911 71837 1912
rect 72643 1952 72701 1953
rect 72643 1912 72652 1952
rect 72692 1912 72701 1952
rect 72643 1911 72701 1912
rect 73995 1952 74037 1961
rect 73995 1912 73996 1952
rect 74036 1912 74037 1952
rect 73995 1903 74037 1912
rect 74187 1952 74229 1961
rect 74187 1912 74188 1952
rect 74228 1912 74229 1952
rect 74187 1903 74229 1912
rect 74275 1952 74333 1953
rect 74275 1912 74284 1952
rect 74324 1912 74333 1952
rect 74275 1911 74333 1912
rect 74563 1952 74621 1953
rect 74563 1912 74572 1952
rect 74612 1912 74621 1952
rect 74563 1911 74621 1912
rect 74667 1952 74709 1961
rect 74667 1912 74668 1952
rect 74708 1912 74709 1952
rect 74667 1903 74709 1912
rect 74859 1952 74901 1961
rect 74859 1912 74860 1952
rect 74900 1912 74901 1952
rect 74859 1903 74901 1912
rect 75139 1952 75197 1953
rect 75139 1912 75148 1952
rect 75188 1912 75197 1952
rect 75139 1911 75197 1912
rect 75243 1952 75285 1961
rect 75243 1912 75244 1952
rect 75284 1912 75285 1952
rect 75243 1903 75285 1912
rect 75435 1952 75477 1961
rect 75435 1912 75436 1952
rect 75476 1912 75477 1952
rect 75435 1903 75477 1912
rect 75627 1952 75669 1961
rect 75627 1912 75628 1952
rect 75668 1912 75669 1952
rect 75627 1903 75669 1912
rect 76003 1952 76061 1953
rect 76003 1912 76012 1952
rect 76052 1912 76061 1952
rect 76003 1911 76061 1912
rect 76867 1952 76925 1953
rect 76867 1912 76876 1952
rect 76916 1912 76925 1952
rect 76867 1911 76925 1912
rect 78219 1952 78261 1961
rect 78219 1912 78220 1952
rect 78260 1912 78261 1952
rect 78219 1903 78261 1912
rect 78411 1952 78453 1961
rect 78411 1912 78412 1952
rect 78452 1912 78453 1952
rect 78411 1903 78453 1912
rect 78499 1952 78557 1953
rect 78499 1912 78508 1952
rect 78548 1912 78557 1952
rect 78499 1911 78557 1912
rect 78691 1952 78749 1953
rect 78691 1912 78700 1952
rect 78740 1912 78749 1952
rect 78691 1911 78749 1912
rect 78891 1952 78933 1961
rect 78891 1912 78892 1952
rect 78932 1912 78933 1952
rect 78891 1903 78933 1912
rect 68611 1784 68669 1785
rect 68611 1744 68620 1784
rect 68660 1744 68669 1784
rect 68611 1743 68669 1744
rect 74859 1784 74901 1793
rect 74859 1744 74860 1784
rect 74900 1744 74901 1784
rect 74859 1735 74901 1744
rect 75435 1784 75477 1793
rect 75435 1744 75436 1784
rect 75476 1744 75477 1784
rect 75435 1735 75477 1744
rect 78795 1784 78837 1793
rect 78795 1744 78796 1784
rect 78836 1744 78837 1784
rect 78795 1735 78837 1744
rect 55939 1700 55997 1701
rect 55939 1660 55948 1700
rect 55988 1660 55997 1700
rect 55939 1659 55997 1660
rect 56235 1700 56277 1709
rect 56235 1660 56236 1700
rect 56276 1660 56277 1700
rect 56235 1651 56277 1660
rect 58915 1700 58973 1701
rect 58915 1660 58924 1700
rect 58964 1660 58973 1700
rect 58915 1659 58973 1660
rect 61507 1700 61565 1701
rect 61507 1660 61516 1700
rect 61556 1660 61565 1700
rect 61507 1659 61565 1660
rect 64099 1700 64157 1701
rect 64099 1660 64108 1700
rect 64148 1660 64157 1700
rect 64099 1659 64157 1660
rect 67371 1700 67413 1709
rect 67371 1660 67372 1700
rect 67412 1660 67413 1700
rect 67371 1651 67413 1660
rect 73995 1700 74037 1709
rect 73995 1660 73996 1700
rect 74036 1660 74037 1700
rect 73995 1651 74037 1660
rect 78219 1700 78261 1709
rect 78219 1660 78220 1700
rect 78260 1660 78261 1700
rect 78219 1651 78261 1660
rect 576 1532 79584 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79584 1532
rect 576 1468 79584 1492
rect 55371 1364 55413 1373
rect 55371 1324 55372 1364
rect 55412 1324 55413 1364
rect 55371 1315 55413 1324
rect 55939 1364 55997 1365
rect 55939 1324 55948 1364
rect 55988 1324 55997 1364
rect 55939 1323 55997 1324
rect 59019 1364 59061 1373
rect 59019 1324 59020 1364
rect 59060 1324 59061 1364
rect 59019 1315 59061 1324
rect 62571 1364 62613 1373
rect 62571 1324 62572 1364
rect 62612 1324 62613 1364
rect 62571 1315 62613 1324
rect 68419 1364 68477 1365
rect 68419 1324 68428 1364
rect 68468 1324 68477 1364
rect 68419 1323 68477 1324
rect 68907 1364 68949 1373
rect 68907 1324 68908 1364
rect 68948 1324 68949 1364
rect 68907 1315 68949 1324
rect 70443 1364 70485 1373
rect 70443 1324 70444 1364
rect 70484 1324 70485 1364
rect 70443 1315 70485 1324
rect 72459 1364 72501 1373
rect 72459 1324 72460 1364
rect 72500 1324 72501 1364
rect 72459 1315 72501 1324
rect 77059 1364 77117 1365
rect 77059 1324 77068 1364
rect 77108 1324 77117 1364
rect 77059 1323 77117 1324
rect 57483 1280 57525 1289
rect 57483 1240 57484 1280
rect 57524 1240 57525 1280
rect 57483 1231 57525 1240
rect 60747 1280 60789 1289
rect 60747 1240 60748 1280
rect 60788 1240 60789 1280
rect 60747 1231 60789 1240
rect 61995 1280 62037 1289
rect 61995 1240 61996 1280
rect 62036 1240 62037 1280
rect 61995 1231 62037 1240
rect 64387 1280 64445 1281
rect 64387 1240 64396 1280
rect 64436 1240 64445 1280
rect 64387 1239 64445 1240
rect 64683 1280 64725 1289
rect 64683 1240 64684 1280
rect 64724 1240 64725 1280
rect 64683 1231 64725 1240
rect 64971 1280 65013 1289
rect 64971 1240 64972 1280
rect 65012 1240 65013 1280
rect 64971 1231 65013 1240
rect 69291 1280 69333 1289
rect 69291 1240 69292 1280
rect 69332 1240 69333 1280
rect 69291 1231 69333 1240
rect 60459 1196 60501 1205
rect 60459 1156 60460 1196
rect 60500 1156 60501 1196
rect 60459 1147 60501 1156
rect 55371 1112 55413 1121
rect 55371 1072 55372 1112
rect 55412 1072 55413 1112
rect 55371 1063 55413 1072
rect 55563 1112 55605 1121
rect 55563 1072 55564 1112
rect 55604 1072 55605 1112
rect 55563 1063 55605 1072
rect 55651 1112 55709 1113
rect 55651 1072 55660 1112
rect 55700 1072 55709 1112
rect 55651 1071 55709 1072
rect 56235 1112 56277 1121
rect 56235 1072 56236 1112
rect 56276 1072 56277 1112
rect 56235 1063 56277 1072
rect 56331 1112 56373 1121
rect 56331 1072 56332 1112
rect 56372 1072 56373 1112
rect 56331 1063 56373 1072
rect 56611 1112 56669 1113
rect 56611 1072 56620 1112
rect 56660 1072 56669 1112
rect 56611 1071 56669 1072
rect 57187 1112 57245 1113
rect 57187 1072 57196 1112
rect 57236 1072 57245 1112
rect 57187 1071 57245 1072
rect 57291 1112 57333 1121
rect 57291 1072 57292 1112
rect 57332 1072 57333 1112
rect 57291 1063 57333 1072
rect 57483 1112 57525 1121
rect 57483 1072 57484 1112
rect 57524 1072 57525 1112
rect 57483 1063 57525 1072
rect 58635 1112 58677 1121
rect 58635 1072 58636 1112
rect 58676 1072 58677 1112
rect 58635 1063 58677 1072
rect 58731 1112 58773 1121
rect 58731 1072 58732 1112
rect 58772 1072 58773 1112
rect 58731 1063 58773 1072
rect 58827 1112 58869 1121
rect 58827 1072 58828 1112
rect 58868 1072 58869 1112
rect 58827 1063 58869 1072
rect 59019 1112 59061 1121
rect 59019 1072 59020 1112
rect 59060 1072 59061 1112
rect 59019 1063 59061 1072
rect 59211 1112 59253 1121
rect 59211 1072 59212 1112
rect 59252 1072 59253 1112
rect 59211 1063 59253 1072
rect 59299 1112 59357 1113
rect 59299 1072 59308 1112
rect 59348 1072 59357 1112
rect 59299 1071 59357 1072
rect 59587 1112 59645 1113
rect 59587 1072 59596 1112
rect 59636 1072 59645 1112
rect 59587 1071 59645 1072
rect 61699 1112 61757 1113
rect 61699 1072 61708 1112
rect 61748 1072 61757 1112
rect 61699 1071 61757 1072
rect 61803 1112 61845 1121
rect 61803 1072 61804 1112
rect 61844 1072 61845 1112
rect 61803 1063 61845 1072
rect 61995 1112 62037 1121
rect 61995 1072 61996 1112
rect 62036 1072 62037 1112
rect 61995 1063 62037 1072
rect 62275 1112 62333 1113
rect 62275 1072 62284 1112
rect 62324 1072 62333 1112
rect 62275 1071 62333 1072
rect 62379 1112 62421 1121
rect 62379 1072 62380 1112
rect 62420 1072 62421 1112
rect 62379 1063 62421 1072
rect 62571 1112 62613 1121
rect 62571 1072 62572 1112
rect 62612 1072 62613 1112
rect 62571 1063 62613 1072
rect 62763 1112 62805 1121
rect 62763 1072 62764 1112
rect 62804 1072 62805 1112
rect 62763 1063 62805 1072
rect 62859 1112 62901 1121
rect 62859 1072 62860 1112
rect 62900 1072 62901 1112
rect 62859 1063 62901 1072
rect 62955 1112 62997 1121
rect 62955 1072 62956 1112
rect 62996 1072 62997 1112
rect 62955 1063 62997 1072
rect 63051 1112 63093 1121
rect 63051 1072 63052 1112
rect 63092 1072 63093 1112
rect 63051 1063 63093 1072
rect 63715 1112 63773 1113
rect 63715 1072 63724 1112
rect 63764 1072 63773 1112
rect 63715 1071 63773 1072
rect 64011 1112 64053 1121
rect 64011 1072 64012 1112
rect 64052 1072 64053 1112
rect 64011 1063 64053 1072
rect 64107 1112 64149 1121
rect 64107 1072 64108 1112
rect 64148 1072 64149 1112
rect 64107 1063 64149 1072
rect 64587 1112 64629 1121
rect 64587 1072 64588 1112
rect 64628 1072 64629 1112
rect 64587 1063 64629 1072
rect 64771 1112 64829 1113
rect 64771 1072 64780 1112
rect 64820 1072 64829 1112
rect 64771 1071 64829 1072
rect 66027 1112 66069 1121
rect 66027 1072 66028 1112
rect 66068 1072 66069 1112
rect 66027 1063 66069 1072
rect 66403 1112 66461 1113
rect 66403 1072 66412 1112
rect 66452 1072 66461 1112
rect 66403 1071 66461 1072
rect 67267 1112 67325 1113
rect 67267 1072 67276 1112
rect 67316 1072 67325 1112
rect 67267 1071 67325 1072
rect 68611 1112 68669 1113
rect 68611 1072 68620 1112
rect 68660 1072 68669 1112
rect 68611 1071 68669 1072
rect 68715 1112 68757 1121
rect 68715 1072 68716 1112
rect 68756 1072 68757 1112
rect 68715 1063 68757 1072
rect 68907 1112 68949 1121
rect 68907 1072 68908 1112
rect 68948 1072 68949 1112
rect 68907 1063 68949 1072
rect 69763 1112 69821 1113
rect 69763 1072 69772 1112
rect 69812 1072 69821 1112
rect 69763 1071 69821 1072
rect 70915 1112 70973 1113
rect 70915 1072 70924 1112
rect 70964 1072 70973 1112
rect 70915 1071 70973 1072
rect 71203 1112 71261 1113
rect 71203 1072 71212 1112
rect 71252 1072 71261 1112
rect 71203 1071 71261 1072
rect 72075 1112 72117 1121
rect 72075 1072 72076 1112
rect 72116 1072 72117 1112
rect 72075 1063 72117 1072
rect 72459 1112 72501 1121
rect 72459 1072 72460 1112
rect 72500 1072 72501 1112
rect 72459 1063 72501 1072
rect 72651 1112 72693 1121
rect 72651 1072 72652 1112
rect 72692 1072 72693 1112
rect 72651 1063 72693 1072
rect 72739 1112 72797 1113
rect 72739 1072 72748 1112
rect 72788 1072 72797 1112
rect 72739 1071 72797 1072
rect 74371 1112 74429 1113
rect 74371 1072 74380 1112
rect 74420 1072 74429 1112
rect 74371 1071 74429 1072
rect 75235 1112 75293 1113
rect 75235 1072 75244 1112
rect 75284 1072 75293 1112
rect 75235 1071 75293 1072
rect 75627 1112 75669 1121
rect 75627 1072 75628 1112
rect 75668 1072 75669 1112
rect 75627 1063 75669 1072
rect 75915 1112 75957 1121
rect 75915 1072 75916 1112
rect 75956 1072 75957 1112
rect 75915 1063 75957 1072
rect 76011 1112 76053 1121
rect 76011 1072 76012 1112
rect 76052 1072 76053 1112
rect 76011 1063 76053 1072
rect 76107 1112 76149 1121
rect 76107 1072 76108 1112
rect 76148 1072 76149 1112
rect 76107 1063 76149 1072
rect 76203 1112 76245 1121
rect 76203 1072 76204 1112
rect 76244 1072 76245 1112
rect 76203 1063 76245 1072
rect 78211 1112 78269 1113
rect 78211 1072 78220 1112
rect 78260 1072 78269 1112
rect 78211 1071 78269 1072
rect 79075 1112 79133 1113
rect 79075 1072 79084 1112
rect 79124 1072 79133 1112
rect 79075 1071 79133 1072
rect 79467 1112 79509 1121
rect 79467 1072 79468 1112
rect 79508 1072 79509 1112
rect 79467 1063 79509 1072
rect 58531 944 58589 945
rect 58531 904 58540 944
rect 58580 904 58589 944
rect 58531 903 58589 904
rect 73219 944 73277 945
rect 73219 904 73228 944
rect 73268 904 73277 944
rect 73219 903 73277 904
rect 576 776 79584 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79584 776
rect 576 712 79584 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 63436 38284 63476 38324
rect 63340 38189 63380 38229
rect 63532 38200 63572 38240
rect 63628 38200 63668 38240
rect 67468 38200 67508 38240
rect 67660 38200 67700 38240
rect 67756 38200 67796 38240
rect 67948 38200 67988 38240
rect 68044 38200 68084 38240
rect 68140 38200 68180 38240
rect 68236 38200 68276 38240
rect 69292 38200 69332 38240
rect 70636 38200 70676 38240
rect 71020 38200 71060 38240
rect 71212 38200 71252 38240
rect 74284 38200 74324 38240
rect 75244 38200 75284 38240
rect 76972 38200 77012 38240
rect 77260 38200 77300 38240
rect 77356 38200 77396 38240
rect 652 38116 692 38156
rect 58348 38116 58388 38156
rect 58924 38116 58964 38156
rect 59308 38116 59348 38156
rect 67084 38116 67124 38156
rect 56908 38032 56948 38072
rect 58540 38032 58580 38072
rect 61612 38032 61652 38072
rect 64204 38032 64244 38072
rect 66508 38032 66548 38072
rect 71404 38032 71444 38072
rect 71980 38032 72020 38072
rect 75916 38032 75956 38072
rect 844 37948 884 37988
rect 58732 37948 58772 37988
rect 59116 37948 59156 37988
rect 67276 37948 67316 37988
rect 67468 37948 67508 37988
rect 69100 37948 69140 37988
rect 70060 37948 70100 37988
rect 71116 37948 71156 37988
rect 77644 37948 77684 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 55180 37528 55220 37568
rect 59788 37528 59828 37568
rect 74284 37528 74324 37568
rect 78412 37528 78452 37568
rect 55756 37360 55796 37400
rect 55948 37360 55988 37400
rect 56044 37360 56084 37400
rect 57388 37360 57428 37400
rect 58252 37360 58292 37400
rect 58828 37360 58868 37400
rect 58924 37360 58964 37400
rect 59020 37360 59060 37400
rect 59116 37360 59156 37400
rect 59308 37360 59348 37400
rect 59500 37360 59540 37400
rect 59596 37360 59636 37400
rect 60172 37360 60212 37400
rect 60364 37360 60404 37400
rect 60460 37362 60500 37402
rect 61516 37360 61556 37400
rect 62380 37360 62420 37400
rect 63724 37360 63764 37400
rect 64108 37360 64148 37400
rect 64972 37360 65012 37400
rect 66316 37360 66356 37400
rect 66700 37360 66740 37400
rect 67564 37360 67604 37400
rect 69580 37360 69620 37400
rect 70444 37360 70484 37400
rect 72844 37360 72884 37400
rect 72940 37360 72980 37400
rect 73036 37360 73076 37400
rect 73132 37360 73172 37400
rect 73324 37360 73364 37400
rect 73516 37360 73556 37400
rect 73612 37360 73652 37400
rect 73804 37360 73844 37400
rect 73996 37360 74036 37400
rect 74092 37360 74132 37400
rect 74284 37360 74324 37400
rect 74476 37360 74516 37400
rect 74572 37360 74612 37400
rect 74956 37360 74996 37400
rect 75052 37360 75092 37400
rect 75148 37360 75188 37400
rect 75820 37360 75860 37400
rect 76684 37360 76724 37400
rect 78028 37360 78068 37400
rect 78220 37360 78260 37400
rect 58636 37276 58676 37316
rect 59404 37276 59444 37316
rect 60268 37276 60308 37316
rect 61132 37276 61172 37316
rect 69196 37276 69236 37316
rect 75436 37276 75476 37316
rect 78124 37276 78164 37316
rect 55852 37192 55892 37232
rect 56236 37192 56276 37232
rect 63532 37192 63572 37232
rect 66124 37192 66164 37232
rect 68716 37192 68756 37232
rect 71596 37192 71636 37232
rect 73420 37192 73460 37232
rect 73900 37192 73940 37232
rect 75244 37192 75284 37232
rect 77836 37192 77876 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 62284 36856 62324 36896
rect 67948 36856 67988 36896
rect 79468 36856 79508 36896
rect 54700 36772 54740 36812
rect 58444 36772 58484 36812
rect 63340 36772 63380 36812
rect 63916 36772 63956 36812
rect 64300 36772 64340 36812
rect 73324 36772 73364 36812
rect 73516 36772 73556 36812
rect 55084 36688 55124 36728
rect 55948 36688 55988 36728
rect 57292 36688 57332 36728
rect 57484 36688 57524 36728
rect 57580 36688 57620 36728
rect 58540 36688 58580 36728
rect 58828 36688 58868 36728
rect 59116 36688 59156 36728
rect 59500 36688 59540 36728
rect 60364 36688 60404 36728
rect 61708 36688 61748 36728
rect 61804 36688 61844 36728
rect 61900 36688 61940 36728
rect 61996 36688 62036 36728
rect 62188 36688 62228 36728
rect 62380 36688 62420 36728
rect 62476 36688 62516 36728
rect 62956 36688 62996 36728
rect 63244 36688 63284 36728
rect 63820 36688 63860 36728
rect 64012 36688 64052 36728
rect 64204 36688 64244 36728
rect 64396 36688 64436 36728
rect 66508 36688 66548 36728
rect 66700 36688 66740 36728
rect 66796 36688 66836 36728
rect 67180 36688 67220 36728
rect 67372 36688 67412 36728
rect 67468 36688 67508 36728
rect 68236 36688 68276 36728
rect 68524 36688 68564 36728
rect 68620 36688 68660 36728
rect 69100 36688 69140 36728
rect 69292 36688 69332 36728
rect 69388 36688 69428 36728
rect 69580 36688 69620 36728
rect 69772 36688 69812 36728
rect 72076 36688 72116 36728
rect 72940 36688 72980 36728
rect 73900 36688 73940 36728
rect 74764 36688 74804 36728
rect 76108 36688 76148 36728
rect 76300 36688 76340 36728
rect 76396 36688 76436 36728
rect 76588 36688 76628 36728
rect 76780 36688 76820 36728
rect 76876 36688 76916 36728
rect 77068 36688 77108 36728
rect 77452 36688 77492 36728
rect 78316 36688 78356 36728
rect 67756 36604 67796 36644
rect 52492 36520 52532 36560
rect 57292 36520 57332 36560
rect 63628 36520 63668 36560
rect 67180 36520 67220 36560
rect 68908 36520 68948 36560
rect 69676 36520 69716 36560
rect 76108 36520 76148 36560
rect 76588 36520 76628 36560
rect 57100 36436 57140 36476
rect 58156 36436 58196 36476
rect 61516 36436 61556 36476
rect 66508 36436 66548 36476
rect 67948 36436 67988 36476
rect 69100 36436 69140 36476
rect 70924 36436 70964 36476
rect 75916 36436 75956 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 62284 36100 62324 36140
rect 73804 36100 73844 36140
rect 77548 36100 77588 36140
rect 49228 36016 49268 36056
rect 60364 36016 60404 36056
rect 69484 36016 69524 36056
rect 73516 36016 73556 36056
rect 74092 36016 74132 36056
rect 77836 36016 77876 36056
rect 50956 35932 50996 35972
rect 57100 35932 57140 35972
rect 51340 35848 51380 35888
rect 51532 35848 51572 35888
rect 52396 35848 52436 35888
rect 53285 35848 53325 35888
rect 55564 35848 55604 35888
rect 55660 35848 55700 35888
rect 55852 35848 55892 35888
rect 56044 35848 56084 35888
rect 56140 35848 56180 35888
rect 56236 35848 56276 35888
rect 56332 35848 56372 35888
rect 56524 35848 56564 35888
rect 56620 35848 56660 35888
rect 56716 35848 56756 35888
rect 58540 35848 58580 35888
rect 58636 35848 58676 35888
rect 58732 35848 58772 35888
rect 58924 35848 58964 35888
rect 59116 35848 59156 35888
rect 59212 35848 59252 35888
rect 59404 35848 59444 35888
rect 59596 35848 59636 35888
rect 61996 35848 62036 35888
rect 62092 35848 62132 35888
rect 62284 35848 62324 35888
rect 64396 35848 64436 35888
rect 64780 35848 64820 35888
rect 65644 35848 65684 35888
rect 66988 35848 67028 35888
rect 67084 35848 67124 35888
rect 67180 35848 67220 35888
rect 67276 35848 67316 35888
rect 69676 35848 69716 35888
rect 69868 35848 69908 35888
rect 69964 35848 70004 35888
rect 71500 35848 71540 35888
rect 71692 35848 71732 35888
rect 71884 35848 71924 35888
rect 72076 35848 72116 35888
rect 72172 35848 72212 35888
rect 72844 35848 72884 35888
rect 73132 35848 73172 35888
rect 73228 35848 73268 35888
rect 73708 35848 73748 35888
rect 73900 35848 73940 35888
rect 76204 35848 76244 35888
rect 76396 35848 76436 35888
rect 76492 35848 76532 35888
rect 77068 35848 77108 35888
rect 77260 35848 77300 35888
rect 77452 35848 77492 35888
rect 77644 35848 77684 35888
rect 51436 35764 51476 35804
rect 52012 35764 52052 35804
rect 59020 35764 59060 35804
rect 59500 35764 59540 35804
rect 69772 35764 69812 35804
rect 71596 35764 71636 35804
rect 76300 35764 76340 35804
rect 77164 35764 77204 35804
rect 50764 35680 50804 35720
rect 54412 35680 54452 35720
rect 55756 35680 55796 35720
rect 56908 35680 56948 35720
rect 66796 35680 66836 35720
rect 71980 35680 72020 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 52204 35344 52244 35384
rect 76588 35344 76628 35384
rect 52684 35260 52724 35300
rect 54892 35260 54932 35300
rect 55180 35260 55220 35300
rect 66028 35260 66068 35300
rect 71308 35260 71348 35300
rect 73420 35260 73460 35300
rect 49708 35176 49748 35216
rect 50572 35176 50612 35216
rect 50956 35176 50996 35216
rect 51436 35176 51476 35216
rect 51532 35176 51572 35216
rect 51820 35176 51860 35216
rect 52108 35176 52148 35216
rect 52300 35176 52340 35216
rect 52396 35176 52436 35216
rect 52588 35176 52628 35216
rect 52780 35176 52820 35216
rect 54796 35176 54836 35216
rect 54988 35176 55028 35216
rect 55564 35176 55604 35216
rect 56428 35176 56468 35216
rect 57772 35176 57812 35216
rect 57964 35176 58004 35216
rect 58060 35176 58100 35216
rect 59884 35176 59924 35216
rect 60268 35176 60308 35216
rect 61132 35176 61172 35216
rect 62764 35176 62804 35216
rect 62860 35176 62900 35216
rect 63148 35176 63188 35216
rect 65932 35176 65972 35216
rect 66124 35176 66164 35216
rect 66604 35176 66644 35216
rect 66700 35176 66740 35216
rect 66988 35176 67028 35216
rect 67276 35176 67316 35216
rect 67660 35176 67700 35216
rect 68524 35176 68564 35216
rect 70348 35176 70388 35216
rect 70444 35176 70484 35216
rect 70540 35176 70580 35216
rect 70636 35176 70676 35216
rect 70924 35176 70964 35216
rect 71212 35176 71252 35216
rect 71788 35176 71828 35216
rect 71980 35176 72020 35216
rect 72076 35176 72116 35216
rect 73324 35176 73364 35216
rect 73516 35176 73556 35216
rect 74188 35176 74228 35216
rect 74572 35176 74612 35216
rect 75436 35176 75476 35216
rect 77068 35176 77108 35216
rect 77452 35176 77492 35216
rect 78316 35176 78356 35216
rect 47116 35008 47156 35048
rect 51148 35008 51188 35048
rect 58444 35008 58484 35048
rect 63628 35008 63668 35048
rect 64876 35008 64916 35048
rect 66316 35008 66356 35048
rect 71596 35008 71636 35048
rect 72556 35008 72596 35048
rect 48556 34924 48596 34964
rect 57580 34924 57620 34964
rect 57772 34924 57812 34964
rect 62284 34924 62324 34964
rect 62476 34924 62516 34964
rect 69676 34924 69716 34964
rect 71788 34924 71828 34964
rect 76588 34924 76628 34964
rect 79468 34924 79508 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 50956 34588 50996 34628
rect 56524 34588 56564 34628
rect 66892 34588 66932 34628
rect 68812 34588 68852 34628
rect 77260 34588 77300 34628
rect 46444 34504 46484 34544
rect 49228 34504 49268 34544
rect 52012 34504 52052 34544
rect 52204 34504 52244 34544
rect 55564 34504 55604 34544
rect 57772 34504 57812 34544
rect 61996 34504 62036 34544
rect 67468 34504 67508 34544
rect 67756 34504 67796 34544
rect 71884 34504 71924 34544
rect 74668 34504 74708 34544
rect 76012 34504 76052 34544
rect 77452 34504 77492 34544
rect 46156 34336 46196 34376
rect 46252 34336 46292 34376
rect 46444 34336 46484 34376
rect 46636 34336 46676 34376
rect 47020 34336 47060 34376
rect 47884 34336 47924 34376
rect 49228 34336 49268 34376
rect 49420 34336 49460 34376
rect 49516 34336 49556 34376
rect 50476 34336 50516 34376
rect 50572 34336 50612 34376
rect 50668 34336 50708 34376
rect 50764 34336 50804 34376
rect 50956 34336 50996 34376
rect 51148 34336 51188 34376
rect 51244 34336 51284 34376
rect 52204 34336 52244 34376
rect 52396 34336 52436 34376
rect 52492 34336 52532 34376
rect 53836 34336 53876 34376
rect 54028 34336 54068 34376
rect 54124 34336 54164 34376
rect 55852 34336 55892 34376
rect 56140 34336 56180 34376
rect 57484 34336 57524 34376
rect 57580 34336 57620 34376
rect 57772 34336 57812 34376
rect 57964 34336 58004 34376
rect 58348 34336 58388 34376
rect 59212 34336 59252 34376
rect 61516 34336 61556 34376
rect 61612 34336 61652 34376
rect 61708 34336 61748 34376
rect 61804 34336 61844 34376
rect 61996 34336 62036 34376
rect 62188 34336 62228 34376
rect 62284 34336 62324 34376
rect 62668 34336 62708 34376
rect 62860 34336 62900 34376
rect 62956 34336 62996 34376
rect 63532 34336 63572 34376
rect 64396 34336 64436 34376
rect 66124 34336 66164 34376
rect 66316 34336 66356 34376
rect 66412 34336 66452 34376
rect 66892 34336 66932 34376
rect 67084 34336 67124 34376
rect 67180 34336 67220 34376
rect 67372 34336 67412 34376
rect 67564 34336 67604 34376
rect 69964 34336 70004 34376
rect 70828 34336 70868 34376
rect 71212 34336 71252 34376
rect 71596 34336 71636 34376
rect 71692 34336 71732 34376
rect 71884 34336 71924 34376
rect 72076 34336 72116 34376
rect 72460 34336 72500 34376
rect 73324 34336 73364 34376
rect 75628 34336 75668 34376
rect 75724 34336 75764 34376
rect 75820 34336 75860 34376
rect 76012 34336 76052 34376
rect 76204 34336 76244 34376
rect 76300 34336 76340 34376
rect 76588 34336 76628 34376
rect 76876 34336 76916 34376
rect 76972 34336 77012 34376
rect 77452 34336 77492 34376
rect 77644 34336 77684 34376
rect 77740 34336 77780 34376
rect 77932 34336 77972 34376
rect 78124 34336 78164 34376
rect 56236 34252 56276 34292
rect 62764 34252 62804 34292
rect 63148 34252 63188 34292
rect 78028 34252 78068 34292
rect 49036 34168 49076 34208
rect 53932 34168 53972 34208
rect 60364 34168 60404 34208
rect 65548 34168 65588 34208
rect 66220 34168 66260 34208
rect 74476 34168 74516 34208
rect 75532 34168 75572 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 46732 33832 46772 33872
rect 58348 33832 58388 33872
rect 62284 33832 62324 33872
rect 51628 33748 51668 33788
rect 62764 33748 62804 33788
rect 63148 33748 63188 33788
rect 66220 33748 66260 33788
rect 71692 33748 71732 33788
rect 46828 33664 46868 33704
rect 46924 33664 46964 33704
rect 47020 33664 47060 33704
rect 49228 33664 49268 33704
rect 49420 33664 49460 33704
rect 49516 33664 49556 33704
rect 52012 33664 52052 33704
rect 52876 33664 52916 33704
rect 54316 33664 54356 33704
rect 54604 33664 54644 33704
rect 54700 33664 54740 33704
rect 55180 33664 55220 33704
rect 55276 33664 55316 33704
rect 55372 33664 55412 33704
rect 58444 33664 58484 33704
rect 58540 33664 58580 33704
rect 58636 33664 58676 33704
rect 58828 33664 58868 33704
rect 59020 33664 59060 33704
rect 62188 33664 62228 33704
rect 62380 33664 62420 33704
rect 62476 33664 62516 33704
rect 62668 33664 62708 33704
rect 62860 33664 62900 33704
rect 63052 33664 63092 33704
rect 63244 33664 63284 33704
rect 66124 33664 66164 33704
rect 66316 33664 66356 33704
rect 66412 33664 66452 33704
rect 66604 33664 66644 33704
rect 66796 33664 66836 33704
rect 71596 33664 71636 33704
rect 71788 33664 71828 33704
rect 71980 33664 72020 33704
rect 72172 33664 72212 33704
rect 72268 33664 72308 33704
rect 72460 33664 72500 33704
rect 72556 33664 72596 33704
rect 72652 33664 72692 33704
rect 75724 33664 75764 33704
rect 75820 33664 75860 33704
rect 76012 33664 76052 33704
rect 76204 33664 76244 33704
rect 76300 33664 76340 33704
rect 76396 33664 76436 33704
rect 76492 33664 76532 33704
rect 76684 33664 76724 33704
rect 76876 33664 76916 33704
rect 76972 33664 77012 33704
rect 77260 33664 77300 33704
rect 77452 33664 77492 33704
rect 77548 33664 77588 33704
rect 54028 33580 54068 33620
rect 48844 33496 48884 33536
rect 54988 33496 55028 33536
rect 55852 33496 55892 33536
rect 59212 33496 59252 33536
rect 63724 33496 63764 33536
rect 66988 33496 67028 33536
rect 69868 33496 69908 33536
rect 72844 33496 72884 33536
rect 75148 33496 75188 33536
rect 77836 33496 77876 33536
rect 49228 33412 49268 33452
rect 58924 33412 58964 33452
rect 66700 33412 66740 33452
rect 71980 33412 72020 33452
rect 76012 33412 76052 33452
rect 76684 33412 76724 33452
rect 77260 33412 77300 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 60940 33076 60980 33116
rect 77164 33076 77204 33116
rect 78412 33076 78452 33116
rect 43852 32992 43892 33032
rect 47116 32992 47156 33032
rect 47308 32992 47348 33032
rect 52300 32992 52340 33032
rect 55084 32992 55124 33032
rect 61132 32992 61172 33032
rect 78124 32992 78164 33032
rect 42700 32908 42740 32948
rect 47788 32908 47828 32948
rect 45868 32824 45908 32864
rect 46060 32824 46100 32864
rect 46156 32824 46196 32864
rect 46444 32824 46484 32864
rect 46732 32824 46772 32864
rect 46828 32824 46868 32864
rect 47692 32824 47732 32864
rect 47884 32824 47924 32864
rect 48460 32824 48500 32864
rect 48844 32824 48884 32864
rect 49708 32824 49748 32864
rect 51052 32824 51092 32864
rect 51244 32824 51284 32864
rect 52588 32824 52628 32864
rect 53452 32824 53492 32864
rect 53548 32824 53588 32864
rect 53644 32824 53684 32864
rect 53740 32824 53780 32864
rect 54412 32824 54452 32864
rect 54508 32824 54548 32864
rect 54604 32824 54644 32864
rect 54796 32824 54836 32864
rect 54892 32824 54932 32864
rect 55084 32824 55124 32864
rect 55276 32824 55316 32864
rect 55660 32824 55700 32864
rect 56524 32824 56564 32864
rect 58060 32824 58100 32864
rect 58252 32824 58292 32864
rect 58348 32824 58388 32864
rect 58924 32824 58964 32864
rect 59788 32824 59828 32864
rect 62476 32824 62516 32864
rect 62572 32824 62612 32864
rect 62668 32824 62708 32864
rect 62860 32824 62900 32864
rect 63052 32824 63092 32864
rect 63628 32824 63668 32864
rect 64492 32824 64532 32864
rect 65836 32824 65876 32864
rect 65932 32824 65972 32864
rect 66028 32824 66068 32864
rect 66124 32824 66164 32864
rect 66316 32824 66356 32864
rect 66700 32824 66740 32864
rect 67564 32824 67604 32864
rect 68908 32824 68948 32864
rect 69004 32824 69044 32864
rect 69196 32835 69236 32875
rect 69772 32824 69812 32864
rect 70636 32824 70676 32864
rect 72172 32824 72212 32864
rect 72556 32824 72596 32864
rect 73420 32824 73460 32864
rect 74764 32824 74804 32864
rect 75148 32824 75188 32864
rect 76012 32824 76052 32864
rect 77452 32824 77492 32864
rect 77740 32824 77780 32864
rect 77836 32824 77876 32864
rect 78316 32824 78356 32864
rect 78508 32824 78548 32864
rect 51148 32740 51188 32780
rect 58156 32740 58196 32780
rect 58540 32740 58580 32780
rect 62956 32740 62996 32780
rect 63244 32740 63284 32780
rect 69388 32740 69428 32780
rect 42892 32656 42932 32696
rect 45964 32656 46004 32696
rect 50860 32656 50900 32696
rect 57676 32656 57716 32696
rect 60940 32656 60980 32696
rect 62380 32656 62420 32696
rect 65644 32656 65684 32696
rect 68716 32656 68756 32696
rect 69100 32656 69140 32696
rect 71788 32656 71828 32696
rect 74572 32656 74612 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 48652 32320 48692 32360
rect 66508 32362 66548 32402
rect 49612 32320 49652 32360
rect 53548 32320 53588 32360
rect 62764 32320 62804 32360
rect 64012 32320 64052 32360
rect 75916 32320 75956 32360
rect 46060 32236 46100 32276
rect 50476 32236 50516 32276
rect 58732 32236 58772 32276
rect 66220 32236 66260 32276
rect 72076 32236 72116 32276
rect 77068 32236 77108 32276
rect 42316 32152 42356 32192
rect 42412 32152 42452 32192
rect 42508 32152 42548 32192
rect 42604 32152 42644 32192
rect 42892 32152 42932 32192
rect 43084 32152 43124 32192
rect 43372 32152 43412 32192
rect 43756 32152 43796 32192
rect 44620 32152 44660 32192
rect 46444 32152 46484 32192
rect 47308 32152 47348 32192
rect 48748 32152 48788 32192
rect 48844 32152 48884 32192
rect 48940 32152 48980 32192
rect 49132 32152 49172 32192
rect 50092 32152 50132 32192
rect 50380 32152 50420 32192
rect 50572 32152 50612 32192
rect 51148 32152 51188 32192
rect 51532 32152 51572 32192
rect 52396 32152 52436 32192
rect 54220 32152 54260 32192
rect 54412 32152 54452 32192
rect 54508 32152 54548 32192
rect 54700 32152 54740 32192
rect 54796 32152 54836 32192
rect 54892 32152 54932 32192
rect 54988 32152 55028 32192
rect 55660 32152 55700 32192
rect 55852 32152 55892 32192
rect 58348 32152 58388 32192
rect 58636 32152 58676 32192
rect 59212 32152 59252 32192
rect 59404 32152 59444 32192
rect 59596 32152 59636 32192
rect 59692 32152 59732 32192
rect 59884 32152 59924 32192
rect 60364 32152 60404 32192
rect 60748 32152 60788 32192
rect 61612 32152 61652 32192
rect 63244 32152 63284 32192
rect 63340 32179 63380 32219
rect 63628 32152 63668 32192
rect 63916 32152 63956 32192
rect 64108 32152 64148 32192
rect 64204 32152 64244 32192
rect 64396 32152 64436 32192
rect 64588 32152 64628 32192
rect 65836 32152 65876 32192
rect 66124 32152 66164 32192
rect 66700 32152 66740 32192
rect 67084 32152 67124 32192
rect 67948 32152 67988 32192
rect 69772 32152 69812 32192
rect 69868 32152 69908 32192
rect 70060 32152 70100 32192
rect 70252 32152 70292 32192
rect 70348 32152 70388 32192
rect 70444 32152 70484 32192
rect 70540 32152 70580 32192
rect 70732 32152 70772 32192
rect 70924 32152 70964 32192
rect 71020 32152 71060 32192
rect 71692 32152 71732 32192
rect 71980 32152 72020 32192
rect 72556 32152 72596 32192
rect 72748 32152 72788 32192
rect 75820 32152 75860 32192
rect 76012 32152 76052 32192
rect 76108 32152 76148 32192
rect 77452 32152 77492 32192
rect 78316 32152 78356 32192
rect 40684 31984 40724 32024
rect 54220 31984 54260 32024
rect 59020 31984 59060 32024
rect 59308 31984 59348 32024
rect 62956 31984 62996 32024
rect 64492 31984 64532 32024
rect 70060 31984 70100 32024
rect 72364 31984 72404 32024
rect 74092 31984 74132 32024
rect 42988 31900 43028 31940
rect 45772 31900 45812 31940
rect 48460 31900 48500 31940
rect 53548 31900 53588 31940
rect 55756 31900 55796 31940
rect 59884 31900 59924 31940
rect 69100 31900 69140 31940
rect 70732 31900 70772 31940
rect 72652 31900 72692 31940
rect 79468 31900 79508 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 42796 31564 42836 31604
rect 44044 31564 44084 31604
rect 46732 31564 46772 31604
rect 49228 31564 49268 31604
rect 50188 31564 50228 31604
rect 51436 31564 51476 31604
rect 55276 31564 55316 31604
rect 60268 31564 60308 31604
rect 60844 31564 60884 31604
rect 66316 31564 66356 31604
rect 71404 31564 71444 31604
rect 72076 31564 72116 31604
rect 76012 31564 76052 31604
rect 77932 31564 77972 31604
rect 51628 31480 51668 31520
rect 63052 31480 63092 31520
rect 63532 31480 63572 31520
rect 66892 31480 66932 31520
rect 67180 31480 67220 31520
rect 68716 31480 68756 31520
rect 71116 31480 71156 31520
rect 72268 31480 72308 31520
rect 60076 31396 60116 31436
rect 60652 31396 60692 31436
rect 71884 31396 71924 31436
rect 40588 31312 40628 31352
rect 41452 31312 41492 31352
rect 43180 31285 43220 31325
rect 43468 31312 43508 31352
rect 43756 31312 43796 31352
rect 43852 31312 43892 31352
rect 44044 31312 44084 31352
rect 46636 31312 46676 31352
rect 46828 31312 46868 31352
rect 48556 31312 48596 31352
rect 48940 31312 48980 31352
rect 49036 31312 49076 31352
rect 49228 31312 49268 31352
rect 49708 31312 49748 31352
rect 49900 31312 49940 31352
rect 49996 31312 50036 31352
rect 50476 31312 50516 31352
rect 50572 31312 50612 31352
rect 50860 31312 50900 31352
rect 51148 31312 51188 31352
rect 51244 31312 51284 31352
rect 51436 31312 51476 31352
rect 53260 31299 53300 31339
rect 54124 31312 54164 31352
rect 55660 31312 55700 31352
rect 55852 31312 55892 31352
rect 55948 31312 55988 31352
rect 56524 31312 56564 31352
rect 57388 31312 57428 31352
rect 59596 31312 59636 31352
rect 59692 31312 59732 31352
rect 59788 31312 59828 31352
rect 62476 31312 62516 31352
rect 62668 31312 62708 31352
rect 62764 31312 62804 31352
rect 40204 31228 40244 31268
rect 43084 31228 43124 31268
rect 52876 31228 52916 31268
rect 56140 31228 56180 31268
rect 62572 31228 62612 31268
rect 63052 31274 63092 31314
rect 63244 31312 63284 31352
rect 63340 31297 63380 31337
rect 66316 31312 66356 31352
rect 66508 31312 66548 31352
rect 66604 31312 66644 31352
rect 66796 31312 66836 31352
rect 66988 31312 67028 31352
rect 70540 31312 70580 31352
rect 70732 31312 70772 31352
rect 70828 31312 70868 31352
rect 71020 31312 71060 31352
rect 71212 31312 71252 31352
rect 71404 31312 71444 31352
rect 71596 31312 71636 31352
rect 71692 31297 71732 31337
rect 73996 31312 74036 31352
rect 74860 31312 74900 31352
rect 76972 31312 77012 31352
rect 77164 31312 77204 31352
rect 77452 31312 77492 31352
rect 77644 31312 77684 31352
rect 77836 31312 77876 31352
rect 78028 31312 78068 31352
rect 73612 31228 73652 31268
rect 77068 31228 77108 31268
rect 77548 31228 77588 31268
rect 42604 31144 42644 31184
rect 49804 31144 49844 31184
rect 55276 31144 55316 31184
rect 55756 31144 55796 31184
rect 58540 31144 58580 31184
rect 59884 31144 59924 31184
rect 60268 31144 60308 31184
rect 60844 31144 60884 31184
rect 70636 31144 70676 31184
rect 76012 31144 76052 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 42508 30808 42548 30848
rect 42796 30808 42836 30848
rect 49228 30808 49268 30848
rect 50380 30808 50420 30848
rect 51532 30808 51572 30848
rect 57964 30808 58004 30848
rect 70828 30808 70868 30848
rect 76876 30850 76916 30890
rect 71500 30808 71540 30848
rect 74860 30808 74900 30848
rect 75436 30808 75476 30848
rect 79468 30808 79508 30848
rect 43276 30724 43316 30764
rect 55564 30724 55604 30764
rect 56140 30724 56180 30764
rect 68236 30724 68276 30764
rect 71692 30724 71732 30764
rect 41452 30640 41492 30680
rect 41644 30640 41684 30680
rect 41740 30640 41780 30680
rect 42700 30640 42740 30680
rect 42892 30640 42932 30680
rect 42988 30640 43028 30680
rect 43179 30661 43219 30701
rect 43372 30640 43412 30680
rect 43756 30640 43796 30680
rect 43948 30640 43988 30680
rect 44044 30640 44084 30680
rect 44620 30640 44660 30680
rect 44716 30640 44756 30680
rect 44812 30640 44852 30680
rect 44908 30640 44948 30680
rect 46060 30640 46100 30680
rect 46252 30640 46292 30680
rect 46348 30640 46388 30680
rect 49612 30640 49652 30680
rect 49708 30640 49748 30680
rect 49804 30640 49844 30680
rect 49900 30640 49940 30680
rect 50572 30640 50612 30680
rect 50764 30640 50804 30680
rect 50956 30640 50996 30680
rect 51159 30661 51199 30701
rect 54604 30640 54644 30680
rect 54796 30640 54836 30680
rect 54892 30640 54932 30680
rect 55180 30640 55220 30680
rect 55468 30640 55508 30680
rect 56044 30617 56084 30657
rect 56236 30640 56276 30680
rect 59116 30640 59156 30680
rect 59980 30640 60020 30680
rect 60364 30640 60404 30680
rect 60556 30640 60596 30680
rect 60748 30640 60788 30680
rect 60844 30640 60884 30680
rect 61036 30640 61076 30680
rect 61228 30640 61268 30680
rect 63052 30640 63092 30680
rect 63436 30640 63476 30680
rect 64300 30640 64340 30680
rect 65644 30661 65684 30701
rect 65836 30640 65876 30680
rect 66028 30640 66068 30680
rect 66220 30640 66260 30680
rect 68620 30640 68660 30680
rect 69484 30640 69524 30680
rect 70924 30640 70964 30680
rect 71020 30640 71060 30680
rect 71116 30640 71156 30680
rect 72076 30640 72116 30680
rect 72940 30640 72980 30680
rect 74956 30640 74996 30680
rect 75052 30640 75092 30680
rect 75148 30640 75188 30680
rect 75340 30640 75380 30680
rect 75532 30640 75572 30680
rect 75628 30640 75668 30680
rect 76204 30640 76244 30680
rect 76492 30640 76532 30680
rect 76588 30640 76628 30680
rect 77068 30640 77108 30680
rect 77452 30640 77492 30680
rect 78316 30640 78356 30680
rect 40876 30556 40916 30596
rect 42316 30556 42356 30596
rect 49420 30556 49460 30596
rect 50188 30556 50228 30596
rect 51340 30556 51380 30596
rect 71308 30556 71348 30596
rect 43756 30472 43796 30512
rect 44236 30472 44276 30512
rect 46828 30472 46868 30512
rect 48268 30472 48308 30512
rect 51724 30472 51764 30512
rect 53356 30472 53396 30512
rect 54604 30472 54644 30512
rect 55852 30472 55892 30512
rect 56620 30472 56660 30512
rect 60556 30472 60596 30512
rect 61420 30472 61460 30512
rect 66508 30472 66548 30512
rect 40684 30388 40724 30428
rect 41452 30388 41492 30428
rect 42508 30388 42548 30428
rect 46060 30388 46100 30428
rect 50380 30388 50420 30428
rect 50668 30388 50708 30428
rect 51052 30388 51092 30428
rect 61132 30388 61172 30428
rect 65452 30388 65492 30428
rect 65740 30388 65780 30428
rect 66124 30388 66164 30428
rect 70636 30388 70676 30428
rect 71500 30388 71540 30428
rect 74092 30388 74132 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 40204 30052 40244 30092
rect 45868 30052 45908 30092
rect 47116 30052 47156 30092
rect 50188 30052 50228 30092
rect 54892 30052 54932 30092
rect 62956 30052 62996 30092
rect 63628 30052 63668 30092
rect 65836 30052 65876 30092
rect 69292 30052 69332 30092
rect 70732 30052 70772 30092
rect 71692 30052 71732 30092
rect 72172 30052 72212 30092
rect 75724 30052 75764 30092
rect 77068 30052 77108 30092
rect 38860 29968 38900 30008
rect 40012 29968 40052 30008
rect 46060 29968 46100 30008
rect 54700 29968 54740 30008
rect 55564 29968 55604 30008
rect 58636 29968 58676 30008
rect 58828 29968 58868 30008
rect 60364 29968 60404 30008
rect 73900 29968 73940 30008
rect 77644 29968 77684 30008
rect 39820 29884 39860 29924
rect 40396 29884 40436 29924
rect 50380 29884 50420 29924
rect 54508 29884 54548 29924
rect 59020 29884 59060 29924
rect 59404 29884 59444 29924
rect 69100 29884 69140 29924
rect 71884 29884 71924 29924
rect 75052 29884 75092 29924
rect 40588 29800 40628 29840
rect 40684 29800 40724 29840
rect 40780 29800 40820 29840
rect 41356 29800 41396 29840
rect 41548 29800 41588 29840
rect 43852 29800 43892 29840
rect 44716 29800 44756 29840
rect 46348 29800 46388 29840
rect 46444 29800 46484 29840
rect 46732 29800 46772 29840
rect 47020 29800 47060 29840
rect 47212 29787 47252 29827
rect 48172 29800 48212 29840
rect 49036 29800 49076 29840
rect 50764 29800 50804 29840
rect 41452 29716 41492 29756
rect 43468 29716 43508 29756
rect 47788 29716 47828 29756
rect 50860 29758 50900 29798
rect 51052 29800 51092 29840
rect 51628 29800 51668 29840
rect 52492 29800 52532 29840
rect 54892 29800 54932 29840
rect 55084 29800 55124 29840
rect 55180 29800 55220 29840
rect 55468 29800 55508 29840
rect 55660 29800 55700 29840
rect 55852 29800 55892 29840
rect 56044 29800 56084 29840
rect 56140 29800 56180 29840
rect 59692 29800 59732 29840
rect 59980 29800 60020 29840
rect 60076 29800 60116 29840
rect 60940 29800 60980 29840
rect 61804 29800 61844 29840
rect 63244 29800 63284 29840
rect 63340 29779 63380 29819
rect 63436 29800 63476 29840
rect 63628 29800 63668 29840
rect 63820 29800 63860 29840
rect 63916 29800 63956 29840
rect 65164 29800 65204 29840
rect 65452 29800 65492 29840
rect 65548 29800 65588 29840
rect 66412 29800 66452 29840
rect 67276 29800 67316 29840
rect 69484 29800 69524 29840
rect 69676 29800 69716 29840
rect 69772 29800 69812 29840
rect 69964 29800 70004 29840
rect 70060 29800 70100 29840
rect 70252 29800 70292 29840
rect 71020 29800 71060 29840
rect 71116 29800 71156 29840
rect 71404 29800 71444 29840
rect 72076 29800 72116 29840
rect 72268 29800 72308 29840
rect 75340 29800 75380 29840
rect 75436 29800 75476 29840
rect 75532 29800 75572 29840
rect 75724 29800 75764 29840
rect 75916 29800 75956 29840
rect 76012 29800 76052 29840
rect 76492 29800 76532 29840
rect 76684 29800 76724 29840
rect 77068 29800 77108 29840
rect 77260 29800 77300 29840
rect 77356 29800 77396 29840
rect 51244 29716 51284 29756
rect 60556 29716 60596 29756
rect 63148 29716 63188 29756
rect 66028 29716 66068 29756
rect 69580 29716 69620 29756
rect 76588 29716 76628 29756
rect 40876 29632 40916 29672
rect 50188 29632 50228 29672
rect 50572 29632 50612 29672
rect 50956 29632 50996 29672
rect 53644 29632 53684 29672
rect 55948 29632 55988 29672
rect 59212 29632 59252 29672
rect 62956 29632 62996 29672
rect 68428 29632 68468 29672
rect 70156 29632 70196 29672
rect 74860 29632 74900 29672
rect 75244 29632 75284 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 45004 29296 45044 29336
rect 55372 29296 55412 29336
rect 59308 29296 59348 29336
rect 60460 29296 60500 29336
rect 61132 29296 61172 29336
rect 63436 29296 63476 29336
rect 70348 29296 70388 29336
rect 70828 29296 70868 29336
rect 71692 29296 71732 29336
rect 75820 29296 75860 29336
rect 46060 29212 46100 29252
rect 46348 29212 46388 29252
rect 50476 29212 50516 29252
rect 56332 29212 56372 29252
rect 60844 29212 60884 29252
rect 65740 29212 65780 29252
rect 67756 29212 67796 29252
rect 76492 29212 76532 29252
rect 38380 29128 38420 29168
rect 38764 29128 38804 29168
rect 39628 29128 39668 29168
rect 41068 29128 41108 29168
rect 41356 29128 41396 29168
rect 41452 29128 41492 29168
rect 41932 29128 41972 29168
rect 42028 29128 42068 29168
rect 42220 29128 42260 29168
rect 44908 29128 44948 29168
rect 45100 29128 45140 29168
rect 45196 29128 45236 29168
rect 45964 29128 46004 29168
rect 46156 29128 46196 29168
rect 46732 29128 46772 29168
rect 47596 29128 47636 29168
rect 49516 29128 49556 29168
rect 49708 29128 49748 29168
rect 49804 29128 49844 29168
rect 50092 29128 50132 29168
rect 50380 29128 50420 29168
rect 51820 29128 51860 29168
rect 52972 29128 53012 29168
rect 53356 29128 53396 29168
rect 54220 29128 54260 29168
rect 55564 29128 55604 29168
rect 55660 29128 55700 29168
rect 55756 29128 55796 29168
rect 55852 29128 55892 29168
rect 56716 29128 56756 29168
rect 57580 29128 57620 29168
rect 59500 29128 59540 29168
rect 59692 29128 59732 29168
rect 59788 29128 59828 29168
rect 60268 29128 60308 29168
rect 60364 29128 60404 29168
rect 60556 29128 60596 29168
rect 60748 29128 60788 29168
rect 60940 29128 60980 29168
rect 63340 29117 63380 29157
rect 63532 29128 63572 29168
rect 63628 29128 63668 29168
rect 63820 29128 63860 29168
rect 63916 29128 63956 29168
rect 64012 29128 64052 29168
rect 64108 29128 64148 29168
rect 64972 29128 65012 29168
rect 65164 29128 65204 29168
rect 65644 29128 65684 29168
rect 65836 29128 65876 29168
rect 65932 29128 65972 29168
rect 68140 29128 68180 29168
rect 69004 29128 69044 29168
rect 70444 29128 70484 29168
rect 70540 29128 70580 29168
rect 70636 29128 70676 29168
rect 71308 29128 71348 29168
rect 71500 29128 71540 29168
rect 73804 29128 73844 29168
rect 74668 29128 74708 29168
rect 76108 29128 76148 29168
rect 76396 29128 76436 29168
rect 51148 29044 51188 29084
rect 51532 29044 51572 29084
rect 59116 29044 59156 29084
rect 61324 29044 61364 29084
rect 73420 29086 73460 29126
rect 77068 29128 77108 29168
rect 77452 29128 77492 29168
rect 78316 29128 78356 29168
rect 70156 29044 70196 29084
rect 71020 29044 71060 29084
rect 71884 29044 71924 29084
rect 41740 28960 41780 29000
rect 42412 28960 42452 29000
rect 49516 28960 49556 29000
rect 50764 28960 50804 29000
rect 62380 28960 62420 29000
rect 76780 28960 76820 29000
rect 40780 28876 40820 28916
rect 42220 28876 42260 28916
rect 48748 28876 48788 28916
rect 50956 28876 50996 28916
rect 51340 28876 51380 28916
rect 58732 28876 58772 28916
rect 59500 28876 59540 28916
rect 65068 28876 65108 28916
rect 70828 28876 70868 28916
rect 71404 28876 71444 28916
rect 71692 28876 71732 28916
rect 79468 28876 79508 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 39628 28540 39668 28580
rect 41452 28540 41492 28580
rect 45292 28540 45332 28580
rect 51244 28540 51284 28580
rect 55276 28540 55316 28580
rect 59020 28540 59060 28580
rect 65260 28540 65300 28580
rect 73804 28540 73844 28580
rect 76684 28540 76724 28580
rect 38188 28456 38228 28496
rect 44332 28456 44372 28496
rect 47500 28456 47540 28496
rect 49228 28456 49268 28496
rect 52492 28456 52532 28496
rect 56812 28456 56852 28496
rect 58636 28456 58676 28496
rect 59788 28456 59828 28496
rect 68332 28456 68372 28496
rect 71020 28456 71060 28496
rect 77548 28456 77588 28496
rect 39436 28372 39476 28412
rect 40012 28372 40052 28412
rect 51052 28372 51092 28412
rect 54412 28372 54452 28412
rect 58444 28372 58484 28412
rect 58828 28372 58868 28412
rect 60940 28372 60980 28412
rect 70060 28372 70100 28412
rect 40204 28288 40244 28328
rect 40396 28288 40436 28328
rect 40492 28288 40532 28328
rect 40876 28288 40916 28328
rect 41068 28288 41108 28328
rect 41164 28288 41204 28328
rect 41356 28288 41396 28328
rect 41548 28288 41588 28328
rect 41740 28288 41780 28328
rect 42124 28288 42164 28328
rect 42988 28288 43028 28328
rect 45004 28288 45044 28328
rect 45100 28288 45140 28328
rect 45292 28288 45332 28328
rect 45484 28288 45524 28328
rect 45676 28288 45716 28328
rect 45772 28288 45812 28328
rect 49420 28288 49460 28328
rect 49612 28288 49652 28328
rect 49708 28288 49748 28328
rect 49900 28288 49940 28328
rect 49996 28288 50036 28328
rect 50188 28288 50228 28328
rect 50476 28288 50516 28328
rect 50572 28288 50612 28328
rect 50668 28288 50708 28328
rect 51724 28288 51764 28328
rect 51820 28288 51860 28328
rect 51916 28288 51956 28328
rect 52108 28288 52148 28328
rect 52300 28288 52340 28328
rect 53068 28288 53108 28328
rect 55564 28288 55604 28328
rect 55660 28288 55700 28328
rect 55948 28288 55988 28328
rect 56236 28288 56276 28328
rect 56428 28288 56468 28328
rect 59212 28288 59252 28328
rect 59404 28288 59444 28328
rect 59500 28288 59540 28328
rect 59692 28288 59732 28328
rect 59884 28288 59924 28328
rect 60076 28288 60116 28328
rect 60268 28288 60308 28328
rect 60364 28288 60404 28328
rect 60556 28288 60596 28328
rect 60652 28288 60692 28328
rect 60748 28288 60788 28328
rect 62284 28288 62324 28328
rect 63148 28288 63188 28328
rect 64588 28288 64628 28328
rect 64876 28288 64916 28328
rect 66124 28288 66164 28328
rect 66988 28288 67028 28328
rect 70348 28288 70388 28328
rect 70636 28288 70676 28328
rect 70732 28288 70772 28328
rect 71788 28288 71828 28328
rect 72652 28288 72692 28328
rect 75244 28288 75284 28328
rect 75436 28288 75476 28328
rect 75532 28288 75572 28328
rect 76684 28288 76724 28328
rect 76876 28288 76916 28328
rect 76972 28288 77012 28328
rect 77164 28288 77204 28328
rect 77356 28288 77396 28328
rect 40972 28204 41012 28244
rect 52204 28204 52244 28244
rect 56332 28204 56372 28244
rect 61900 28204 61940 28244
rect 64972 28204 65012 28244
rect 65740 28204 65780 28244
rect 71404 28204 71444 28244
rect 75340 28204 75380 28244
rect 77260 28204 77300 28244
rect 39820 28120 39860 28160
rect 40300 28120 40340 28160
rect 44140 28120 44180 28160
rect 45580 28120 45620 28160
rect 49516 28120 49556 28160
rect 50092 28120 50132 28160
rect 50380 28120 50420 28160
rect 51244 28120 51284 28160
rect 59020 28120 59060 28160
rect 59308 28120 59348 28160
rect 60172 28120 60212 28160
rect 61132 28120 61172 28160
rect 64300 28120 64340 28160
rect 68140 28120 68180 28160
rect 69868 28120 69908 28160
rect 73804 28120 73844 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 45964 27784 46004 27824
rect 51244 27784 51284 27824
rect 54508 27784 54548 27824
rect 54796 27784 54836 27824
rect 59692 27784 59732 27824
rect 64012 27784 64052 27824
rect 68620 27784 68660 27824
rect 75532 27784 75572 27824
rect 37708 27700 37748 27740
rect 40396 27700 40436 27740
rect 43564 27700 43604 27740
rect 46444 27700 46484 27740
rect 48844 27700 48884 27740
rect 51724 27700 51764 27740
rect 52108 27700 52148 27740
rect 57100 27700 57140 27740
rect 60460 27700 60500 27740
rect 65260 27700 65300 27740
rect 70732 27700 70772 27740
rect 71116 27700 71156 27740
rect 38092 27616 38132 27656
rect 38956 27616 38996 27656
rect 40300 27616 40340 27656
rect 40492 27616 40532 27656
rect 40588 27616 40628 27656
rect 40972 27616 41012 27656
rect 41164 27616 41204 27656
rect 43948 27616 43988 27656
rect 44812 27616 44852 27656
rect 46540 27616 46580 27656
rect 46828 27616 46868 27656
rect 47116 27616 47156 27656
rect 47308 27616 47348 27656
rect 47404 27616 47444 27656
rect 47596 27616 47636 27656
rect 47692 27616 47732 27656
rect 47788 27616 47828 27656
rect 49228 27616 49268 27656
rect 50092 27616 50132 27656
rect 51628 27616 51668 27656
rect 51820 27616 51860 27656
rect 51916 27616 51956 27656
rect 52492 27616 52532 27656
rect 53356 27616 53396 27656
rect 54700 27616 54740 27656
rect 54892 27616 54932 27656
rect 54988 27616 55028 27656
rect 55180 27616 55220 27656
rect 55372 27616 55412 27656
rect 55468 27616 55508 27656
rect 55660 27616 55700 27656
rect 55756 27616 55796 27656
rect 55852 27616 55892 27656
rect 55948 27616 55988 27656
rect 57484 27616 57524 27656
rect 58348 27616 58388 27656
rect 59788 27616 59828 27656
rect 59884 27616 59924 27656
rect 59980 27616 60020 27656
rect 60844 27616 60884 27656
rect 61708 27616 61748 27656
rect 63820 27616 63860 27656
rect 63916 27616 63956 27656
rect 64108 27616 64148 27656
rect 65164 27616 65204 27656
rect 65356 27616 65396 27656
rect 65452 27616 65492 27656
rect 65644 27616 65684 27656
rect 65836 27616 65876 27656
rect 69580 27616 69620 27656
rect 69772 27616 69812 27656
rect 69868 27616 69908 27656
rect 70060 27616 70100 27656
rect 70252 27616 70292 27656
rect 70348 27616 70388 27656
rect 70636 27616 70676 27656
rect 70828 27616 70868 27656
rect 71020 27616 71060 27656
rect 71212 27616 71252 27656
rect 71308 27616 71348 27656
rect 74860 27616 74900 27656
rect 75052 27616 75092 27656
rect 75148 27616 75188 27656
rect 75436 27616 75476 27656
rect 75628 27616 75668 27656
rect 75724 27616 75764 27656
rect 76780 27616 76820 27656
rect 76876 27616 76916 27656
rect 76972 27616 77012 27656
rect 77164 27616 77204 27656
rect 77356 27616 77396 27656
rect 41548 27532 41588 27572
rect 65740 27532 65780 27572
rect 67564 27532 67604 27572
rect 68428 27532 68468 27572
rect 36460 27448 36500 27488
rect 41356 27448 41396 27488
rect 55180 27448 55220 27488
rect 66220 27448 66260 27488
rect 69388 27448 69428 27488
rect 70060 27448 70100 27488
rect 71884 27448 71924 27488
rect 73516 27448 73556 27488
rect 77548 27448 77588 27488
rect 40108 27364 40148 27404
rect 41068 27364 41108 27404
rect 46156 27364 46196 27404
rect 47116 27364 47156 27404
rect 51244 27364 51284 27404
rect 59500 27364 59540 27404
rect 62860 27364 62900 27404
rect 67372 27364 67412 27404
rect 69580 27364 69620 27404
rect 74860 27364 74900 27404
rect 77260 27364 77300 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 41068 27028 41108 27068
rect 44908 27028 44948 27068
rect 45868 27028 45908 27068
rect 46348 27028 46388 27068
rect 49420 27028 49460 27068
rect 51916 27028 51956 27068
rect 54220 27028 54260 27068
rect 58444 27028 58484 27068
rect 59404 27028 59444 27068
rect 60748 27028 60788 27068
rect 63820 27028 63860 27068
rect 71884 27028 71924 27068
rect 72076 27028 72116 27068
rect 76876 27028 76916 27068
rect 33004 26944 33044 26984
rect 35308 26944 35348 26984
rect 38860 26944 38900 26984
rect 53452 26944 53492 26984
rect 57580 26944 57620 26984
rect 61132 26944 61172 26984
rect 62092 26944 62132 26984
rect 35596 26860 35636 26900
rect 38668 26860 38708 26900
rect 39052 26860 39092 26900
rect 39436 26860 39476 26900
rect 44716 26860 44756 26900
rect 52108 26860 52148 26900
rect 58252 26860 58292 26900
rect 59020 26860 59060 26900
rect 60364 26860 60404 26900
rect 60940 26860 60980 26900
rect 71692 26860 71732 26900
rect 72268 26860 72308 26900
rect 75436 26860 75476 26900
rect 4300 26776 4340 26816
rect 35212 26776 35252 26816
rect 35404 26776 35444 26816
rect 36364 26776 36404 26816
rect 37228 26776 37268 26816
rect 39820 26776 39860 26816
rect 39916 26776 39956 26816
rect 40012 26776 40052 26816
rect 40108 26776 40148 26816
rect 40396 26776 40436 26816
rect 40684 26776 40724 26816
rect 40780 26776 40820 26816
rect 41260 26776 41300 26816
rect 41356 26776 41396 26816
rect 41452 26776 41492 26816
rect 42028 26776 42068 26816
rect 42892 26776 42932 26816
rect 45100 26776 45140 26816
rect 45196 26776 45236 26816
rect 45292 26776 45332 26816
rect 45388 26776 45428 26816
rect 45580 26776 45620 26816
rect 45676 26776 45716 26816
rect 45868 26776 45908 26816
rect 46243 26763 46283 26803
rect 46444 26776 46484 26816
rect 46636 26776 46676 26816
rect 46828 26776 46868 26816
rect 47020 26776 47060 26816
rect 47404 26776 47444 26816
rect 48268 26776 48308 26816
rect 50092 26776 50132 26816
rect 50284 26776 50324 26816
rect 50380 26776 50420 26816
rect 50572 26776 50612 26816
rect 50668 26776 50708 26816
rect 50860 26776 50900 26816
rect 51244 26776 51284 26816
rect 51532 26776 51572 26816
rect 51628 26776 51668 26816
rect 55372 26776 55412 26816
rect 56236 26776 56276 26816
rect 59788 26776 59828 26816
rect 60076 26776 60116 26816
rect 63820 26776 63860 26816
rect 64012 26776 64052 26816
rect 64108 26776 64148 26816
rect 66892 26776 66932 26816
rect 67756 26776 67796 26816
rect 68332 26776 68372 26816
rect 68524 26776 68564 26816
rect 68620 26776 68660 26816
rect 69100 26776 69140 26816
rect 69484 26776 69524 26816
rect 70348 26776 70388 26816
rect 73036 26776 73076 26816
rect 73420 26812 73460 26852
rect 74284 26776 74324 26816
rect 75628 26776 75668 26816
rect 75724 26776 75764 26816
rect 75820 26755 75860 26795
rect 75916 26776 75956 26816
rect 76204 26776 76244 26816
rect 76492 26776 76532 26816
rect 76588 26776 76628 26816
rect 77452 26776 77492 26816
rect 78316 26776 78356 26816
rect 35980 26692 36020 26732
rect 41644 26692 41684 26732
rect 46732 26692 46772 26732
rect 50188 26692 50228 26732
rect 56620 26692 56660 26732
rect 59692 26692 59732 26732
rect 68140 26692 68180 26732
rect 77068 26692 77108 26732
rect 4204 26608 4244 26648
rect 35788 26608 35828 26648
rect 38380 26608 38420 26648
rect 39244 26608 39284 26648
rect 39628 26608 39668 26648
rect 44044 26608 44084 26648
rect 44908 26608 44948 26648
rect 49420 26608 49460 26648
rect 50764 26608 50804 26648
rect 52300 26608 52340 26648
rect 58828 26608 58868 26648
rect 60556 26608 60596 26648
rect 60748 26608 60788 26648
rect 65740 26608 65780 26648
rect 68428 26608 68468 26648
rect 71500 26608 71540 26648
rect 71884 26608 71924 26648
rect 79468 26608 79508 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 35884 26272 35924 26312
rect 39148 26272 39188 26312
rect 56428 26272 56468 26312
rect 57676 26272 57716 26312
rect 61228 26272 61268 26312
rect 67756 26272 67796 26312
rect 69580 26272 69620 26312
rect 75244 26272 75284 26312
rect 76972 26272 77012 26312
rect 36364 26188 36404 26228
rect 33388 26104 33428 26144
rect 34252 26104 34292 26144
rect 34636 26104 34676 26144
rect 34924 26104 34964 26144
rect 35212 26104 35252 26144
rect 35308 26104 35348 26144
rect 35788 26104 35828 26144
rect 35980 26104 36020 26144
rect 36076 26104 36116 26144
rect 36268 26104 36308 26144
rect 36460 26104 36500 26144
rect 39340 26104 39380 26144
rect 39820 26146 39860 26186
rect 48748 26188 48788 26228
rect 52108 26188 52148 26228
rect 55852 26188 55892 26228
rect 61612 26188 61652 26228
rect 64780 26188 64820 26228
rect 71308 26188 71348 26228
rect 71884 26188 71924 26228
rect 39532 26104 39572 26144
rect 39628 26104 39668 26144
rect 40012 26090 40052 26130
rect 40108 26104 40148 26144
rect 41164 26104 41204 26144
rect 41260 26104 41300 26144
rect 41452 26104 41492 26144
rect 43660 26104 43700 26144
rect 44044 26104 44084 26144
rect 44908 26104 44948 26144
rect 47212 26104 47252 26144
rect 47980 26104 48020 26144
rect 48172 26104 48212 26144
rect 49132 26104 49172 26144
rect 49996 26104 50036 26144
rect 52012 26104 52052 26144
rect 52204 26104 52244 26144
rect 52396 26104 52436 26144
rect 52588 26104 52628 26144
rect 55468 26104 55508 26144
rect 55756 26104 55796 26144
rect 56332 26104 56372 26144
rect 56524 26104 56564 26144
rect 56620 26104 56660 26144
rect 56812 26104 56852 26144
rect 57004 26104 57044 26144
rect 57100 26104 57140 26144
rect 58348 26104 58388 26144
rect 58540 26104 58580 26144
rect 58636 26104 58676 26144
rect 58828 26104 58868 26144
rect 59020 26104 59060 26144
rect 59116 26104 59156 26144
rect 59404 26104 59444 26144
rect 59500 26104 59540 26144
rect 59596 26104 59636 26144
rect 59788 26104 59828 26144
rect 59884 26104 59924 26144
rect 60076 26104 60116 26144
rect 61996 26104 62036 26144
rect 62860 26104 62900 26144
rect 64204 26104 64244 26144
rect 64300 26104 64340 26144
rect 64396 26104 64436 26144
rect 64492 26104 64532 26144
rect 64684 26093 64724 26133
rect 64876 26104 64916 26144
rect 64972 26104 65012 26144
rect 65452 26104 65492 26144
rect 65644 26104 65684 26144
rect 65740 26104 65780 26144
rect 67180 26104 67220 26144
rect 67276 26104 67316 26144
rect 67372 26104 67412 26144
rect 67468 26104 67508 26144
rect 67660 26104 67700 26144
rect 67852 26104 67892 26144
rect 67948 26104 67988 26144
rect 68140 26104 68180 26144
rect 68332 26104 68372 26144
rect 69292 26104 69332 26144
rect 69388 26104 69428 26144
rect 69484 26104 69524 26144
rect 70924 26104 70964 26144
rect 71212 26104 71252 26144
rect 71788 26104 71828 26144
rect 71980 26104 72020 26144
rect 74188 26104 74228 26144
rect 74284 26104 74324 26144
rect 74476 26104 74516 26144
rect 74668 26104 74708 26144
rect 74764 26104 74804 26144
rect 74860 26104 74900 26144
rect 74956 26104 74996 26144
rect 75148 26104 75188 26144
rect 75340 26104 75380 26144
rect 75436 26104 75476 26144
rect 76876 26104 76916 26144
rect 77068 26104 77108 26144
rect 77164 26104 77204 26144
rect 652 26020 692 26060
rect 38956 26020 38996 26060
rect 40492 26020 40532 26060
rect 48076 26020 48116 26060
rect 51532 26020 51572 26060
rect 57484 26020 57524 26060
rect 60268 26020 60308 26060
rect 60652 26020 60692 26060
rect 61036 26020 61076 26060
rect 68812 26020 68852 26060
rect 70444 26020 70484 26060
rect 844 25936 884 25976
rect 32236 25936 32276 25976
rect 35596 25936 35636 25976
rect 39820 25936 39860 25976
rect 40684 25936 40724 25976
rect 41452 25936 41492 25976
rect 42124 25936 42164 25976
rect 47020 25936 47060 25976
rect 47596 25936 47636 25976
rect 48556 25936 48596 25976
rect 51724 25936 51764 25976
rect 52780 25936 52820 25976
rect 54892 25936 54932 25976
rect 56812 25936 56852 25976
rect 57868 25936 57908 25976
rect 58348 25936 58388 25976
rect 58828 25936 58868 25976
rect 60460 25936 60500 25976
rect 60844 25936 60884 25976
rect 65452 25936 65492 25976
rect 66412 25936 66452 25976
rect 68620 25936 68660 25976
rect 71596 25936 71636 25976
rect 39148 25852 39188 25892
rect 39340 25852 39380 25892
rect 46060 25852 46100 25892
rect 51148 25852 51188 25892
rect 52492 25852 52532 25892
rect 56140 25852 56180 25892
rect 60076 25852 60116 25892
rect 64012 25852 64052 25892
rect 68236 25852 68276 25892
rect 70636 25852 70676 25892
rect 73420 25894 73460 25934
rect 74476 25936 74516 25976
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 34924 25516 34964 25556
rect 40396 25516 40436 25556
rect 45100 25516 45140 25556
rect 46828 25516 46868 25556
rect 52108 25516 52148 25556
rect 56236 25516 56276 25556
rect 67756 25516 67796 25556
rect 75628 25516 75668 25556
rect 75916 25516 75956 25556
rect 35692 25432 35732 25472
rect 44140 25432 44180 25472
rect 55756 25432 55796 25472
rect 63820 25432 63860 25472
rect 76492 25432 76532 25472
rect 652 25348 692 25388
rect 40588 25347 40628 25387
rect 54700 25348 54740 25388
rect 30124 25264 30164 25304
rect 30988 25264 31028 25304
rect 32812 25264 32852 25304
rect 29740 25180 29780 25220
rect 33100 25222 33140 25262
rect 33292 25264 33332 25304
rect 33388 25264 33428 25304
rect 34444 25264 34484 25304
rect 34540 25264 34580 25304
rect 34636 25264 34676 25304
rect 34732 25264 34772 25304
rect 34924 25264 34964 25304
rect 35116 25264 35156 25304
rect 35212 25264 35252 25304
rect 35692 25264 35732 25304
rect 35884 25264 35924 25304
rect 35980 25264 36020 25304
rect 37228 25264 37268 25304
rect 37612 25264 37652 25304
rect 38476 25264 38516 25304
rect 39820 25264 39860 25304
rect 39916 25264 39956 25304
rect 40012 25264 40052 25304
rect 40108 25264 40148 25304
rect 41260 25264 41300 25304
rect 42124 25264 42164 25304
rect 44812 25264 44852 25304
rect 44908 25264 44948 25304
rect 45100 25264 45140 25304
rect 45292 25264 45332 25304
rect 45388 25264 45428 25304
rect 45484 25264 45524 25304
rect 45580 25264 45620 25304
rect 45772 25264 45812 25304
rect 46156 25264 46196 25304
rect 46444 25264 46484 25304
rect 46540 25264 46580 25304
rect 47404 25264 47444 25304
rect 48268 25264 48308 25304
rect 50572 25264 50612 25304
rect 50668 25264 50708 25304
rect 50764 25264 50804 25304
rect 50860 25264 50900 25304
rect 51436 25264 51476 25304
rect 51724 25264 51764 25304
rect 52684 25264 52724 25304
rect 53548 25264 53588 25304
rect 55276 25264 55316 25304
rect 55468 25264 55508 25304
rect 55564 25264 55604 25304
rect 56140 25264 56180 25304
rect 56332 25264 56372 25304
rect 57388 25264 57428 25304
rect 57772 25264 57812 25304
rect 58636 25264 58676 25304
rect 60268 25264 60308 25304
rect 60652 25264 60692 25304
rect 61516 25264 61556 25304
rect 63148 25264 63188 25304
rect 63436 25264 63476 25304
rect 63532 25264 63572 25304
rect 64396 25264 64436 25304
rect 65260 25264 65300 25304
rect 67084 25264 67124 25304
rect 67372 25264 67412 25304
rect 67468 25264 67508 25304
rect 68332 25264 68372 25304
rect 69196 25264 69236 25304
rect 71020 25264 71060 25304
rect 71884 25264 71924 25304
rect 73228 25264 73268 25304
rect 73612 25264 73652 25304
rect 74476 25264 74516 25304
rect 75820 25264 75860 25304
rect 76005 25279 76045 25319
rect 76204 25264 76244 25304
rect 76300 25264 76340 25304
rect 76492 25264 76532 25304
rect 76684 25264 76724 25304
rect 77068 25264 77108 25304
rect 77932 25264 77972 25304
rect 40876 25180 40916 25220
rect 47020 25180 47060 25220
rect 51820 25180 51860 25220
rect 52300 25180 52340 25220
rect 64012 25180 64052 25220
rect 67948 25180 67988 25220
rect 70636 25180 70676 25220
rect 844 25096 884 25136
rect 32140 25096 32180 25136
rect 33196 25096 33236 25136
rect 39628 25096 39668 25136
rect 43276 25096 43316 25136
rect 49420 25096 49460 25136
rect 55372 25096 55412 25136
rect 59788 25096 59828 25136
rect 62668 25096 62708 25136
rect 66412 25096 66452 25136
rect 70348 25096 70388 25136
rect 73036 25096 73076 25136
rect 75628 25096 75668 25136
rect 79084 25096 79124 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 32236 24760 32276 24800
rect 39148 24760 39188 24800
rect 40588 24760 40628 24800
rect 45004 24760 45044 24800
rect 46828 24760 46868 24800
rect 50188 24760 50228 24800
rect 51436 24760 51476 24800
rect 52204 24760 52244 24800
rect 58348 24760 58388 24800
rect 59020 24760 59060 24800
rect 64012 24760 64052 24800
rect 67756 24760 67796 24800
rect 74380 24760 74420 24800
rect 34924 24676 34964 24716
rect 40012 24676 40052 24716
rect 54892 24676 54932 24716
rect 59500 24676 59540 24716
rect 60268 24676 60308 24716
rect 64492 24676 64532 24716
rect 64876 24676 64916 24716
rect 68236 24676 68276 24716
rect 75820 24676 75860 24716
rect 76492 24676 76532 24716
rect 31660 24592 31700 24632
rect 31756 24592 31796 24632
rect 31852 24592 31892 24632
rect 31948 24592 31988 24632
rect 32140 24592 32180 24632
rect 32332 24592 32372 24632
rect 32428 24592 32468 24632
rect 32716 24592 32756 24632
rect 32908 24592 32948 24632
rect 34156 24592 34196 24632
rect 35308 24592 35348 24632
rect 36172 24592 36212 24632
rect 39628 24592 39668 24632
rect 39916 24592 39956 24632
rect 40492 24592 40532 24632
rect 40684 24592 40724 24632
rect 40780 24592 40820 24632
rect 40972 24592 41012 24632
rect 41164 24592 41204 24632
rect 42316 24592 42356 24632
rect 42700 24592 42740 24632
rect 43564 24592 43604 24632
rect 44908 24592 44948 24632
rect 45100 24592 45140 24632
rect 45196 24592 45236 24632
rect 46732 24592 46772 24632
rect 46924 24592 46964 24632
rect 47020 24592 47060 24632
rect 50380 24592 50420 24632
rect 50572 24592 50612 24632
rect 50668 24592 50708 24632
rect 50860 24592 50900 24632
rect 51052 24592 51092 24632
rect 52108 24592 52148 24632
rect 52300 24592 52340 24632
rect 52396 24592 52436 24632
rect 55276 24592 55316 24632
rect 56140 24592 56180 24632
rect 58060 24592 58100 24632
rect 58156 24592 58196 24632
rect 58252 24592 58292 24632
rect 59596 24592 59636 24632
rect 59884 24592 59924 24632
rect 60172 24592 60212 24632
rect 60364 24592 60404 24632
rect 63916 24592 63956 24632
rect 64108 24592 64148 24632
rect 64204 24592 64244 24632
rect 64396 24592 64436 24632
rect 64588 24592 64628 24632
rect 64780 24592 64820 24632
rect 64972 24592 65012 24632
rect 67660 24592 67700 24632
rect 67852 24592 67892 24632
rect 67948 24592 67988 24632
rect 68140 24592 68180 24632
rect 68332 24592 68372 24632
rect 70732 24592 70772 24632
rect 70924 24592 70964 24632
rect 71020 24592 71060 24632
rect 71212 24592 71252 24632
rect 71308 24592 71348 24632
rect 71404 24592 71444 24632
rect 74284 24592 74324 24632
rect 74476 24592 74516 24632
rect 74572 24592 74612 24632
rect 75436 24592 75476 24632
rect 75724 24592 75764 24632
rect 76396 24592 76436 24632
rect 76588 24592 76628 24632
rect 652 24508 692 24548
rect 39340 24508 39380 24548
rect 41068 24508 41108 24548
rect 49996 24508 50036 24548
rect 51244 24508 51284 24548
rect 57292 24508 57332 24548
rect 58828 24508 58868 24548
rect 60748 24508 60788 24548
rect 30220 24424 30260 24464
rect 33868 24424 33908 24464
rect 37708 24424 37748 24464
rect 41356 24424 41396 24464
rect 48556 24424 48596 24464
rect 52588 24424 52628 24464
rect 59212 24424 59252 24464
rect 60940 24424 60980 24464
rect 65164 24424 65204 24464
rect 68524 24424 68564 24464
rect 70732 24424 70772 24464
rect 71596 24424 71636 24464
rect 76108 24424 76148 24464
rect 77164 24424 77204 24464
rect 844 24340 884 24380
rect 32812 24340 32852 24380
rect 37324 24340 37364 24380
rect 40300 24340 40340 24380
rect 44716 24340 44756 24380
rect 50188 24340 50228 24380
rect 50380 24340 50420 24380
rect 50956 24340 50996 24380
rect 60556 24340 60596 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 36556 24004 36596 24044
rect 40204 24004 40244 24044
rect 41452 24004 41492 24044
rect 44428 24004 44468 24044
rect 55756 24004 55796 24044
rect 28876 23920 28916 23960
rect 32524 23920 32564 23960
rect 35500 23920 35540 23960
rect 40684 23920 40724 23960
rect 42796 23920 42836 23960
rect 45676 23920 45716 23960
rect 46924 23920 46964 23960
rect 51436 23920 51476 23960
rect 652 23836 692 23876
rect 1804 23836 1844 23876
rect 1996 23836 2036 23876
rect 30892 23836 30932 23876
rect 40492 23836 40532 23876
rect 41260 23836 41300 23876
rect 31276 23752 31316 23792
rect 31468 23752 31508 23792
rect 31564 23752 31604 23792
rect 31852 23752 31892 23792
rect 32140 23752 32180 23792
rect 32236 23752 32276 23792
rect 33292 23752 33332 23792
rect 34156 23752 34196 23792
rect 36076 23752 36116 23792
rect 36172 23752 36212 23792
rect 36268 23752 36308 23792
rect 36364 23752 36404 23792
rect 36556 23752 36596 23792
rect 36748 23752 36788 23792
rect 36844 23752 36884 23792
rect 38764 23752 38804 23792
rect 38860 23752 38900 23792
rect 38956 23752 38996 23792
rect 39244 23752 39284 23792
rect 39436 23752 39476 23792
rect 39532 23752 39572 23792
rect 40108 23752 40148 23792
rect 40300 23752 40340 23792
rect 40876 23752 40916 23792
rect 41068 23752 41108 23792
rect 44044 23752 44084 23792
rect 44140 23752 44180 23792
rect 44236 23752 44276 23792
rect 44428 23752 44468 23792
rect 44620 23752 44660 23792
rect 44716 23752 44756 23792
rect 45004 23752 45044 23792
rect 45292 23752 45332 23792
rect 45388 23752 45428 23792
rect 45868 23752 45908 23792
rect 45964 23752 46004 23792
rect 46060 23752 46100 23792
rect 48460 23752 48500 23792
rect 49324 23752 49364 23792
rect 50668 23752 50708 23792
rect 50860 23752 50900 23792
rect 50956 23752 50996 23792
rect 51148 23752 51188 23792
rect 51244 23766 51284 23806
rect 51436 23752 51476 23792
rect 51724 23752 51764 23792
rect 52108 23752 52148 23792
rect 52972 23752 53012 23792
rect 54796 23752 54836 23792
rect 55180 23752 55220 23792
rect 55660 23752 55700 23792
rect 55852 23752 55892 23792
rect 56140 23752 56180 23792
rect 56428 23752 56468 23792
rect 56620 23752 56660 23792
rect 56908 23752 56948 23792
rect 57292 23752 57332 23792
rect 57676 23752 57716 23792
rect 58060 23752 58100 23792
rect 58444 23752 58484 23792
rect 58828 23752 58868 23792
rect 59308 23752 59348 23792
rect 59692 23752 59732 23792
rect 60076 23752 60116 23792
rect 60460 23752 60500 23792
rect 60844 23752 60884 23792
rect 61324 23752 61364 23792
rect 61708 23752 61748 23792
rect 62092 23752 62132 23792
rect 62476 23752 62516 23792
rect 62860 23752 62900 23792
rect 63244 23752 63284 23792
rect 63628 23752 63668 23792
rect 64108 23752 64148 23792
rect 64492 23752 64532 23792
rect 64876 23752 64916 23792
rect 65260 23752 65300 23792
rect 65740 23752 65780 23792
rect 66124 23752 66164 23792
rect 66508 23752 66548 23792
rect 66892 23752 66932 23792
rect 67276 23752 67316 23792
rect 67660 23752 67700 23792
rect 68140 23752 68180 23792
rect 68524 23752 68564 23792
rect 68908 23752 68948 23792
rect 69292 23752 69332 23792
rect 69676 23752 69716 23792
rect 70156 23752 70196 23792
rect 70540 23752 70580 23792
rect 70924 23752 70964 23792
rect 71308 23752 71348 23792
rect 71692 23752 71732 23792
rect 72076 23752 72116 23792
rect 72460 23752 72500 23792
rect 72844 23752 72884 23792
rect 73324 23752 73364 23792
rect 73708 23752 73748 23792
rect 74092 23752 74132 23792
rect 74476 23752 74516 23792
rect 74860 23752 74900 23792
rect 75244 23752 75284 23792
rect 75628 23752 75668 23792
rect 76108 23752 76148 23792
rect 76972 23752 77012 23792
rect 77260 23752 77300 23792
rect 77548 23752 77588 23792
rect 77740 23752 77780 23792
rect 78124 23752 78164 23792
rect 78508 23752 78548 23792
rect 78796 23752 78836 23792
rect 79084 23752 79124 23792
rect 79372 23752 79412 23792
rect 32908 23668 32948 23708
rect 39052 23668 39092 23708
rect 40972 23668 41012 23708
rect 48076 23668 48116 23708
rect 50764 23668 50804 23708
rect 844 23584 884 23624
rect 1612 23584 1652 23624
rect 2188 23584 2228 23624
rect 31084 23584 31124 23624
rect 31372 23584 31412 23624
rect 35308 23584 35348 23624
rect 39340 23584 39380 23624
rect 41452 23584 41492 23624
rect 43948 23584 43988 23624
rect 50476 23584 50516 23624
rect 54124 23584 54164 23624
rect 54892 23584 54932 23624
rect 55276 23584 55316 23624
rect 56044 23584 56084 23624
rect 56332 23584 56372 23624
rect 56716 23584 56756 23624
rect 57004 23584 57044 23624
rect 57388 23584 57428 23624
rect 57772 23584 57812 23624
rect 58156 23584 58196 23624
rect 58540 23584 58580 23624
rect 58924 23584 58964 23624
rect 59404 23584 59444 23624
rect 59788 23584 59828 23624
rect 60172 23584 60212 23624
rect 60556 23584 60596 23624
rect 60940 23584 60980 23624
rect 61420 23584 61460 23624
rect 61804 23584 61844 23624
rect 62188 23584 62228 23624
rect 62572 23584 62612 23624
rect 62956 23584 62996 23624
rect 63340 23584 63380 23624
rect 63724 23584 63764 23624
rect 64204 23584 64244 23624
rect 64588 23584 64628 23624
rect 64972 23584 65012 23624
rect 65356 23584 65396 23624
rect 65836 23584 65876 23624
rect 66220 23584 66260 23624
rect 66604 23584 66644 23624
rect 66988 23584 67028 23624
rect 67372 23584 67412 23624
rect 67756 23584 67796 23624
rect 68236 23584 68276 23624
rect 68620 23584 68660 23624
rect 69004 23584 69044 23624
rect 69388 23584 69428 23624
rect 69772 23584 69812 23624
rect 70252 23584 70292 23624
rect 70636 23584 70676 23624
rect 71020 23584 71060 23624
rect 71404 23584 71444 23624
rect 71788 23584 71828 23624
rect 72172 23584 72212 23624
rect 72556 23584 72596 23624
rect 72940 23584 72980 23624
rect 73420 23584 73460 23624
rect 73804 23584 73844 23624
rect 74188 23584 74228 23624
rect 74572 23584 74612 23624
rect 74956 23584 74996 23624
rect 75340 23584 75380 23624
rect 75724 23584 75764 23624
rect 76204 23584 76244 23624
rect 76876 23584 76916 23624
rect 77164 23584 77204 23624
rect 77452 23584 77492 23624
rect 77836 23584 77876 23624
rect 78220 23584 78260 23624
rect 78604 23584 78644 23624
rect 78892 23584 78932 23624
rect 79180 23584 79220 23624
rect 79468 23584 79508 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 41068 23290 41108 23330
rect 32620 23248 32660 23288
rect 37900 23248 37940 23288
rect 40876 23248 40916 23288
rect 44716 23248 44756 23288
rect 48748 23248 48788 23288
rect 51052 23290 51092 23330
rect 49612 23248 49652 23288
rect 50092 23248 50132 23288
rect 32236 23164 32276 23204
rect 36652 23164 36692 23204
rect 41356 23164 41396 23204
rect 45580 23164 45620 23204
rect 50764 23164 50804 23204
rect 51340 23164 51380 23204
rect 1516 23080 1556 23120
rect 1900 23080 1940 23120
rect 2092 23080 2132 23120
rect 28396 23080 28436 23120
rect 28780 23080 28820 23120
rect 29644 23080 29684 23120
rect 30988 23080 31028 23120
rect 31180 23080 31220 23120
rect 31276 23080 31316 23120
rect 31756 23080 31796 23120
rect 31948 23080 31988 23120
rect 32140 23080 32180 23120
rect 32332 23080 32372 23120
rect 32524 23080 32564 23120
rect 32716 23080 32756 23120
rect 32812 23080 32852 23120
rect 36268 23080 36308 23120
rect 36556 23080 36596 23120
rect 37132 23080 37172 23120
rect 37228 23080 37268 23120
rect 37324 23080 37364 23120
rect 37804 23080 37844 23120
rect 37996 23080 38036 23120
rect 38092 23080 38132 23120
rect 38476 23080 38516 23120
rect 38860 23080 38900 23120
rect 39724 23080 39764 23120
rect 41452 23080 41492 23120
rect 41740 23080 41780 23120
rect 44620 23080 44660 23120
rect 44812 23080 44852 23120
rect 44908 23080 44948 23120
rect 45484 23080 45524 23120
rect 45676 23080 45716 23120
rect 45868 23080 45908 23120
rect 45964 23080 46004 23120
rect 46156 23080 46196 23120
rect 46348 23080 46388 23120
rect 46732 23080 46772 23120
rect 47596 23080 47636 23120
rect 652 22996 692 23036
rect 49420 22996 49460 23036
rect 49804 23035 49844 23075
rect 49900 23080 49940 23120
rect 49996 23080 50036 23120
rect 50380 23080 50420 23120
rect 50668 23080 50708 23120
rect 51244 23101 51284 23141
rect 51436 23080 51476 23120
rect 52492 23080 52532 23120
rect 51724 22996 51764 23036
rect 1516 22912 1556 22952
rect 30988 22912 31028 22952
rect 33388 22912 33428 22952
rect 35980 22912 36020 22952
rect 36940 22912 36980 22952
rect 42028 22912 42068 22952
rect 42892 22912 42932 22952
rect 46156 22912 46196 22952
rect 52300 22912 52340 22952
rect 844 22828 884 22868
rect 1708 22828 1748 22868
rect 1900 22828 1940 22868
rect 30796 22828 30836 22868
rect 31852 22828 31892 22868
rect 49612 22828 49652 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 28300 22492 28340 22532
rect 31852 22492 31892 22532
rect 35212 22492 35252 22532
rect 39052 22492 39092 22532
rect 43564 22492 43604 22532
rect 50380 22492 50420 22532
rect 52012 22492 52052 22532
rect 52396 22492 52436 22532
rect 52684 22492 52724 22532
rect 652 22408 692 22448
rect 27916 22408 27956 22448
rect 38860 22408 38900 22448
rect 40972 22408 41012 22448
rect 44908 22408 44948 22448
rect 46444 22408 46484 22448
rect 48172 22408 48212 22448
rect 27724 22324 27764 22364
rect 28108 22324 28148 22364
rect 50188 22324 50228 22364
rect 28492 22240 28532 22280
rect 28684 22240 28724 22280
rect 28876 22240 28916 22280
rect 29068 22240 29108 22280
rect 29548 22240 29588 22280
rect 29740 22240 29780 22280
rect 29836 22240 29876 22280
rect 30604 22240 30644 22280
rect 30700 22240 30740 22280
rect 30796 22240 30836 22280
rect 30892 22240 30932 22280
rect 31180 22240 31220 22280
rect 31468 22240 31508 22280
rect 31564 22240 31604 22280
rect 28588 22156 28628 22196
rect 28972 22156 29012 22196
rect 32140 22198 32180 22238
rect 32332 22240 32372 22280
rect 32428 22240 32468 22280
rect 33196 22240 33236 22280
rect 34060 22240 34100 22280
rect 36076 22240 36116 22280
rect 36940 22240 36980 22280
rect 39052 22240 39092 22280
rect 39244 22240 39284 22280
rect 39340 22240 39380 22280
rect 40684 22240 40724 22280
rect 40780 22240 40820 22280
rect 40972 22240 41012 22280
rect 41164 22240 41204 22280
rect 41548 22240 41588 22280
rect 42412 22240 42452 22280
rect 44812 22240 44852 22280
rect 45004 22240 45044 22280
rect 45196 22240 45236 22280
rect 45388 22240 45428 22280
rect 45484 22240 45524 22280
rect 45676 22240 45716 22280
rect 45868 22240 45908 22280
rect 48556 22240 48596 22280
rect 48652 22240 48692 22280
rect 48748 22240 48788 22280
rect 49420 22240 49460 22280
rect 49612 22240 49652 22280
rect 49708 22240 49748 22280
rect 50572 22240 50612 22280
rect 50764 22240 50804 22280
rect 51628 22240 51668 22280
rect 52108 22229 52148 22269
rect 52300 22240 52340 22280
rect 52588 22240 52628 22280
rect 32236 22156 32276 22196
rect 32812 22156 32852 22196
rect 35692 22156 35732 22196
rect 45772 22156 45812 22196
rect 50668 22156 50708 22196
rect 28300 22072 28340 22112
rect 29644 22072 29684 22112
rect 35212 22072 35252 22112
rect 38092 22072 38132 22112
rect 43564 22072 43604 22112
rect 45292 22072 45332 22112
rect 48844 22072 48884 22112
rect 49516 22072 49556 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 36172 21736 36212 21776
rect 44812 21736 44852 21776
rect 32428 21652 32468 21692
rect 41260 21652 41300 21692
rect 42412 21652 42452 21692
rect 51052 21652 51092 21692
rect 26668 21568 26708 21608
rect 27532 21568 27572 21608
rect 27916 21568 27956 21608
rect 28204 21568 28244 21608
rect 28492 21568 28532 21608
rect 28588 21568 28628 21608
rect 29356 21568 29396 21608
rect 29740 21568 29780 21608
rect 30604 21568 30644 21608
rect 32332 21568 32372 21608
rect 32524 21568 32564 21608
rect 36076 21568 36116 21608
rect 36268 21568 36308 21608
rect 36364 21568 36404 21608
rect 36556 21568 36596 21608
rect 36748 21568 36788 21608
rect 38956 21568 38996 21608
rect 39052 21568 39092 21608
rect 39148 21568 39188 21608
rect 39244 21568 39284 21608
rect 41164 21568 41204 21608
rect 41356 21568 41396 21608
rect 42796 21568 42836 21608
rect 43660 21568 43700 21608
rect 45292 21568 45332 21608
rect 45388 21568 45428 21608
rect 45676 21568 45716 21608
rect 45964 21568 46004 21608
rect 46348 21568 46388 21608
rect 47212 21568 47252 21608
rect 48844 21568 48884 21608
rect 49036 21568 49076 21608
rect 49132 21568 49172 21608
rect 49516 21568 49556 21608
rect 49612 21568 49652 21608
rect 49708 21568 49748 21608
rect 50188 21568 50228 21608
rect 50284 21568 50324 21608
rect 50572 21568 50612 21608
rect 50860 21568 50900 21608
rect 50956 21568 50996 21608
rect 51148 21568 51188 21608
rect 52300 21568 52340 21608
rect 52396 21568 52436 21608
rect 52588 21568 52628 21608
rect 52684 21568 52724 21608
rect 3052 21484 3092 21524
rect 3628 21484 3668 21524
rect 4012 21484 4052 21524
rect 4204 21484 4244 21524
rect 3244 21400 3284 21440
rect 28876 21400 28916 21440
rect 31756 21400 31796 21440
rect 32716 21400 32756 21440
rect 33292 21400 33332 21440
rect 35692 21400 35732 21440
rect 36652 21400 36692 21440
rect 39436 21400 39476 21440
rect 45004 21400 45044 21440
rect 49900 21400 49940 21440
rect 51340 21400 51380 21440
rect 3436 21316 3476 21356
rect 3820 21316 3860 21356
rect 4396 21316 4436 21356
rect 25516 21316 25556 21356
rect 48364 21316 48404 21356
rect 48844 21316 48884 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 26956 20980 26996 21020
rect 28300 20980 28340 21020
rect 29068 20980 29108 21020
rect 43852 20980 43892 21020
rect 46348 20980 46388 21020
rect 50092 20980 50132 21020
rect 52684 20980 52724 21020
rect 652 20896 692 20936
rect 26188 20896 26228 20936
rect 29836 20896 29876 20936
rect 38476 20896 38516 20936
rect 41932 20896 41972 20936
rect 5068 20812 5108 20852
rect 23212 20812 23252 20852
rect 26380 20812 26420 20852
rect 26764 20812 26804 20852
rect 27148 20812 27188 20852
rect 42892 20812 42932 20852
rect 43468 20812 43508 20852
rect 43660 20812 43700 20852
rect 44044 20812 44084 20852
rect 44620 20812 44660 20852
rect 3532 20728 3572 20768
rect 3628 20728 3668 20768
rect 3820 20728 3860 20768
rect 27820 20728 27860 20768
rect 27916 20728 27956 20768
rect 28012 20728 28052 20768
rect 28108 20728 28148 20768
rect 28300 20728 28340 20768
rect 28492 20728 28532 20768
rect 28588 20728 28628 20768
rect 28780 20728 28820 20768
rect 28876 20728 28916 20768
rect 29068 20728 29108 20768
rect 32620 20728 32660 20768
rect 33484 20728 33524 20768
rect 35692 20728 35732 20768
rect 36556 20728 36596 20768
rect 38188 20728 38228 20768
rect 38284 20728 38324 20768
rect 38476 20728 38516 20768
rect 38668 20728 38708 20768
rect 39052 20728 39092 20768
rect 39916 20728 39956 20768
rect 42412 20728 42452 20768
rect 42508 20728 42548 20768
rect 42604 20728 42644 20768
rect 44812 20728 44852 20768
rect 44908 20728 44948 20768
rect 45004 20728 45044 20768
rect 45100 20728 45140 20768
rect 45484 20728 45524 20768
rect 45676 20728 45716 20768
rect 45772 20728 45812 20768
rect 46348 20728 46388 20768
rect 46540 20728 46580 20768
rect 46636 20728 46676 20768
rect 47692 20728 47732 20768
rect 48076 20728 48116 20768
rect 48940 20728 48980 20768
rect 50284 20728 50324 20768
rect 50668 20728 50708 20768
rect 51532 20728 51572 20768
rect 32236 20644 32276 20684
rect 35308 20644 35348 20684
rect 3724 20560 3764 20600
rect 5260 20560 5300 20600
rect 23020 20560 23060 20600
rect 26572 20560 26612 20600
rect 26956 20560 26996 20600
rect 27340 20560 27380 20600
rect 34636 20560 34676 20600
rect 37708 20560 37748 20600
rect 41068 20560 41108 20600
rect 42316 20560 42356 20600
rect 43084 20560 43124 20600
rect 43276 20560 43316 20600
rect 44236 20560 44276 20600
rect 44428 20560 44468 20600
rect 45580 20560 45620 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 23500 20224 23540 20264
rect 32332 20224 32372 20264
rect 35692 20224 35732 20264
rect 37996 20224 38036 20264
rect 4684 20056 4724 20096
rect 10924 20056 10964 20096
rect 11020 20077 11060 20117
rect 11116 20056 11156 20096
rect 11212 20056 11252 20096
rect 11404 20056 11444 20096
rect 11596 20056 11636 20096
rect 11692 20056 11732 20096
rect 22540 20056 22580 20096
rect 22732 20056 22772 20096
rect 22828 20056 22868 20096
rect 26476 20056 26516 20096
rect 26668 20056 26708 20096
rect 26764 20056 26804 20096
rect 29932 20056 29972 20096
rect 30028 20056 30068 20096
rect 30124 20056 30164 20096
rect 30220 20056 30260 20096
rect 32140 20056 32180 20096
rect 32236 20056 32276 20096
rect 32428 20056 32468 20096
rect 32620 20056 32660 20096
rect 32716 20056 32756 20096
rect 32812 20056 32852 20096
rect 32908 20056 32948 20096
rect 34828 20056 34868 20096
rect 34924 20056 34964 20096
rect 35116 20056 35156 20096
rect 35500 20056 35540 20096
rect 35596 20056 35636 20096
rect 35788 20056 35828 20096
rect 35980 20056 36020 20096
rect 36076 20056 36116 20096
rect 36172 20056 36212 20096
rect 36268 20056 36308 20096
rect 37804 20056 37844 20096
rect 37900 20056 37940 20096
rect 38092 20056 38132 20096
rect 38284 20056 38324 20096
rect 38476 20056 38516 20096
rect 38668 20056 38708 20096
rect 38860 20056 38900 20096
rect 39148 20056 39188 20096
rect 41452 20056 41492 20096
rect 41836 20056 41876 20096
rect 42700 20056 42740 20096
rect 49132 20056 49172 20096
rect 49324 20056 49364 20096
rect 5068 19972 5108 20012
rect 23692 19972 23732 20012
rect 31756 19972 31796 20012
rect 43852 19972 43892 20012
rect 44524 19972 44564 20012
rect 45292 19972 45332 20012
rect 45676 19972 45716 20012
rect 47500 19972 47540 20012
rect 47884 19972 47924 20012
rect 652 19888 692 19928
rect 9580 19888 9620 19928
rect 12748 19888 12788 19928
rect 23116 19888 23156 19928
rect 26476 19888 26516 19928
rect 26956 19888 26996 19928
rect 29740 19888 29780 19928
rect 33388 19888 33428 19928
rect 35116 19888 35156 19928
rect 40780 19888 40820 19928
rect 44716 19888 44756 19928
rect 46732 19888 46772 19928
rect 50092 19888 50132 19928
rect 4588 19804 4628 19844
rect 4876 19804 4916 19844
rect 11404 19804 11444 19844
rect 22540 19804 22580 19844
rect 31948 19804 31988 19844
rect 38380 19804 38420 19844
rect 38764 19804 38804 19844
rect 44332 19804 44372 19844
rect 45100 19804 45140 19844
rect 45484 19804 45524 19844
rect 47308 19804 47348 19844
rect 47692 19804 47732 19844
rect 49228 19804 49268 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 14668 19468 14708 19508
rect 32140 19468 32180 19508
rect 35788 19468 35828 19508
rect 39052 19468 39092 19508
rect 40588 19468 40628 19508
rect 48940 19468 48980 19508
rect 652 19384 692 19424
rect 29068 19384 29108 19424
rect 33580 19384 33620 19424
rect 36076 19384 36116 19424
rect 37036 19384 37076 19424
rect 38380 19384 38420 19424
rect 40396 19384 40436 19424
rect 41260 19384 41300 19424
rect 43468 19384 43508 19424
rect 21772 19300 21812 19340
rect 31660 19300 31700 19340
rect 10060 19216 10100 19256
rect 10924 19216 10964 19256
rect 11308 19216 11348 19256
rect 11788 19216 11828 19256
rect 11980 19216 12020 19256
rect 12076 19216 12116 19256
rect 12652 19216 12692 19256
rect 13516 19216 13556 19256
rect 22156 19216 22196 19256
rect 22252 19216 22292 19256
rect 22348 19216 22388 19256
rect 22444 19216 22484 19256
rect 22636 19216 22676 19256
rect 23020 19252 23060 19292
rect 40204 19300 40244 19340
rect 40780 19311 40820 19351
rect 41548 19300 41588 19340
rect 23884 19216 23924 19256
rect 25228 19216 25268 19256
rect 25324 19216 25364 19256
rect 25516 19216 25556 19256
rect 25804 19216 25844 19256
rect 25900 19216 25940 19256
rect 25996 19216 26036 19256
rect 26572 19216 26612 19256
rect 27436 19216 27476 19256
rect 28780 19216 28820 19256
rect 28876 19216 28916 19256
rect 29068 19216 29108 19256
rect 29260 19216 29300 19256
rect 29644 19216 29684 19256
rect 30508 19216 30548 19256
rect 31852 19216 31892 19256
rect 31948 19216 31988 19256
rect 32140 19216 32180 19256
rect 32908 19216 32948 19256
rect 33196 19216 33236 19256
rect 33292 19216 33332 19256
rect 33772 19216 33812 19256
rect 33964 19216 34004 19256
rect 35692 19216 35732 19256
rect 35884 19216 35924 19256
rect 36364 19216 36404 19256
rect 36460 19216 36500 19256
rect 36748 19216 36788 19256
rect 38572 19216 38612 19256
rect 38764 19216 38804 19256
rect 38860 19216 38900 19256
rect 39340 19216 39380 19256
rect 39436 19216 39476 19256
rect 39724 19216 39764 19256
rect 40972 19216 41012 19256
rect 41068 19216 41108 19256
rect 41260 19216 41300 19256
rect 41932 19216 41972 19256
rect 42028 19216 42068 19256
rect 42220 19216 42260 19256
rect 42796 19216 42836 19256
rect 43180 19258 43220 19298
rect 43084 19216 43124 19256
rect 44044 19216 44084 19256
rect 44908 19216 44948 19256
rect 46636 19216 46676 19256
rect 47500 19216 47540 19256
rect 48940 19216 48980 19256
rect 49132 19216 49172 19256
rect 49228 19216 49268 19256
rect 49612 19216 49652 19256
rect 49996 19216 50036 19256
rect 50860 19216 50900 19256
rect 11884 19132 11924 19172
rect 12268 19132 12308 19172
rect 26188 19132 26228 19172
rect 33868 19132 33908 19172
rect 42124 19132 42164 19172
rect 43660 19132 43700 19172
rect 46252 19132 46292 19172
rect 8908 19048 8948 19088
rect 14668 19048 14708 19088
rect 21964 19048 22004 19088
rect 25036 19048 25076 19088
rect 25420 19048 25460 19088
rect 25708 19048 25748 19088
rect 28588 19048 28628 19088
rect 38668 19048 38708 19088
rect 41740 19048 41780 19088
rect 46060 19048 46100 19088
rect 48652 19048 48692 19088
rect 52012 19048 52052 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 22540 18712 22580 18752
rect 26284 18712 26324 18752
rect 41164 18712 41204 18752
rect 44044 18712 44084 18752
rect 11020 18628 11060 18668
rect 11596 18628 11636 18668
rect 12172 18628 12212 18668
rect 23020 18628 23060 18668
rect 27244 18628 27284 18668
rect 28876 18628 28916 18668
rect 29740 18628 29780 18668
rect 30316 18628 30356 18668
rect 32524 18628 32564 18668
rect 32908 18628 32948 18668
rect 35788 18628 35828 18668
rect 36172 18628 36212 18668
rect 38764 18628 38804 18668
rect 43660 18628 43700 18668
rect 49324 18628 49364 18668
rect 10636 18544 10676 18584
rect 10924 18544 10964 18584
rect 11500 18544 11540 18584
rect 11692 18544 11732 18584
rect 12076 18544 12116 18584
rect 12268 18544 12308 18584
rect 23116 18544 23156 18584
rect 23404 18544 23444 18584
rect 26188 18544 26228 18584
rect 26380 18544 26420 18584
rect 26476 18544 26516 18584
rect 26860 18544 26900 18584
rect 27148 18544 27188 18584
rect 27724 18544 27764 18584
rect 27820 18544 27860 18584
rect 27916 18544 27956 18584
rect 28684 18544 28724 18584
rect 28780 18544 28820 18584
rect 28972 18544 29012 18584
rect 29644 18544 29684 18584
rect 29836 18544 29876 18584
rect 30412 18544 30452 18584
rect 30700 18544 30740 18584
rect 31180 18544 31220 18584
rect 32428 18544 32468 18584
rect 32620 18544 32660 18584
rect 32716 18544 32756 18584
rect 33292 18544 33332 18584
rect 34156 18544 34196 18584
rect 35692 18544 35732 18584
rect 35884 18544 35924 18584
rect 35980 18544 36020 18584
rect 36556 18544 36596 18584
rect 37420 18544 37460 18584
rect 39148 18544 39188 18584
rect 40012 18544 40052 18584
rect 41932 18544 41972 18584
rect 42124 18544 42164 18584
rect 42220 18544 42260 18584
rect 42412 18544 42452 18584
rect 42604 18544 42644 18584
rect 42700 18544 42740 18584
rect 43564 18544 43604 18584
rect 43756 18544 43796 18584
rect 43948 18544 43988 18584
rect 44140 18544 44180 18584
rect 44236 18544 44276 18584
rect 44428 18544 44468 18584
rect 44620 18544 44660 18584
rect 46732 18544 46772 18584
rect 46828 18544 46868 18584
rect 47020 18544 47060 18584
rect 47404 18544 47444 18584
rect 47500 18544 47540 18584
rect 47596 18544 47636 18584
rect 47692 18544 47732 18584
rect 48364 18544 48404 18584
rect 48652 18544 48692 18584
rect 48748 18544 48788 18584
rect 49228 18565 49268 18605
rect 49420 18544 49460 18584
rect 52300 18544 52340 18584
rect 52684 18544 52724 18584
rect 1708 18460 1748 18500
rect 21964 18460 22004 18500
rect 22348 18460 22388 18500
rect 23692 18460 23732 18500
rect 24076 18460 24116 18500
rect 24460 18460 24500 18500
rect 24844 18460 24884 18500
rect 25708 18460 25748 18500
rect 35308 18460 35348 18500
rect 41740 18460 41780 18500
rect 43084 18460 43124 18500
rect 49804 18460 49844 18500
rect 50476 18460 50516 18500
rect 51340 18460 51380 18500
rect 51532 18460 51572 18500
rect 652 18376 692 18416
rect 11308 18376 11348 18416
rect 22156 18376 22196 18416
rect 25516 18376 25556 18416
rect 27532 18376 27572 18416
rect 30028 18376 30068 18416
rect 41548 18376 41588 18416
rect 44524 18376 44564 18416
rect 47020 18376 47060 18416
rect 49036 18376 49076 18416
rect 50764 18376 50804 18416
rect 1516 18292 1556 18332
rect 22732 18292 22772 18332
rect 23884 18292 23924 18332
rect 24268 18292 24308 18332
rect 24652 18292 24692 18332
rect 25036 18292 25076 18332
rect 31564 18292 31604 18332
rect 38572 18292 38612 18332
rect 41164 18292 41204 18332
rect 41932 18292 41972 18332
rect 42412 18292 42452 18332
rect 42892 18292 42932 18332
rect 49996 18292 50036 18332
rect 50284 18292 50324 18332
rect 51148 18292 51188 18332
rect 51724 18292 51764 18332
rect 52396 18292 52436 18332
rect 52588 18292 52628 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 33388 17956 33428 17996
rect 36556 17956 36596 17996
rect 37036 17956 37076 17996
rect 46444 17956 46484 17996
rect 50092 17956 50132 17996
rect 652 17872 692 17912
rect 23212 17872 23252 17912
rect 34828 17872 34868 17912
rect 37900 17872 37940 17912
rect 39436 17872 39476 17912
rect 22636 17788 22676 17828
rect 34348 17788 34388 17828
rect 36844 17788 36884 17828
rect 46828 17788 46868 17828
rect 49516 17788 49556 17828
rect 22540 17704 22580 17744
rect 22732 17704 22772 17744
rect 22924 17704 22964 17744
rect 23020 17718 23060 17758
rect 23212 17704 23252 17744
rect 23404 17704 23444 17744
rect 23788 17704 23828 17744
rect 24652 17704 24692 17744
rect 26668 17704 26708 17744
rect 26860 17704 26900 17744
rect 26956 17704 26996 17744
rect 27532 17704 27572 17744
rect 28396 17704 28436 17744
rect 29836 17704 29876 17744
rect 30028 17704 30068 17744
rect 30124 17704 30164 17744
rect 30700 17704 30740 17744
rect 31564 17704 31604 17744
rect 33292 17704 33332 17744
rect 33484 17704 33524 17744
rect 36460 17704 36500 17744
rect 36652 17704 36692 17744
rect 39820 17704 39860 17744
rect 40204 17704 40244 17744
rect 41068 17704 41108 17744
rect 42604 17704 42644 17744
rect 42796 17704 42836 17744
rect 42892 17704 42932 17744
rect 43468 17704 43508 17744
rect 44332 17704 44372 17744
rect 45772 17704 45812 17744
rect 45964 17704 46004 17744
rect 46156 17704 46196 17744
rect 46252 17704 46292 17744
rect 46444 17704 46484 17744
rect 48652 17704 48692 17744
rect 48748 17704 48788 17744
rect 48940 17704 48980 17744
rect 49420 17704 49460 17744
rect 49612 17704 49652 17744
rect 49804 17704 49844 17744
rect 49900 17704 49940 17744
rect 50092 17704 50132 17744
rect 50284 17704 50324 17744
rect 50668 17704 50708 17744
rect 51532 17704 51572 17744
rect 27148 17620 27188 17660
rect 29932 17620 29972 17660
rect 30316 17620 30356 17660
rect 42700 17620 42740 17660
rect 43084 17620 43124 17660
rect 45868 17620 45908 17660
rect 25804 17536 25844 17576
rect 26764 17536 26804 17576
rect 29548 17536 29588 17576
rect 32716 17536 32756 17576
rect 34156 17536 34196 17576
rect 37036 17536 37076 17576
rect 42220 17536 42260 17576
rect 45484 17536 45524 17576
rect 46636 17536 46676 17576
rect 48844 17536 48884 17576
rect 52684 17536 52724 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 23212 17200 23252 17240
rect 41644 17200 41684 17240
rect 51436 17200 51476 17240
rect 52684 17200 52724 17240
rect 23692 17116 23732 17156
rect 27340 17116 27380 17156
rect 30508 17116 30548 17156
rect 42604 17116 42644 17156
rect 44044 17116 44084 17156
rect 45772 17116 45812 17156
rect 51724 17116 51764 17156
rect 4204 17032 4244 17072
rect 4396 17032 4436 17072
rect 23596 17032 23636 17072
rect 23788 17032 23828 17072
rect 27244 17032 27284 17072
rect 27436 17032 27476 17072
rect 30412 17032 30452 17072
rect 30604 17032 30644 17072
rect 33388 17032 33428 17072
rect 33580 17032 33620 17072
rect 33772 17032 33812 17072
rect 33868 17032 33908 17072
rect 34060 17032 34100 17072
rect 34252 17032 34292 17072
rect 34636 17032 34676 17072
rect 35500 17032 35540 17072
rect 36940 17032 36980 17072
rect 37132 17032 37172 17072
rect 37324 17032 37364 17072
rect 37708 17032 37748 17072
rect 38572 17032 38612 17072
rect 41740 17032 41780 17072
rect 41836 17032 41876 17072
rect 41932 17032 41972 17072
rect 42220 17032 42260 17072
rect 42508 17032 42548 17072
rect 43948 17032 43988 17072
rect 44140 17032 44180 17072
rect 45388 17032 45428 17072
rect 45676 17032 45716 17072
rect 46252 17032 46292 17072
rect 46636 17032 46676 17072
rect 47500 17032 47540 17072
rect 49132 17032 49172 17072
rect 49228 17032 49268 17072
rect 49420 17032 49460 17072
rect 49708 17032 49748 17072
rect 49804 17032 49844 17072
rect 49900 17032 49940 17072
rect 49996 17032 50036 17072
rect 50380 17032 50420 17072
rect 50668 17032 50708 17072
rect 50764 17032 50804 17072
rect 51628 17032 51668 17072
rect 51820 17032 51860 17072
rect 52300 17032 52340 17072
rect 52588 17032 52628 17072
rect 2764 16948 2804 16988
rect 3148 16948 3188 16988
rect 4780 16948 4820 16988
rect 23404 16948 23444 16988
rect 40876 16948 40916 16988
rect 41452 16948 41492 16988
rect 43276 16948 43316 16988
rect 44524 16948 44564 16988
rect 44908 16948 44948 16988
rect 48652 16948 48692 16988
rect 51244 16948 51284 16988
rect 652 16864 692 16904
rect 2956 16864 2996 16904
rect 3340 16864 3380 16904
rect 4588 16864 4628 16904
rect 23980 16864 24020 16904
rect 27628 16864 27668 16904
rect 30796 16864 30836 16904
rect 31564 16864 31604 16904
rect 33484 16864 33524 16904
rect 34060 16864 34100 16904
rect 39724 16864 39764 16904
rect 41068 16864 41108 16904
rect 42892 16864 42932 16904
rect 43084 16864 43124 16904
rect 43564 16864 43604 16904
rect 44716 16864 44756 16904
rect 51052 16864 51092 16904
rect 4300 16780 4340 16820
rect 36652 16780 36692 16820
rect 37036 16780 37076 16820
rect 41260 16780 41300 16820
rect 45100 16780 45140 16820
rect 46060 16780 46100 16820
rect 49420 16780 49460 16820
rect 51436 16780 51476 16820
rect 52396 16780 52436 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 1996 16444 2036 16484
rect 2572 16444 2612 16484
rect 4012 16444 4052 16484
rect 6988 16444 7028 16484
rect 34732 16444 34772 16484
rect 37996 16444 38036 16484
rect 45772 16444 45812 16484
rect 46252 16444 46292 16484
rect 51052 16444 51092 16484
rect 54796 16444 54836 16484
rect 55084 16444 55124 16484
rect 55372 16444 55412 16484
rect 55756 16444 55796 16484
rect 56620 16444 56660 16484
rect 57388 16444 57428 16484
rect 58060 16444 58100 16484
rect 58348 16444 58388 16484
rect 58636 16444 58676 16484
rect 59020 16444 59060 16484
rect 60172 16444 60212 16484
rect 60556 16444 60596 16484
rect 60844 16444 60884 16484
rect 61516 16444 61556 16484
rect 62188 16444 62228 16484
rect 62476 16444 62516 16484
rect 62764 16444 62804 16484
rect 63052 16444 63092 16484
rect 63436 16444 63476 16484
rect 64588 16444 64628 16484
rect 65068 16444 65108 16484
rect 65452 16444 65492 16484
rect 65836 16444 65876 16484
rect 66604 16444 66644 16484
rect 67084 16444 67124 16484
rect 67468 16444 67508 16484
rect 67852 16444 67892 16484
rect 68236 16444 68276 16484
rect 69004 16444 69044 16484
rect 69484 16444 69524 16484
rect 69868 16444 69908 16484
rect 70252 16444 70292 16484
rect 70636 16444 70676 16484
rect 71020 16444 71060 16484
rect 71404 16444 71444 16484
rect 71884 16444 71924 16484
rect 72268 16444 72308 16484
rect 72652 16444 72692 16484
rect 73036 16444 73076 16484
rect 73420 16444 73460 16484
rect 74284 16444 74324 16484
rect 74668 16444 74708 16484
rect 75052 16444 75092 16484
rect 75436 16444 75476 16484
rect 76492 16444 76532 16484
rect 76876 16444 76916 16484
rect 77260 16444 77300 16484
rect 77644 16444 77684 16484
rect 78028 16444 78068 16484
rect 78316 16444 78356 16484
rect 78700 16444 78740 16484
rect 78988 16444 79028 16484
rect 79276 16444 79316 16484
rect 652 16360 692 16400
rect 1804 16360 1844 16400
rect 4204 16360 4244 16400
rect 34444 16360 34484 16400
rect 37516 16360 37556 16400
rect 43084 16360 43124 16400
rect 46732 16360 46772 16400
rect 52108 16360 52148 16400
rect 53644 16360 53684 16400
rect 53932 16360 53972 16400
rect 54316 16360 54356 16400
rect 57580 16360 57620 16400
rect 61036 16360 61076 16400
rect 2188 16276 2228 16316
rect 2380 16276 2420 16316
rect 3436 16276 3476 16316
rect 3820 16276 3860 16316
rect 4396 16276 4436 16316
rect 61708 16276 61748 16316
rect 2764 16192 2804 16232
rect 2956 16192 2996 16232
rect 3052 16192 3092 16232
rect 4972 16192 5012 16232
rect 5836 16192 5876 16232
rect 31468 16192 31508 16232
rect 32332 16192 32372 16232
rect 33772 16192 33812 16232
rect 34060 16192 34100 16232
rect 34636 16192 34676 16232
rect 34828 16192 34868 16232
rect 36844 16209 36884 16249
rect 37132 16192 37172 16232
rect 37708 16192 37748 16232
rect 37804 16192 37844 16232
rect 37996 16192 38036 16232
rect 39820 16192 39860 16232
rect 40012 16192 40052 16232
rect 40588 16192 40628 16232
rect 41452 16192 41492 16232
rect 42988 16192 43028 16232
rect 43173 16207 43213 16247
rect 43756 16192 43796 16232
rect 44620 16192 44660 16232
rect 45964 16192 46004 16232
rect 46060 16192 46100 16232
rect 46252 16192 46292 16232
rect 47116 16192 47156 16232
rect 47212 16192 47252 16232
rect 47308 16192 47348 16232
rect 48652 16192 48692 16232
rect 49036 16192 49076 16232
rect 49900 16192 49940 16232
rect 51628 16192 51668 16232
rect 51724 16192 51764 16232
rect 51820 16192 51860 16232
rect 52396 16192 52436 16232
rect 52492 16192 52532 16232
rect 52780 16192 52820 16232
rect 53068 16178 53108 16218
rect 53356 16192 53396 16232
rect 53548 16192 53588 16232
rect 53740 16192 53780 16232
rect 4588 16108 4628 16148
rect 31084 16108 31124 16148
rect 34156 16108 34196 16148
rect 37228 16108 37268 16148
rect 39916 16108 39956 16148
rect 40204 16108 40244 16148
rect 43372 16108 43412 16148
rect 53260 16150 53300 16190
rect 54700 16192 54740 16232
rect 54988 16192 55028 16232
rect 55276 16192 55316 16232
rect 55660 16192 55700 16232
rect 56044 16192 56084 16232
rect 56524 16192 56564 16232
rect 56908 16192 56948 16232
rect 57292 16192 57332 16232
rect 57964 16192 58004 16232
rect 58252 16192 58292 16232
rect 58540 16192 58580 16232
rect 58924 16192 58964 16232
rect 59308 16192 59348 16232
rect 59692 16192 59732 16232
rect 60076 16192 60116 16232
rect 60460 16192 60500 16232
rect 60748 16192 60788 16232
rect 61420 16192 61460 16232
rect 62092 16192 62132 16232
rect 62380 16192 62420 16232
rect 62668 16192 62708 16232
rect 62956 16192 62996 16232
rect 63327 16181 63367 16221
rect 63724 16192 63764 16232
rect 64108 16192 64148 16232
rect 64492 16192 64532 16232
rect 64972 16192 65012 16232
rect 65356 16192 65396 16232
rect 65740 16192 65780 16232
rect 66124 16192 66164 16232
rect 66508 16192 66548 16232
rect 66988 16192 67028 16232
rect 67372 16192 67412 16232
rect 67756 16192 67796 16232
rect 68140 16192 68180 16232
rect 68524 16192 68564 16232
rect 68908 16192 68948 16232
rect 69388 16192 69428 16232
rect 69772 16192 69812 16232
rect 70156 16192 70196 16232
rect 70540 16192 70580 16232
rect 70924 16192 70964 16232
rect 71308 16192 71348 16232
rect 71788 16192 71828 16232
rect 72172 16192 72212 16232
rect 72556 16192 72596 16232
rect 72940 16192 72980 16232
rect 73324 16192 73364 16232
rect 73708 16192 73748 16232
rect 74188 16192 74228 16232
rect 74572 16192 74612 16232
rect 74956 16192 74996 16232
rect 75340 16192 75380 16232
rect 75724 16192 75764 16232
rect 76588 16192 76628 16232
rect 76972 16192 77012 16232
rect 77164 16192 77204 16232
rect 77548 16192 77588 16232
rect 77932 16192 77972 16232
rect 78220 16192 78260 16232
rect 78604 16192 78644 16232
rect 78892 16192 78932 16232
rect 79180 16192 79220 16232
rect 63820 16108 63860 16148
rect 1996 16024 2036 16064
rect 2860 16024 2900 16064
rect 3628 16024 3668 16064
rect 33484 16024 33524 16064
rect 42604 16024 42644 16064
rect 45772 16024 45812 16064
rect 51532 16024 51572 16064
rect 53164 16024 53204 16064
rect 56140 16024 56180 16064
rect 57004 16024 57044 16064
rect 59404 16024 59444 16064
rect 59788 16024 59828 16064
rect 61900 16024 61940 16064
rect 64204 16024 64244 16064
rect 66220 16024 66260 16064
rect 68620 16024 68660 16064
rect 73804 16024 73844 16064
rect 75820 16024 75860 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 4492 15688 4532 15728
rect 33964 15688 34004 15728
rect 40492 15688 40532 15728
rect 46060 15688 46100 15728
rect 50188 15688 50228 15728
rect 55468 15688 55508 15728
rect 59500 15688 59540 15728
rect 62956 15688 62996 15728
rect 67852 15688 67892 15728
rect 79468 15688 79508 15728
rect 3532 15604 3572 15644
rect 3820 15604 3860 15644
rect 32140 15604 32180 15644
rect 38380 15604 38420 15644
rect 53068 15604 53108 15644
rect 2284 15520 2324 15560
rect 3148 15520 3188 15560
rect 3724 15520 3764 15560
rect 3916 15520 3956 15560
rect 4300 15520 4340 15560
rect 4396 15520 4436 15560
rect 4588 15520 4628 15560
rect 31564 15520 31604 15560
rect 31756 15520 31796 15560
rect 31852 15520 31892 15560
rect 32044 15520 32084 15560
rect 32236 15520 32276 15560
rect 33388 15520 33428 15560
rect 33484 15520 33524 15560
rect 33580 15520 33620 15560
rect 33676 15520 33716 15560
rect 33868 15520 33908 15560
rect 34060 15520 34100 15560
rect 34156 15520 34196 15560
rect 34924 15520 34964 15560
rect 35116 15520 35156 15560
rect 35212 15520 35252 15560
rect 36268 15520 36308 15560
rect 36364 15520 36404 15560
rect 36460 15520 36500 15560
rect 36556 15520 36596 15560
rect 36748 15520 36788 15560
rect 36940 15520 36980 15560
rect 37036 15520 37076 15560
rect 37516 15520 37556 15560
rect 38284 15520 38324 15560
rect 38476 15520 38516 15560
rect 39052 15520 39092 15560
rect 39148 15520 39188 15560
rect 39244 15520 39284 15560
rect 39724 15520 39764 15560
rect 39820 15520 39860 15560
rect 40108 15520 40148 15560
rect 40396 15520 40436 15560
rect 40588 15520 40628 15560
rect 40684 15520 40724 15560
rect 41836 15520 41876 15560
rect 42028 15520 42068 15560
rect 42124 15520 42164 15560
rect 45484 15520 45524 15560
rect 45580 15520 45620 15560
rect 45676 15520 45716 15560
rect 45772 15520 45812 15560
rect 45964 15520 46004 15560
rect 46156 15520 46196 15560
rect 46252 15520 46292 15560
rect 47500 15520 47540 15560
rect 47692 15520 47732 15560
rect 47884 15520 47924 15560
rect 48076 15520 48116 15560
rect 50764 15520 50804 15560
rect 50860 15520 50900 15560
rect 51052 15520 51092 15560
rect 51244 15520 51284 15560
rect 51724 15520 51764 15560
rect 52684 15520 52724 15560
rect 53452 15520 53492 15560
rect 54316 15520 54356 15560
rect 57100 15520 57140 15560
rect 57484 15520 57524 15560
rect 58348 15520 58388 15560
rect 60556 15520 60596 15560
rect 60940 15520 60980 15560
rect 61804 15520 61844 15560
rect 64876 15520 64916 15560
rect 65068 15520 65108 15560
rect 65452 15520 65492 15560
rect 65836 15520 65876 15560
rect 66700 15520 66740 15560
rect 70060 15520 70100 15560
rect 70156 15520 70196 15560
rect 70348 15520 70388 15560
rect 70924 15520 70964 15560
rect 71020 15520 71060 15560
rect 71116 15520 71156 15560
rect 75148 15520 75188 15560
rect 75340 15520 75380 15560
rect 79372 15520 79412 15560
rect 844 15436 884 15476
rect 49996 15436 50036 15476
rect 50380 15436 50420 15476
rect 60364 15436 60404 15476
rect 68716 15436 68756 15476
rect 69868 15436 69908 15476
rect 70732 15436 70772 15476
rect 5068 15352 5108 15392
rect 31564 15352 31604 15392
rect 34924 15352 34964 15392
rect 35692 15352 35732 15392
rect 38092 15352 38132 15392
rect 40876 15352 40916 15392
rect 43852 15352 43892 15392
rect 48460 15352 48500 15392
rect 49132 15352 49172 15392
rect 52012 15352 52052 15392
rect 60172 15352 60212 15392
rect 68044 15352 68084 15392
rect 71308 15352 71348 15392
rect 72652 15352 72692 15392
rect 76684 15352 76724 15392
rect 652 15268 692 15308
rect 1132 15268 1172 15308
rect 36748 15268 36788 15308
rect 39436 15268 39476 15308
rect 41836 15268 41876 15308
rect 47596 15268 47636 15308
rect 47980 15268 48020 15308
rect 50188 15268 50228 15308
rect 50572 15268 50612 15308
rect 51052 15268 51092 15308
rect 59500 15268 59540 15308
rect 64972 15268 65012 15308
rect 68908 15268 68948 15308
rect 69676 15268 69716 15308
rect 70348 15268 70388 15308
rect 70540 15268 70580 15308
rect 75244 15268 75284 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 1516 14932 1556 14972
rect 3628 14932 3668 14972
rect 32908 14932 32948 14972
rect 34828 14932 34868 14972
rect 46348 14932 46388 14972
rect 47692 14932 47732 14972
rect 50380 14932 50420 14972
rect 53164 14932 53204 14972
rect 56908 14932 56948 14972
rect 60556 14932 60596 14972
rect 65452 14932 65492 14972
rect 72748 14932 72788 14972
rect 75340 14932 75380 14972
rect 1996 14848 2036 14888
rect 40012 14848 40052 14888
rect 45100 14848 45140 14888
rect 56716 14848 56756 14888
rect 57484 14848 57524 14888
rect 58636 14848 58676 14888
rect 60172 14848 60212 14888
rect 61804 14848 61844 14888
rect 64204 14848 64244 14888
rect 65932 14848 65972 14888
rect 75532 14848 75572 14888
rect 844 14764 884 14804
rect 1324 14764 1364 14804
rect 1708 14764 1748 14804
rect 2188 14764 2228 14804
rect 60364 14764 60404 14804
rect 62188 14764 62228 14804
rect 62956 14764 62996 14804
rect 63916 14764 63956 14804
rect 67180 14764 67220 14804
rect 2380 14680 2420 14720
rect 2476 14680 2516 14720
rect 2572 14680 2612 14720
rect 2668 14680 2708 14720
rect 2956 14680 2996 14720
rect 3244 14680 3284 14720
rect 3340 14680 3380 14720
rect 30220 14680 30260 14720
rect 30604 14680 30644 14720
rect 31468 14680 31508 14720
rect 32812 14680 32852 14720
rect 33004 14680 33044 14720
rect 33196 14680 33236 14720
rect 33388 14680 33428 14720
rect 33484 14680 33524 14720
rect 35980 14680 36020 14720
rect 36844 14680 36884 14720
rect 37228 14680 37268 14720
rect 38572 14680 38612 14720
rect 39436 14680 39476 14720
rect 39820 14680 39860 14720
rect 40012 14680 40052 14720
rect 40204 14680 40244 14720
rect 40300 14680 40340 14720
rect 41164 14680 41204 14720
rect 41260 14680 41300 14720
rect 41356 14680 41396 14720
rect 42700 14680 42740 14720
rect 42892 14680 42932 14720
rect 42988 14680 43028 14720
rect 43180 14680 43220 14720
rect 43276 14680 43316 14720
rect 43372 14680 43412 14720
rect 46060 14680 46100 14720
rect 46156 14680 46196 14720
rect 46348 14680 46388 14720
rect 47020 14680 47060 14720
rect 47308 14680 47348 14720
rect 48364 14680 48404 14720
rect 49228 14680 49268 14720
rect 51148 14680 51188 14720
rect 52012 14680 52052 14720
rect 53452 14680 53492 14720
rect 54892 14680 54932 14720
rect 56044 14680 56084 14720
rect 56332 14680 56372 14720
rect 56908 14680 56948 14720
rect 57100 14680 57140 14720
rect 57196 14680 57236 14720
rect 57388 14680 57428 14720
rect 57580 14680 57620 14720
rect 60556 14680 60596 14720
rect 60748 14680 60788 14720
rect 60844 14680 60884 14720
rect 61132 14680 61172 14720
rect 61420 14680 61460 14720
rect 62380 14680 62420 14720
rect 62476 14680 62516 14720
rect 62572 14680 62612 14720
rect 63820 14680 63860 14720
rect 64012 14680 64052 14720
rect 64588 14680 64628 14720
rect 64876 14680 64916 14720
rect 65164 14680 65204 14720
rect 65260 14680 65300 14720
rect 65452 14680 65492 14720
rect 67948 14680 67988 14720
rect 68812 14680 68852 14720
rect 70348 14680 70388 14720
rect 70732 14680 70772 14720
rect 71596 14680 71636 14720
rect 73612 14680 73652 14720
rect 73804 14680 73844 14720
rect 73900 14680 73940 14720
rect 74092 14680 74132 14720
rect 74188 14680 74228 14720
rect 74284 14680 74324 14720
rect 74380 14680 74420 14720
rect 74668 14680 74708 14720
rect 74956 14680 74996 14720
rect 47404 14596 47444 14636
rect 47980 14596 48020 14636
rect 50764 14596 50804 14636
rect 56428 14596 56468 14636
rect 61516 14596 61556 14636
rect 64492 14596 64532 14636
rect 67564 14596 67604 14636
rect 75052 14596 75092 14636
rect 75532 14638 75572 14678
rect 75724 14680 75764 14720
rect 75820 14680 75860 14720
rect 76204 14680 76244 14720
rect 76588 14680 76628 14720
rect 77452 14680 77492 14720
rect 652 14512 692 14552
rect 1132 14512 1172 14552
rect 32620 14512 32660 14552
rect 33292 14512 33332 14552
rect 37420 14512 37460 14552
rect 41452 14512 41492 14552
rect 42796 14512 42836 14552
rect 53164 14512 53204 14552
rect 61996 14512 62036 14552
rect 62764 14512 62804 14552
rect 67372 14512 67412 14552
rect 69964 14512 70004 14552
rect 73708 14512 73748 14552
rect 78604 14512 78644 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 1324 14176 1364 14216
rect 2860 14176 2900 14216
rect 7276 14176 7316 14216
rect 38572 14176 38612 14216
rect 39436 14176 39476 14216
rect 40012 14176 40052 14216
rect 42700 14176 42740 14216
rect 47020 14176 47060 14216
rect 56140 14176 56180 14216
rect 60556 14176 60596 14216
rect 61036 14176 61076 14216
rect 66988 14176 67028 14216
rect 69004 14176 69044 14216
rect 70732 14176 70772 14216
rect 71116 14176 71156 14216
rect 79372 14176 79412 14216
rect 43180 14092 43220 14132
rect 47692 14092 47732 14132
rect 52588 14092 52628 14132
rect 67468 14092 67508 14132
rect 70060 14092 70100 14132
rect 72172 14092 72212 14132
rect 75916 14092 75956 14132
rect 2092 14008 2132 14048
rect 2188 14008 2228 14048
rect 2284 14008 2324 14048
rect 2380 14008 2420 14048
rect 2668 14008 2708 14048
rect 2764 14008 2804 14048
rect 2956 14008 2996 14048
rect 3244 14008 3284 14048
rect 3532 14008 3572 14048
rect 3628 14008 3668 14048
rect 4396 14008 4436 14048
rect 4492 14008 4532 14048
rect 4684 14008 4724 14048
rect 4876 14008 4916 14048
rect 5260 14008 5300 14048
rect 6124 14008 6164 14048
rect 31660 14008 31700 14048
rect 31756 14008 31796 14048
rect 31852 14008 31892 14048
rect 31948 14008 31988 14048
rect 32236 14008 32276 14048
rect 32524 14008 32564 14048
rect 32620 14008 32660 14048
rect 33484 14008 33524 14048
rect 34348 14008 34388 14048
rect 37324 14008 37364 14048
rect 38284 14008 38324 14048
rect 38476 14008 38516 14048
rect 33100 13966 33140 14006
rect 38668 14008 38708 14048
rect 38764 14008 38804 14048
rect 39148 14008 39188 14048
rect 39244 14008 39284 14048
rect 39340 14008 39380 14048
rect 39820 14008 39860 14048
rect 39916 14008 39956 14048
rect 40108 14008 40148 14048
rect 40300 14008 40340 14048
rect 40684 14008 40724 14048
rect 41548 14008 41588 14048
rect 43276 14008 43316 14048
rect 43564 14008 43604 14048
rect 44620 14008 44660 14048
rect 45004 14008 45044 14048
rect 45868 14008 45908 14048
rect 47212 14008 47252 14048
rect 47596 14008 47636 14048
rect 47788 14008 47828 14048
rect 47884 14008 47924 14048
rect 51148 14008 51188 14048
rect 51244 14008 51284 14048
rect 51436 14008 51476 14048
rect 52492 14008 52532 14048
rect 52684 14008 52724 14048
rect 53250 14023 53290 14063
rect 53356 14008 53396 14048
rect 53548 14008 53588 14048
rect 53740 14008 53780 14048
rect 54124 14008 54164 14048
rect 54988 14008 55028 14048
rect 56428 14008 56468 14048
rect 56620 14008 56660 14048
rect 57772 14029 57812 14069
rect 57964 14008 58004 14048
rect 58156 14008 58196 14048
rect 58540 14008 58580 14048
rect 59404 14008 59444 14048
rect 61228 14008 61268 14048
rect 61612 14008 61652 14048
rect 62476 14008 62516 14048
rect 63820 14008 63860 14048
rect 63916 14008 63956 14048
rect 64108 14008 64148 14048
rect 64588 14008 64628 14048
rect 64972 14008 65012 14048
rect 65836 14008 65876 14048
rect 67276 14008 67316 14048
rect 67372 14008 67412 14048
rect 67564 14008 67604 14048
rect 68044 14008 68084 14048
rect 68140 14008 68180 14048
rect 68332 14008 68372 14048
rect 68524 14008 68564 14048
rect 68620 14008 68660 14048
rect 68716 14008 68756 14048
rect 68812 14008 68852 14048
rect 69676 14008 69716 14048
rect 69964 14008 70004 14048
rect 72556 14008 72596 14048
rect 73445 14008 73485 14048
rect 74764 14008 74804 14048
rect 74956 14008 74996 14048
rect 75052 14008 75092 14048
rect 75820 14008 75860 14048
rect 76012 14008 76052 14048
rect 76972 14008 77012 14048
rect 77356 14008 77396 14048
rect 78220 14008 78260 14048
rect 1516 13924 1556 13964
rect 60844 13924 60884 13964
rect 63628 13924 63668 13964
rect 69196 13924 69236 13964
rect 70540 13924 70580 13964
rect 70924 13924 70964 13964
rect 1900 13840 1940 13880
rect 4684 13840 4724 13880
rect 30700 13840 30740 13880
rect 32908 13840 32948 13880
rect 43852 13840 43892 13880
rect 51628 13840 51668 13880
rect 74764 13840 74804 13880
rect 3916 13756 3956 13796
rect 35500 13756 35540 13796
rect 42892 13756 42932 13796
rect 51436 13756 51476 13796
rect 53548 13756 53588 13796
rect 56140 13756 56180 13796
rect 56524 13756 56564 13796
rect 57868 13756 57908 13796
rect 61036 13756 61076 13796
rect 64108 13756 64148 13796
rect 68332 13756 68372 13796
rect 70348 13756 70388 13796
rect 70732 13756 70772 13796
rect 71116 13756 71156 13796
rect 74572 13756 74612 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 3820 13420 3860 13460
rect 4300 13420 4340 13460
rect 32812 13420 32852 13460
rect 42796 13420 42836 13460
rect 45484 13420 45524 13460
rect 46156 13420 46196 13460
rect 47212 13420 47252 13460
rect 51628 13420 51668 13460
rect 58924 13420 58964 13460
rect 61132 13420 61172 13460
rect 61900 13420 61940 13460
rect 1036 13336 1076 13376
rect 5548 13336 5588 13376
rect 33580 13336 33620 13376
rect 39340 13336 39380 13376
rect 40780 13336 40820 13376
rect 47404 13336 47444 13376
rect 52492 13336 52532 13376
rect 62188 13378 62228 13418
rect 64492 13420 64532 13460
rect 70156 13420 70196 13460
rect 76492 13420 76532 13460
rect 56332 13336 56372 13376
rect 58444 13336 58484 13376
rect 65164 13336 65204 13376
rect 70924 13336 70964 13376
rect 72076 13336 72116 13376
rect 76108 13336 76148 13376
rect 77068 13336 77108 13376
rect 77452 13336 77492 13376
rect 844 13252 884 13292
rect 1228 13252 1268 13292
rect 1804 13168 1844 13208
rect 2668 13168 2708 13208
rect 4204 13168 4244 13208
rect 4396 13168 4436 13208
rect 4972 13168 5012 13208
rect 32812 13168 32852 13208
rect 33004 13168 33044 13208
rect 33118 13179 33158 13219
rect 34924 13168 34964 13208
rect 35020 13168 35060 13208
rect 35212 13168 35252 13208
rect 36556 13168 36596 13208
rect 36748 13168 36788 13208
rect 37324 13168 37364 13208
rect 38188 13168 38228 13208
rect 41452 13168 41492 13208
rect 41644 13168 41684 13208
rect 41740 13168 41780 13208
rect 42700 13168 42740 13208
rect 42892 13168 42932 13208
rect 43084 13168 43124 13208
rect 43468 13168 43508 13208
rect 44332 13168 44372 13208
rect 45676 13168 45716 13208
rect 45772 13168 45812 13208
rect 45868 13168 45908 13208
rect 45964 13168 46004 13208
rect 46156 13168 46196 13208
rect 46348 13168 46388 13208
rect 46444 13168 46484 13208
rect 46828 13168 46868 13208
rect 47884 13168 47924 13208
rect 48076 13168 48116 13208
rect 48172 13168 48212 13208
rect 48556 13168 48596 13208
rect 48748 13168 48788 13208
rect 49612 13168 49652 13208
rect 50476 13168 50516 13208
rect 51916 13168 51956 13208
rect 52108 13168 52148 13208
rect 54412 13168 54452 13208
rect 54508 13168 54548 13208
rect 54700 13168 54740 13208
rect 55084 13168 55124 13208
rect 55180 13168 55220 13208
rect 55276 13168 55316 13208
rect 55372 13168 55412 13208
rect 56044 13168 56084 13208
rect 56140 13168 56180 13208
rect 56332 13168 56372 13208
rect 56524 13168 56564 13208
rect 56716 13154 56756 13194
rect 56812 13168 56852 13208
rect 57772 13168 57812 13208
rect 58060 13168 58100 13208
rect 58636 13168 58676 13208
rect 58732 13168 58772 13208
rect 58924 13168 58964 13208
rect 60844 13168 60884 13208
rect 60940 13168 60980 13208
rect 61132 13168 61172 13208
rect 61324 13168 61364 13208
rect 61420 13168 61460 13208
rect 61516 13205 61556 13245
rect 74668 13252 74708 13292
rect 61612 13168 61652 13208
rect 61804 13168 61844 13208
rect 61996 13168 62036 13208
rect 64204 13168 64244 13208
rect 64300 13168 64340 13208
rect 64492 13168 64532 13208
rect 64684 13168 64724 13208
rect 64780 13168 64820 13208
rect 64876 13168 64916 13208
rect 64972 13168 65012 13208
rect 68620 13168 68660 13208
rect 68716 13168 68756 13208
rect 68812 13168 68852 13208
rect 69004 13168 69044 13208
rect 69100 13168 69140 13208
rect 69292 13168 69332 13208
rect 69676 13168 69716 13208
rect 69868 13168 69908 13208
rect 70060 13168 70100 13208
rect 70252 13168 70292 13208
rect 72652 13168 72692 13208
rect 73516 13168 73556 13208
rect 74956 13168 74996 13208
rect 75052 13168 75092 13208
rect 75148 13168 75188 13208
rect 75436 13168 75476 13208
rect 75724 13168 75764 13208
rect 75820 13168 75860 13208
rect 76492 13168 76532 13208
rect 76684 13168 76724 13208
rect 76780 13168 76820 13208
rect 76972 13168 77012 13208
rect 77164 13168 77204 13208
rect 1420 13084 1460 13124
rect 36652 13084 36692 13124
rect 36940 13084 36980 13124
rect 41548 13084 41588 13124
rect 47980 13084 48020 13124
rect 48652 13084 48692 13124
rect 49228 13084 49268 13124
rect 52012 13084 52052 13124
rect 54604 13084 54644 13124
rect 58156 13084 58196 13124
rect 69772 13084 69812 13124
rect 72268 13084 72308 13124
rect 652 13000 692 13040
rect 35116 13000 35156 13040
rect 51628 13000 51668 13040
rect 56620 13000 56660 13040
rect 68524 13000 68564 13040
rect 69196 13000 69236 13040
rect 74860 13000 74900 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 2380 12664 2420 12704
rect 47692 12664 47732 12704
rect 48940 12664 48980 12704
rect 54412 12664 54452 12704
rect 57196 12664 57236 12704
rect 57964 12664 58004 12704
rect 62092 12664 62132 12704
rect 67180 12664 67220 12704
rect 72844 12664 72884 12704
rect 74380 12664 74420 12704
rect 4108 12580 4148 12620
rect 48364 12580 48404 12620
rect 54796 12580 54836 12620
rect 2284 12496 2324 12536
rect 2476 12496 2516 12536
rect 2572 12496 2612 12536
rect 2764 12496 2804 12536
rect 2956 12496 2996 12536
rect 3052 12496 3092 12536
rect 4012 12496 4052 12536
rect 4204 12496 4244 12536
rect 4780 12496 4820 12536
rect 5644 12496 5684 12536
rect 29932 12496 29972 12536
rect 31372 12496 31412 12536
rect 33868 12496 33908 12536
rect 34252 12496 34292 12536
rect 35116 12496 35156 12536
rect 36748 12496 36788 12536
rect 36844 12496 36884 12536
rect 37132 12496 37172 12536
rect 39148 12496 39188 12536
rect 39532 12496 39572 12536
rect 40396 12496 40436 12536
rect 41932 12496 41972 12536
rect 42028 12496 42068 12536
rect 42220 12496 42260 12536
rect 42412 12496 42452 12536
rect 42508 12496 42548 12536
rect 42604 12496 42644 12536
rect 45292 12496 45332 12536
rect 45676 12496 45716 12536
rect 46540 12496 46580 12536
rect 47980 12496 48020 12536
rect 48268 12496 48308 12536
rect 48844 12496 48884 12536
rect 49036 12496 49076 12536
rect 49132 12496 49172 12536
rect 49324 12496 49364 12536
rect 49516 12496 49556 12536
rect 52012 12496 52052 12536
rect 52396 12496 52436 12536
rect 53293 12496 53333 12536
rect 55180 12496 55220 12536
rect 56044 12496 56084 12536
rect 58156 12496 58196 12536
rect 58348 12496 58388 12536
rect 59308 12496 59348 12536
rect 59509 12509 59549 12549
rect 61996 12496 62036 12536
rect 62188 12496 62228 12536
rect 62284 12496 62324 12536
rect 63296 12496 63336 12536
rect 63628 12496 63668 12536
rect 63724 12496 63764 12536
rect 64396 12496 64436 12536
rect 64588 12496 64628 12536
rect 64780 12496 64820 12536
rect 65164 12496 65204 12536
rect 66028 12496 66068 12536
rect 67372 12496 67412 12536
rect 67756 12496 67796 12536
rect 68620 12496 68660 12536
rect 69964 12496 70004 12536
rect 70060 12496 70100 12536
rect 70252 12538 70292 12578
rect 76108 12580 76148 12620
rect 70444 12496 70484 12536
rect 70828 12496 70868 12536
rect 71692 12496 71732 12536
rect 74284 12496 74324 12536
rect 74476 12496 74516 12536
rect 74572 12496 74612 12536
rect 74764 12496 74804 12536
rect 74956 12496 74996 12536
rect 75052 12496 75092 12536
rect 76012 12496 76052 12536
rect 76204 12496 76244 12536
rect 76876 12496 76916 12536
rect 77260 12496 77300 12536
rect 78124 12496 78164 12536
rect 844 12412 884 12452
rect 1324 12412 1364 12452
rect 1708 12412 1748 12452
rect 49420 12412 49460 12452
rect 50284 12412 50324 12452
rect 51148 12412 51188 12452
rect 51628 12412 51668 12452
rect 57772 12412 57812 12452
rect 652 12328 692 12368
rect 1132 12328 1172 12368
rect 1900 12328 1940 12368
rect 2764 12328 2804 12368
rect 4972 12328 5012 12368
rect 5836 12328 5876 12368
rect 36268 12328 36308 12368
rect 37420 12328 37460 12368
rect 41548 12328 41588 12368
rect 42892 12328 42932 12368
rect 48652 12328 48692 12368
rect 49708 12328 49748 12368
rect 58252 12328 58292 12368
rect 59788 12328 59828 12368
rect 70252 12328 70292 12368
rect 74764 12328 74804 12368
rect 1516 12244 1556 12284
rect 36460 12244 36500 12284
rect 42220 12244 42260 12284
rect 47692 12244 47732 12284
rect 50092 12244 50132 12284
rect 50956 12244 50996 12284
rect 51820 12244 51860 12284
rect 57964 12244 58004 12284
rect 59404 12244 59444 12284
rect 64012 12244 64052 12284
rect 64492 12244 64532 12284
rect 69772 12244 69812 12284
rect 79276 12244 79316 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 7372 11908 7412 11948
rect 34828 11908 34868 11948
rect 36844 11908 36884 11948
rect 38860 11908 38900 11948
rect 44812 11908 44852 11948
rect 48268 11908 48308 11948
rect 51724 11908 51764 11948
rect 61708 11908 61748 11948
rect 64204 11908 64244 11948
rect 68908 11908 68948 11948
rect 70156 11908 70196 11948
rect 70540 11908 70580 11948
rect 74956 11908 74996 11948
rect 76492 11908 76532 11948
rect 34348 11824 34388 11864
rect 36268 11824 36308 11864
rect 37036 11824 37076 11864
rect 39436 11824 39476 11864
rect 39724 11824 39764 11864
rect 42220 11824 42260 11864
rect 45004 11824 45044 11864
rect 45772 11824 45812 11864
rect 48940 11824 48980 11864
rect 49228 11824 49268 11864
rect 51532 11824 51572 11864
rect 55276 11824 55316 11864
rect 56332 11824 56372 11864
rect 57292 11824 57332 11864
rect 62092 11824 62132 11864
rect 65260 11824 65300 11864
rect 67468 11824 67508 11864
rect 76012 11824 76052 11864
rect 77356 11824 77396 11864
rect 1132 11740 1172 11780
rect 57484 11740 57524 11780
rect 1708 11656 1748 11696
rect 2572 11656 2612 11696
rect 3916 11656 3956 11696
rect 4108 11656 4148 11696
rect 4492 11656 4532 11696
rect 4684 11656 4724 11696
rect 4780 11656 4820 11696
rect 4972 11656 5012 11696
rect 5356 11656 5396 11696
rect 6220 11656 6260 11696
rect 34828 11656 34868 11696
rect 35020 11656 35060 11696
rect 35116 11656 35156 11696
rect 35308 11656 35348 11696
rect 35404 11656 35444 11696
rect 35500 11656 35540 11696
rect 35596 11656 35636 11696
rect 36172 11656 36212 11696
rect 36364 11656 36404 11696
rect 36556 11656 36596 11696
rect 36652 11656 36692 11696
rect 36844 11656 36884 11696
rect 38860 11656 38900 11696
rect 39052 11656 39092 11696
rect 39148 11656 39188 11696
rect 39340 11656 39380 11696
rect 39532 11656 39572 11696
rect 41548 11656 41588 11696
rect 41836 11656 41876 11696
rect 42412 11656 42452 11696
rect 42796 11656 42836 11696
rect 43660 11656 43700 11696
rect 47788 11656 47828 11696
rect 47884 11656 47924 11696
rect 47980 11656 48020 11696
rect 48076 11656 48116 11696
rect 48268 11656 48308 11696
rect 48460 11656 48500 11696
rect 48556 11656 48596 11696
rect 49228 11656 49268 11696
rect 49420 11656 49460 11696
rect 49516 11656 49556 11696
rect 50860 11656 50900 11696
rect 51148 11656 51188 11696
rect 51724 11656 51764 11696
rect 51916 11656 51956 11696
rect 52012 11656 52052 11696
rect 52204 11656 52244 11696
rect 52396 11656 52436 11696
rect 56524 11656 56564 11696
rect 56620 11656 56660 11696
rect 56716 11656 56756 11696
rect 56812 11656 56852 11696
rect 57676 11656 57716 11696
rect 57868 11656 57908 11696
rect 57964 11656 58004 11696
rect 58252 11656 58292 11696
rect 58348 11656 58388 11696
rect 58444 11656 58484 11696
rect 58828 11656 58868 11696
rect 59020 11656 59060 11696
rect 59116 11656 59156 11696
rect 59692 11656 59732 11696
rect 60556 11656 60596 11696
rect 62764 11656 62804 11696
rect 62860 11656 62900 11696
rect 62956 11656 62996 11696
rect 63052 11656 63092 11696
rect 63244 11656 63284 11696
rect 63436 11656 63476 11696
rect 63532 11656 63572 11696
rect 63820 11656 63860 11696
rect 63916 11656 63956 11696
rect 64012 11656 64052 11696
rect 64204 11656 64244 11696
rect 64396 11656 64436 11696
rect 64492 11656 64532 11696
rect 68908 11656 68948 11696
rect 69100 11656 69140 11696
rect 69196 11656 69236 11696
rect 69484 11656 69524 11696
rect 69772 11656 69812 11696
rect 70444 11656 70484 11696
rect 70636 11656 70676 11696
rect 72940 11656 72980 11696
rect 73804 11656 73844 11696
rect 75340 11656 75380 11696
rect 75628 11656 75668 11696
rect 75724 11656 75764 11696
rect 76492 11656 76532 11696
rect 76684 11656 76724 11696
rect 76780 11656 76820 11696
rect 76972 11656 77012 11696
rect 77164 11656 77204 11696
rect 1324 11572 1364 11612
rect 4012 11572 4052 11612
rect 4588 11572 4628 11612
rect 41932 11572 41972 11612
rect 51244 11572 51284 11612
rect 52300 11572 52340 11612
rect 58924 11572 58964 11612
rect 59308 11572 59348 11612
rect 69868 11572 69908 11612
rect 72556 11572 72596 11612
rect 77068 11572 77108 11612
rect 940 11488 980 11528
rect 3724 11488 3764 11528
rect 7372 11488 7412 11528
rect 57772 11488 57812 11528
rect 58156 11488 58196 11528
rect 63340 11488 63380 11528
rect 74956 11488 74996 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 652 11152 692 11192
rect 42604 11152 42644 11192
rect 46732 11152 46772 11192
rect 48172 11152 48212 11192
rect 56332 11152 56372 11192
rect 58924 11152 58964 11192
rect 60940 11152 60980 11192
rect 75244 11152 75284 11192
rect 3532 11068 3572 11108
rect 4972 11068 5012 11108
rect 59404 11068 59444 11108
rect 63340 11068 63380 11108
rect 76204 11068 76244 11108
rect 1804 10984 1844 11024
rect 1900 10984 1940 11024
rect 1996 10984 2036 11024
rect 2092 10984 2132 11024
rect 2284 10984 2324 11024
rect 2476 10984 2516 11024
rect 2572 10984 2612 11024
rect 3148 10984 3188 11024
rect 3436 10984 3476 11024
rect 4876 10984 4916 11024
rect 5068 10984 5108 11024
rect 36460 10984 36500 11024
rect 36556 10984 36596 11024
rect 36748 10984 36788 11024
rect 36940 10984 36980 11024
rect 37036 10984 37076 11024
rect 37228 10984 37268 11024
rect 37420 10984 37460 11024
rect 37516 10984 37556 11024
rect 37612 10984 37652 11024
rect 37708 10984 37748 11024
rect 38572 10984 38612 11024
rect 38860 10984 38900 11024
rect 38956 10984 38996 11024
rect 39436 10984 39476 11024
rect 39628 10984 39668 11024
rect 40684 10984 40724 11024
rect 42892 10984 42932 11024
rect 43084 10984 43124 11024
rect 43948 10984 43988 11024
rect 44140 10984 44180 11024
rect 44332 10984 44372 11024
rect 44716 10984 44756 11024
rect 45580 10984 45620 11024
rect 46924 10984 46964 11024
rect 47116 10984 47156 11024
rect 49324 10984 49364 11024
rect 50188 10984 50228 11024
rect 50572 10984 50612 11024
rect 50764 10984 50804 11024
rect 50860 10984 50900 11024
rect 50956 10984 50996 11024
rect 51052 10984 51092 11024
rect 51244 10984 51284 11024
rect 51436 10984 51476 11024
rect 51532 10984 51572 11024
rect 52492 10984 52532 11024
rect 52684 10984 52724 11024
rect 52780 10984 52820 11024
rect 53068 10984 53108 11024
rect 53164 10984 53204 11024
rect 53260 10961 53300 11001
rect 53452 10984 53492 11024
rect 53548 10984 53588 11024
rect 53740 10984 53780 11024
rect 53932 10984 53972 11024
rect 54316 10984 54356 11024
rect 55180 10984 55220 11024
rect 56524 10984 56564 11024
rect 56908 10984 56948 11024
rect 57772 10984 57812 11024
rect 59500 10984 59540 11024
rect 59788 10984 59828 11024
rect 62092 10984 62132 11024
rect 62956 10984 62996 11024
rect 64492 10984 64532 11024
rect 64684 10984 64724 11024
rect 64876 10984 64916 11024
rect 65068 10984 65108 11024
rect 65164 10984 65204 11024
rect 68908 10984 68948 11024
rect 69100 10984 69140 11024
rect 69196 10984 69236 11024
rect 74668 10984 74708 11024
rect 74764 10984 74804 11024
rect 74860 10984 74900 11024
rect 74956 10984 74996 11024
rect 75148 10984 75188 11024
rect 75340 10984 75380 11024
rect 75436 10984 75476 11024
rect 75628 10984 75668 11024
rect 75820 10984 75860 11024
rect 75916 10984 75956 11024
rect 76108 10984 76148 11024
rect 76311 10983 76351 11023
rect 77068 10984 77108 11024
rect 77260 10984 77300 11024
rect 844 10900 884 10940
rect 1228 10900 1268 10940
rect 1612 10900 1652 10940
rect 39532 10900 39572 10940
rect 51916 10900 51956 10940
rect 64588 10900 64628 10940
rect 69580 10900 69620 10940
rect 69964 10900 70004 10940
rect 70348 10900 70388 10940
rect 70540 10900 70580 10940
rect 71116 10900 71156 10940
rect 76492 10889 76532 10929
rect 1420 10816 1460 10856
rect 2284 10816 2324 10856
rect 3820 10816 3860 10856
rect 36748 10816 36788 10856
rect 39244 10816 39284 10856
rect 40012 10816 40052 10856
rect 51244 10816 51284 10856
rect 53740 10816 53780 10856
rect 65740 10816 65780 10856
rect 71308 10816 71348 10856
rect 73036 10816 73076 10856
rect 75628 10816 75668 10856
rect 77644 10816 77684 10856
rect 1036 10732 1076 10772
rect 37228 10732 37268 10772
rect 42988 10732 43028 10772
rect 44044 10732 44084 10772
rect 47020 10732 47060 10772
rect 51724 10732 51764 10772
rect 52492 10732 52532 10772
rect 59116 10732 59156 10772
rect 64876 10732 64916 10772
rect 68908 10732 68948 10772
rect 69388 10732 69428 10772
rect 69772 10732 69812 10772
rect 70156 10732 70196 10772
rect 70732 10732 70772 10772
rect 70924 10732 70964 10772
rect 76684 10732 76724 10772
rect 77164 10732 77204 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 2572 10396 2612 10436
rect 38860 10396 38900 10436
rect 41836 10396 41876 10436
rect 42316 10396 42356 10436
rect 44812 10396 44852 10436
rect 49228 10396 49268 10436
rect 53740 10396 53780 10436
rect 58060 10396 58100 10436
rect 63436 10396 63476 10436
rect 64204 10396 64244 10436
rect 67660 10396 67700 10436
rect 72940 10396 72980 10436
rect 75916 10396 75956 10436
rect 76876 10396 76916 10436
rect 1516 10312 1556 10352
rect 3052 10312 3092 10352
rect 43564 10312 43604 10352
rect 53452 10312 53492 10352
rect 54412 10312 54452 10352
rect 57580 10312 57620 10352
rect 58732 10312 58772 10352
rect 62380 10312 62420 10352
rect 67852 10312 67892 10352
rect 69964 10312 70004 10352
rect 70348 10312 70388 10352
rect 844 10228 884 10268
rect 1708 10228 1748 10268
rect 3244 10228 3284 10268
rect 7180 10228 7220 10268
rect 42124 10228 42164 10268
rect 57388 10228 57428 10268
rect 58924 10228 58964 10268
rect 70156 10228 70196 10268
rect 79468 10228 79508 10268
rect 2572 10144 2612 10184
rect 2764 10144 2804 10184
rect 2870 10129 2910 10169
rect 5164 10144 5204 10184
rect 6028 10144 6068 10184
rect 36460 10144 36500 10184
rect 36844 10144 36884 10184
rect 37708 10144 37748 10184
rect 39820 10144 39860 10184
rect 40684 10144 40724 10184
rect 43948 10144 43988 10184
rect 44236 10144 44276 10184
rect 44524 10144 44564 10184
rect 44620 10144 44660 10184
rect 44812 10144 44852 10184
rect 46348 10144 46388 10184
rect 46540 10144 46580 10184
rect 46636 10144 46676 10184
rect 46828 10144 46868 10184
rect 47212 10144 47252 10184
rect 48076 10144 48116 10184
rect 49804 10144 49844 10184
rect 50188 10144 50228 10184
rect 51052 10144 51092 10184
rect 52780 10144 52820 10184
rect 53068 10144 53108 10184
rect 53644 10144 53684 10184
rect 53836 10144 53876 10184
rect 57772 10144 57812 10184
rect 57868 10144 57908 10184
rect 58060 10144 58100 10184
rect 58252 10144 58292 10184
rect 58444 10144 58484 10184
rect 58540 10144 58580 10184
rect 59116 10144 59156 10184
rect 59308 10144 59348 10184
rect 59500 10144 59540 10184
rect 59692 10144 59732 10184
rect 63436 10144 63476 10184
rect 63628 10144 63668 10184
rect 63724 10144 63764 10184
rect 64588 10144 64628 10184
rect 64876 10144 64916 10184
rect 65260 10144 65300 10184
rect 65644 10144 65684 10184
rect 66508 10144 66548 10184
rect 68332 10144 68372 10184
rect 68428 10144 68468 10184
rect 68524 10144 68564 10184
rect 68716 10144 68756 10184
rect 68908 10144 68948 10184
rect 69004 10144 69044 10184
rect 69292 10144 69332 10184
rect 69580 10144 69620 10184
rect 69676 10144 69716 10184
rect 70924 10144 70964 10184
rect 71788 10144 71828 10184
rect 73900 10144 73940 10184
rect 74764 10144 74804 10184
rect 76204 10144 76244 10184
rect 76492 10144 76532 10184
rect 76588 10144 76628 10184
rect 77452 10144 77492 10184
rect 78316 10144 78356 10184
rect 4780 10060 4820 10100
rect 39436 10060 39476 10100
rect 43852 10060 43892 10100
rect 46444 10060 46484 10100
rect 53164 10060 53204 10100
rect 59212 10060 59252 10100
rect 59596 10060 59636 10100
rect 64492 10060 64532 10100
rect 68236 10060 68276 10100
rect 68812 10060 68852 10100
rect 70540 10060 70580 10100
rect 73516 10060 73556 10100
rect 77068 10060 77108 10100
rect 652 9976 692 10016
rect 52204 9976 52244 10016
rect 58348 9976 58388 10016
rect 75916 9976 75956 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 652 9640 692 9680
rect 3436 9640 3476 9680
rect 4492 9640 4532 9680
rect 40204 9640 40244 9680
rect 42796 9640 42836 9680
rect 51532 9640 51572 9680
rect 52492 9640 52532 9680
rect 52780 9640 52820 9680
rect 61996 9640 62036 9680
rect 64588 9640 64628 9680
rect 69292 9640 69332 9680
rect 70636 9640 70676 9680
rect 75532 9640 75572 9680
rect 77164 9640 77204 9680
rect 62188 9556 62228 9596
rect 64876 9556 64916 9596
rect 65356 9556 65396 9596
rect 66892 9556 66932 9596
rect 1036 9472 1076 9512
rect 1420 9472 1460 9512
rect 2284 9472 2324 9512
rect 3628 9472 3668 9512
rect 3820 9472 3860 9512
rect 4396 9472 4436 9512
rect 4588 9472 4628 9512
rect 4684 9472 4724 9512
rect 4876 9472 4916 9512
rect 5068 9472 5108 9512
rect 39244 9472 39284 9512
rect 39340 9472 39380 9512
rect 39532 9472 39572 9512
rect 40012 9472 40052 9512
rect 40108 9472 40148 9512
rect 40300 9472 40340 9512
rect 40684 9472 40724 9512
rect 40780 9472 40820 9512
rect 40876 9472 40916 9512
rect 40972 9472 41012 9512
rect 41740 9472 41780 9512
rect 41836 9472 41876 9512
rect 42028 9472 42068 9512
rect 42220 9472 42260 9512
rect 42316 9472 42356 9512
rect 42508 9472 42548 9512
rect 42892 9472 42932 9512
rect 42988 9472 43028 9512
rect 43084 9472 43124 9512
rect 43948 9472 43988 9512
rect 44140 9472 44180 9512
rect 46636 9472 46676 9512
rect 46732 9472 46772 9512
rect 47020 9472 47060 9512
rect 51436 9472 51476 9512
rect 51628 9472 51668 9512
rect 51724 9472 51764 9512
rect 52204 9472 52244 9512
rect 52300 9472 52340 9512
rect 52396 9472 52436 9512
rect 52684 9472 52724 9512
rect 52876 9472 52916 9512
rect 52972 9472 53012 9512
rect 53644 9472 53684 9512
rect 53836 9472 53876 9512
rect 54124 9472 54164 9512
rect 54316 9472 54356 9512
rect 57772 9472 57812 9512
rect 57964 9472 58004 9512
rect 58060 9472 58100 9512
rect 58348 9472 58388 9512
rect 58636 9472 58676 9512
rect 58732 9472 58772 9512
rect 59596 9472 59636 9512
rect 59980 9472 60020 9512
rect 60844 9472 60884 9512
rect 62572 9472 62612 9512
rect 63436 9472 63476 9512
rect 64780 9472 64820 9512
rect 64972 9472 65012 9512
rect 65068 9472 65108 9512
rect 65260 9472 65300 9512
rect 65452 9472 65492 9512
rect 67276 9472 67316 9512
rect 68140 9472 68180 9512
rect 69484 9472 69524 9512
rect 69580 9472 69620 9512
rect 69772 9472 69812 9512
rect 69964 9472 70004 9512
rect 70156 9472 70196 9512
rect 70252 9472 70292 9512
rect 70828 9472 70868 9512
rect 70924 9472 70964 9512
rect 71020 9472 71060 9512
rect 71308 9472 71348 9512
rect 71500 9472 71540 9512
rect 71692 9472 71732 9512
rect 71884 9472 71924 9512
rect 75628 9472 75668 9512
rect 75724 9472 75764 9512
rect 75820 9472 75860 9512
rect 76012 9472 76052 9512
rect 76204 9458 76244 9498
rect 76300 9472 76340 9512
rect 77068 9472 77108 9512
rect 77260 9472 77300 9512
rect 77356 9472 77396 9512
rect 77548 9472 77588 9512
rect 77644 9472 77684 9512
rect 77740 9472 77780 9512
rect 844 9388 884 9428
rect 57388 9388 57428 9428
rect 59404 9388 59444 9428
rect 70444 9388 70484 9428
rect 76492 9388 76532 9428
rect 4972 9304 5012 9344
rect 5260 9304 5300 9344
rect 39532 9304 39572 9344
rect 41548 9304 41588 9344
rect 42028 9304 42068 9344
rect 44620 9304 44660 9344
rect 47308 9304 47348 9344
rect 50380 9304 50420 9344
rect 54796 9304 54836 9344
rect 56428 9304 56468 9344
rect 69964 9304 70004 9344
rect 72172 9304 72212 9344
rect 73996 9304 74036 9344
rect 76684 9304 76724 9344
rect 3724 9220 3764 9260
rect 42508 9220 42548 9260
rect 44044 9220 44084 9260
rect 46348 9220 46388 9260
rect 53740 9220 53780 9260
rect 54220 9220 54260 9260
rect 57580 9220 57620 9260
rect 57772 9220 57812 9260
rect 59020 9220 59060 9260
rect 59212 9220 59252 9260
rect 64588 9220 64628 9260
rect 69772 9220 69812 9260
rect 70636 9220 70676 9260
rect 71404 9220 71444 9260
rect 71788 9220 71828 9260
rect 76012 9220 76052 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 652 8884 692 8924
rect 3436 8884 3476 8924
rect 43948 8884 43988 8924
rect 46540 8884 46580 8924
rect 53836 8884 53876 8924
rect 56716 8884 56756 8924
rect 59500 8884 59540 8924
rect 68428 8884 68468 8924
rect 69868 8884 69908 8924
rect 71500 8884 71540 8924
rect 74092 8884 74132 8924
rect 75916 8884 75956 8924
rect 79468 8884 79508 8924
rect 1516 8800 1556 8840
rect 5260 8800 5300 8840
rect 49324 8800 49364 8840
rect 50956 8800 50996 8840
rect 60076 8800 60116 8840
rect 64972 8800 65012 8840
rect 70156 8800 70196 8840
rect 74284 8800 74324 8840
rect 76876 8800 76916 8840
rect 844 8716 884 8756
rect 58252 8716 58292 8756
rect 58732 8716 58772 8756
rect 59692 8716 59732 8756
rect 64780 8716 64820 8756
rect 68908 8716 68948 8756
rect 1708 8632 1748 8672
rect 1804 8632 1844 8672
rect 1900 8632 1940 8672
rect 2188 8632 2228 8672
rect 2380 8632 2420 8672
rect 2476 8632 2516 8672
rect 2764 8632 2804 8672
rect 3052 8632 3092 8672
rect 3148 8632 3188 8672
rect 41932 8632 41972 8672
rect 42796 8632 42836 8672
rect 44524 8632 44564 8672
rect 45388 8632 45428 8672
rect 46732 8632 46772 8672
rect 46924 8632 46964 8672
rect 48460 8632 48500 8672
rect 48652 8632 48692 8672
rect 48844 8632 48884 8672
rect 49036 8632 49076 8672
rect 49132 8632 49172 8672
rect 53164 8632 53204 8672
rect 53452 8632 53492 8672
rect 54700 8632 54740 8672
rect 55564 8632 55604 8672
rect 57772 8632 57812 8672
rect 57868 8632 57908 8672
rect 57964 8632 58004 8672
rect 58060 8632 58100 8672
rect 58636 8632 58676 8672
rect 58828 8632 58868 8672
rect 59020 8632 59060 8672
rect 59212 8632 59252 8672
rect 59308 8632 59348 8672
rect 60460 8632 60500 8672
rect 60652 8632 60692 8672
rect 63820 8632 63860 8672
rect 63916 8632 63956 8672
rect 64012 8632 64052 8672
rect 64108 8632 64148 8672
rect 64300 8632 64340 8672
rect 64492 8632 64532 8672
rect 64588 8632 64628 8672
rect 66412 8632 66452 8672
rect 67276 8632 67316 8672
rect 69292 8632 69332 8672
rect 69484 8632 69524 8672
rect 69580 8632 69620 8672
rect 69772 8632 69812 8672
rect 69964 8632 70004 8672
rect 70828 8632 70868 8672
rect 71116 8632 71156 8672
rect 72076 8632 72116 8672
rect 72940 8632 72980 8672
rect 75628 8632 75668 8672
rect 75724 8632 75764 8672
rect 75916 8632 75956 8672
rect 76204 8632 76244 8672
rect 76492 8632 76532 8672
rect 77452 8632 77492 8672
rect 78316 8632 78356 8672
rect 1996 8548 2036 8588
rect 2284 8548 2324 8588
rect 41548 8548 41588 8588
rect 44140 8548 44180 8588
rect 46828 8548 46868 8588
rect 48556 8548 48596 8588
rect 53548 8548 53588 8588
rect 54316 8548 54356 8588
rect 60556 8548 60596 8588
rect 64396 8548 64436 8588
rect 66028 8548 66068 8588
rect 71212 8548 71252 8588
rect 71692 8548 71732 8588
rect 76588 8548 76628 8588
rect 77068 8548 77108 8588
rect 43948 8464 43988 8504
rect 46540 8464 46580 8504
rect 48940 8464 48980 8504
rect 58444 8464 58484 8504
rect 59116 8464 59156 8504
rect 68428 8464 68468 8504
rect 69100 8464 69140 8504
rect 69388 8464 69428 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 652 8128 692 8168
rect 4396 8128 4436 8168
rect 7180 8128 7220 8168
rect 44908 8128 44948 8168
rect 52876 8128 52916 8168
rect 62860 8128 62900 8168
rect 64108 8128 64148 8168
rect 65644 8128 65684 8168
rect 70732 8128 70772 8168
rect 71500 8128 71540 8168
rect 77068 8128 77108 8168
rect 4780 8044 4820 8084
rect 54028 8044 54068 8084
rect 55948 8044 55988 8084
rect 68332 8044 68372 8084
rect 73612 8044 73652 8084
rect 76300 8044 76340 8084
rect 1996 7960 2036 8000
rect 2092 7960 2132 8000
rect 2188 7960 2228 8000
rect 2284 7960 2324 8000
rect 2572 7960 2612 8000
rect 2764 7960 2804 8000
rect 2878 7960 2918 8000
rect 3340 7960 3380 8000
rect 3628 7960 3668 8000
rect 3724 7960 3764 8000
rect 4300 7960 4340 8000
rect 4492 7960 4532 8000
rect 4588 7960 4628 8000
rect 5164 7960 5204 8000
rect 6028 7960 6068 8000
rect 44140 7960 44180 8000
rect 44236 7960 44276 8000
rect 44428 7960 44468 8000
rect 44716 7960 44756 8000
rect 44812 7960 44852 8000
rect 45004 7960 45044 8000
rect 45388 7960 45428 8000
rect 45484 7960 45524 8000
rect 45580 7960 45620 8000
rect 45676 7960 45716 8000
rect 46732 7960 46772 8000
rect 46828 7960 46868 8000
rect 47020 7960 47060 8000
rect 47212 7960 47252 8000
rect 47308 7960 47348 8000
rect 47500 7960 47540 8000
rect 47980 7960 48020 8000
rect 48268 7960 48308 8000
rect 48364 7960 48404 8000
rect 48844 7973 48884 8013
rect 49036 7960 49076 8000
rect 49420 7960 49460 8000
rect 50476 7960 50516 8000
rect 50860 7960 50900 8000
rect 51724 7960 51764 8000
rect 53068 7960 53108 8000
rect 53164 7960 53204 8000
rect 53260 7981 53300 8021
rect 53356 7960 53396 8000
rect 53932 7960 53972 8000
rect 54124 7960 54164 8000
rect 54220 7960 54260 8000
rect 56332 7960 56372 8000
rect 57196 7960 57236 8000
rect 58540 7960 58580 8000
rect 58636 7960 58676 8000
rect 58828 7960 58868 8000
rect 60460 7960 60500 8000
rect 60844 7960 60884 8000
rect 61708 7960 61748 8000
rect 63628 7960 63668 8000
rect 63820 7960 63860 8000
rect 63916 7960 63956 8000
rect 64204 7960 64244 8000
rect 64300 7960 64340 8000
rect 64396 7960 64436 8000
rect 64684 7960 64724 8000
rect 64972 7960 65012 8000
rect 65068 7960 65108 8000
rect 65548 7960 65588 8000
rect 65740 7960 65780 8000
rect 65836 7960 65876 8000
rect 66028 7960 66068 8000
rect 66220 7960 66260 8000
rect 68716 7960 68756 8000
rect 69580 7960 69620 8000
rect 71404 7960 71444 8000
rect 71596 7960 71636 8000
rect 71692 7960 71732 8000
rect 73996 7960 74036 8000
rect 74860 7960 74900 8000
rect 76204 7960 76244 8000
rect 76396 7960 76436 8000
rect 76492 7960 76532 8000
rect 76972 7960 77012 8000
rect 77164 7960 77204 8000
rect 77260 7960 77300 8000
rect 77452 7960 77492 8000
rect 77548 7960 77588 8000
rect 77644 7960 77684 8000
rect 844 7876 884 7916
rect 1708 7876 1748 7916
rect 58348 7876 58388 7916
rect 59884 7876 59924 7916
rect 60268 7876 60308 7916
rect 1324 7792 1364 7832
rect 44428 7792 44468 7832
rect 45964 7792 46004 7832
rect 47020 7792 47060 7832
rect 48652 7792 48692 7832
rect 48940 7792 48980 7832
rect 63052 7792 63092 7832
rect 66124 7792 66164 7832
rect 66508 7792 66548 7832
rect 77836 7792 77876 7832
rect 1516 7708 1556 7748
rect 2572 7708 2612 7748
rect 4012 7708 4052 7748
rect 7180 7708 7220 7748
rect 47500 7708 47540 7748
rect 49612 7708 49652 7748
rect 58828 7708 58868 7748
rect 59692 7708 59732 7748
rect 60076 7708 60116 7748
rect 63628 7708 63668 7748
rect 65356 7708 65396 7748
rect 70732 7708 70772 7748
rect 76012 7708 76052 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 3724 7372 3764 7412
rect 4876 7372 4916 7412
rect 47788 7372 47828 7412
rect 51148 7372 51188 7412
rect 64588 7372 64628 7412
rect 65356 7372 65396 7412
rect 77452 7372 77492 7412
rect 652 7288 692 7328
rect 51916 7288 51956 7328
rect 55276 7288 55316 7328
rect 61036 7288 61076 7328
rect 69388 7288 69428 7328
rect 72364 7288 72404 7328
rect 77836 7288 77876 7328
rect 844 7204 884 7244
rect 54892 7204 54932 7244
rect 1708 7120 1748 7160
rect 2572 7120 2612 7160
rect 4012 7120 4052 7160
rect 4204 7120 4244 7160
rect 4780 7120 4820 7160
rect 4972 7120 5012 7160
rect 45388 7120 45428 7160
rect 45772 7120 45812 7160
rect 46636 7120 46676 7160
rect 48364 7120 48404 7160
rect 48748 7120 48788 7160
rect 49132 7120 49172 7160
rect 49996 7120 50036 7160
rect 52780 7120 52820 7160
rect 52972 7120 53012 7160
rect 53068 7120 53108 7160
rect 1324 7036 1364 7076
rect 4108 7036 4148 7076
rect 52876 7036 52916 7076
rect 53260 7078 53300 7118
rect 53452 7120 53492 7160
rect 53548 7120 53588 7160
rect 54220 7120 54260 7160
rect 54412 7120 54452 7160
rect 57292 7120 57332 7160
rect 58156 7120 58196 7160
rect 59692 7120 59732 7160
rect 59980 7120 60020 7160
rect 60556 7120 60596 7160
rect 60652 7120 60692 7160
rect 60844 7120 60884 7160
rect 62188 7120 62228 7160
rect 62572 7120 62612 7160
rect 63436 7120 63476 7160
rect 64780 7120 64820 7160
rect 64972 7120 65012 7160
rect 65068 7120 65108 7160
rect 65260 7120 65300 7160
rect 65452 7120 65492 7160
rect 66220 7120 66260 7160
rect 66412 7120 66452 7160
rect 66700 7120 66740 7160
rect 66892 7120 66932 7160
rect 69676 7120 69716 7160
rect 69772 7120 69812 7160
rect 69868 7120 69908 7160
rect 70060 7120 70100 7160
rect 70252 7120 70292 7160
rect 70348 7139 70388 7179
rect 71212 7120 71252 7160
rect 71404 7120 71444 7160
rect 71596 7120 71636 7160
rect 71788 7120 71828 7160
rect 71884 7120 71924 7160
rect 75436 7120 75476 7160
rect 75532 7120 75572 7160
rect 75628 7120 75668 7160
rect 75724 7120 75764 7160
rect 75916 7120 75956 7160
rect 76108 7120 76148 7160
rect 76204 7120 76244 7160
rect 76876 7120 76916 7160
rect 77068 7120 77108 7160
rect 77356 7120 77396 7160
rect 77548 7120 77588 7160
rect 53356 7036 53396 7076
rect 54316 7036 54356 7076
rect 56908 7036 56948 7076
rect 60076 7036 60116 7076
rect 64876 7036 64916 7076
rect 66316 7036 66356 7076
rect 66796 7036 66836 7076
rect 71308 7036 71348 7076
rect 76012 7036 76052 7076
rect 76972 7036 77012 7076
rect 55084 6952 55124 6992
rect 59308 6952 59348 6992
rect 60748 6952 60788 6992
rect 69580 6952 69620 6992
rect 70156 6952 70196 6992
rect 71692 6952 71732 6992
rect 60364 6910 60404 6950
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 47212 6616 47252 6656
rect 57004 6616 57044 6656
rect 69100 6616 69140 6656
rect 74284 6616 74324 6656
rect 2188 6448 2228 6488
rect 2380 6448 2420 6488
rect 2476 6448 2516 6488
rect 2668 6448 2708 6488
rect 2860 6490 2900 6530
rect 54220 6532 54260 6572
rect 54604 6532 54644 6572
rect 58540 6532 58580 6572
rect 66124 6532 66164 6572
rect 71884 6532 71924 6572
rect 2956 6448 2996 6488
rect 4108 6448 4148 6488
rect 4204 6448 4244 6488
rect 4492 6448 4532 6488
rect 4876 6448 4916 6488
rect 5068 6448 5108 6488
rect 47308 6448 47348 6488
rect 47404 6448 47444 6488
rect 47500 6448 47540 6488
rect 47692 6448 47732 6488
rect 47884 6448 47924 6488
rect 47980 6448 48020 6488
rect 48844 6448 48884 6488
rect 49228 6448 49268 6488
rect 50092 6448 50132 6488
rect 51436 6448 51476 6488
rect 51820 6448 51860 6488
rect 52684 6448 52724 6488
rect 54124 6448 54164 6488
rect 54316 6448 54356 6488
rect 54412 6448 54452 6488
rect 54988 6448 55028 6488
rect 55852 6448 55892 6488
rect 58060 6448 58100 6488
rect 58252 6448 58292 6488
rect 58348 6448 58388 6488
rect 58636 6448 58676 6488
rect 58732 6448 58772 6488
rect 58828 6448 58868 6488
rect 59212 6448 59252 6488
rect 59308 6448 59348 6488
rect 59500 6448 59540 6488
rect 60172 6448 60212 6488
rect 60364 6448 60404 6488
rect 61420 6448 61460 6488
rect 61612 6448 61652 6488
rect 65740 6448 65780 6488
rect 66028 6448 66068 6488
rect 66700 6448 66740 6488
rect 67084 6448 67124 6488
rect 67948 6448 67988 6488
rect 69292 6448 69332 6488
rect 69676 6448 69716 6488
rect 70540 6448 70580 6488
rect 72268 6448 72308 6488
rect 73132 6448 73172 6488
rect 75628 6448 75668 6488
rect 75724 6448 75764 6488
rect 75820 6448 75860 6488
rect 75916 6411 75956 6451
rect 76204 6448 76244 6488
rect 76492 6448 76532 6488
rect 76588 6448 76628 6488
rect 77068 6448 77108 6488
rect 77452 6448 77492 6488
rect 78316 6448 78356 6488
rect 844 6364 884 6404
rect 652 6280 692 6320
rect 1708 6280 1748 6320
rect 2188 6280 2228 6320
rect 2668 6280 2708 6320
rect 5452 6280 5492 6320
rect 57388 6280 57428 6320
rect 58060 6280 58100 6320
rect 60268 6280 60308 6320
rect 63628 6280 63668 6320
rect 66412 6280 66452 6320
rect 74476 6280 74516 6320
rect 76876 6280 76916 6320
rect 3820 6196 3860 6236
rect 4972 6196 5012 6236
rect 47692 6196 47732 6236
rect 51244 6196 51284 6236
rect 53836 6196 53876 6236
rect 57004 6196 57044 6236
rect 59500 6196 59540 6236
rect 61516 6196 61556 6236
rect 71692 6196 71732 6236
rect 74284 6196 74324 6236
rect 79468 6196 79508 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 7372 5860 7412 5900
rect 49036 5860 49076 5900
rect 54508 5860 54548 5900
rect 66412 5860 66452 5900
rect 69772 5860 69812 5900
rect 71116 5860 71156 5900
rect 76012 5860 76052 5900
rect 77068 5860 77108 5900
rect 46348 5776 46388 5816
rect 48844 5776 48884 5816
rect 49516 5776 49556 5816
rect 56620 5776 56660 5816
rect 59692 5776 59732 5816
rect 67180 5776 67220 5816
rect 1036 5692 1076 5732
rect 3628 5692 3668 5732
rect 54796 5692 54836 5732
rect 63724 5692 63764 5732
rect 72172 5692 72212 5732
rect 1612 5608 1652 5648
rect 2476 5608 2516 5648
rect 4108 5608 4148 5648
rect 5356 5608 5396 5648
rect 6220 5608 6260 5648
rect 47212 5608 47252 5648
rect 47404 5608 47444 5648
rect 47500 5608 47540 5648
rect 48172 5608 48212 5648
rect 48460 5608 48500 5648
rect 49036 5608 49076 5648
rect 49228 5608 49268 5648
rect 49324 5608 49364 5648
rect 49900 5608 49940 5648
rect 50092 5608 50132 5648
rect 52300 5608 52340 5648
rect 52396 5608 52436 5648
rect 52588 5608 52628 5648
rect 52780 5608 52820 5648
rect 52876 5608 52916 5648
rect 52972 5608 53012 5648
rect 53068 5608 53108 5648
rect 53836 5608 53876 5648
rect 54124 5608 54164 5648
rect 54220 5608 54260 5648
rect 54700 5608 54740 5648
rect 54892 5608 54932 5648
rect 56236 5608 56276 5648
rect 56428 5608 56468 5648
rect 59212 5608 59252 5648
rect 59404 5608 59444 5648
rect 59500 5608 59540 5648
rect 60844 5608 60884 5648
rect 61036 5608 61076 5648
rect 61132 5608 61172 5648
rect 61708 5608 61748 5648
rect 62572 5608 62612 5648
rect 64588 5608 64628 5648
rect 64780 5608 64820 5648
rect 64876 5608 64916 5648
rect 65068 5608 65108 5648
rect 65164 5608 65204 5648
rect 65260 5608 65300 5648
rect 65356 5608 65396 5648
rect 66412 5608 66452 5648
rect 66604 5608 66644 5648
rect 66700 5608 66740 5648
rect 69292 5608 69332 5648
rect 69388 5608 69428 5648
rect 69484 5608 69524 5648
rect 69580 5608 69620 5648
rect 69772 5608 69812 5648
rect 69964 5608 70004 5648
rect 70060 5608 70100 5648
rect 71404 5608 71444 5648
rect 71500 5608 71540 5648
rect 71788 5608 71828 5648
rect 72076 5608 72116 5648
rect 72268 5608 72308 5648
rect 73996 5608 74036 5648
rect 74860 5608 74900 5648
rect 76204 5608 76244 5648
rect 76396 5608 76436 5648
rect 76492 5608 76532 5648
rect 77068 5608 77108 5648
rect 77260 5608 77300 5648
rect 77356 5608 77396 5648
rect 77548 5608 77588 5648
rect 77740 5608 77780 5648
rect 1228 5524 1268 5564
rect 4972 5524 5012 5564
rect 48556 5524 48596 5564
rect 49996 5524 50036 5564
rect 52492 5524 52532 5564
rect 56332 5524 56372 5564
rect 61324 5524 61364 5564
rect 73612 5524 73652 5564
rect 76300 5524 76340 5564
rect 77644 5524 77684 5564
rect 844 5440 884 5480
rect 7372 5440 7412 5480
rect 47308 5440 47348 5480
rect 59308 5440 59348 5480
rect 60940 5440 60980 5480
rect 64684 5440 64724 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 652 5104 692 5144
rect 2284 5104 2324 5144
rect 52204 5104 52244 5144
rect 55756 5104 55796 5144
rect 65548 5104 65588 5144
rect 65836 5104 65876 5144
rect 71692 5104 71732 5144
rect 76108 5104 76148 5144
rect 1996 5020 2036 5060
rect 1708 4936 1748 4976
rect 1804 4936 1844 4976
rect 1900 4936 1940 4976
rect 2188 4978 2228 5018
rect 45868 5020 45908 5060
rect 56140 5020 56180 5060
rect 58924 5020 58964 5060
rect 62284 5020 62324 5060
rect 63148 5020 63188 5060
rect 66316 5020 66356 5060
rect 2380 4936 2420 4976
rect 2476 4936 2516 4976
rect 3724 4936 3764 4976
rect 3916 4936 3956 4976
rect 4108 4936 4148 4976
rect 5068 4936 5108 4976
rect 46252 4936 46292 4976
rect 47116 4936 47156 4976
rect 48460 4936 48500 4976
rect 48652 4936 48692 4976
rect 48844 4936 48884 4976
rect 48940 4936 48980 4976
rect 49132 4936 49172 4976
rect 51532 4936 51572 4976
rect 51628 4936 51668 4976
rect 51820 4936 51860 4976
rect 52012 4936 52052 4976
rect 52108 4936 52148 4976
rect 52300 4936 52340 4976
rect 52492 4936 52532 4976
rect 52684 4936 52724 4976
rect 55660 4936 55700 4976
rect 55852 4936 55892 4976
rect 55948 4936 55988 4976
rect 56524 4936 56564 4976
rect 57388 4936 57428 4976
rect 59308 4936 59348 4976
rect 60172 4936 60212 4976
rect 62188 4936 62228 4976
rect 62380 4936 62420 4976
rect 63532 4936 63572 4976
rect 64396 4936 64436 4976
rect 65740 4936 65780 4976
rect 65932 4936 65972 4976
rect 66028 4936 66068 4976
rect 66220 4936 66260 4976
rect 66412 4936 66452 4976
rect 68908 4936 68948 4976
rect 69100 4936 69140 4976
rect 69196 4936 69236 4976
rect 71596 4936 71636 4976
rect 71788 4936 71828 4976
rect 71884 4936 71924 4976
rect 72076 4936 72116 4976
rect 72172 4936 72212 4976
rect 72268 4936 72308 4976
rect 75916 4936 75956 4976
rect 76012 4936 76052 4976
rect 76204 4936 76244 4976
rect 76963 4949 77003 4989
rect 77164 4936 77204 4976
rect 77452 4936 77492 4976
rect 77644 4949 77684 4989
rect 844 4852 884 4892
rect 1516 4852 1556 4892
rect 3820 4768 3860 4808
rect 5548 4768 5588 4808
rect 48556 4768 48596 4808
rect 50188 4768 50228 4808
rect 52876 4768 52916 4808
rect 58540 4768 58580 4808
rect 61804 4768 61844 4808
rect 66892 4768 66932 4808
rect 69388 4768 69428 4808
rect 72460 4768 72500 4808
rect 74284 4768 74324 4808
rect 77836 4768 77876 4808
rect 1324 4684 1364 4724
rect 48268 4684 48308 4724
rect 49132 4684 49172 4724
rect 51820 4684 51860 4724
rect 52588 4684 52628 4724
rect 61324 4684 61364 4724
rect 68908 4684 68948 4724
rect 77068 4684 77108 4724
rect 77548 4684 77588 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 2572 4348 2612 4388
rect 52012 4348 52052 4388
rect 61516 4348 61556 4388
rect 66220 4348 66260 4388
rect 76876 4348 76916 4388
rect 652 4264 692 4304
rect 1900 4264 1940 4304
rect 4204 4264 4244 4304
rect 7468 4264 7508 4304
rect 55180 4264 55220 4304
rect 56908 4264 56948 4304
rect 57964 4264 58004 4304
rect 60172 4264 60212 4304
rect 68812 4264 68852 4304
rect 74380 4264 74420 4304
rect 844 4180 884 4220
rect 1228 4180 1268 4220
rect 79468 4180 79508 4220
rect 2092 4096 2132 4136
rect 2188 4096 2228 4136
rect 2284 4096 2324 4136
rect 2572 4096 2612 4136
rect 2764 4096 2804 4136
rect 2878 4096 2918 4136
rect 3532 4096 3572 4136
rect 3820 4096 3860 4136
rect 4588 4096 4628 4136
rect 4780 4096 4820 4136
rect 4876 4096 4916 4136
rect 5452 4096 5492 4136
rect 6316 4096 6356 4136
rect 47404 4096 47444 4136
rect 47500 4096 47540 4136
rect 47596 4096 47636 4136
rect 47692 4096 47732 4136
rect 49996 4096 50036 4136
rect 50860 4096 50900 4136
rect 52396 4096 52436 4136
rect 52780 4096 52820 4136
rect 53644 4096 53684 4136
rect 55660 4096 55700 4136
rect 55756 4096 55796 4136
rect 55852 4096 55892 4136
rect 55948 4096 55988 4136
rect 56236 4096 56276 4136
rect 56524 4096 56564 4136
rect 57100 4096 57140 4136
rect 57292 4096 57332 4136
rect 57388 4096 57428 4136
rect 57964 4096 58004 4136
rect 58156 4096 58196 4136
rect 58252 4096 58292 4136
rect 59020 4096 59060 4136
rect 59116 4096 59156 4136
rect 59212 4096 59252 4136
rect 59308 4096 59348 4136
rect 60844 4096 60884 4136
rect 61132 4096 61172 4136
rect 61228 4096 61268 4136
rect 63244 4096 63284 4136
rect 64108 4096 64148 4136
rect 65548 4096 65588 4136
rect 65836 4096 65876 4136
rect 66796 4096 66836 4136
rect 67660 4096 67700 4136
rect 69388 4096 69428 4136
rect 70252 4096 70292 4136
rect 71596 4096 71636 4136
rect 71788 4096 71828 4136
rect 71980 4096 72020 4136
rect 72364 4096 72404 4136
rect 73228 4096 73268 4136
rect 75148 4096 75188 4136
rect 75340 4096 75380 4136
rect 75436 4096 75476 4136
rect 75628 4096 75668 4136
rect 75724 4096 75764 4136
rect 75820 4096 75860 4136
rect 75916 4096 75956 4136
rect 76204 4096 76244 4136
rect 76492 4096 76532 4136
rect 76588 4096 76628 4136
rect 77452 4096 77492 4136
rect 78316 4096 78356 4136
rect 3916 4012 3956 4052
rect 5068 4012 5108 4052
rect 49612 4012 49652 4052
rect 56620 4012 56660 4052
rect 62860 4012 62900 4052
rect 65932 4012 65972 4052
rect 66412 4012 66452 4052
rect 69004 4012 69044 4052
rect 71692 4012 71732 4052
rect 77068 4012 77108 4052
rect 1036 3928 1076 3968
rect 2380 3928 2420 3968
rect 4684 3928 4724 3968
rect 52012 3928 52052 3968
rect 54796 3928 54836 3968
rect 57196 3928 57236 3968
rect 65260 3928 65300 3968
rect 71404 3928 71444 3968
rect 75244 3928 75284 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 3820 3592 3860 3632
rect 4684 3592 4724 3632
rect 50284 3592 50324 3632
rect 53932 3592 53972 3632
rect 62092 3592 62132 3632
rect 64012 3592 64052 3632
rect 66220 3592 66260 3632
rect 69388 3592 69428 3632
rect 76204 3592 76244 3632
rect 76492 3592 76532 3632
rect 77260 3592 77300 3632
rect 52108 3508 52148 3548
rect 52684 3508 52724 3548
rect 56332 3508 56372 3548
rect 56812 3508 56852 3548
rect 73804 3508 73844 3548
rect 1420 3424 1460 3464
rect 1804 3424 1844 3464
rect 2668 3424 2708 3464
rect 4204 3424 4244 3464
rect 4396 3424 4436 3464
rect 4588 3413 4628 3453
rect 4780 3424 4820 3464
rect 4876 3424 4916 3464
rect 5068 3424 5108 3464
rect 5260 3424 5300 3464
rect 50092 3424 50132 3464
rect 50188 3424 50228 3464
rect 50380 3424 50420 3464
rect 50668 3424 50708 3464
rect 50764 3424 50804 3464
rect 50860 3424 50900 3464
rect 50956 3424 50996 3464
rect 51724 3424 51764 3464
rect 52012 3424 52052 3464
rect 52588 3424 52628 3464
rect 52780 3424 52820 3464
rect 55084 3424 55124 3464
rect 55948 3424 55988 3464
rect 56716 3424 56756 3464
rect 56908 3424 56948 3464
rect 59308 3424 59348 3464
rect 59500 3424 59540 3464
rect 59692 3424 59732 3464
rect 60076 3424 60116 3464
rect 60940 3424 60980 3464
rect 63820 3424 63860 3464
rect 63916 3424 63956 3464
rect 64108 3424 64148 3464
rect 64300 3424 64340 3464
rect 64396 3424 64436 3464
rect 64492 3424 64532 3464
rect 64588 3424 64628 3464
rect 66124 3424 66164 3464
rect 66316 3424 66356 3464
rect 66412 3424 66452 3464
rect 66604 3424 66644 3464
rect 66796 3424 66836 3464
rect 68620 3424 68660 3464
rect 68716 3424 68756 3464
rect 68908 3424 68948 3464
rect 69196 3424 69236 3464
rect 69292 3424 69332 3464
rect 69484 3424 69524 3464
rect 69772 3424 69812 3464
rect 69868 3424 69908 3464
rect 69964 3424 70004 3464
rect 70060 3424 70100 3464
rect 71212 3424 71252 3464
rect 71500 3424 71540 3464
rect 71596 3424 71636 3464
rect 72076 3424 72116 3464
rect 72172 3424 72212 3464
rect 72364 3424 72404 3464
rect 74188 3424 74228 3464
rect 75052 3424 75092 3464
rect 76396 3424 76436 3464
rect 76588 3424 76628 3464
rect 76684 3424 76724 3464
rect 77164 3424 77204 3464
rect 77356 3424 77396 3464
rect 77452 3424 77492 3464
rect 844 3340 884 3380
rect 1228 3340 1268 3380
rect 1036 3256 1076 3296
rect 63340 3298 63380 3338
rect 5164 3256 5204 3296
rect 52396 3256 52436 3296
rect 66700 3256 66740 3296
rect 68908 3256 68948 3296
rect 71884 3256 71924 3296
rect 652 3172 692 3212
rect 4300 3172 4340 3212
rect 59404 3172 59444 3212
rect 72364 3172 72404 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 59116 2836 59156 2876
rect 64012 2836 64052 2876
rect 73516 2836 73556 2876
rect 1516 2752 1556 2792
rect 54028 2752 54068 2792
rect 56812 2752 56852 2792
rect 57100 2752 57140 2792
rect 60076 2752 60116 2792
rect 62188 2752 62228 2792
rect 66508 2752 66548 2792
rect 68716 2752 68756 2792
rect 71500 2752 71540 2792
rect 72940 2752 72980 2792
rect 74956 2752 74996 2792
rect 76108 2752 76148 2792
rect 77452 2752 77492 2792
rect 78220 2752 78260 2792
rect 844 2668 884 2708
rect 1708 2668 1748 2708
rect 64780 2668 64820 2708
rect 2380 2584 2420 2624
rect 2572 2584 2612 2624
rect 2668 2584 2708 2624
rect 2860 2584 2900 2624
rect 3052 2584 3092 2624
rect 3148 2584 3188 2624
rect 55372 2584 55412 2624
rect 55468 2584 55508 2624
rect 55564 2584 55604 2624
rect 55756 2584 55796 2624
rect 55948 2584 55988 2624
rect 56044 2584 56084 2624
rect 56236 2584 56276 2624
rect 56428 2584 56468 2624
rect 56524 2584 56564 2624
rect 56716 2584 56756 2624
rect 56908 2584 56948 2624
rect 58828 2584 58868 2624
rect 58924 2584 58964 2624
rect 59116 2584 59156 2624
rect 59404 2584 59444 2624
rect 59692 2584 59732 2624
rect 60268 2584 60308 2624
rect 60364 2584 60404 2624
rect 60460 2584 60500 2624
rect 63724 2584 63764 2624
rect 63820 2584 63860 2624
rect 64012 2584 64052 2624
rect 64204 2584 64244 2624
rect 64396 2584 64436 2624
rect 64492 2584 64532 2624
rect 64684 2584 64724 2624
rect 64876 2584 64916 2624
rect 68236 2584 68276 2624
rect 68332 2584 68372 2624
rect 68428 2584 68468 2624
rect 68620 2584 68660 2624
rect 68812 2584 68852 2624
rect 69004 2584 69044 2624
rect 69196 2584 69236 2624
rect 71788 2584 71828 2624
rect 71884 2584 71924 2624
rect 71980 2584 72020 2624
rect 72268 2584 72308 2624
rect 72556 2584 72596 2624
rect 72652 2584 72692 2624
rect 73228 2584 73268 2624
rect 74188 2584 74228 2624
rect 74380 2584 74420 2624
rect 74572 2584 74612 2624
rect 75148 2584 75188 2624
rect 75340 2584 75380 2624
rect 76780 2584 76820 2624
rect 77068 2584 77108 2624
rect 77644 2584 77684 2624
rect 77836 2584 77876 2624
rect 2476 2500 2516 2540
rect 59788 2500 59828 2540
rect 69100 2500 69140 2540
rect 74476 2500 74516 2540
rect 75244 2500 75284 2540
rect 77164 2500 77204 2540
rect 77740 2500 77780 2540
rect 652 2416 692 2456
rect 2956 2416 2996 2456
rect 55276 2416 55316 2456
rect 55852 2416 55892 2456
rect 56332 2416 56372 2456
rect 64300 2416 64340 2456
rect 68140 2416 68180 2456
rect 71692 2416 71732 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 55948 2080 55988 2120
rect 58924 2080 58964 2120
rect 61516 2080 61556 2120
rect 64108 2080 64148 2120
rect 66892 2080 66932 2120
rect 71212 2080 71252 2120
rect 73804 2080 73844 2120
rect 78028 2080 78068 2120
rect 56524 1996 56564 2036
rect 53548 1912 53588 1952
rect 53932 1912 53972 1952
rect 54796 1912 54836 1952
rect 56140 1912 56180 1952
rect 56332 1912 56372 1952
rect 56908 1912 56948 1952
rect 57772 1912 57812 1952
rect 59116 1912 59156 1952
rect 59500 1912 59540 1952
rect 60364 1912 60404 1952
rect 61708 1912 61748 1952
rect 62092 1912 62132 1952
rect 62956 1912 62996 1952
rect 64492 1912 64532 1952
rect 64876 1912 64916 1952
rect 65740 1912 65780 1952
rect 67372 1912 67412 1952
rect 67564 1912 67604 1952
rect 67660 1912 67700 1952
rect 67948 1912 67988 1952
rect 68236 1912 68276 1952
rect 68332 1912 68372 1952
rect 68812 1912 68852 1952
rect 69196 1912 69236 1952
rect 70060 1912 70100 1952
rect 71404 1912 71444 1952
rect 71788 1912 71828 1952
rect 72652 1912 72692 1952
rect 73996 1912 74036 1952
rect 74188 1912 74228 1952
rect 74284 1912 74324 1952
rect 74572 1912 74612 1952
rect 74668 1912 74708 1952
rect 74860 1912 74900 1952
rect 75148 1912 75188 1952
rect 75244 1912 75284 1952
rect 75436 1912 75476 1952
rect 75628 1912 75668 1952
rect 76012 1912 76052 1952
rect 76876 1912 76916 1952
rect 78220 1912 78260 1952
rect 78412 1912 78452 1952
rect 78508 1912 78548 1952
rect 78700 1912 78740 1952
rect 78892 1912 78932 1952
rect 68620 1744 68660 1784
rect 74860 1744 74900 1784
rect 75436 1744 75476 1784
rect 78796 1744 78836 1784
rect 55948 1660 55988 1700
rect 56236 1660 56276 1700
rect 58924 1660 58964 1700
rect 61516 1660 61556 1700
rect 64108 1660 64148 1700
rect 67372 1660 67412 1700
rect 73996 1660 74036 1700
rect 78220 1660 78260 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 55372 1324 55412 1364
rect 55948 1324 55988 1364
rect 59020 1324 59060 1364
rect 62572 1324 62612 1364
rect 68428 1324 68468 1364
rect 68908 1324 68948 1364
rect 70444 1324 70484 1364
rect 72460 1324 72500 1364
rect 77068 1324 77108 1364
rect 57484 1240 57524 1280
rect 60748 1240 60788 1280
rect 61996 1240 62036 1280
rect 64396 1240 64436 1280
rect 64684 1240 64724 1280
rect 64972 1240 65012 1280
rect 69292 1240 69332 1280
rect 60460 1156 60500 1196
rect 55372 1072 55412 1112
rect 55564 1072 55604 1112
rect 55660 1072 55700 1112
rect 56236 1072 56276 1112
rect 56332 1072 56372 1112
rect 56620 1072 56660 1112
rect 57196 1072 57236 1112
rect 57292 1072 57332 1112
rect 57484 1072 57524 1112
rect 58636 1072 58676 1112
rect 58732 1072 58772 1112
rect 58828 1072 58868 1112
rect 59020 1072 59060 1112
rect 59212 1072 59252 1112
rect 59308 1072 59348 1112
rect 59596 1072 59636 1112
rect 61708 1072 61748 1112
rect 61804 1072 61844 1112
rect 61996 1072 62036 1112
rect 62284 1072 62324 1112
rect 62380 1072 62420 1112
rect 62572 1072 62612 1112
rect 62764 1072 62804 1112
rect 62860 1072 62900 1112
rect 62956 1072 62996 1112
rect 63052 1072 63092 1112
rect 63724 1072 63764 1112
rect 64012 1072 64052 1112
rect 64108 1072 64148 1112
rect 64588 1072 64628 1112
rect 64780 1072 64820 1112
rect 66028 1072 66068 1112
rect 66412 1072 66452 1112
rect 67276 1072 67316 1112
rect 68620 1072 68660 1112
rect 68716 1072 68756 1112
rect 68908 1072 68948 1112
rect 69772 1072 69812 1112
rect 70924 1072 70964 1112
rect 71212 1072 71252 1112
rect 72076 1072 72116 1112
rect 72460 1072 72500 1112
rect 72652 1072 72692 1112
rect 72748 1072 72788 1112
rect 74380 1072 74420 1112
rect 75244 1072 75284 1112
rect 75628 1072 75668 1112
rect 75916 1072 75956 1112
rect 76012 1072 76052 1112
rect 76108 1072 76148 1112
rect 76204 1072 76244 1112
rect 78220 1072 78260 1112
rect 79084 1072 79124 1112
rect 79468 1072 79508 1112
rect 58540 904 58580 944
rect 73228 904 73268 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 63436 38324 63476 38333
rect 63340 38229 63380 38238
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 58348 38156 58388 38165
rect 56907 38072 56949 38081
rect 56907 38032 56908 38072
rect 56948 38032 56949 38072
rect 56907 38023 56949 38032
rect 58251 38072 58293 38081
rect 58251 38032 58252 38072
rect 58292 38032 58293 38072
rect 58251 38023 58293 38032
rect 844 37988 884 37997
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 844 37460 884 37948
rect 56908 37938 56948 38023
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 55180 37568 55220 37577
rect 844 37420 980 37460
rect 652 26060 692 26069
rect 652 25817 692 26020
rect 843 25976 885 25985
rect 843 25936 844 25976
rect 884 25936 885 25976
rect 843 25927 885 25936
rect 844 25842 884 25927
rect 651 25808 693 25817
rect 651 25768 652 25808
rect 692 25768 693 25808
rect 651 25759 693 25768
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 844 25002 884 25087
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 844 24380 884 24389
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 844 23885 884 24340
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 843 23876 885 23885
rect 843 23836 844 23876
rect 884 23836 885 23876
rect 843 23827 885 23836
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 844 23490 884 23575
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 23036 692 23045
rect 556 22996 652 23036
rect 556 22457 596 22996
rect 652 22987 692 22996
rect 844 22868 884 22877
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 844 20777 884 22828
rect 940 20861 980 37420
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 54699 36812 54741 36821
rect 54699 36772 54700 36812
rect 54740 36772 54741 36812
rect 54699 36763 54741 36772
rect 54700 36678 54740 36763
rect 55084 36728 55124 36737
rect 55180 36728 55220 37528
rect 55659 37400 55701 37409
rect 55659 37360 55660 37400
rect 55700 37360 55701 37400
rect 55659 37351 55701 37360
rect 55756 37400 55796 37409
rect 55124 36688 55220 36728
rect 55084 36679 55124 36688
rect 52492 36560 52532 36569
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 49227 36056 49269 36065
rect 49227 36016 49228 36056
rect 49268 36016 49269 36056
rect 49227 36007 49269 36016
rect 50571 36056 50613 36065
rect 50571 36016 50572 36056
rect 50612 36016 50613 36056
rect 50571 36007 50613 36016
rect 49228 35922 49268 36007
rect 50379 35972 50421 35981
rect 50379 35932 50380 35972
rect 50420 35932 50421 35972
rect 50379 35923 50421 35932
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 49707 35216 49749 35225
rect 49612 35176 49708 35216
rect 49748 35176 49749 35216
rect 47116 35048 47156 35057
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 46155 34544 46197 34553
rect 46155 34504 46156 34544
rect 46196 34504 46197 34544
rect 46155 34495 46197 34504
rect 46444 34544 46484 34553
rect 46484 34504 46676 34544
rect 46444 34495 46484 34504
rect 46156 34376 46196 34495
rect 46156 34327 46196 34336
rect 46252 34376 46292 34385
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 43852 33032 43892 33041
rect 42219 32948 42261 32957
rect 42219 32908 42220 32948
rect 42260 32908 42261 32948
rect 42219 32899 42261 32908
rect 42699 32948 42741 32957
rect 42699 32908 42700 32948
rect 42740 32908 42741 32948
rect 42699 32899 42741 32908
rect 42123 32696 42165 32705
rect 42123 32656 42124 32696
rect 42164 32656 42165 32696
rect 42123 32647 42165 32656
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 40684 32024 40724 32033
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 40588 31352 40628 31361
rect 40684 31352 40724 31984
rect 40628 31312 40724 31352
rect 41451 31352 41493 31361
rect 41451 31312 41452 31352
rect 41492 31312 41493 31352
rect 40588 31303 40628 31312
rect 41451 31303 41493 31312
rect 40204 31268 40244 31277
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 40204 30857 40244 31228
rect 41452 31218 41492 31303
rect 41067 31100 41109 31109
rect 41067 31060 41068 31100
rect 41108 31060 41109 31100
rect 41067 31051 41109 31060
rect 40203 30848 40245 30857
rect 40203 30808 40204 30848
rect 40244 30808 40245 30848
rect 40203 30799 40245 30808
rect 40203 30680 40245 30689
rect 40203 30640 40204 30680
rect 40244 30640 40245 30680
rect 40203 30631 40245 30640
rect 40204 30269 40244 30631
rect 40875 30596 40917 30605
rect 40875 30556 40876 30596
rect 40916 30556 40917 30596
rect 40875 30547 40917 30556
rect 40876 30462 40916 30547
rect 40684 30428 40724 30437
rect 40396 30388 40684 30428
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 39723 30260 39765 30269
rect 39723 30220 39724 30260
rect 39764 30220 39765 30260
rect 39723 30211 39765 30220
rect 40203 30260 40245 30269
rect 40203 30220 40204 30260
rect 40244 30220 40245 30260
rect 40203 30211 40245 30220
rect 38860 30008 38900 30017
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 38380 29168 38420 29177
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 38188 28496 38228 28505
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 37707 27740 37749 27749
rect 37707 27700 37708 27740
rect 37748 27700 37749 27740
rect 37707 27691 37749 27700
rect 37708 27606 37748 27691
rect 38092 27656 38132 27665
rect 38188 27656 38228 28456
rect 38380 28253 38420 29128
rect 38764 29168 38804 29177
rect 38860 29168 38900 29968
rect 39628 29168 39668 29177
rect 38804 29128 38900 29168
rect 38956 29128 39628 29168
rect 38764 29119 38804 29128
rect 38379 28244 38421 28253
rect 38379 28204 38380 28244
rect 38420 28204 38421 28244
rect 38379 28195 38421 28204
rect 38667 27908 38709 27917
rect 38667 27868 38668 27908
rect 38708 27868 38709 27908
rect 38667 27859 38709 27868
rect 38132 27616 38228 27656
rect 38092 27607 38132 27616
rect 36460 27488 36500 27497
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 33003 26984 33045 26993
rect 33003 26944 33004 26984
rect 33044 26944 33045 26984
rect 33003 26935 33045 26944
rect 34251 26984 34293 26993
rect 35308 26984 35348 26993
rect 34251 26944 34252 26984
rect 34292 26944 34293 26984
rect 34251 26935 34293 26944
rect 35116 26944 35308 26984
rect 33004 26850 33044 26935
rect 4300 26816 4340 26825
rect 4340 26776 4820 26816
rect 4300 26767 4340 26776
rect 4204 26648 4244 26657
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3915 25136 3957 25145
rect 3915 25096 3916 25136
rect 3956 25096 3957 25136
rect 3915 25087 3957 25096
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 1804 23876 1844 23885
rect 1804 23633 1844 23836
rect 1995 23876 2037 23885
rect 1995 23836 1996 23876
rect 2036 23836 2037 23876
rect 1995 23827 2037 23836
rect 1996 23742 2036 23827
rect 1419 23624 1461 23633
rect 1419 23584 1420 23624
rect 1460 23584 1461 23624
rect 1419 23575 1461 23584
rect 1612 23624 1652 23633
rect 1420 23129 1460 23575
rect 1515 23204 1557 23213
rect 1612 23204 1652 23584
rect 1803 23624 1845 23633
rect 1803 23584 1804 23624
rect 1844 23584 1845 23624
rect 1803 23575 1845 23584
rect 2187 23624 2229 23633
rect 2187 23584 2188 23624
rect 2228 23584 2229 23624
rect 2187 23575 2229 23584
rect 2188 23490 2228 23575
rect 1515 23164 1516 23204
rect 1556 23164 1652 23204
rect 1515 23155 1557 23164
rect 1419 23120 1461 23129
rect 1419 23080 1420 23120
rect 1460 23080 1461 23120
rect 1419 23071 1461 23080
rect 1516 23120 1556 23155
rect 1420 22952 1460 23071
rect 1516 23069 1556 23080
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 1941 23120
rect 1899 23071 1941 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 1900 22986 1940 23071
rect 2092 22986 2132 23071
rect 1516 22952 1556 22961
rect 1420 22912 1516 22952
rect 1516 22903 1556 22912
rect 1707 22868 1749 22877
rect 1707 22828 1708 22868
rect 1748 22828 1749 22868
rect 1707 22819 1749 22828
rect 1900 22868 1940 22877
rect 1708 22734 1748 22819
rect 1900 21533 1940 22828
rect 2763 22868 2805 22877
rect 2763 22828 2764 22868
rect 2804 22828 2805 22868
rect 2763 22819 2805 22828
rect 1899 21524 1941 21533
rect 1899 21484 1900 21524
rect 1940 21484 1941 21524
rect 1899 21475 1941 21484
rect 939 20852 981 20861
rect 939 20812 940 20852
rect 980 20812 981 20852
rect 939 20803 981 20812
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 843 20768 885 20777
rect 843 20728 844 20768
rect 884 20728 885 20768
rect 843 20719 885 20728
rect 2667 20096 2709 20105
rect 2667 20056 2668 20096
rect 2708 20056 2709 20096
rect 2667 20047 2709 20056
rect 1995 20012 2037 20021
rect 1995 19972 1996 20012
rect 2036 19972 2037 20012
rect 1995 19963 2037 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 1707 18500 1749 18509
rect 1707 18460 1708 18500
rect 1748 18460 1749 18500
rect 1707 18451 1749 18460
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 1708 18366 1748 18451
rect 1516 18332 1556 18341
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 1516 17300 1556 18292
rect 1516 17260 1652 17300
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 652 15737 692 16360
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 844 15476 884 15485
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 844 14981 884 15436
rect 1132 15308 1172 15317
rect 1172 15268 1364 15308
rect 1132 15259 1172 15268
rect 843 14972 885 14981
rect 843 14932 844 14972
rect 884 14932 885 14972
rect 843 14923 885 14932
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 844 14804 884 14813
rect 1324 14804 1364 15268
rect 1515 14972 1557 14981
rect 1515 14932 1516 14972
rect 1556 14932 1557 14972
rect 1515 14923 1557 14932
rect 1516 14838 1556 14923
rect 884 14764 1268 14804
rect 844 14755 884 14764
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 1132 14552 1172 14561
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 1036 13376 1076 13385
rect 844 13336 1036 13376
rect 844 13292 884 13336
rect 1036 13327 1076 13336
rect 844 13243 884 13252
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 1132 12980 1172 14512
rect 1228 14216 1268 14764
rect 1324 14729 1364 14764
rect 1323 14720 1365 14729
rect 1323 14680 1324 14720
rect 1364 14680 1365 14720
rect 1323 14671 1365 14680
rect 1324 14640 1364 14671
rect 1324 14216 1364 14225
rect 1228 14176 1324 14216
rect 1324 14167 1364 14176
rect 1515 14216 1557 14225
rect 1515 14176 1516 14216
rect 1556 14176 1557 14216
rect 1515 14167 1557 14176
rect 1516 13964 1556 14167
rect 1516 13915 1556 13924
rect 1227 13292 1269 13301
rect 1227 13252 1228 13292
rect 1268 13252 1269 13292
rect 1227 13243 1269 13252
rect 1228 13158 1268 13243
rect 1420 13124 1460 13133
rect 1132 12940 1268 12980
rect 844 12452 884 12461
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 844 12368 884 12412
rect 1132 12368 1172 12377
rect 844 12328 1132 12368
rect 651 12319 693 12328
rect 1132 12319 1172 12328
rect 555 12284 597 12293
rect 555 12244 556 12284
rect 596 12244 597 12284
rect 555 12235 597 12244
rect 556 7253 596 12235
rect 652 12234 692 12319
rect 1131 11780 1173 11789
rect 1131 11740 1132 11780
rect 1172 11740 1173 11780
rect 1131 11731 1173 11740
rect 1132 11646 1172 11731
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 940 11528 980 11537
rect 1228 11528 1268 12940
rect 1420 12713 1460 13084
rect 1419 12704 1461 12713
rect 1419 12664 1420 12704
rect 1460 12664 1461 12704
rect 1419 12655 1461 12664
rect 1323 12452 1365 12461
rect 1323 12412 1324 12452
rect 1364 12412 1365 12452
rect 1323 12403 1365 12412
rect 1324 12318 1364 12403
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 1516 12150 1556 12235
rect 652 11192 692 11479
rect 652 11143 692 11152
rect 844 10940 884 10949
rect 940 10940 980 11488
rect 884 10900 980 10940
rect 1132 11488 1268 11528
rect 1324 11612 1364 11621
rect 844 10891 884 10900
rect 1035 10772 1077 10781
rect 1035 10732 1036 10772
rect 1076 10732 1077 10772
rect 1035 10723 1077 10732
rect 1036 10638 1076 10723
rect 844 10268 884 10277
rect 748 10228 844 10268
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9689
rect 748 9680 788 10228
rect 844 10219 884 10228
rect 843 10100 885 10109
rect 843 10060 844 10100
rect 884 10060 885 10100
rect 843 10051 885 10060
rect 692 9640 788 9680
rect 652 9631 692 9640
rect 844 9596 884 10051
rect 748 9556 884 9596
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8924 692 8959
rect 652 8873 692 8884
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 8034 692 8119
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 555 7244 597 7253
rect 555 7204 556 7244
rect 596 7204 597 7244
rect 555 7195 597 7204
rect 652 7194 692 7279
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 652 6320 692 6439
rect 748 6404 788 9556
rect 1036 9512 1076 9521
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 843 9176 885 9185
rect 843 9136 844 9176
rect 884 9136 885 9176
rect 843 9127 885 9136
rect 844 8756 884 9127
rect 844 8707 884 8716
rect 1036 8597 1076 9472
rect 1035 8588 1077 8597
rect 1035 8548 1036 8588
rect 1076 8548 1077 8588
rect 1035 8539 1077 8548
rect 844 7916 884 7925
rect 1132 7916 1172 11488
rect 1324 11033 1364 11572
rect 1612 11108 1652 17260
rect 1996 16484 2036 19963
rect 2379 17156 2421 17165
rect 2379 17116 2380 17156
rect 2420 17116 2421 17156
rect 2379 17107 2421 17116
rect 2187 16904 2229 16913
rect 2187 16864 2188 16904
rect 2228 16864 2229 16904
rect 2187 16855 2229 16864
rect 1996 16435 2036 16444
rect 1804 16400 1844 16409
rect 1804 15569 1844 16360
rect 2188 16316 2228 16855
rect 2188 16267 2228 16276
rect 2380 16316 2420 17107
rect 2571 16568 2613 16577
rect 2571 16528 2572 16568
rect 2612 16528 2613 16568
rect 2571 16519 2613 16528
rect 2572 16484 2612 16519
rect 2572 16433 2612 16444
rect 2380 16267 2420 16276
rect 1996 16064 2036 16073
rect 2036 16024 2516 16064
rect 1996 16015 2036 16024
rect 1803 15560 1845 15569
rect 1803 15520 1804 15560
rect 1844 15520 1845 15560
rect 1803 15511 1845 15520
rect 2284 15560 2324 15569
rect 1995 14888 2037 14897
rect 1995 14848 1996 14888
rect 2036 14848 2037 14888
rect 1995 14839 2037 14848
rect 1708 14804 1748 14813
rect 1708 14645 1748 14764
rect 1996 14754 2036 14839
rect 2187 14804 2229 14813
rect 2187 14764 2188 14804
rect 2228 14764 2229 14804
rect 2187 14755 2229 14764
rect 2188 14670 2228 14755
rect 1707 14636 1749 14645
rect 1707 14596 1708 14636
rect 1748 14596 1749 14636
rect 1707 14587 1749 14596
rect 2187 14384 2229 14393
rect 2187 14344 2188 14384
rect 2228 14344 2229 14384
rect 2187 14335 2229 14344
rect 1707 14048 1749 14057
rect 1707 14008 1708 14048
rect 1748 14008 1749 14048
rect 1707 13999 1749 14008
rect 2091 14048 2133 14057
rect 2091 14008 2092 14048
rect 2132 14008 2133 14048
rect 2091 13999 2133 14008
rect 2188 14048 2228 14335
rect 2284 14216 2324 15520
rect 2379 14720 2421 14729
rect 2379 14680 2380 14720
rect 2420 14680 2421 14720
rect 2379 14671 2421 14680
rect 2476 14720 2516 16024
rect 2571 14888 2613 14897
rect 2668 14888 2708 20047
rect 2764 16988 2804 22819
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3051 21524 3093 21533
rect 3051 21484 3052 21524
rect 3092 21484 3093 21524
rect 3051 21475 3093 21484
rect 3052 21390 3092 21475
rect 3244 21449 3284 21534
rect 3628 21524 3668 21535
rect 3628 21449 3668 21484
rect 3243 21440 3285 21449
rect 3243 21400 3244 21440
rect 3284 21400 3285 21440
rect 3243 21391 3285 21400
rect 3627 21440 3669 21449
rect 3627 21400 3628 21440
rect 3668 21400 3669 21440
rect 3627 21391 3669 21400
rect 3436 21356 3476 21365
rect 3820 21356 3860 21365
rect 3476 21316 3572 21356
rect 3436 21307 3476 21316
rect 3532 21272 3572 21316
rect 3532 21232 3764 21272
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3627 21104 3669 21113
rect 3627 21064 3628 21104
rect 3668 21064 3669 21104
rect 3627 21055 3669 21064
rect 3531 20768 3573 20777
rect 3531 20728 3532 20768
rect 3572 20728 3573 20768
rect 3531 20719 3573 20728
rect 3628 20768 3668 21055
rect 3724 20768 3764 21232
rect 3820 21113 3860 21316
rect 3819 21104 3861 21113
rect 3819 21064 3820 21104
rect 3860 21064 3861 21104
rect 3819 21055 3861 21064
rect 3820 20768 3860 20777
rect 3724 20728 3820 20768
rect 3532 20634 3572 20719
rect 3628 20525 3668 20728
rect 3723 20600 3765 20609
rect 3723 20560 3724 20600
rect 3764 20560 3765 20600
rect 3723 20551 3765 20560
rect 3627 20516 3669 20525
rect 3627 20476 3628 20516
rect 3668 20476 3669 20516
rect 3627 20467 3669 20476
rect 3724 20466 3764 20551
rect 3820 19844 3860 20728
rect 2956 19804 3860 19844
rect 2956 17300 2996 19804
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3916 17300 3956 25087
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4011 21524 4053 21533
rect 4011 21484 4012 21524
rect 4052 21484 4053 21524
rect 4011 21475 4053 21484
rect 4012 21390 4052 21475
rect 4108 18425 4148 23071
rect 4204 21524 4244 26608
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 4780 23129 4820 26776
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 33388 26144 33428 26153
rect 32235 25976 32277 25985
rect 32235 25936 32236 25976
rect 32276 25936 32277 25976
rect 32235 25927 32277 25936
rect 33195 25976 33237 25985
rect 33195 25936 33196 25976
rect 33236 25936 33237 25976
rect 33195 25927 33237 25936
rect 32236 25842 32276 25927
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33196 25556 33236 25927
rect 33388 25901 33428 26104
rect 34252 26144 34292 26935
rect 35019 26900 35061 26909
rect 35019 26860 35020 26900
rect 35060 26860 35061 26900
rect 35019 26851 35061 26860
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34923 26312 34965 26321
rect 34923 26272 34924 26312
rect 34964 26272 34965 26312
rect 34923 26263 34965 26272
rect 34252 26095 34292 26104
rect 34443 26144 34485 26153
rect 34443 26104 34444 26144
rect 34484 26104 34485 26144
rect 34443 26095 34485 26104
rect 34636 26144 34676 26153
rect 34924 26144 34964 26263
rect 34676 26104 34868 26144
rect 34636 26095 34676 26104
rect 34444 25985 34484 26095
rect 34443 25976 34485 25985
rect 34443 25936 34444 25976
rect 34484 25936 34485 25976
rect 34443 25927 34485 25936
rect 33387 25892 33429 25901
rect 33387 25852 33388 25892
rect 33428 25852 33429 25892
rect 33387 25843 33429 25852
rect 33867 25892 33909 25901
rect 33867 25852 33868 25892
rect 33908 25852 33909 25892
rect 33867 25843 33909 25852
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 33196 25516 33428 25556
rect 31755 25388 31797 25397
rect 31755 25348 31756 25388
rect 31796 25348 31797 25388
rect 31755 25339 31797 25348
rect 30124 25304 30164 25313
rect 30987 25304 31029 25313
rect 30164 25264 30260 25304
rect 30124 25255 30164 25264
rect 29740 25220 29780 25229
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 29740 24809 29780 25180
rect 29739 24800 29781 24809
rect 29739 24760 29740 24800
rect 29780 24760 29781 24800
rect 29739 24751 29781 24760
rect 7467 24716 7509 24725
rect 7467 24676 7468 24716
rect 7508 24676 7509 24716
rect 7467 24667 7509 24676
rect 4779 23120 4821 23129
rect 4779 23080 4780 23120
rect 4820 23080 4821 23120
rect 4779 23071 4821 23080
rect 6987 22028 7029 22037
rect 6987 21988 6988 22028
rect 7028 21988 7029 22028
rect 6987 21979 7029 21988
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4204 21475 4244 21484
rect 4395 21524 4437 21533
rect 4395 21484 4396 21524
rect 4436 21484 4437 21524
rect 4395 21475 4437 21484
rect 4396 21356 4436 21475
rect 4396 20693 4436 21316
rect 5067 20852 5109 20861
rect 5067 20812 5068 20852
rect 5108 20812 5109 20852
rect 5067 20803 5109 20812
rect 5068 20718 5108 20803
rect 4395 20684 4437 20693
rect 4395 20644 4396 20684
rect 4436 20644 4437 20684
rect 4395 20635 4437 20644
rect 5260 20600 5300 20609
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4684 20096 4724 20105
rect 4724 20056 4916 20096
rect 4684 20047 4724 20056
rect 4876 19853 4916 20056
rect 5068 20012 5108 20021
rect 5260 20012 5300 20560
rect 5355 20516 5397 20525
rect 5355 20476 5356 20516
rect 5396 20476 5397 20516
rect 5355 20467 5397 20476
rect 5108 19972 5300 20012
rect 4588 19844 4628 19853
rect 4875 19844 4917 19853
rect 4628 19804 4820 19844
rect 4588 19795 4628 19804
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4107 18416 4149 18425
rect 4107 18376 4108 18416
rect 4148 18376 4149 18416
rect 4107 18367 4149 18376
rect 2764 16939 2804 16948
rect 2860 17260 2996 17300
rect 3148 17260 3956 17300
rect 2860 16400 2900 17260
rect 3148 16988 3188 17260
rect 3339 17156 3381 17165
rect 3339 17116 3340 17156
rect 3380 17116 3381 17156
rect 3339 17107 3381 17116
rect 3148 16939 3188 16948
rect 2955 16904 2997 16913
rect 2955 16864 2956 16904
rect 2996 16864 2997 16904
rect 2955 16855 2997 16864
rect 3340 16904 3380 17107
rect 4108 16904 4148 18367
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4780 17300 4820 19804
rect 4875 19804 4876 19844
rect 4916 19804 5012 19844
rect 4875 19795 4917 19804
rect 4876 19710 4916 19795
rect 4875 18584 4917 18593
rect 4875 18544 4876 18584
rect 4916 18544 4917 18584
rect 4875 18535 4917 18544
rect 4492 17260 4820 17300
rect 4203 17072 4245 17081
rect 4203 17032 4204 17072
rect 4244 17032 4245 17072
rect 4203 17023 4245 17032
rect 4396 17072 4436 17081
rect 4204 16938 4244 17023
rect 3340 16855 3380 16864
rect 3724 16864 4148 16904
rect 2956 16770 2996 16855
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 3339 16484 3381 16493
rect 3339 16444 3340 16484
rect 3380 16444 3381 16484
rect 3339 16435 3381 16444
rect 2860 16360 3284 16400
rect 2571 14848 2572 14888
rect 2612 14848 2708 14888
rect 2764 16232 2804 16241
rect 2571 14839 2613 14848
rect 2380 14586 2420 14671
rect 2476 14393 2516 14680
rect 2572 14720 2612 14839
rect 2475 14384 2517 14393
rect 2475 14344 2476 14384
rect 2516 14344 2517 14384
rect 2475 14335 2517 14344
rect 2284 14176 2516 14216
rect 1708 12452 1748 13999
rect 1995 13964 2037 13973
rect 1995 13924 1996 13964
rect 2036 13924 2037 13964
rect 1995 13915 2037 13924
rect 1900 13880 1940 13889
rect 1804 13840 1900 13880
rect 1804 13208 1844 13840
rect 1900 13831 1940 13840
rect 1804 13159 1844 13168
rect 1708 12403 1748 12412
rect 1900 12368 1940 12377
rect 1708 11696 1748 11705
rect 1900 11696 1940 12328
rect 1748 11656 1940 11696
rect 1708 11647 1748 11656
rect 1899 11192 1941 11201
rect 1899 11152 1900 11192
rect 1940 11152 1941 11192
rect 1899 11143 1941 11152
rect 1516 11068 1652 11108
rect 1803 11108 1845 11117
rect 1803 11068 1804 11108
rect 1844 11068 1845 11108
rect 1323 11024 1365 11033
rect 1323 10984 1324 11024
rect 1364 10984 1365 11024
rect 1323 10975 1365 10984
rect 1228 10940 1268 10949
rect 1228 10856 1268 10900
rect 1420 10856 1460 10865
rect 1228 10816 1420 10856
rect 1420 10807 1460 10816
rect 1516 10772 1556 11068
rect 1803 11059 1845 11068
rect 1804 11024 1844 11059
rect 1612 10940 1652 10949
rect 1652 10900 1748 10940
rect 1612 10891 1652 10900
rect 1516 10732 1652 10772
rect 1516 10352 1556 10361
rect 1516 10109 1556 10312
rect 1515 10100 1557 10109
rect 1515 10060 1516 10100
rect 1556 10060 1557 10100
rect 1515 10051 1557 10060
rect 1420 9512 1460 9521
rect 1420 8840 1460 9472
rect 1612 9185 1652 10732
rect 1708 10445 1748 10900
rect 1707 10436 1749 10445
rect 1707 10396 1708 10436
rect 1748 10396 1749 10436
rect 1707 10387 1749 10396
rect 1708 10268 1748 10277
rect 1804 10268 1844 10984
rect 1748 10228 1844 10268
rect 1900 11024 1940 11143
rect 1708 10219 1748 10228
rect 1900 10100 1940 10984
rect 1804 10060 1940 10100
rect 1996 11024 2036 13915
rect 2092 13914 2132 13999
rect 2188 11201 2228 14008
rect 2284 14048 2324 14059
rect 2284 13973 2324 14008
rect 2380 14048 2420 14057
rect 2283 13964 2325 13973
rect 2283 13924 2284 13964
rect 2324 13924 2325 13964
rect 2283 13915 2325 13924
rect 2380 12980 2420 14008
rect 2476 13208 2516 14176
rect 2572 13973 2612 14680
rect 2668 14720 2708 14729
rect 2764 14720 2804 16192
rect 2956 16232 2996 16241
rect 2860 16064 2900 16073
rect 2860 15653 2900 16024
rect 2956 15737 2996 16192
rect 3052 16232 3092 16241
rect 2955 15728 2997 15737
rect 2955 15688 2956 15728
rect 2996 15688 2997 15728
rect 2955 15679 2997 15688
rect 2859 15644 2901 15653
rect 2859 15604 2860 15644
rect 2900 15604 2901 15644
rect 2859 15595 2901 15604
rect 3052 15392 3092 16192
rect 3147 15560 3189 15569
rect 3147 15520 3148 15560
rect 3188 15520 3189 15560
rect 3147 15511 3189 15520
rect 3148 15426 3188 15511
rect 2708 14680 2804 14720
rect 2860 15352 3092 15392
rect 2668 14671 2708 14680
rect 2860 14216 2900 15352
rect 3244 15308 3284 16360
rect 3043 15268 3284 15308
rect 3340 15308 3380 16435
rect 3436 16316 3476 16325
rect 3724 16316 3764 16864
rect 4300 16820 4340 16829
rect 4108 16780 4300 16820
rect 4011 16652 4053 16661
rect 4011 16612 4012 16652
rect 4052 16612 4053 16652
rect 4011 16603 4053 16612
rect 4012 16484 4052 16603
rect 4012 16435 4052 16444
rect 3476 16276 3764 16316
rect 3819 16316 3861 16325
rect 3819 16276 3820 16316
rect 3860 16276 3861 16316
rect 3436 16267 3476 16276
rect 3819 16267 3861 16276
rect 3820 16182 3860 16267
rect 3627 16064 3669 16073
rect 3627 16024 3628 16064
rect 3668 16024 3669 16064
rect 3627 16015 3669 16024
rect 3915 16064 3957 16073
rect 3915 16024 3916 16064
rect 3956 16024 3957 16064
rect 3915 16015 3957 16024
rect 3628 15930 3668 16015
rect 3819 15728 3861 15737
rect 3819 15688 3820 15728
rect 3860 15688 3861 15728
rect 3819 15679 3861 15688
rect 3531 15644 3573 15653
rect 3531 15604 3532 15644
rect 3572 15604 3573 15644
rect 3531 15595 3573 15604
rect 3820 15644 3860 15679
rect 3532 15510 3572 15595
rect 3820 15593 3860 15604
rect 3724 15560 3764 15569
rect 3628 15520 3724 15560
rect 3340 15268 3572 15308
rect 3043 15224 3083 15268
rect 2956 15184 3083 15224
rect 2956 14888 2996 15184
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 2956 14848 3092 14888
rect 2956 14720 2996 14729
rect 2956 14477 2996 14680
rect 2955 14468 2997 14477
rect 2955 14428 2956 14468
rect 2996 14428 2997 14468
rect 2955 14419 2997 14428
rect 2860 14167 2900 14176
rect 2667 14048 2709 14057
rect 2667 14008 2668 14048
rect 2708 14008 2709 14048
rect 2667 13999 2709 14008
rect 2764 14048 2804 14057
rect 2956 14048 2996 14057
rect 3052 14048 3092 14848
rect 3244 14720 3284 14731
rect 3244 14645 3284 14680
rect 3339 14720 3381 14729
rect 3339 14680 3340 14720
rect 3380 14680 3381 14720
rect 3339 14671 3381 14680
rect 3243 14636 3285 14645
rect 3243 14596 3244 14636
rect 3284 14596 3285 14636
rect 3243 14587 3285 14596
rect 3340 14586 3380 14671
rect 3243 14468 3285 14477
rect 3243 14428 3244 14468
rect 3284 14428 3285 14468
rect 3243 14419 3285 14428
rect 2571 13964 2613 13973
rect 2571 13924 2572 13964
rect 2612 13924 2613 13964
rect 2571 13915 2613 13924
rect 2668 13914 2708 13999
rect 2764 13217 2804 14008
rect 2860 14008 2956 14048
rect 2996 14008 3092 14048
rect 3244 14048 3284 14419
rect 3532 14384 3572 15268
rect 3628 14972 3668 15520
rect 3724 15511 3764 15520
rect 3916 15560 3956 16015
rect 4011 15812 4053 15821
rect 4011 15772 4012 15812
rect 4052 15772 4053 15812
rect 4011 15763 4053 15772
rect 3628 14923 3668 14932
rect 3436 14344 3572 14384
rect 3436 14048 3476 14344
rect 3531 14216 3573 14225
rect 3531 14176 3532 14216
rect 3572 14176 3573 14216
rect 3531 14167 3573 14176
rect 3284 14008 3476 14048
rect 2668 13208 2708 13217
rect 2476 13168 2668 13208
rect 2284 12940 2420 12980
rect 2284 12536 2324 12940
rect 2475 12872 2517 12881
rect 2475 12832 2476 12872
rect 2516 12832 2517 12872
rect 2475 12823 2517 12832
rect 2379 12704 2421 12713
rect 2379 12664 2380 12704
rect 2420 12664 2421 12704
rect 2379 12655 2421 12664
rect 2380 12570 2420 12655
rect 2284 12487 2324 12496
rect 2476 12536 2516 12823
rect 2668 12797 2708 13168
rect 2763 13208 2805 13217
rect 2763 13168 2764 13208
rect 2804 13168 2805 13208
rect 2763 13159 2805 13168
rect 2860 12980 2900 14008
rect 2956 13999 2996 14008
rect 3244 13999 3284 14008
rect 3436 13796 3476 14008
rect 3532 14048 3572 14167
rect 3532 13999 3572 14008
rect 3627 14048 3669 14057
rect 3627 14008 3628 14048
rect 3668 14008 3669 14048
rect 3627 13999 3669 14008
rect 3819 14048 3861 14057
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 3628 13914 3668 13999
rect 3436 13756 3668 13796
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3531 13292 3573 13301
rect 3531 13252 3532 13292
rect 3572 13252 3573 13292
rect 3531 13243 3573 13252
rect 2955 13208 2997 13217
rect 2955 13168 2956 13208
rect 2996 13168 2997 13208
rect 2955 13159 2997 13168
rect 2764 12940 2900 12980
rect 2667 12788 2709 12797
rect 2667 12748 2668 12788
rect 2708 12748 2709 12788
rect 2667 12739 2709 12748
rect 2476 12487 2516 12496
rect 2572 12536 2612 12545
rect 2572 12377 2612 12496
rect 2571 12368 2613 12377
rect 2571 12328 2572 12368
rect 2612 12328 2613 12368
rect 2571 12319 2613 12328
rect 2572 11696 2612 11705
rect 2668 11696 2708 12739
rect 2764 12536 2804 12940
rect 2956 12536 2996 13159
rect 2804 12496 2891 12536
rect 2764 12487 2804 12496
rect 2763 12368 2805 12377
rect 2763 12328 2764 12368
rect 2804 12328 2805 12368
rect 2763 12319 2805 12328
rect 2764 12234 2804 12319
rect 2851 12116 2891 12496
rect 2956 12487 2996 12496
rect 3052 12536 3092 12545
rect 3052 12284 3092 12496
rect 2380 11656 2572 11696
rect 2612 11656 2708 11696
rect 2764 12076 2891 12116
rect 2956 12244 3092 12284
rect 2187 11192 2229 11201
rect 2187 11152 2188 11192
rect 2228 11152 2229 11192
rect 2187 11143 2229 11152
rect 1611 9176 1653 9185
rect 1611 9136 1612 9176
rect 1652 9136 1653 9176
rect 1611 9127 1653 9136
rect 1516 8840 1556 8849
rect 1420 8800 1516 8840
rect 1516 8791 1556 8800
rect 1707 8756 1749 8765
rect 1707 8716 1708 8756
rect 1748 8716 1749 8756
rect 1707 8707 1749 8716
rect 884 7876 1172 7916
rect 1708 8672 1748 8707
rect 1708 7916 1748 8632
rect 1804 8672 1844 10060
rect 1996 8840 2036 10984
rect 2092 11024 2132 11033
rect 2284 11024 2324 11033
rect 2132 10984 2284 11024
rect 2092 10975 2132 10984
rect 2284 10975 2324 10984
rect 2283 10856 2325 10865
rect 2283 10816 2284 10856
rect 2324 10816 2325 10856
rect 2283 10807 2325 10816
rect 2284 10722 2324 10807
rect 2284 9512 2324 9521
rect 2380 9512 2420 11656
rect 2572 11647 2612 11656
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2572 11024 2612 11033
rect 2476 10890 2516 10975
rect 2475 10436 2517 10445
rect 2475 10396 2476 10436
rect 2516 10396 2517 10436
rect 2475 10387 2517 10396
rect 2572 10436 2612 10984
rect 2764 10436 2804 12076
rect 2956 11537 2996 12244
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3532 11948 3572 13243
rect 3628 12620 3668 13756
rect 3820 13460 3860 13999
rect 3916 13964 3956 15520
rect 4012 14645 4052 15763
rect 4108 15560 4148 16780
rect 4300 16771 4340 16780
rect 4396 16493 4436 17032
rect 4395 16484 4437 16493
rect 4300 16444 4396 16484
rect 4436 16444 4437 16484
rect 4204 16400 4244 16411
rect 4204 16325 4244 16360
rect 4203 16316 4245 16325
rect 4203 16276 4204 16316
rect 4244 16276 4245 16316
rect 4203 16267 4245 16276
rect 4300 16064 4340 16444
rect 4395 16435 4437 16444
rect 4396 16316 4436 16325
rect 4492 16316 4532 17260
rect 4587 17072 4629 17081
rect 4587 17032 4588 17072
rect 4628 17032 4629 17072
rect 4587 17023 4629 17032
rect 4588 16904 4628 17023
rect 4780 16988 4820 16997
rect 4876 16988 4916 18535
rect 4820 16948 4916 16988
rect 4780 16939 4820 16948
rect 4588 16855 4628 16864
rect 4972 16400 5012 19804
rect 5068 19769 5108 19972
rect 5067 19760 5109 19769
rect 5067 19720 5068 19760
rect 5108 19720 5109 19760
rect 5067 19711 5109 19720
rect 5356 18593 5396 20467
rect 5355 18584 5397 18593
rect 5355 18544 5356 18584
rect 5396 18544 5397 18584
rect 5355 18535 5397 18544
rect 5163 17072 5205 17081
rect 5163 17032 5164 17072
rect 5204 17032 5205 17072
rect 5163 17023 5205 17032
rect 5067 16652 5109 16661
rect 5067 16612 5068 16652
rect 5108 16612 5109 16652
rect 5067 16603 5109 16612
rect 4436 16276 4532 16316
rect 4876 16360 5012 16400
rect 4396 16267 4436 16276
rect 4588 16148 4628 16157
rect 4628 16108 4820 16148
rect 4588 16099 4628 16108
rect 4204 16024 4340 16064
rect 4204 15821 4244 16024
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4203 15812 4245 15821
rect 4203 15772 4204 15812
rect 4244 15772 4245 15812
rect 4203 15763 4245 15772
rect 4395 15728 4437 15737
rect 4395 15688 4396 15728
rect 4436 15688 4437 15728
rect 4395 15679 4437 15688
rect 4492 15728 4532 15737
rect 4780 15728 4820 16108
rect 4532 15688 4820 15728
rect 4492 15679 4532 15688
rect 4300 15560 4340 15569
rect 4108 15520 4300 15560
rect 4300 15511 4340 15520
rect 4396 15560 4436 15679
rect 4396 15511 4436 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4779 15560 4821 15569
rect 4779 15520 4780 15560
rect 4820 15520 4821 15560
rect 4779 15511 4821 15520
rect 4588 15426 4628 15511
rect 4011 14636 4053 14645
rect 4011 14596 4012 14636
rect 4052 14596 4053 14636
rect 4011 14587 4053 14596
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4203 14216 4245 14225
rect 4203 14176 4204 14216
rect 4244 14176 4245 14216
rect 4203 14167 4245 14176
rect 3916 13924 4148 13964
rect 3916 13796 3956 13805
rect 3956 13756 4052 13796
rect 3916 13747 3956 13756
rect 3820 13411 3860 13420
rect 3627 12580 3668 12620
rect 3627 12452 3667 12580
rect 4012 12536 4052 13756
rect 4108 13040 4148 13924
rect 4204 13208 4244 14167
rect 4396 14048 4436 14057
rect 4300 13460 4340 13469
rect 4396 13460 4436 14008
rect 4340 13420 4436 13460
rect 4492 14048 4532 14057
rect 4684 14048 4724 14057
rect 4780 14048 4820 15511
rect 4876 14813 4916 16360
rect 4972 16232 5012 16241
rect 4972 15392 5012 16192
rect 5068 15569 5108 16603
rect 5067 15560 5109 15569
rect 5067 15520 5068 15560
rect 5108 15520 5109 15560
rect 5067 15511 5109 15520
rect 5068 15392 5108 15401
rect 4972 15352 5068 15392
rect 5068 15343 5108 15352
rect 4875 14804 4917 14813
rect 4875 14764 4876 14804
rect 4916 14764 4917 14804
rect 4875 14755 4917 14764
rect 4300 13411 4340 13420
rect 4396 13217 4436 13302
rect 4204 13159 4244 13168
rect 4395 13208 4437 13217
rect 4395 13168 4396 13208
rect 4436 13168 4437 13208
rect 4395 13159 4437 13168
rect 4492 13049 4532 14008
rect 4588 14008 4684 14048
rect 4724 14008 4820 14048
rect 4876 14048 4916 14057
rect 4491 13040 4533 13049
rect 4108 13000 4244 13040
rect 4107 12872 4149 12881
rect 4107 12832 4108 12872
rect 4148 12832 4149 12872
rect 4107 12823 4149 12832
rect 4108 12620 4148 12823
rect 4108 12571 4148 12580
rect 4012 12487 4052 12496
rect 4204 12536 4244 13000
rect 4491 13000 4492 13040
rect 4532 13000 4533 13040
rect 4588 13040 4628 14008
rect 4684 13999 4724 14008
rect 4684 13880 4724 13889
rect 4876 13880 4916 14008
rect 4724 13840 4916 13880
rect 4684 13831 4724 13840
rect 5164 13217 5204 17023
rect 6988 16493 7028 21979
rect 6987 16484 7029 16493
rect 6987 16444 6988 16484
rect 7028 16444 7029 16484
rect 6987 16435 7029 16444
rect 6988 16350 7028 16435
rect 5836 16232 5876 16241
rect 5260 14048 5300 14057
rect 5836 14048 5876 16192
rect 7371 15308 7413 15317
rect 7371 15268 7372 15308
rect 7412 15268 7413 15308
rect 7371 15259 7413 15268
rect 7275 14216 7317 14225
rect 7275 14176 7276 14216
rect 7316 14176 7317 14216
rect 7275 14167 7317 14176
rect 7276 14082 7316 14167
rect 6124 14048 6164 14057
rect 5300 14008 5588 14048
rect 5836 14008 6124 14048
rect 6164 14008 6260 14048
rect 5260 13999 5300 14008
rect 5548 13376 5588 14008
rect 6124 13999 6164 14008
rect 5548 13327 5588 13336
rect 4972 13208 5012 13217
rect 4588 13000 4820 13040
rect 4491 12991 4533 13000
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4780 12704 4820 13000
rect 4972 12797 5012 13168
rect 5163 13208 5205 13217
rect 5163 13168 5164 13208
rect 5204 13168 5205 13208
rect 5163 13159 5205 13168
rect 4971 12788 5013 12797
rect 4971 12748 4972 12788
rect 5012 12748 5013 12788
rect 4971 12739 5013 12748
rect 3627 12412 3668 12452
rect 3436 11908 3572 11948
rect 2955 11528 2997 11537
rect 2955 11488 2956 11528
rect 2996 11488 2997 11528
rect 2955 11479 2997 11488
rect 3436 11201 3476 11908
rect 3531 11528 3573 11537
rect 3531 11488 3532 11528
rect 3572 11488 3573 11528
rect 3531 11479 3573 11488
rect 3435 11192 3477 11201
rect 3435 11152 3436 11192
rect 3476 11152 3477 11192
rect 3435 11143 3477 11152
rect 3148 11024 3188 11033
rect 3148 10772 3188 10984
rect 3436 11024 3476 11143
rect 3532 11117 3572 11479
rect 3531 11108 3573 11117
rect 3531 11068 3532 11108
rect 3572 11068 3573 11108
rect 3531 11059 3573 11068
rect 3436 10975 3476 10984
rect 3532 10974 3572 11059
rect 3628 10772 3668 12412
rect 3916 11696 3956 11705
rect 3723 11528 3765 11537
rect 3723 11488 3724 11528
rect 3764 11488 3765 11528
rect 3723 11479 3765 11488
rect 3724 11394 3764 11479
rect 3820 10856 3860 10865
rect 3916 10856 3956 11656
rect 4108 11696 4148 11705
rect 4204 11696 4244 12496
rect 4148 11656 4244 11696
rect 4492 12664 4820 12704
rect 4492 11696 4532 12664
rect 4779 12536 4821 12545
rect 4779 12496 4780 12536
rect 4820 12496 4821 12536
rect 4779 12487 4821 12496
rect 4780 12402 4820 12487
rect 4972 12368 5012 12739
rect 4972 12319 5012 12328
rect 4012 11612 4052 11621
rect 4012 11537 4052 11572
rect 4011 11528 4053 11537
rect 4011 11488 4012 11528
rect 4052 11488 4053 11528
rect 4011 11479 4053 11488
rect 4012 11033 4052 11479
rect 4011 11024 4053 11033
rect 4011 10984 4012 11024
rect 4052 10984 4053 11024
rect 4011 10975 4053 10984
rect 3860 10816 3956 10856
rect 3820 10807 3860 10816
rect 3148 10732 3668 10772
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 2572 10387 2612 10396
rect 2668 10396 2804 10436
rect 2324 9472 2420 9512
rect 2284 9463 2324 9472
rect 1804 8168 1844 8632
rect 1900 8800 2036 8840
rect 2476 8840 2516 10387
rect 2668 10268 2708 10396
rect 3052 10361 3092 10446
rect 2859 10352 2901 10361
rect 2572 10228 2708 10268
rect 2764 10312 2860 10352
rect 2900 10312 2901 10352
rect 2572 10184 2612 10228
rect 2764 10184 2804 10312
rect 2859 10303 2901 10312
rect 3051 10352 3093 10361
rect 3051 10312 3052 10352
rect 3092 10312 3093 10352
rect 3051 10303 3093 10312
rect 2860 10284 2900 10303
rect 3243 10268 3285 10277
rect 3243 10228 3244 10268
rect 3284 10228 3285 10268
rect 3243 10219 3285 10228
rect 2572 9017 2612 10144
rect 2668 10144 2764 10184
rect 2571 9008 2613 9017
rect 2571 8968 2572 9008
rect 2612 8968 2613 9008
rect 2571 8959 2613 8968
rect 2476 8800 2612 8840
rect 1900 8672 1940 8800
rect 2188 8672 2228 8681
rect 1900 8420 1940 8632
rect 1996 8632 2188 8672
rect 1996 8588 2036 8632
rect 2188 8623 2228 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2476 8672 2516 8681
rect 1996 8539 2036 8548
rect 2283 8588 2325 8597
rect 2283 8548 2284 8588
rect 2324 8548 2325 8588
rect 2283 8539 2325 8548
rect 2284 8454 2324 8539
rect 2380 8538 2420 8623
rect 1900 8380 2228 8420
rect 1804 8128 2132 8168
rect 844 7867 884 7876
rect 1708 7867 1748 7876
rect 1996 8000 2036 8009
rect 1324 7832 1364 7841
rect 1364 7792 1460 7832
rect 1324 7783 1364 7792
rect 939 7748 981 7757
rect 939 7708 940 7748
rect 980 7708 981 7748
rect 939 7699 981 7708
rect 843 7244 885 7253
rect 843 7204 844 7244
rect 884 7204 885 7244
rect 843 7195 885 7204
rect 844 7110 884 7195
rect 844 6404 884 6413
rect 748 6364 844 6404
rect 844 6355 884 6364
rect 652 6271 692 6280
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5144 692 5599
rect 844 5480 884 5489
rect 652 5095 692 5104
rect 748 5440 844 5480
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4304 692 4759
rect 652 4255 692 4264
rect 748 4220 788 5440
rect 844 5431 884 5440
rect 844 4892 884 4901
rect 940 4892 980 7699
rect 1035 7664 1077 7673
rect 1035 7624 1036 7664
rect 1076 7624 1077 7664
rect 1035 7615 1077 7624
rect 1036 5732 1076 7615
rect 1420 7160 1460 7792
rect 1515 7748 1557 7757
rect 1515 7708 1516 7748
rect 1556 7708 1557 7748
rect 1515 7699 1557 7708
rect 1516 7614 1556 7699
rect 1996 7673 2036 7960
rect 2092 8000 2132 8128
rect 1995 7664 2037 7673
rect 1995 7624 1996 7664
rect 2036 7624 2037 7664
rect 1995 7615 2037 7624
rect 2092 7244 2132 7960
rect 1996 7204 2132 7244
rect 2188 8000 2228 8380
rect 1708 7160 1748 7169
rect 1420 7120 1708 7160
rect 1708 7111 1748 7120
rect 1324 7076 1364 7085
rect 1324 6329 1364 7036
rect 1323 6320 1365 6329
rect 1323 6280 1324 6320
rect 1364 6280 1365 6320
rect 1323 6271 1365 6280
rect 1708 6320 1748 6329
rect 1036 5683 1076 5692
rect 1612 5648 1652 5657
rect 1708 5648 1748 6280
rect 1803 5732 1845 5741
rect 1803 5692 1804 5732
rect 1844 5692 1845 5732
rect 1803 5683 1845 5692
rect 1652 5608 1748 5648
rect 1612 5599 1652 5608
rect 1228 5564 1268 5573
rect 1804 5564 1844 5683
rect 1228 5153 1268 5524
rect 1708 5524 1844 5564
rect 1227 5144 1269 5153
rect 1227 5104 1228 5144
rect 1268 5104 1269 5144
rect 1227 5095 1269 5104
rect 1708 4976 1748 5524
rect 1996 5480 2036 7204
rect 2188 7160 2228 7960
rect 884 4852 980 4892
rect 1516 4892 1556 4901
rect 1708 4892 1748 4936
rect 1804 5440 2036 5480
rect 2092 7120 2228 7160
rect 2284 8000 2324 8009
rect 1804 4976 1844 5440
rect 2092 5228 2132 7120
rect 2188 6488 2228 6497
rect 2284 6488 2324 7960
rect 2476 7748 2516 8632
rect 2572 8336 2612 8800
rect 2668 8513 2708 10144
rect 2764 10135 2804 10144
rect 2870 10169 2910 10178
rect 3244 10134 3284 10219
rect 2870 9857 2910 10129
rect 2869 9848 2911 9857
rect 3435 9848 3477 9857
rect 2869 9808 2870 9848
rect 2910 9808 2996 9848
rect 2869 9799 2911 9808
rect 2763 9344 2805 9353
rect 2763 9304 2764 9344
rect 2804 9304 2805 9344
rect 2763 9295 2805 9304
rect 2764 8933 2804 9295
rect 2763 8924 2805 8933
rect 2763 8884 2764 8924
rect 2804 8884 2805 8924
rect 2763 8875 2805 8884
rect 2764 8672 2804 8875
rect 2956 8765 2996 9808
rect 3435 9808 3436 9848
rect 3476 9808 3477 9848
rect 3435 9799 3477 9808
rect 3436 9680 3476 9799
rect 3436 9631 3476 9640
rect 3532 9353 3572 10732
rect 3628 9512 3668 9521
rect 3531 9344 3573 9353
rect 3531 9304 3532 9344
rect 3572 9304 3573 9344
rect 3531 9295 3573 9304
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3339 8924 3381 8933
rect 3339 8884 3340 8924
rect 3380 8884 3381 8924
rect 3339 8875 3381 8884
rect 3436 8924 3476 8933
rect 3628 8924 3668 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 3820 9512 3860 9521
rect 4108 9512 4148 11656
rect 4492 11528 4532 11656
rect 4588 11824 5012 11864
rect 4588 11612 4628 11824
rect 4588 11563 4628 11572
rect 4684 11696 4724 11705
rect 4684 11537 4724 11656
rect 4780 11696 4820 11705
rect 4204 11488 4532 11528
rect 4683 11528 4725 11537
rect 4683 11488 4684 11528
rect 4724 11488 4725 11528
rect 4204 11192 4244 11488
rect 4683 11479 4725 11488
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4780 11192 4820 11656
rect 4972 11696 5012 11824
rect 4972 11647 5012 11656
rect 4204 11152 4340 11192
rect 4780 11152 5012 11192
rect 4300 10100 4340 11152
rect 4972 11108 5012 11152
rect 4972 11059 5012 11068
rect 4876 11024 4916 11033
rect 4876 10772 4916 10984
rect 5067 11024 5109 11033
rect 5067 10984 5068 11024
rect 5108 10984 5109 11024
rect 5067 10975 5109 10984
rect 5068 10890 5108 10975
rect 5164 10772 5204 13159
rect 5451 12536 5493 12545
rect 5451 12496 5452 12536
rect 5492 12496 5493 12536
rect 5451 12487 5493 12496
rect 5644 12536 5684 12545
rect 5355 12368 5397 12377
rect 5355 12328 5356 12368
rect 5396 12328 5397 12368
rect 5355 12319 5397 12328
rect 5356 11696 5396 12319
rect 5356 11647 5396 11656
rect 4876 10732 5204 10772
rect 4876 10277 4916 10732
rect 4875 10268 4917 10277
rect 4875 10228 4876 10268
rect 4916 10228 4917 10268
rect 4875 10219 4917 10228
rect 3860 9472 4148 9512
rect 4204 10060 4340 10100
rect 4780 10100 4820 10109
rect 4204 9512 4244 10060
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4492 9680 4532 9689
rect 4780 9680 4820 10060
rect 4532 9640 4820 9680
rect 4492 9631 4532 9640
rect 4396 9512 4436 9521
rect 4204 9472 4396 9512
rect 3476 8884 3668 8924
rect 3724 9260 3764 9463
rect 3436 8875 3476 8884
rect 3051 8840 3093 8849
rect 3051 8800 3052 8840
rect 3092 8800 3093 8840
rect 3051 8791 3093 8800
rect 2955 8756 2997 8765
rect 2955 8716 2956 8756
rect 2996 8716 2997 8756
rect 2955 8707 2997 8716
rect 2764 8623 2804 8632
rect 3052 8672 3092 8791
rect 3147 8756 3189 8765
rect 3147 8716 3148 8756
rect 3188 8716 3189 8756
rect 3147 8707 3189 8716
rect 3052 8623 3092 8632
rect 3148 8672 3188 8707
rect 3148 8621 3188 8632
rect 2667 8504 2709 8513
rect 2667 8464 2668 8504
rect 2708 8464 2709 8504
rect 2667 8455 2709 8464
rect 2572 8296 2891 8336
rect 2851 8252 2891 8296
rect 2851 8212 3092 8252
rect 2764 8093 2804 8124
rect 2763 8084 2805 8093
rect 2763 8044 2764 8084
rect 2804 8044 2805 8084
rect 2763 8035 2805 8044
rect 2571 8000 2613 8009
rect 2764 8000 2804 8035
rect 2571 7960 2572 8000
rect 2612 7960 2708 8000
rect 2571 7951 2613 7960
rect 2572 7866 2612 7951
rect 2572 7748 2612 7757
rect 2476 7708 2572 7748
rect 2572 7699 2612 7708
rect 2572 7160 2612 7169
rect 2379 7076 2421 7085
rect 2379 7036 2380 7076
rect 2420 7036 2421 7076
rect 2379 7027 2421 7036
rect 2228 6448 2324 6488
rect 2380 6488 2420 7027
rect 2188 6439 2228 6448
rect 2380 6439 2420 6448
rect 2476 6488 2516 6497
rect 2476 6329 2516 6448
rect 2187 6320 2229 6329
rect 2187 6280 2188 6320
rect 2228 6280 2229 6320
rect 2187 6271 2229 6280
rect 2475 6320 2517 6329
rect 2475 6280 2476 6320
rect 2516 6280 2517 6320
rect 2475 6271 2517 6280
rect 2188 6186 2228 6271
rect 2475 5648 2517 5657
rect 2572 5648 2612 7120
rect 2668 6497 2708 7960
rect 2667 6488 2709 6497
rect 2667 6448 2668 6488
rect 2708 6448 2709 6488
rect 2667 6439 2709 6448
rect 2764 6404 2804 7960
rect 2877 8000 2919 8009
rect 2877 7960 2878 8000
rect 2918 7960 2919 8000
rect 2877 7951 2919 7960
rect 2878 7673 2918 7951
rect 3052 7748 3092 8212
rect 3340 8000 3380 8875
rect 3724 8681 3764 9220
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 3628 8000 3668 8009
rect 3380 7960 3572 8000
rect 3340 7951 3380 7960
rect 2974 7708 3092 7748
rect 2877 7664 2919 7673
rect 2877 7624 2878 7664
rect 2918 7624 2919 7664
rect 2877 7615 2919 7624
rect 2974 7580 3014 7708
rect 2956 7540 3014 7580
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 2956 7412 2996 7540
rect 3112 7531 3480 7540
rect 2956 7372 3092 7412
rect 2859 6740 2901 6749
rect 2859 6700 2860 6740
rect 2900 6700 2901 6740
rect 2859 6691 2901 6700
rect 2860 6530 2900 6691
rect 3052 6497 3092 7372
rect 3532 6581 3572 7960
rect 3628 7757 3668 7960
rect 3723 8000 3765 8009
rect 3723 7960 3724 8000
rect 3764 7960 3765 8000
rect 3723 7951 3765 7960
rect 3627 7748 3669 7757
rect 3627 7708 3628 7748
rect 3668 7708 3669 7748
rect 3627 7699 3669 7708
rect 3724 7412 3764 7951
rect 3724 7363 3764 7372
rect 3820 6824 3860 9472
rect 4107 9344 4149 9353
rect 4107 9304 4108 9344
rect 4148 9304 4149 9344
rect 4107 9295 4149 9304
rect 4108 8513 4148 9295
rect 4107 8504 4149 8513
rect 4396 8504 4436 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4684 9512 4724 9521
rect 4588 9378 4628 9463
rect 4684 9344 4724 9472
rect 4876 9512 4916 10219
rect 5164 10184 5204 10193
rect 5204 10144 5300 10184
rect 5164 10135 5204 10144
rect 5067 10016 5109 10025
rect 5067 9976 5068 10016
rect 5108 9976 5109 10016
rect 5067 9967 5109 9976
rect 4876 9463 4916 9472
rect 5068 9512 5108 9967
rect 4972 9344 5012 9353
rect 4684 9304 4972 9344
rect 4972 9295 5012 9304
rect 5068 8849 5108 9472
rect 5260 9344 5300 10144
rect 5260 9295 5300 9304
rect 5067 8840 5109 8849
rect 5067 8800 5068 8840
rect 5108 8800 5109 8840
rect 5067 8791 5109 8800
rect 5260 8840 5300 8849
rect 4107 8464 4108 8504
rect 4148 8464 4149 8504
rect 4107 8455 4149 8464
rect 4204 8464 4436 8504
rect 4204 8000 4244 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4396 8168 4436 8177
rect 4436 8128 4820 8168
rect 4396 8119 4436 8128
rect 4780 8084 4820 8128
rect 4780 8035 4820 8044
rect 4299 8000 4341 8009
rect 4204 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4492 8000 4532 8009
rect 4300 7866 4340 7951
rect 4012 7748 4052 7757
rect 4012 7160 4052 7708
rect 4012 7111 4052 7120
rect 4204 7160 4244 7169
rect 4107 7076 4149 7085
rect 4107 7036 4108 7076
rect 4148 7036 4149 7076
rect 4107 7027 4149 7036
rect 4108 6942 4148 7027
rect 4204 6824 4244 7120
rect 4492 7085 4532 7960
rect 4588 8000 4628 8009
rect 4588 7412 4628 7960
rect 5164 8000 5204 8009
rect 5260 8000 5300 8800
rect 5204 7960 5300 8000
rect 5164 7951 5204 7960
rect 4971 7748 5013 7757
rect 4971 7708 4972 7748
rect 5012 7708 5013 7748
rect 4971 7699 5013 7708
rect 4876 7412 4916 7421
rect 4588 7372 4876 7412
rect 4876 7363 4916 7372
rect 4780 7160 4820 7169
rect 4972 7160 5012 7699
rect 4820 7120 4916 7160
rect 4780 7111 4820 7120
rect 4491 7076 4533 7085
rect 4491 7036 4492 7076
rect 4532 7036 4533 7076
rect 4491 7027 4533 7036
rect 3820 6784 4244 6824
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 3531 6572 3573 6581
rect 3531 6532 3532 6572
rect 3572 6532 3580 6572
rect 3531 6523 3580 6532
rect 2860 6404 2900 6490
rect 2764 6364 2900 6404
rect 2956 6488 2996 6497
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 2668 6186 2708 6271
rect 2667 6068 2709 6077
rect 2667 6028 2668 6068
rect 2708 6028 2709 6068
rect 2667 6019 2709 6028
rect 2475 5608 2476 5648
rect 2516 5608 2612 5648
rect 2475 5599 2517 5608
rect 1804 4901 1844 4936
rect 1900 5188 2132 5228
rect 1900 4976 1940 5188
rect 2476 5153 2516 5599
rect 2283 5144 2325 5153
rect 1996 5104 2228 5144
rect 1996 5060 2036 5104
rect 1996 5011 2036 5020
rect 2188 5018 2228 5104
rect 2283 5104 2284 5144
rect 2324 5104 2325 5144
rect 2283 5095 2325 5104
rect 2475 5144 2517 5153
rect 2475 5104 2476 5144
rect 2516 5104 2517 5144
rect 2475 5095 2517 5104
rect 2284 5010 2324 5095
rect 2188 4969 2228 4978
rect 2380 4976 2420 4985
rect 1556 4852 1748 4892
rect 1803 4892 1845 4901
rect 1803 4852 1804 4892
rect 1844 4852 1845 4892
rect 844 4843 884 4852
rect 1516 4843 1556 4852
rect 1803 4843 1845 4852
rect 1324 4724 1364 4733
rect 1228 4684 1324 4724
rect 844 4220 884 4229
rect 748 4180 844 4220
rect 844 4171 884 4180
rect 1228 4220 1268 4684
rect 1324 4675 1364 4684
rect 1900 4649 1940 4936
rect 2187 4892 2229 4901
rect 2187 4852 2188 4892
rect 2228 4852 2229 4892
rect 2187 4843 2229 4852
rect 1899 4640 1941 4649
rect 1899 4600 1900 4640
rect 1940 4600 1941 4640
rect 1899 4591 1941 4600
rect 1900 4304 1940 4313
rect 1228 4171 1268 4180
rect 1804 4264 1900 4304
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 1036 3834 1076 3919
rect 1420 3464 1460 3473
rect 844 3380 884 3389
rect 844 3296 884 3340
rect 1227 3380 1269 3389
rect 1227 3340 1228 3380
rect 1268 3340 1269 3380
rect 1227 3331 1269 3340
rect 1036 3296 1076 3305
rect 844 3256 1036 3296
rect 1036 3247 1076 3256
rect 1228 3246 1268 3331
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 843 2792 885 2801
rect 843 2752 844 2792
rect 884 2752 885 2792
rect 843 2743 885 2752
rect 844 2708 884 2743
rect 844 2657 884 2668
rect 1420 2549 1460 3424
rect 1804 3464 1844 4264
rect 1900 4255 1940 4264
rect 2091 4136 2133 4145
rect 2091 4096 2092 4136
rect 2132 4096 2133 4136
rect 2091 4087 2133 4096
rect 2188 4136 2228 4843
rect 2380 4817 2420 4936
rect 2476 4976 2516 4985
rect 2516 4936 2549 4976
rect 2476 4927 2549 4936
rect 2509 4892 2549 4927
rect 2509 4852 2612 4892
rect 2379 4808 2421 4817
rect 2379 4768 2380 4808
rect 2420 4768 2421 4808
rect 2379 4759 2421 4768
rect 2475 4724 2517 4733
rect 2475 4684 2476 4724
rect 2516 4684 2517 4724
rect 2475 4675 2517 4684
rect 2283 4640 2325 4649
rect 2283 4600 2284 4640
rect 2324 4600 2325 4640
rect 2283 4591 2325 4600
rect 2188 4087 2228 4096
rect 2284 4136 2324 4591
rect 2284 4087 2324 4096
rect 1804 3415 1844 3424
rect 2092 3389 2132 4087
rect 2380 3968 2420 3977
rect 2091 3380 2133 3389
rect 2091 3340 2092 3380
rect 2132 3340 2133 3380
rect 2091 3331 2133 3340
rect 1515 2792 1557 2801
rect 1515 2752 1516 2792
rect 1556 2752 1557 2792
rect 1515 2743 1557 2752
rect 1516 2658 1556 2743
rect 1707 2708 1749 2717
rect 1707 2668 1708 2708
rect 1748 2668 1749 2708
rect 1707 2659 1749 2668
rect 1708 2574 1748 2659
rect 2380 2624 2420 3928
rect 2476 3464 2516 4675
rect 2572 4388 2612 4852
rect 2572 4339 2612 4348
rect 2572 4136 2612 4145
rect 2572 3884 2612 4096
rect 2668 3884 2708 6019
rect 2764 4388 2804 6364
rect 2956 5741 2996 6448
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3540 6404 3580 6523
rect 3532 6364 3580 6404
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 2955 5732 2997 5741
rect 2955 5692 2956 5732
rect 2996 5692 2997 5732
rect 2955 5683 2997 5692
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 2764 4348 2996 4388
rect 2956 4304 2996 4348
rect 2956 4264 3006 4304
rect 2878 4145 2918 4230
rect 2764 4136 2804 4145
rect 2764 3968 2804 4096
rect 2877 4136 2919 4145
rect 2877 4096 2878 4136
rect 2918 4096 2919 4136
rect 2877 4087 2919 4096
rect 2966 4052 3006 4264
rect 3532 4136 3572 6364
rect 3820 6236 3860 6245
rect 3724 6196 3820 6236
rect 3627 5732 3669 5741
rect 3627 5692 3628 5732
rect 3668 5692 3669 5732
rect 3627 5683 3669 5692
rect 3628 5598 3668 5683
rect 3724 4976 3764 6196
rect 3820 6187 3860 6196
rect 3724 4927 3764 4936
rect 3916 4976 3956 4985
rect 4012 4976 4052 6784
rect 4352 6775 4720 6784
rect 4876 6749 4916 7120
rect 4972 7111 5012 7120
rect 4875 6740 4917 6749
rect 4875 6700 4876 6740
rect 4916 6700 4917 6740
rect 4875 6691 4917 6700
rect 4491 6572 4533 6581
rect 4491 6532 4492 6572
rect 4532 6532 4533 6572
rect 4491 6523 4533 6532
rect 4108 6488 4148 6497
rect 4108 5825 4148 6448
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 4492 6488 4532 6523
rect 4204 6354 4244 6439
rect 4492 6437 4532 6448
rect 4876 6488 4916 6691
rect 4876 6439 4916 6448
rect 5067 6488 5109 6497
rect 5452 6488 5492 12487
rect 5644 11705 5684 12496
rect 5835 12368 5877 12377
rect 5835 12328 5836 12368
rect 5876 12328 5877 12368
rect 5835 12319 5877 12328
rect 5836 12234 5876 12319
rect 6220 11705 6260 14008
rect 7372 11948 7412 15259
rect 7372 11899 7412 11908
rect 5643 11696 5685 11705
rect 5643 11656 5644 11696
rect 5684 11656 5685 11696
rect 5643 11647 5685 11656
rect 6219 11696 6261 11705
rect 6219 11656 6220 11696
rect 6260 11656 6261 11696
rect 6219 11647 6261 11656
rect 6028 10184 6068 10193
rect 6220 10184 6260 11647
rect 7372 11528 7412 11537
rect 7372 11033 7412 11488
rect 7371 11024 7413 11033
rect 7371 10984 7372 11024
rect 7412 10984 7413 11024
rect 7371 10975 7413 10984
rect 6068 10144 6260 10184
rect 7180 10268 7220 10277
rect 6028 8000 6068 10144
rect 7180 10025 7220 10228
rect 7179 10016 7221 10025
rect 7179 9976 7180 10016
rect 7220 9976 7221 10016
rect 7179 9967 7221 9976
rect 7468 9512 7508 24667
rect 30220 24464 30260 25264
rect 30987 25264 30988 25304
rect 31028 25264 31029 25304
rect 30987 25255 31029 25264
rect 30220 24415 30260 24424
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 28876 23960 28916 23969
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 28395 23120 28437 23129
rect 28395 23080 28396 23120
rect 28436 23080 28437 23120
rect 28395 23071 28437 23080
rect 28780 23120 28820 23129
rect 28876 23120 28916 23920
rect 29547 23960 29589 23969
rect 29547 23920 29548 23960
rect 29588 23920 29589 23960
rect 29547 23911 29589 23920
rect 30891 23960 30933 23969
rect 30891 23920 30892 23960
rect 30932 23920 30933 23960
rect 30891 23911 30933 23920
rect 29548 23213 29588 23911
rect 30892 23876 30932 23911
rect 30892 23825 30932 23836
rect 30988 23456 31028 25255
rect 31659 25136 31701 25145
rect 31659 25096 31660 25136
rect 31700 25096 31701 25136
rect 31659 25087 31701 25096
rect 31660 24632 31700 25087
rect 31276 23792 31316 23801
rect 31180 23752 31276 23792
rect 31083 23708 31125 23717
rect 31083 23668 31084 23708
rect 31124 23668 31125 23708
rect 31083 23659 31125 23668
rect 31084 23624 31124 23659
rect 31084 23573 31124 23584
rect 31180 23465 31220 23752
rect 31276 23743 31316 23752
rect 31468 23792 31508 23803
rect 31660 23801 31700 24592
rect 31756 24632 31796 25339
rect 32811 25304 32853 25313
rect 32811 25264 32812 25304
rect 32852 25264 32853 25304
rect 33292 25304 33332 25313
rect 32811 25255 32853 25264
rect 33100 25262 33140 25271
rect 32812 25170 32852 25255
rect 33003 25220 33045 25229
rect 33003 25180 33004 25220
rect 33044 25180 33045 25220
rect 33003 25171 33045 25180
rect 32139 25136 32181 25145
rect 32139 25096 32140 25136
rect 32180 25096 32181 25136
rect 32139 25087 32181 25096
rect 32140 25002 32180 25087
rect 31851 24884 31893 24893
rect 31851 24844 31852 24884
rect 31892 24844 31893 24884
rect 31851 24835 31893 24844
rect 31468 23717 31508 23752
rect 31564 23792 31604 23801
rect 31659 23792 31701 23801
rect 31604 23752 31660 23792
rect 31700 23752 31701 23792
rect 31564 23743 31604 23752
rect 31659 23743 31701 23752
rect 31467 23708 31509 23717
rect 31467 23668 31468 23708
rect 31508 23668 31509 23708
rect 31467 23659 31509 23668
rect 31660 23658 31700 23743
rect 31372 23624 31412 23633
rect 31276 23584 31372 23624
rect 31179 23456 31221 23465
rect 30988 23416 31124 23456
rect 28971 23204 29013 23213
rect 28971 23164 28972 23204
rect 29012 23164 29013 23204
rect 28971 23155 29013 23164
rect 29547 23204 29589 23213
rect 29547 23164 29548 23204
rect 29588 23164 29589 23204
rect 29547 23155 29589 23164
rect 28820 23080 28916 23120
rect 28780 23071 28820 23080
rect 28396 22986 28436 23071
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 28299 22532 28341 22541
rect 28299 22492 28300 22532
rect 28340 22492 28341 22532
rect 28299 22483 28341 22492
rect 27627 22448 27669 22457
rect 27627 22408 27628 22448
rect 27668 22408 27669 22448
rect 27627 22399 27669 22408
rect 27915 22448 27957 22457
rect 27915 22408 27916 22448
rect 27956 22408 27957 22448
rect 27915 22399 27957 22408
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 23211 21692 23253 21701
rect 23211 21652 23212 21692
rect 23252 21652 23253 21692
rect 23211 21643 23253 21652
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 23212 20852 23252 21643
rect 26668 21608 26708 21617
rect 27532 21608 27572 21617
rect 26708 21568 26900 21608
rect 26668 21559 26708 21568
rect 25516 21356 25556 21365
rect 23252 20812 23540 20852
rect 23212 20803 23252 20812
rect 22827 20600 22869 20609
rect 23020 20600 23060 20609
rect 22827 20560 22828 20600
rect 22868 20560 22869 20600
rect 22827 20551 22869 20560
rect 22924 20560 23020 20600
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 10828 20224 11060 20264
rect 10828 20021 10868 20224
rect 11020 20117 11060 20224
rect 10924 20096 10964 20105
rect 11020 20068 11060 20077
rect 11115 20096 11157 20105
rect 10827 20012 10869 20021
rect 10827 19972 10828 20012
rect 10868 19972 10869 20012
rect 10924 20012 10964 20056
rect 11115 20056 11116 20096
rect 11156 20056 11157 20096
rect 11115 20047 11157 20056
rect 11212 20096 11252 20105
rect 11404 20096 11444 20105
rect 11252 20056 11404 20096
rect 11212 20047 11252 20056
rect 11404 20047 11444 20056
rect 11596 20096 11636 20105
rect 10924 19972 11060 20012
rect 10827 19963 10869 19972
rect 9580 19928 9620 19937
rect 9580 19601 9620 19888
rect 9579 19592 9621 19601
rect 9579 19552 9580 19592
rect 9620 19552 9621 19592
rect 9579 19543 9621 19552
rect 10923 19592 10965 19601
rect 10923 19552 10924 19592
rect 10964 19552 10965 19592
rect 10923 19543 10965 19552
rect 10059 19256 10101 19265
rect 10059 19216 10060 19256
rect 10100 19216 10101 19256
rect 10059 19207 10101 19216
rect 10924 19256 10964 19543
rect 10924 19207 10964 19216
rect 10060 19122 10100 19207
rect 8908 19088 8948 19097
rect 8908 18761 8948 19048
rect 11020 18761 11060 19972
rect 11116 19962 11156 20047
rect 11404 19844 11444 19853
rect 11308 19256 11348 19265
rect 11404 19256 11444 19804
rect 11348 19216 11444 19256
rect 11596 19424 11636 20056
rect 11691 20096 11733 20105
rect 22540 20096 22580 20105
rect 11691 20056 11692 20096
rect 11732 20056 11733 20096
rect 11691 20047 11733 20056
rect 22156 20056 22540 20096
rect 11692 19962 11732 20047
rect 12748 19928 12788 19937
rect 12652 19888 12748 19928
rect 11596 19384 12020 19424
rect 11308 19207 11348 19216
rect 8907 18752 8949 18761
rect 8907 18712 8908 18752
rect 8948 18712 8949 18752
rect 8907 18703 8949 18712
rect 11019 18752 11061 18761
rect 11019 18712 11020 18752
rect 11060 18712 11061 18752
rect 11019 18703 11061 18712
rect 8619 15224 8661 15233
rect 8619 15184 8620 15224
rect 8660 15184 8661 15224
rect 8619 15175 8661 15184
rect 8620 14225 8660 15175
rect 8619 14216 8661 14225
rect 8619 14176 8620 14216
rect 8660 14176 8661 14216
rect 8619 14167 8661 14176
rect 7180 9472 7508 9512
rect 7180 8168 7220 9472
rect 7467 8504 7509 8513
rect 7467 8464 7468 8504
rect 7508 8464 7509 8504
rect 7467 8455 7509 8464
rect 7180 8119 7220 8128
rect 6028 7951 6068 7960
rect 7179 7748 7221 7757
rect 7179 7708 7180 7748
rect 7220 7708 7221 7748
rect 7179 7699 7221 7708
rect 7180 7614 7220 7699
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5164 6448 5492 6488
rect 7371 6488 7413 6497
rect 7371 6448 7372 6488
rect 7412 6448 7413 6488
rect 5068 6354 5108 6439
rect 4972 6236 5012 6245
rect 4876 6196 4972 6236
rect 4107 5816 4149 5825
rect 4107 5776 4108 5816
rect 4148 5776 4149 5816
rect 4107 5767 4149 5776
rect 4107 5648 4149 5657
rect 4107 5608 4108 5648
rect 4148 5608 4149 5648
rect 4107 5599 4149 5608
rect 3956 4936 4052 4976
rect 3916 4927 3956 4936
rect 3819 4808 3861 4817
rect 3819 4768 3820 4808
rect 3860 4768 3861 4808
rect 3819 4759 3861 4768
rect 3820 4674 3860 4759
rect 3532 4087 3572 4096
rect 3820 4136 3860 4147
rect 3916 4145 3956 4176
rect 3820 4061 3860 4096
rect 3915 4136 3957 4145
rect 3915 4096 3916 4136
rect 3956 4096 3957 4136
rect 3915 4087 3957 4096
rect 2956 4012 3006 4052
rect 3819 4052 3861 4061
rect 3819 4012 3820 4052
rect 3860 4012 3861 4052
rect 2956 3968 2996 4012
rect 3819 4003 3861 4012
rect 3916 4052 3956 4087
rect 2764 3928 2996 3968
rect 2572 3844 2804 3884
rect 2668 3464 2708 3473
rect 2476 3424 2668 3464
rect 2668 3415 2708 3424
rect 2380 2575 2420 2584
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2668 2624 2708 2633
rect 2764 2624 2804 3844
rect 2956 3473 2996 3928
rect 3820 3632 3860 3641
rect 3916 3632 3956 4012
rect 4012 3641 4052 4936
rect 4108 4976 4148 5599
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4108 4927 4148 4936
rect 4779 4808 4821 4817
rect 4779 4768 4780 4808
rect 4820 4768 4821 4808
rect 4779 4759 4821 4768
rect 4204 4304 4244 4313
rect 3860 3592 3956 3632
rect 4011 3632 4053 3641
rect 4011 3592 4012 3632
rect 4052 3592 4053 3632
rect 3820 3583 3860 3592
rect 4011 3583 4053 3592
rect 2955 3464 2997 3473
rect 2955 3424 2956 3464
rect 2996 3424 2997 3464
rect 2955 3415 2997 3424
rect 4204 3464 4244 4264
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4780 4136 4820 4759
rect 4780 4087 4820 4096
rect 4876 4136 4916 6196
rect 4972 6187 5012 6196
rect 4876 4087 4916 4096
rect 4972 5564 5012 5573
rect 4588 4002 4628 4087
rect 4684 3968 4724 3977
rect 4972 3968 5012 5524
rect 5068 4976 5108 4985
rect 5164 4976 5204 6448
rect 7371 6439 7413 6448
rect 5452 6320 5492 6329
rect 5356 6280 5452 6320
rect 5356 5648 5396 6280
rect 5452 6271 5492 6280
rect 7372 5900 7412 6439
rect 7372 5851 7412 5860
rect 5356 5599 5396 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6356 5648
rect 6219 5599 6261 5608
rect 6220 5514 6260 5599
rect 5108 4936 5204 4976
rect 5068 4927 5108 4936
rect 5548 4808 5588 4817
rect 5452 4768 5548 4808
rect 5452 4136 5492 4768
rect 5548 4759 5588 4768
rect 5452 4087 5492 4096
rect 6316 4136 6356 5608
rect 7371 5480 7413 5489
rect 7371 5440 7372 5480
rect 7412 5440 7413 5480
rect 7371 5431 7413 5440
rect 7372 5346 7412 5431
rect 6316 4087 6356 4096
rect 7468 4304 7508 8455
rect 4724 3928 5012 3968
rect 5068 4052 5108 4061
rect 4684 3919 4724 3928
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 5068 3716 5108 4012
rect 5259 4052 5301 4061
rect 5259 4012 5260 4052
rect 5300 4012 5301 4052
rect 5259 4003 5301 4012
rect 4972 3676 5108 3716
rect 4395 3632 4437 3641
rect 4395 3592 4396 3632
rect 4436 3592 4437 3632
rect 4395 3583 4437 3592
rect 4684 3632 4724 3641
rect 4972 3632 5012 3676
rect 4724 3592 5012 3632
rect 4684 3583 4724 3592
rect 4204 3415 4244 3424
rect 4396 3464 4436 3583
rect 5068 3473 5108 3558
rect 5260 3473 5300 4003
rect 7468 3473 7508 4264
rect 4780 3464 4820 3473
rect 4396 3415 4436 3424
rect 4588 3453 4628 3462
rect 2860 2624 2900 2633
rect 2764 2584 2860 2624
rect 2956 2624 2996 3415
rect 4588 3305 4628 3413
rect 4587 3296 4629 3305
rect 4587 3256 4588 3296
rect 4628 3256 4629 3296
rect 4587 3247 4629 3256
rect 4300 3212 4340 3221
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 3147 2708 3189 2717
rect 3147 2668 3148 2708
rect 3188 2668 3189 2708
rect 3147 2659 3189 2668
rect 3052 2624 3092 2633
rect 2956 2584 3052 2624
rect 1419 2540 1461 2549
rect 1419 2500 1420 2540
rect 1460 2500 1461 2540
rect 1419 2491 1461 2500
rect 2475 2540 2517 2549
rect 2475 2500 2476 2540
rect 2516 2500 2517 2540
rect 2475 2491 2517 2500
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 2476 2406 2516 2491
rect 2572 2490 2612 2575
rect 2668 2456 2708 2584
rect 2860 2575 2900 2584
rect 3052 2575 3092 2584
rect 3148 2624 3188 2659
rect 4300 2633 4340 3172
rect 4780 2633 4820 3424
rect 4876 3464 4916 3473
rect 4876 3296 4916 3424
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 5259 3464 5301 3473
rect 5259 3424 5260 3464
rect 5300 3424 5301 3464
rect 5259 3415 5301 3424
rect 7467 3464 7509 3473
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 5260 3330 5300 3415
rect 5164 3296 5204 3305
rect 4876 3256 5164 3296
rect 5164 3247 5204 3256
rect 8908 2717 8948 18703
rect 11020 18668 11060 18703
rect 11020 18617 11060 18628
rect 11596 18668 11636 19384
rect 11596 18619 11636 18628
rect 11788 19256 11828 19265
rect 10636 18584 10676 18593
rect 10636 16577 10676 18544
rect 10924 18584 10964 18595
rect 10924 18509 10964 18544
rect 11500 18584 11540 18593
rect 10923 18500 10965 18509
rect 10923 18460 10924 18500
rect 10964 18460 10965 18500
rect 10923 18451 10965 18460
rect 11308 18416 11348 18425
rect 11500 18416 11540 18544
rect 11348 18376 11540 18416
rect 11692 18584 11732 18593
rect 11308 18367 11348 18376
rect 10635 16568 10677 16577
rect 10635 16528 10636 16568
rect 10676 16528 10677 16568
rect 10635 16519 10677 16528
rect 11692 16073 11732 18544
rect 11788 16661 11828 19216
rect 11980 19256 12020 19384
rect 11980 19207 12020 19216
rect 12076 19256 12116 19265
rect 12652 19256 12692 19888
rect 12748 19879 12788 19888
rect 21771 19844 21813 19853
rect 21771 19804 21772 19844
rect 21812 19804 21813 19844
rect 21771 19795 21813 19804
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 14667 19508 14709 19517
rect 14667 19468 14668 19508
rect 14708 19468 14709 19508
rect 14667 19459 14709 19468
rect 14668 19374 14708 19459
rect 21772 19349 21812 19795
rect 21771 19340 21813 19349
rect 21771 19300 21772 19340
rect 21812 19300 21813 19340
rect 21771 19291 21813 19300
rect 12116 19216 12212 19256
rect 12076 19207 12116 19216
rect 11883 19172 11925 19181
rect 11883 19132 11884 19172
rect 11924 19132 11925 19172
rect 11883 19123 11925 19132
rect 11884 19038 11924 19123
rect 12075 18668 12117 18677
rect 12075 18628 12076 18668
rect 12116 18628 12117 18668
rect 12075 18619 12117 18628
rect 12172 18668 12212 19216
rect 12652 19207 12692 19216
rect 13515 19256 13557 19265
rect 13515 19216 13516 19256
rect 13556 19216 13557 19256
rect 13515 19207 13557 19216
rect 12267 19172 12309 19181
rect 12267 19132 12268 19172
rect 12308 19132 12309 19172
rect 12267 19123 12309 19132
rect 12268 19038 12308 19123
rect 13516 19122 13556 19207
rect 21772 19206 21812 19291
rect 22156 19256 22196 20056
rect 22540 20047 22580 20056
rect 22732 20096 22772 20105
rect 22540 19844 22580 19853
rect 22156 19207 22196 19216
rect 22252 19256 22292 19265
rect 14668 19088 14708 19097
rect 12172 18619 12212 18628
rect 12076 18584 12116 18619
rect 12076 18533 12116 18544
rect 12268 18584 12308 18595
rect 12268 18509 12308 18544
rect 14668 18509 14708 19048
rect 21964 19088 22004 19099
rect 21964 19013 22004 19048
rect 22252 19013 22292 19216
rect 22348 19256 22388 19267
rect 22348 19181 22388 19216
rect 22444 19256 22484 19265
rect 22540 19256 22580 19804
rect 22636 19256 22676 19265
rect 22540 19216 22636 19256
rect 22347 19172 22389 19181
rect 22347 19132 22348 19172
rect 22388 19132 22389 19172
rect 22347 19123 22389 19132
rect 21963 19004 22005 19013
rect 21963 18964 21964 19004
rect 22004 18964 22005 19004
rect 21963 18955 22005 18964
rect 22251 19004 22293 19013
rect 22251 18964 22252 19004
rect 22292 18964 22293 19004
rect 22251 18955 22293 18964
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 22444 18761 22484 19216
rect 22636 19207 22676 19216
rect 22539 19088 22581 19097
rect 22539 19048 22540 19088
rect 22580 19048 22581 19088
rect 22539 19039 22581 19048
rect 22443 18752 22485 18761
rect 22443 18712 22444 18752
rect 22484 18712 22485 18752
rect 22443 18703 22485 18712
rect 22540 18752 22580 19039
rect 22540 18703 22580 18712
rect 22155 18584 22197 18593
rect 22155 18544 22156 18584
rect 22196 18544 22197 18584
rect 22155 18535 22197 18544
rect 12267 18500 12309 18509
rect 12267 18460 12268 18500
rect 12308 18460 12309 18500
rect 12267 18451 12309 18460
rect 14667 18500 14709 18509
rect 14667 18460 14668 18500
rect 14708 18460 14709 18500
rect 14667 18451 14709 18460
rect 21964 18500 22004 18509
rect 21964 18341 22004 18460
rect 22156 18416 22196 18535
rect 22347 18500 22389 18509
rect 22347 18460 22348 18500
rect 22388 18460 22389 18500
rect 22732 18500 22772 20056
rect 22828 20096 22868 20551
rect 22828 20047 22868 20056
rect 22732 18460 22868 18500
rect 22347 18451 22389 18460
rect 22156 18367 22196 18376
rect 22348 18366 22388 18451
rect 21963 18332 22005 18341
rect 22732 18332 22772 18341
rect 21963 18292 21964 18332
rect 22004 18292 22005 18332
rect 21963 18283 22005 18292
rect 22636 18292 22732 18332
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 21964 17417 22004 18283
rect 22636 17996 22676 18292
rect 22732 18283 22772 18292
rect 22540 17956 22676 17996
rect 22540 17744 22580 17956
rect 22828 17912 22868 18460
rect 22924 18341 22964 20560
rect 23020 20532 23060 20560
rect 23500 20264 23540 20812
rect 23500 20215 23540 20224
rect 25516 20189 25556 21316
rect 26187 20936 26229 20945
rect 26187 20896 26188 20936
rect 26228 20896 26229 20936
rect 26187 20887 26229 20896
rect 25899 20852 25941 20861
rect 25899 20812 25900 20852
rect 25940 20812 25941 20852
rect 25899 20803 25941 20812
rect 25515 20180 25557 20189
rect 25515 20140 25516 20180
rect 25556 20140 25557 20180
rect 25515 20131 25557 20140
rect 23692 20012 23732 20021
rect 23116 19928 23156 19937
rect 23116 19592 23156 19888
rect 23692 19853 23732 19972
rect 23499 19844 23541 19853
rect 23499 19804 23500 19844
rect 23540 19804 23541 19844
rect 23499 19795 23541 19804
rect 23691 19844 23733 19853
rect 23691 19804 23692 19844
rect 23732 19804 23733 19844
rect 23691 19795 23733 19804
rect 23020 19552 23156 19592
rect 23020 19292 23060 19552
rect 23020 19243 23060 19252
rect 23019 18752 23061 18761
rect 23019 18712 23020 18752
rect 23060 18712 23061 18752
rect 23019 18703 23061 18712
rect 23020 18668 23060 18703
rect 23020 18617 23060 18628
rect 23116 18584 23156 18593
rect 22923 18332 22965 18341
rect 22923 18292 22924 18332
rect 22964 18292 22965 18332
rect 22923 18283 22965 18292
rect 22636 17872 23060 17912
rect 22636 17828 22676 17872
rect 22636 17779 22676 17788
rect 23020 17758 23060 17872
rect 22540 17695 22580 17704
rect 22731 17744 22773 17753
rect 22731 17704 22732 17744
rect 22772 17704 22773 17744
rect 22731 17695 22773 17704
rect 22923 17744 22965 17753
rect 22923 17704 22924 17744
rect 22964 17704 22965 17744
rect 23020 17709 23060 17718
rect 22923 17695 22965 17704
rect 22732 17610 22772 17695
rect 22924 17610 22964 17695
rect 23116 17585 23156 18544
rect 23403 18584 23445 18593
rect 23403 18544 23404 18584
rect 23444 18544 23445 18584
rect 23403 18535 23445 18544
rect 23404 18450 23444 18535
rect 23212 17912 23252 17921
rect 23252 17872 23444 17912
rect 23212 17863 23252 17872
rect 23212 17744 23252 17753
rect 23212 17669 23252 17704
rect 23404 17744 23444 17872
rect 23404 17695 23444 17704
rect 23211 17660 23253 17669
rect 23211 17620 23212 17660
rect 23252 17620 23253 17660
rect 23211 17611 23253 17620
rect 23115 17576 23157 17585
rect 23115 17536 23116 17576
rect 23156 17536 23157 17576
rect 23115 17527 23157 17536
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 21963 17408 22005 17417
rect 21963 17368 21964 17408
rect 22004 17368 22005 17408
rect 21963 17359 22005 17368
rect 23212 17240 23252 17611
rect 23212 17191 23252 17200
rect 23500 17165 23540 19795
rect 25900 19424 25940 20803
rect 26188 20802 26228 20887
rect 26379 20852 26421 20861
rect 26764 20852 26804 20861
rect 26379 20812 26380 20852
rect 26420 20812 26421 20852
rect 26379 20803 26421 20812
rect 26476 20812 26764 20852
rect 26380 20718 26420 20803
rect 26476 20264 26516 20812
rect 26764 20803 26804 20812
rect 25612 19384 25940 19424
rect 26092 20224 26516 20264
rect 26572 20600 26612 20609
rect 23884 19256 23924 19265
rect 25228 19256 25268 19265
rect 23924 19216 24020 19256
rect 23884 19207 23924 19216
rect 23691 18500 23733 18509
rect 23691 18460 23692 18500
rect 23732 18460 23733 18500
rect 23691 18451 23733 18460
rect 23692 18366 23732 18451
rect 23980 18341 24020 19216
rect 25036 19088 25076 19097
rect 25228 19088 25268 19216
rect 25076 19048 25268 19088
rect 25324 19256 25364 19265
rect 24459 18920 24501 18929
rect 24459 18880 24460 18920
rect 24500 18880 24501 18920
rect 24459 18871 24501 18880
rect 24076 18500 24116 18509
rect 23884 18332 23924 18341
rect 23884 18173 23924 18292
rect 23979 18332 24021 18341
rect 23979 18292 23980 18332
rect 24020 18292 24021 18332
rect 23979 18283 24021 18292
rect 24076 18173 24116 18460
rect 24460 18500 24500 18871
rect 25036 18761 25076 19048
rect 25035 18752 25077 18761
rect 25035 18712 25036 18752
rect 25076 18712 25077 18752
rect 25035 18703 25077 18712
rect 24843 18668 24885 18677
rect 24843 18628 24844 18668
rect 24884 18628 24885 18668
rect 24843 18619 24885 18628
rect 24844 18509 24884 18619
rect 24268 18332 24308 18343
rect 24268 18257 24308 18292
rect 24267 18248 24309 18257
rect 24267 18208 24268 18248
rect 24308 18208 24309 18248
rect 24267 18199 24309 18208
rect 23883 18164 23925 18173
rect 23883 18124 23884 18164
rect 23924 18124 23925 18164
rect 23883 18115 23925 18124
rect 24075 18164 24117 18173
rect 24075 18124 24076 18164
rect 24116 18124 24117 18164
rect 24075 18115 24117 18124
rect 24268 17837 24308 18199
rect 24267 17828 24309 17837
rect 24267 17788 24268 17828
rect 24308 17788 24309 17828
rect 24267 17779 24309 17788
rect 23691 17744 23733 17753
rect 23691 17704 23692 17744
rect 23732 17704 23733 17744
rect 23691 17695 23733 17704
rect 23788 17744 23828 17753
rect 23828 17704 24020 17744
rect 23788 17695 23828 17704
rect 23595 17576 23637 17585
rect 23595 17536 23596 17576
rect 23636 17536 23637 17576
rect 23595 17527 23637 17536
rect 23499 17156 23541 17165
rect 23499 17116 23500 17156
rect 23540 17116 23541 17156
rect 23499 17107 23541 17116
rect 23596 17072 23636 17527
rect 23692 17156 23732 17695
rect 23787 17492 23829 17501
rect 23787 17452 23788 17492
rect 23828 17452 23829 17492
rect 23787 17443 23829 17452
rect 23692 17107 23732 17116
rect 23596 17023 23636 17032
rect 23788 17072 23828 17443
rect 23788 17023 23828 17032
rect 23403 16988 23445 16997
rect 23403 16948 23404 16988
rect 23444 16948 23445 16988
rect 23403 16939 23445 16948
rect 23404 16854 23444 16939
rect 23980 16904 24020 17704
rect 23980 16855 24020 16864
rect 11787 16652 11829 16661
rect 11787 16612 11788 16652
rect 11828 16612 11829 16652
rect 11787 16603 11829 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 24460 16325 24500 18460
rect 24843 18500 24885 18509
rect 24843 18460 24844 18500
rect 24884 18460 24885 18500
rect 24843 18451 24885 18460
rect 24844 18366 24884 18451
rect 24652 18332 24692 18341
rect 24556 18292 24652 18332
rect 24556 18089 24596 18292
rect 24652 18283 24692 18292
rect 24747 18332 24789 18341
rect 24747 18292 24748 18332
rect 24788 18292 24789 18332
rect 24747 18283 24789 18292
rect 25036 18332 25076 18341
rect 25324 18332 25364 19216
rect 25516 19256 25556 19265
rect 25419 19088 25461 19097
rect 25419 19048 25420 19088
rect 25460 19048 25461 19088
rect 25419 19039 25461 19048
rect 25420 18954 25460 19039
rect 25516 18425 25556 19216
rect 25612 18500 25652 19384
rect 25804 19256 25844 19265
rect 25708 19088 25748 19097
rect 25708 18761 25748 19048
rect 25804 19013 25844 19216
rect 25900 19256 25940 19267
rect 25900 19181 25940 19216
rect 25996 19256 26036 19265
rect 25899 19172 25941 19181
rect 25899 19132 25900 19172
rect 25940 19132 25941 19172
rect 25899 19123 25941 19132
rect 25803 19004 25845 19013
rect 25803 18964 25804 19004
rect 25844 18964 25845 19004
rect 25803 18955 25845 18964
rect 25996 18845 26036 19216
rect 25995 18836 26037 18845
rect 25995 18796 25996 18836
rect 26036 18796 26037 18836
rect 25995 18787 26037 18796
rect 25707 18752 25749 18761
rect 25707 18712 25708 18752
rect 25748 18712 25749 18752
rect 25707 18703 25749 18712
rect 26092 18509 26132 20224
rect 26476 20096 26516 20124
rect 26572 20105 26612 20560
rect 26667 20600 26709 20609
rect 26667 20560 26668 20600
rect 26708 20560 26709 20600
rect 26667 20551 26709 20560
rect 26571 20096 26613 20105
rect 26516 20056 26572 20096
rect 26612 20056 26613 20096
rect 26476 20047 26516 20056
rect 26571 20047 26613 20056
rect 26668 20096 26708 20551
rect 26763 20180 26805 20189
rect 26763 20140 26764 20180
rect 26804 20140 26805 20180
rect 26763 20131 26805 20140
rect 26668 20047 26708 20056
rect 26764 20096 26804 20131
rect 26764 20045 26804 20056
rect 26379 19928 26421 19937
rect 26476 19928 26516 19937
rect 26379 19888 26380 19928
rect 26420 19888 26476 19928
rect 26379 19879 26421 19888
rect 26476 19879 26516 19888
rect 26571 19928 26613 19937
rect 26571 19888 26572 19928
rect 26612 19888 26613 19928
rect 26571 19879 26613 19888
rect 26572 19256 26612 19879
rect 26860 19256 26900 21568
rect 26955 21524 26997 21533
rect 26955 21484 26956 21524
rect 26996 21484 26997 21524
rect 26955 21475 26997 21484
rect 26956 21020 26996 21475
rect 27147 21440 27189 21449
rect 27147 21400 27148 21440
rect 27188 21400 27189 21440
rect 27147 21391 27189 21400
rect 26956 20971 26996 20980
rect 27148 20861 27188 21391
rect 27532 20945 27572 21568
rect 27531 20936 27573 20945
rect 27531 20896 27532 20936
rect 27572 20896 27573 20936
rect 27531 20887 27573 20896
rect 27147 20852 27189 20861
rect 27147 20812 27148 20852
rect 27188 20812 27189 20852
rect 27147 20803 27189 20812
rect 27148 20718 27188 20803
rect 27628 20777 27668 22399
rect 27723 22364 27765 22373
rect 27723 22324 27724 22364
rect 27764 22324 27765 22364
rect 27723 22315 27765 22324
rect 27724 22230 27764 22315
rect 27916 22314 27956 22399
rect 28300 22398 28340 22483
rect 28108 22364 28148 22373
rect 28012 22324 28108 22364
rect 28012 21776 28052 22324
rect 28108 22315 28148 22324
rect 28203 22364 28245 22373
rect 28972 22364 29012 23155
rect 29548 22952 29588 23155
rect 29644 23120 29684 23129
rect 30988 23120 31028 23129
rect 29684 23080 29972 23120
rect 29644 23071 29684 23080
rect 29548 22912 29780 22952
rect 28203 22324 28204 22364
rect 28244 22324 28245 22364
rect 28203 22315 28245 22324
rect 28876 22324 29012 22364
rect 27724 21736 28052 21776
rect 27339 20768 27381 20777
rect 27339 20728 27340 20768
rect 27380 20728 27381 20768
rect 27339 20719 27381 20728
rect 27627 20768 27669 20777
rect 27627 20728 27628 20768
rect 27668 20728 27669 20768
rect 27627 20719 27669 20728
rect 27340 20609 27380 20719
rect 26955 20600 26997 20609
rect 26955 20560 26956 20600
rect 26996 20560 26997 20600
rect 26955 20551 26997 20560
rect 27339 20600 27381 20609
rect 27339 20560 27340 20600
rect 27380 20560 27381 20600
rect 27339 20551 27381 20560
rect 26956 20466 26996 20551
rect 27340 20466 27380 20551
rect 26955 19928 26997 19937
rect 26955 19888 26956 19928
rect 26996 19888 26997 19928
rect 26955 19879 26997 19888
rect 26956 19794 26996 19879
rect 27724 19349 27764 21736
rect 28204 21701 28244 22315
rect 28491 22280 28533 22289
rect 28491 22240 28492 22280
rect 28532 22240 28533 22280
rect 28491 22231 28533 22240
rect 28684 22280 28724 22289
rect 28876 22280 28916 22324
rect 28724 22240 28820 22280
rect 28684 22231 28724 22240
rect 28492 22146 28532 22231
rect 28588 22196 28628 22205
rect 28300 22112 28340 22121
rect 28203 21692 28245 21701
rect 28203 21652 28204 21692
rect 28244 21652 28245 21692
rect 28203 21643 28245 21652
rect 27819 21608 27861 21617
rect 27819 21568 27820 21608
rect 27860 21568 27861 21608
rect 27819 21559 27861 21568
rect 27916 21608 27956 21617
rect 28204 21608 28244 21643
rect 27956 21568 28148 21608
rect 27916 21559 27956 21568
rect 27820 20768 27860 21559
rect 28011 21188 28053 21197
rect 28011 21148 28012 21188
rect 28052 21148 28053 21188
rect 28011 21139 28053 21148
rect 27820 20189 27860 20728
rect 27915 20768 27957 20777
rect 27915 20728 27916 20768
rect 27956 20728 27957 20768
rect 27915 20719 27957 20728
rect 28012 20768 28052 21139
rect 28108 21020 28148 21568
rect 28204 21558 28244 21568
rect 28300 21197 28340 22072
rect 28588 21776 28628 22156
rect 28683 22112 28725 22121
rect 28683 22072 28684 22112
rect 28724 22072 28725 22112
rect 28683 22063 28725 22072
rect 28396 21736 28628 21776
rect 28299 21188 28341 21197
rect 28299 21148 28300 21188
rect 28340 21148 28341 21188
rect 28299 21139 28341 21148
rect 28300 21020 28340 21029
rect 28108 20980 28300 21020
rect 28300 20971 28340 20980
rect 28012 20719 28052 20728
rect 28108 20768 28148 20777
rect 28300 20768 28340 20777
rect 28148 20728 28300 20768
rect 28396 20768 28436 21736
rect 28492 21608 28532 21617
rect 28492 21449 28532 21568
rect 28587 21608 28629 21617
rect 28587 21568 28588 21608
rect 28628 21568 28629 21608
rect 28587 21559 28629 21568
rect 28588 21474 28628 21559
rect 28491 21440 28533 21449
rect 28491 21400 28492 21440
rect 28532 21400 28533 21440
rect 28491 21391 28533 21400
rect 28491 20768 28533 20777
rect 28396 20728 28492 20768
rect 28532 20728 28533 20768
rect 28108 20719 28148 20728
rect 28300 20719 28340 20728
rect 28491 20719 28533 20728
rect 28588 20768 28628 20777
rect 28684 20768 28724 22063
rect 28780 21440 28820 22240
rect 28876 21617 28916 22240
rect 29068 22280 29108 22289
rect 28972 22196 29012 22205
rect 28875 21608 28917 21617
rect 28875 21568 28876 21608
rect 28916 21568 28917 21608
rect 28875 21559 28917 21568
rect 28876 21440 28916 21449
rect 28780 21400 28876 21440
rect 28876 21391 28916 21400
rect 28972 21272 29012 22156
rect 29068 21785 29108 22240
rect 29548 22280 29588 22289
rect 29067 21776 29109 21785
rect 29067 21736 29068 21776
rect 29108 21736 29109 21776
rect 29067 21727 29109 21736
rect 29356 21608 29396 21617
rect 28628 20728 28724 20768
rect 28780 21232 29012 21272
rect 29068 21568 29356 21608
rect 28780 20768 28820 21232
rect 29068 21020 29108 21568
rect 29356 21559 29396 21568
rect 29451 21608 29493 21617
rect 29451 21568 29452 21608
rect 29492 21568 29493 21608
rect 29451 21559 29493 21568
rect 29068 20971 29108 20980
rect 28971 20852 29013 20861
rect 28971 20812 28972 20852
rect 29012 20812 29013 20852
rect 28971 20803 29013 20812
rect 28588 20719 28628 20728
rect 28780 20719 28820 20728
rect 28875 20768 28917 20777
rect 28875 20728 28876 20768
rect 28916 20728 28917 20768
rect 28875 20719 28917 20728
rect 27916 20634 27956 20719
rect 28492 20634 28532 20719
rect 28876 20634 28916 20719
rect 27819 20180 27861 20189
rect 27819 20140 27820 20180
rect 27860 20140 27861 20180
rect 27819 20131 27861 20140
rect 28972 19853 29012 20803
rect 29068 20768 29108 20777
rect 29452 20768 29492 21559
rect 29108 20728 29492 20768
rect 29068 20719 29108 20728
rect 28971 19844 29013 19853
rect 28971 19804 28972 19844
rect 29012 19804 29013 19844
rect 28971 19795 29013 19804
rect 29068 19433 29108 19518
rect 29067 19424 29109 19433
rect 29067 19384 29068 19424
rect 29108 19384 29109 19424
rect 29067 19375 29109 19384
rect 29259 19424 29301 19433
rect 29259 19384 29260 19424
rect 29300 19384 29301 19424
rect 29259 19375 29301 19384
rect 27723 19340 27765 19349
rect 27723 19300 27724 19340
rect 27764 19300 27765 19340
rect 27723 19291 27765 19300
rect 27436 19256 27476 19265
rect 26860 19216 27436 19256
rect 26572 19207 26612 19216
rect 26188 19172 26228 19181
rect 26228 19132 26324 19172
rect 26188 19123 26228 19132
rect 26187 18752 26229 18761
rect 26187 18712 26188 18752
rect 26228 18712 26229 18752
rect 26187 18703 26229 18712
rect 26284 18752 26324 19132
rect 26475 19088 26517 19097
rect 26475 19048 26476 19088
rect 26516 19048 26517 19088
rect 26475 19039 26517 19048
rect 26284 18703 26324 18712
rect 26188 18584 26228 18703
rect 26188 18535 26228 18544
rect 26379 18584 26421 18593
rect 26379 18544 26380 18584
rect 26420 18544 26421 18584
rect 26379 18535 26421 18544
rect 26476 18584 26516 19039
rect 27243 18836 27285 18845
rect 27243 18796 27244 18836
rect 27284 18796 27285 18836
rect 27243 18787 27285 18796
rect 26859 18668 26901 18677
rect 26859 18628 26860 18668
rect 26900 18628 26901 18668
rect 26859 18619 26901 18628
rect 27244 18668 27284 18787
rect 27244 18619 27284 18628
rect 26476 18535 26516 18544
rect 26763 18584 26805 18593
rect 26763 18544 26764 18584
rect 26804 18544 26805 18584
rect 26763 18535 26805 18544
rect 26860 18584 26900 18619
rect 25708 18500 25748 18509
rect 25612 18460 25708 18500
rect 25708 18451 25748 18460
rect 26091 18500 26133 18509
rect 26091 18460 26092 18500
rect 26132 18460 26133 18500
rect 26091 18451 26133 18460
rect 26380 18450 26420 18535
rect 25515 18416 25557 18425
rect 25515 18376 25516 18416
rect 25556 18376 25557 18416
rect 25515 18367 25557 18376
rect 25076 18292 25364 18332
rect 25036 18283 25076 18292
rect 24555 18080 24597 18089
rect 24555 18040 24556 18080
rect 24596 18040 24597 18080
rect 24555 18031 24597 18040
rect 24556 16997 24596 18031
rect 24652 17744 24692 17753
rect 24748 17744 24788 18283
rect 24692 17704 24788 17744
rect 24652 17695 24692 17704
rect 25324 17501 25364 18292
rect 25516 18282 25556 18367
rect 26668 17744 26708 17755
rect 26764 17744 26804 18535
rect 26860 18533 26900 18544
rect 27148 18584 27188 18593
rect 27148 17912 27188 18544
rect 27436 18341 27476 19216
rect 28780 19256 28820 19265
rect 28588 19088 28628 19097
rect 28588 18845 28628 19048
rect 28587 18836 28629 18845
rect 28587 18796 28588 18836
rect 28628 18796 28724 18836
rect 28587 18787 28629 18796
rect 27724 18584 27764 18593
rect 27532 18416 27572 18425
rect 27724 18416 27764 18544
rect 27819 18584 27861 18593
rect 27819 18544 27820 18584
rect 27860 18544 27861 18584
rect 27819 18535 27861 18544
rect 27916 18584 27956 18593
rect 27820 18450 27860 18535
rect 27572 18376 27764 18416
rect 27532 18367 27572 18376
rect 27435 18332 27477 18341
rect 27435 18292 27436 18332
rect 27476 18292 27477 18332
rect 27435 18283 27477 18292
rect 27916 18257 27956 18544
rect 28684 18584 28724 18796
rect 28780 18752 28820 19216
rect 28876 19256 28916 19265
rect 29068 19256 29108 19267
rect 28916 19216 29012 19256
rect 28876 19207 28916 19216
rect 28972 18761 29012 19216
rect 29068 19181 29108 19216
rect 29260 19256 29300 19375
rect 29260 19207 29300 19216
rect 29067 19172 29109 19181
rect 29067 19132 29068 19172
rect 29108 19132 29109 19172
rect 29067 19123 29109 19132
rect 28971 18752 29013 18761
rect 28780 18712 28916 18752
rect 28876 18668 28916 18712
rect 28971 18712 28972 18752
rect 29012 18712 29013 18752
rect 28971 18703 29013 18712
rect 28876 18619 28916 18628
rect 28684 18535 28724 18544
rect 28780 18584 28820 18593
rect 28395 18332 28437 18341
rect 28395 18292 28396 18332
rect 28436 18292 28437 18332
rect 28395 18283 28437 18292
rect 27915 18248 27957 18257
rect 27915 18208 27916 18248
rect 27956 18208 27957 18248
rect 27915 18199 27957 18208
rect 27148 17872 27476 17912
rect 26956 17788 27380 17828
rect 26860 17744 26900 17753
rect 26764 17704 26860 17744
rect 26668 17669 26708 17704
rect 26860 17695 26900 17704
rect 26956 17744 26996 17788
rect 26956 17695 26996 17704
rect 26667 17660 26709 17669
rect 26667 17620 26668 17660
rect 26708 17620 26709 17660
rect 26667 17611 26709 17620
rect 27148 17660 27188 17669
rect 25803 17576 25845 17585
rect 25803 17536 25804 17576
rect 25844 17536 25845 17576
rect 25803 17527 25845 17536
rect 26764 17576 26804 17585
rect 27148 17576 27188 17620
rect 26804 17536 27188 17576
rect 26764 17527 26804 17536
rect 25323 17492 25365 17501
rect 25323 17452 25324 17492
rect 25364 17452 25365 17492
rect 25323 17443 25365 17452
rect 25804 17442 25844 17527
rect 27243 17492 27285 17501
rect 27243 17452 27244 17492
rect 27284 17452 27285 17492
rect 27243 17443 27285 17452
rect 27244 17072 27284 17443
rect 27340 17156 27380 17788
rect 27436 17585 27476 17872
rect 27532 17744 27572 17753
rect 27435 17576 27477 17585
rect 27435 17536 27436 17576
rect 27476 17536 27477 17576
rect 27435 17527 27477 17536
rect 27340 17107 27380 17116
rect 27244 17023 27284 17032
rect 27436 17072 27476 17527
rect 27436 17023 27476 17032
rect 24555 16988 24597 16997
rect 24555 16948 24556 16988
rect 24596 16948 24597 16988
rect 24555 16939 24597 16948
rect 27532 16904 27572 17704
rect 28396 17744 28436 18283
rect 28396 17695 28436 17704
rect 28780 17501 28820 18544
rect 28972 18584 29012 18595
rect 28972 18509 29012 18544
rect 28971 18500 29013 18509
rect 28971 18460 28972 18500
rect 29012 18460 29013 18500
rect 28971 18451 29013 18460
rect 29356 18089 29396 20728
rect 29548 20105 29588 22240
rect 29740 22280 29780 22912
rect 29740 22231 29780 22240
rect 29835 22280 29877 22289
rect 29835 22240 29836 22280
rect 29876 22240 29877 22280
rect 29835 22231 29877 22240
rect 29836 22146 29876 22231
rect 29643 22112 29685 22121
rect 29643 22072 29644 22112
rect 29684 22072 29685 22112
rect 29643 22063 29685 22072
rect 29644 21978 29684 22063
rect 29740 21608 29780 21617
rect 29932 21608 29972 23080
rect 30892 23080 30988 23120
rect 30796 22868 30836 22877
rect 30604 22828 30796 22868
rect 30604 22289 30644 22828
rect 30796 22819 30836 22828
rect 30795 22532 30837 22541
rect 30795 22492 30796 22532
rect 30836 22492 30837 22532
rect 30795 22483 30837 22492
rect 30699 22448 30741 22457
rect 30699 22408 30700 22448
rect 30740 22408 30741 22448
rect 30699 22399 30741 22408
rect 30603 22280 30645 22289
rect 30603 22240 30604 22280
rect 30644 22240 30645 22280
rect 30603 22231 30645 22240
rect 30700 22280 30740 22399
rect 30700 22231 30740 22240
rect 30796 22280 30836 22483
rect 30604 22146 30644 22231
rect 30027 22112 30069 22121
rect 30027 22072 30028 22112
rect 30068 22072 30069 22112
rect 30027 22063 30069 22072
rect 30028 21953 30068 22063
rect 30027 21944 30069 21953
rect 30027 21904 30028 21944
rect 30068 21904 30069 21944
rect 30027 21895 30069 21904
rect 30604 21608 30644 21617
rect 29932 21568 30604 21608
rect 29740 20936 29780 21568
rect 30315 21020 30357 21029
rect 30315 20980 30316 21020
rect 30356 20980 30357 21020
rect 30315 20971 30357 20980
rect 29836 20936 29876 20945
rect 29740 20896 29836 20936
rect 29836 20887 29876 20896
rect 29547 20096 29589 20105
rect 29547 20056 29548 20096
rect 29588 20056 29589 20096
rect 29547 20047 29589 20056
rect 29932 20096 29972 20105
rect 29548 19853 29588 20047
rect 29740 19928 29780 19937
rect 29547 19844 29589 19853
rect 29547 19804 29548 19844
rect 29588 19804 29589 19844
rect 29547 19795 29589 19804
rect 29644 19256 29684 19265
rect 29740 19256 29780 19888
rect 29684 19216 29780 19256
rect 29644 19207 29684 19216
rect 29932 19181 29972 20056
rect 30028 20096 30068 20105
rect 29931 19172 29973 19181
rect 29931 19132 29932 19172
rect 29972 19132 29973 19172
rect 29931 19123 29973 19132
rect 30028 19013 30068 20056
rect 30124 20096 30164 20105
rect 30124 19097 30164 20056
rect 30220 20096 30260 20105
rect 30220 19349 30260 20056
rect 30219 19340 30261 19349
rect 30219 19300 30220 19340
rect 30260 19300 30261 19340
rect 30219 19291 30261 19300
rect 30123 19088 30165 19097
rect 30123 19048 30124 19088
rect 30164 19048 30165 19088
rect 30123 19039 30165 19048
rect 29451 19004 29493 19013
rect 29451 18964 29452 19004
rect 29492 18964 29493 19004
rect 29451 18955 29493 18964
rect 30027 19004 30069 19013
rect 30027 18964 30028 19004
rect 30068 18964 30069 19004
rect 30027 18955 30069 18964
rect 29355 18080 29397 18089
rect 29355 18040 29356 18080
rect 29396 18040 29397 18080
rect 29355 18031 29397 18040
rect 28779 17492 28821 17501
rect 28779 17452 28780 17492
rect 28820 17452 28821 17492
rect 28779 17443 28821 17452
rect 27628 16904 27668 16913
rect 27532 16864 27628 16904
rect 27628 16855 27668 16864
rect 24459 16316 24501 16325
rect 24459 16276 24460 16316
rect 24500 16276 24501 16316
rect 24459 16267 24501 16276
rect 11691 16064 11733 16073
rect 11691 16024 11692 16064
rect 11732 16024 11733 16064
rect 11691 16015 11733 16024
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 29452 15569 29492 18955
rect 29739 18752 29781 18761
rect 29739 18712 29740 18752
rect 29780 18712 29781 18752
rect 29739 18703 29781 18712
rect 29740 18668 29780 18703
rect 30220 18668 30260 19291
rect 30316 18929 30356 20971
rect 30508 19256 30548 21568
rect 30604 21559 30644 21568
rect 30796 20525 30836 22240
rect 30892 22280 30932 23080
rect 30988 23071 31028 23080
rect 30987 22952 31029 22961
rect 30987 22912 30988 22952
rect 31028 22912 31029 22952
rect 30987 22903 31029 22912
rect 30988 22818 31028 22903
rect 30892 22231 30932 22240
rect 30795 20516 30837 20525
rect 30795 20476 30796 20516
rect 30836 20476 30837 20516
rect 30795 20467 30837 20476
rect 31084 19265 31124 23416
rect 31179 23416 31180 23456
rect 31220 23416 31221 23456
rect 31179 23407 31221 23416
rect 31179 23120 31221 23129
rect 31179 23080 31180 23120
rect 31220 23080 31221 23120
rect 31179 23071 31221 23080
rect 31276 23120 31316 23584
rect 31372 23575 31412 23584
rect 31371 23456 31413 23465
rect 31371 23416 31372 23456
rect 31412 23416 31413 23456
rect 31371 23407 31413 23416
rect 31276 23071 31316 23080
rect 31180 22986 31220 23071
rect 31179 22364 31221 22373
rect 31179 22324 31180 22364
rect 31220 22324 31221 22364
rect 31179 22315 31221 22324
rect 31180 22280 31220 22315
rect 31180 22229 31220 22240
rect 31372 20609 31412 23407
rect 31756 23372 31796 24592
rect 31852 24632 31892 24835
rect 32235 24800 32277 24809
rect 32235 24760 32236 24800
rect 32276 24760 32277 24800
rect 32235 24751 32277 24760
rect 32236 24666 32276 24751
rect 31852 24583 31892 24592
rect 31948 24632 31988 24641
rect 32140 24632 32180 24641
rect 31988 24592 32140 24632
rect 31948 24583 31988 24592
rect 32140 24583 32180 24592
rect 32332 24632 32372 24641
rect 32332 24044 32372 24592
rect 32427 24632 32469 24641
rect 32427 24592 32428 24632
rect 32468 24592 32469 24632
rect 32427 24583 32469 24592
rect 32716 24632 32756 24641
rect 32428 24498 32468 24583
rect 32716 24305 32756 24592
rect 32908 24632 32948 24641
rect 33004 24632 33044 25171
rect 33100 25061 33140 25222
rect 33292 25145 33332 25264
rect 33388 25304 33428 25516
rect 33868 25313 33908 25843
rect 33388 25255 33428 25264
rect 33867 25304 33909 25313
rect 33867 25264 33868 25304
rect 33908 25264 33909 25304
rect 33867 25255 33909 25264
rect 34444 25304 34484 25927
rect 34828 25556 34868 26104
rect 34924 26095 34964 26104
rect 34924 25556 34964 25565
rect 34828 25516 34924 25556
rect 34924 25507 34964 25516
rect 34444 25255 34484 25264
rect 34539 25304 34581 25313
rect 34539 25264 34540 25304
rect 34580 25264 34581 25304
rect 34539 25255 34581 25264
rect 34636 25304 34676 25315
rect 33483 25220 33525 25229
rect 33483 25180 33484 25220
rect 33524 25180 33525 25220
rect 33483 25171 33525 25180
rect 33196 25136 33236 25145
rect 33099 25052 33141 25061
rect 33099 25012 33100 25052
rect 33140 25012 33141 25052
rect 33099 25003 33141 25012
rect 33196 24641 33236 25096
rect 33291 25136 33333 25145
rect 33291 25096 33292 25136
rect 33332 25096 33333 25136
rect 33291 25087 33333 25096
rect 33484 24893 33524 25171
rect 33483 24884 33525 24893
rect 33483 24844 33484 24884
rect 33524 24844 33525 24884
rect 33483 24835 33525 24844
rect 32948 24592 33044 24632
rect 32908 24583 32948 24592
rect 32812 24380 32852 24389
rect 32715 24296 32757 24305
rect 32715 24256 32716 24296
rect 32756 24256 32757 24296
rect 32715 24247 32757 24256
rect 32044 24004 32372 24044
rect 31564 23332 31796 23372
rect 31852 23792 31892 23801
rect 31564 22457 31604 23332
rect 31852 23288 31892 23752
rect 32044 23540 32084 24004
rect 32524 23960 32564 23969
rect 32332 23920 32524 23960
rect 32139 23876 32181 23885
rect 32139 23836 32140 23876
rect 32180 23836 32181 23876
rect 32139 23827 32181 23836
rect 32140 23792 32180 23827
rect 32140 23741 32180 23752
rect 32235 23792 32277 23801
rect 32235 23752 32236 23792
rect 32276 23752 32277 23792
rect 32235 23743 32277 23752
rect 32236 23658 32276 23743
rect 32044 23500 32276 23540
rect 31660 23248 31892 23288
rect 31563 22448 31605 22457
rect 31563 22408 31564 22448
rect 31604 22408 31605 22448
rect 31563 22399 31605 22408
rect 31660 22373 31700 23248
rect 32140 23213 32180 23244
rect 32139 23204 32181 23213
rect 32139 23164 32140 23204
rect 32180 23164 32181 23204
rect 32139 23155 32181 23164
rect 32236 23204 32276 23500
rect 31756 23120 31796 23131
rect 31756 23045 31796 23080
rect 31851 23120 31893 23129
rect 31851 23080 31852 23120
rect 31892 23080 31893 23120
rect 31851 23071 31893 23080
rect 31948 23120 31988 23129
rect 31755 23036 31797 23045
rect 31755 22996 31756 23036
rect 31796 22996 31797 23036
rect 31755 22987 31797 22996
rect 31756 22956 31796 22987
rect 31852 22868 31892 23071
rect 31756 22828 31852 22868
rect 31659 22364 31701 22373
rect 31659 22324 31660 22364
rect 31700 22324 31701 22364
rect 31659 22315 31701 22324
rect 31756 22289 31796 22828
rect 31852 22819 31892 22828
rect 31852 22532 31892 22541
rect 31948 22532 31988 23080
rect 32140 23120 32180 23155
rect 32236 23129 32276 23164
rect 32140 23045 32180 23080
rect 32235 23120 32277 23129
rect 32235 23080 32236 23120
rect 32276 23080 32277 23120
rect 32235 23071 32277 23080
rect 32332 23120 32372 23920
rect 32524 23911 32564 23920
rect 32716 23885 32756 24247
rect 32715 23876 32757 23885
rect 32715 23836 32716 23876
rect 32756 23836 32757 23876
rect 32715 23827 32757 23836
rect 32619 23288 32661 23297
rect 32619 23248 32620 23288
rect 32660 23248 32661 23288
rect 32619 23239 32661 23248
rect 32620 23154 32660 23239
rect 32332 23071 32372 23080
rect 32524 23120 32564 23129
rect 32139 23036 32181 23045
rect 32236 23040 32276 23071
rect 32139 22996 32140 23036
rect 32180 22996 32181 23036
rect 32139 22987 32181 22996
rect 31892 22492 31988 22532
rect 31852 22483 31892 22492
rect 32140 22448 32180 22987
rect 32122 22408 32180 22448
rect 32122 22364 32162 22408
rect 32057 22324 32162 22364
rect 31468 22280 31508 22289
rect 31468 21701 31508 22240
rect 31563 22280 31605 22289
rect 31563 22240 31564 22280
rect 31604 22240 31605 22280
rect 31563 22231 31605 22240
rect 31755 22280 31797 22289
rect 32057 22280 32097 22324
rect 31755 22240 31756 22280
rect 31796 22240 31797 22280
rect 31755 22231 31797 22240
rect 32044 22240 32097 22280
rect 32331 22280 32373 22289
rect 31564 22146 31604 22231
rect 31467 21692 31509 21701
rect 31467 21652 31468 21692
rect 31508 21652 31509 21692
rect 31467 21643 31509 21652
rect 31755 21440 31797 21449
rect 31755 21400 31756 21440
rect 31796 21400 31797 21440
rect 31755 21391 31797 21400
rect 31756 21306 31796 21391
rect 31371 20600 31413 20609
rect 31371 20560 31372 20600
rect 31412 20560 31413 20600
rect 31371 20551 31413 20560
rect 31756 20012 31796 20021
rect 31659 19340 31701 19349
rect 31659 19300 31660 19340
rect 31700 19300 31701 19340
rect 31659 19291 31701 19300
rect 30315 18920 30357 18929
rect 30315 18880 30316 18920
rect 30356 18880 30357 18920
rect 30315 18871 30357 18880
rect 30316 18668 30356 18677
rect 30220 18628 30316 18668
rect 29644 18584 29684 18593
rect 29644 18257 29684 18544
rect 29643 18248 29685 18257
rect 29643 18208 29644 18248
rect 29684 18208 29685 18248
rect 29643 18199 29685 18208
rect 29740 17996 29780 18628
rect 30316 18619 30356 18628
rect 29836 18584 29876 18593
rect 29836 18416 29876 18544
rect 30412 18584 30452 18593
rect 30028 18416 30068 18425
rect 29836 18376 30028 18416
rect 30028 18367 30068 18376
rect 29740 17956 30068 17996
rect 29835 17744 29877 17753
rect 29835 17704 29836 17744
rect 29876 17704 29877 17744
rect 29835 17695 29877 17704
rect 30028 17744 30068 17956
rect 30028 17695 30068 17704
rect 30124 17744 30164 17753
rect 29836 17610 29876 17695
rect 29931 17660 29973 17669
rect 29931 17620 29932 17660
rect 29972 17620 29973 17660
rect 29931 17611 29973 17620
rect 29547 17576 29589 17585
rect 29547 17536 29548 17576
rect 29588 17536 29589 17576
rect 29547 17527 29589 17536
rect 29548 17442 29588 17527
rect 29932 17526 29972 17611
rect 30124 17165 30164 17704
rect 30315 17660 30357 17669
rect 30315 17620 30316 17660
rect 30356 17620 30357 17660
rect 30315 17611 30357 17620
rect 30316 17526 30356 17611
rect 30219 17492 30261 17501
rect 30219 17452 30220 17492
rect 30260 17452 30261 17492
rect 30219 17443 30261 17452
rect 30123 17156 30165 17165
rect 30123 17116 30124 17156
rect 30164 17116 30165 17156
rect 30123 17107 30165 17116
rect 30220 17072 30260 17443
rect 30412 17333 30452 18544
rect 30508 18341 30548 19216
rect 31083 19256 31125 19265
rect 31083 19216 31084 19256
rect 31124 19216 31125 19256
rect 31083 19207 31125 19216
rect 31660 19206 31700 19291
rect 30699 18668 30741 18677
rect 30699 18628 30700 18668
rect 30740 18628 30741 18668
rect 30699 18619 30741 18628
rect 30700 18584 30740 18619
rect 30700 18533 30740 18544
rect 31179 18584 31221 18593
rect 31179 18544 31180 18584
rect 31220 18544 31221 18584
rect 31179 18535 31221 18544
rect 31659 18584 31701 18593
rect 31659 18544 31660 18584
rect 31700 18544 31701 18584
rect 31659 18535 31701 18544
rect 31180 18450 31220 18535
rect 30507 18332 30549 18341
rect 30507 18292 30508 18332
rect 30548 18292 30549 18332
rect 30507 18283 30549 18292
rect 31563 18332 31605 18341
rect 31563 18292 31564 18332
rect 31604 18292 31605 18332
rect 31563 18283 31605 18292
rect 31564 17753 31604 18283
rect 30700 17744 30740 17753
rect 31371 17744 31413 17753
rect 30740 17704 30836 17744
rect 30700 17695 30740 17704
rect 30411 17324 30453 17333
rect 30411 17284 30412 17324
rect 30452 17284 30453 17324
rect 30411 17275 30453 17284
rect 30603 17324 30645 17333
rect 30603 17284 30604 17324
rect 30644 17284 30645 17324
rect 30603 17275 30645 17284
rect 30507 17156 30549 17165
rect 30507 17116 30508 17156
rect 30548 17116 30549 17156
rect 30507 17107 30549 17116
rect 30412 17072 30452 17081
rect 30220 17032 30412 17072
rect 30412 17023 30452 17032
rect 30508 17022 30548 17107
rect 30604 17072 30644 17275
rect 30604 17023 30644 17032
rect 30796 16904 30836 17704
rect 31371 17704 31372 17744
rect 31412 17704 31413 17744
rect 31371 17695 31413 17704
rect 31563 17744 31605 17753
rect 31563 17704 31564 17744
rect 31604 17704 31605 17744
rect 31563 17695 31605 17704
rect 31275 17408 31317 17417
rect 31275 17368 31276 17408
rect 31316 17368 31317 17408
rect 31275 17359 31317 17368
rect 30796 16855 30836 16864
rect 31084 16148 31124 16157
rect 31084 15905 31124 16108
rect 31083 15896 31125 15905
rect 31083 15856 31084 15896
rect 31124 15856 31125 15896
rect 31083 15847 31125 15856
rect 29451 15560 29493 15569
rect 29451 15520 29452 15560
rect 29492 15520 29493 15560
rect 29451 15511 29493 15520
rect 30219 15392 30261 15401
rect 30219 15352 30220 15392
rect 30260 15352 30261 15392
rect 30219 15343 30261 15352
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 30220 14720 30260 15343
rect 30220 14671 30260 14680
rect 30604 14720 30644 14729
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 30219 14048 30261 14057
rect 30219 14008 30220 14048
rect 30260 14008 30261 14048
rect 30219 13999 30261 14008
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 29931 12536 29973 12545
rect 30220 12536 30260 13999
rect 30604 13880 30644 14680
rect 31276 14141 31316 17359
rect 31372 15560 31412 17695
rect 31564 17610 31604 17695
rect 31564 16904 31604 16913
rect 31468 16232 31508 16241
rect 31564 16232 31604 16864
rect 31508 16192 31604 16232
rect 31468 16183 31508 16192
rect 31564 15560 31604 15569
rect 31372 15520 31564 15560
rect 31564 15511 31604 15520
rect 31563 15392 31605 15401
rect 31563 15352 31564 15392
rect 31604 15352 31605 15392
rect 31563 15343 31605 15352
rect 31564 15258 31604 15343
rect 31660 15140 31700 18535
rect 31756 17501 31796 19972
rect 31948 19844 31988 19853
rect 31851 19340 31893 19349
rect 31851 19300 31852 19340
rect 31892 19300 31893 19340
rect 31851 19291 31893 19300
rect 31852 19256 31892 19291
rect 31852 19205 31892 19216
rect 31948 19256 31988 19804
rect 32044 19433 32084 22240
rect 32140 22238 32180 22247
rect 32331 22240 32332 22280
rect 32372 22240 32373 22280
rect 32331 22231 32373 22240
rect 32428 22280 32468 22289
rect 32140 21617 32180 22198
rect 32235 22196 32277 22205
rect 32235 22156 32236 22196
rect 32276 22156 32277 22196
rect 32235 22147 32277 22156
rect 32236 22062 32276 22147
rect 32332 22146 32372 22231
rect 32331 21692 32373 21701
rect 32331 21652 32332 21692
rect 32372 21652 32373 21692
rect 32331 21643 32373 21652
rect 32428 21692 32468 22240
rect 32524 21776 32564 23080
rect 32715 23120 32757 23129
rect 32715 23080 32716 23120
rect 32756 23080 32757 23120
rect 32715 23071 32757 23080
rect 32812 23120 32852 24340
rect 33004 23717 33044 24592
rect 33195 24632 33237 24641
rect 33195 24592 33196 24632
rect 33236 24592 33237 24632
rect 33195 24583 33237 24592
rect 33868 24557 33908 25255
rect 34540 25170 34580 25255
rect 34636 25229 34676 25264
rect 34732 25304 34772 25313
rect 34924 25304 34964 25313
rect 34772 25264 34924 25304
rect 34732 25255 34772 25264
rect 34924 25255 34964 25264
rect 34635 25220 34677 25229
rect 34635 25180 34636 25220
rect 34676 25180 34677 25220
rect 34635 25171 34677 25180
rect 35020 25052 35060 26851
rect 35116 25901 35156 26944
rect 35308 26935 35348 26944
rect 35595 26900 35637 26909
rect 35595 26860 35596 26900
rect 35636 26860 35637 26900
rect 35595 26851 35637 26860
rect 35211 26816 35253 26825
rect 35211 26776 35212 26816
rect 35252 26776 35253 26816
rect 35211 26767 35253 26776
rect 35404 26816 35444 26825
rect 35212 26682 35252 26767
rect 35212 26144 35252 26153
rect 35212 25985 35252 26104
rect 35307 26144 35349 26153
rect 35307 26104 35308 26144
rect 35348 26104 35349 26144
rect 35307 26095 35349 26104
rect 35308 26010 35348 26095
rect 35211 25976 35253 25985
rect 35211 25936 35212 25976
rect 35252 25936 35253 25976
rect 35404 25976 35444 26776
rect 35596 26766 35636 26851
rect 35691 26816 35733 26825
rect 35691 26776 35692 26816
rect 35732 26776 35733 26816
rect 35691 26767 35733 26776
rect 36364 26816 36404 26825
rect 36460 26816 36500 27448
rect 38668 26900 38708 27859
rect 38956 27656 38996 29128
rect 39628 29119 39668 29128
rect 39628 28589 39668 28674
rect 39627 28580 39669 28589
rect 39627 28540 39628 28580
rect 39668 28540 39669 28580
rect 39627 28531 39669 28540
rect 39436 28412 39476 28421
rect 39724 28412 39764 30211
rect 40204 30092 40244 30211
rect 40204 30043 40244 30052
rect 40012 30008 40052 30017
rect 39476 28372 39764 28412
rect 39820 29924 39860 29933
rect 39436 28363 39476 28372
rect 39820 28328 39860 29884
rect 40012 29849 40052 29968
rect 40396 29924 40436 30388
rect 40684 30379 40724 30388
rect 40779 30428 40821 30437
rect 40779 30388 40780 30428
rect 40820 30388 40821 30428
rect 40779 30379 40821 30388
rect 40011 29840 40053 29849
rect 40011 29800 40012 29840
rect 40052 29800 40053 29840
rect 40011 29791 40053 29800
rect 40011 28748 40053 28757
rect 40011 28708 40012 28748
rect 40052 28708 40053 28748
rect 40011 28699 40053 28708
rect 40012 28412 40052 28699
rect 40396 28673 40436 29884
rect 40588 29840 40628 29849
rect 40588 29168 40628 29800
rect 40683 29840 40725 29849
rect 40683 29800 40684 29840
rect 40724 29800 40725 29840
rect 40683 29791 40725 29800
rect 40780 29840 40820 30379
rect 40780 29791 40820 29800
rect 40684 29706 40724 29791
rect 40876 29672 40916 29681
rect 40779 29168 40821 29177
rect 40588 29128 40780 29168
rect 40820 29128 40821 29168
rect 40779 29119 40821 29128
rect 40780 28916 40820 29119
rect 40395 28664 40437 28673
rect 40395 28624 40396 28664
rect 40436 28624 40437 28664
rect 40395 28615 40437 28624
rect 40395 28496 40437 28505
rect 40395 28456 40396 28496
rect 40436 28456 40437 28496
rect 40395 28447 40437 28456
rect 40012 28363 40052 28372
rect 40396 28337 40436 28447
rect 38860 26984 38900 26995
rect 38860 26909 38900 26944
rect 38572 26860 38668 26900
rect 36404 26776 36500 26816
rect 37228 26816 37268 26825
rect 36364 26767 36404 26776
rect 35596 25976 35636 25985
rect 35404 25936 35596 25976
rect 35692 25976 35732 26767
rect 35980 26732 36020 26741
rect 35788 26648 35828 26657
rect 35788 26321 35828 26608
rect 35787 26312 35829 26321
rect 35787 26272 35788 26312
rect 35828 26272 35829 26312
rect 35787 26263 35829 26272
rect 35884 26312 35924 26321
rect 35980 26312 36020 26692
rect 37035 26396 37077 26405
rect 37035 26356 37036 26396
rect 37076 26356 37077 26396
rect 37035 26347 37077 26356
rect 35924 26272 36020 26312
rect 36076 26272 36404 26312
rect 35884 26263 35924 26272
rect 35788 26144 35828 26153
rect 35980 26144 36020 26153
rect 35828 26104 35924 26144
rect 35788 26095 35828 26104
rect 35692 25936 35828 25976
rect 35211 25927 35253 25936
rect 35596 25927 35636 25936
rect 35115 25892 35157 25901
rect 35115 25852 35116 25892
rect 35156 25852 35157 25892
rect 35115 25843 35157 25852
rect 35116 25304 35156 25843
rect 35692 25472 35732 25481
rect 35116 25255 35156 25264
rect 35212 25432 35692 25472
rect 35212 25304 35252 25432
rect 35692 25423 35732 25432
rect 35212 25255 35252 25264
rect 35595 25304 35637 25313
rect 35595 25264 35596 25304
rect 35636 25264 35637 25304
rect 35595 25255 35637 25264
rect 35692 25304 35732 25313
rect 35020 25012 35156 25052
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 35019 24884 35061 24893
rect 35019 24844 35020 24884
rect 35060 24844 35061 24884
rect 35019 24835 35061 24844
rect 34924 24716 34964 24725
rect 35020 24716 35060 24835
rect 34964 24676 35060 24716
rect 34924 24667 34964 24676
rect 34156 24632 34196 24641
rect 34196 24592 34292 24632
rect 34156 24583 34196 24592
rect 33867 24548 33909 24557
rect 33867 24508 33868 24548
rect 33908 24508 33909 24548
rect 33867 24499 33909 24508
rect 33868 24464 33908 24499
rect 33868 24413 33908 24424
rect 34155 24464 34197 24473
rect 34155 24424 34156 24464
rect 34196 24424 34197 24464
rect 34155 24415 34197 24424
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 33292 23792 33332 23801
rect 32908 23708 32948 23717
rect 32908 23297 32948 23668
rect 33003 23708 33045 23717
rect 33003 23668 33004 23708
rect 33044 23668 33045 23708
rect 33003 23659 33045 23668
rect 32907 23288 32949 23297
rect 32907 23248 32908 23288
rect 32948 23248 32949 23288
rect 32907 23239 32949 23248
rect 32812 23071 32852 23080
rect 32716 22986 32756 23071
rect 32907 22448 32949 22457
rect 32907 22408 32908 22448
rect 32948 22408 32949 22448
rect 32907 22399 32949 22408
rect 32811 22196 32853 22205
rect 32811 22156 32812 22196
rect 32852 22156 32853 22196
rect 32811 22147 32853 22156
rect 32812 22062 32852 22147
rect 32908 21869 32948 22399
rect 32907 21860 32949 21869
rect 32907 21820 32908 21860
rect 32948 21820 32949 21860
rect 32907 21811 32949 21820
rect 32524 21736 32660 21776
rect 32428 21643 32468 21652
rect 32139 21608 32181 21617
rect 32139 21568 32140 21608
rect 32180 21568 32181 21608
rect 32139 21559 32181 21568
rect 32332 21608 32372 21643
rect 32620 21617 32660 21736
rect 32332 21557 32372 21568
rect 32524 21608 32564 21617
rect 32236 20684 32276 20693
rect 32236 20264 32276 20644
rect 32524 20273 32564 21568
rect 32619 21608 32661 21617
rect 32619 21568 32620 21608
rect 32660 21568 32661 21608
rect 32619 21559 32661 21568
rect 32716 21440 32756 21449
rect 32620 20768 32660 20777
rect 32716 20768 32756 21400
rect 32660 20728 32756 20768
rect 32620 20719 32660 20728
rect 32908 20600 32948 21811
rect 32812 20560 32948 20600
rect 32715 20516 32757 20525
rect 32715 20476 32716 20516
rect 32756 20476 32757 20516
rect 32715 20467 32757 20476
rect 32332 20264 32372 20273
rect 32236 20224 32332 20264
rect 32332 20215 32372 20224
rect 32523 20264 32565 20273
rect 32523 20224 32524 20264
rect 32564 20224 32565 20264
rect 32523 20215 32565 20224
rect 32140 20096 32180 20105
rect 32140 19508 32180 20056
rect 32140 19459 32180 19468
rect 32236 20096 32276 20105
rect 32043 19424 32085 19433
rect 32043 19384 32044 19424
rect 32084 19384 32085 19424
rect 32043 19375 32085 19384
rect 32140 19256 32180 19265
rect 31988 19216 32084 19256
rect 31948 19207 31988 19216
rect 31947 19088 31989 19097
rect 31947 19048 31948 19088
rect 31988 19048 31989 19088
rect 31947 19039 31989 19048
rect 31851 19004 31893 19013
rect 31851 18964 31852 19004
rect 31892 18964 31893 19004
rect 31851 18955 31893 18964
rect 31852 18173 31892 18955
rect 31851 18164 31893 18173
rect 31851 18124 31852 18164
rect 31892 18124 31893 18164
rect 31851 18115 31893 18124
rect 31755 17492 31797 17501
rect 31755 17452 31756 17492
rect 31796 17452 31797 17492
rect 31755 17443 31797 17452
rect 31851 15644 31893 15653
rect 31851 15604 31852 15644
rect 31892 15604 31893 15644
rect 31851 15595 31893 15604
rect 31564 15100 31700 15140
rect 31756 15560 31796 15569
rect 31467 14720 31509 14729
rect 31467 14680 31468 14720
rect 31508 14680 31509 14720
rect 31467 14671 31509 14680
rect 31468 14586 31508 14671
rect 31275 14132 31317 14141
rect 31275 14092 31276 14132
rect 31316 14092 31317 14132
rect 31275 14083 31317 14092
rect 31564 14057 31604 15100
rect 31756 14981 31796 15520
rect 31852 15560 31892 15595
rect 31852 15509 31892 15520
rect 31948 15308 31988 19039
rect 31852 15268 31988 15308
rect 32044 15560 32084 19216
rect 32140 18509 32180 19216
rect 32236 18761 32276 20056
rect 32428 20096 32468 20105
rect 32620 20096 32660 20105
rect 32468 20056 32620 20096
rect 32428 20047 32468 20056
rect 32620 20047 32660 20056
rect 32716 20096 32756 20467
rect 32716 20047 32756 20056
rect 32812 20096 32852 20560
rect 33004 20189 33044 23659
rect 33292 23060 33332 23752
rect 34156 23792 34196 24415
rect 34156 23060 34196 23752
rect 33292 23020 33428 23060
rect 33388 22952 33428 23020
rect 33388 22903 33428 22912
rect 34060 23020 34196 23060
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 33196 22280 33236 22289
rect 34060 22280 34100 23020
rect 33236 22240 33332 22280
rect 33196 22231 33236 22240
rect 33292 21440 33332 22240
rect 34060 22231 34100 22240
rect 33292 21391 33332 21400
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 33484 20768 33524 20777
rect 33524 20728 34196 20768
rect 33484 20719 33524 20728
rect 33003 20180 33045 20189
rect 33003 20140 33004 20180
rect 33044 20140 33045 20180
rect 33003 20131 33045 20140
rect 32812 20047 32852 20056
rect 32908 20096 32948 20105
rect 32908 19937 32948 20056
rect 32907 19928 32949 19937
rect 32907 19888 32908 19928
rect 32948 19888 32949 19928
rect 32907 19879 32949 19888
rect 32908 19433 32948 19879
rect 33004 19601 33044 20131
rect 33388 19928 33428 19937
rect 33196 19888 33388 19928
rect 33003 19592 33045 19601
rect 33003 19552 33004 19592
rect 33044 19552 33045 19592
rect 33003 19543 33045 19552
rect 33196 19550 33236 19888
rect 33388 19879 33428 19888
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 33196 19510 33428 19550
rect 32907 19424 32949 19433
rect 32907 19384 32908 19424
rect 32948 19384 32949 19424
rect 32907 19375 32949 19384
rect 33291 19424 33333 19433
rect 33291 19384 33292 19424
rect 33332 19384 33333 19424
rect 33291 19375 33333 19384
rect 32908 19256 32948 19265
rect 33196 19256 33236 19265
rect 32948 19216 33044 19256
rect 32908 19207 32948 19216
rect 32524 18880 32852 18920
rect 32235 18752 32277 18761
rect 32235 18712 32236 18752
rect 32276 18712 32277 18752
rect 32235 18703 32277 18712
rect 32524 18668 32564 18880
rect 32619 18752 32661 18761
rect 32619 18712 32620 18752
rect 32660 18712 32661 18752
rect 32619 18703 32661 18712
rect 32524 18619 32564 18628
rect 32428 18584 32468 18593
rect 32139 18500 32181 18509
rect 32139 18460 32140 18500
rect 32180 18460 32181 18500
rect 32139 18451 32181 18460
rect 32331 18500 32373 18509
rect 32331 18460 32332 18500
rect 32372 18460 32373 18500
rect 32331 18451 32373 18460
rect 32140 17669 32180 18451
rect 32332 17753 32372 18451
rect 32428 18425 32468 18544
rect 32620 18584 32660 18703
rect 32812 18668 32852 18880
rect 33004 18677 33044 19216
rect 33196 18677 33236 19216
rect 33292 19256 33332 19375
rect 33292 19207 33332 19216
rect 32908 18668 32948 18677
rect 32812 18628 32908 18668
rect 32908 18619 32948 18628
rect 33003 18668 33045 18677
rect 33003 18628 33004 18668
rect 33044 18628 33045 18668
rect 33003 18619 33045 18628
rect 33195 18668 33237 18677
rect 33195 18628 33196 18668
rect 33236 18628 33237 18668
rect 33195 18619 33237 18628
rect 32620 18535 32660 18544
rect 32716 18584 32756 18593
rect 32427 18416 32469 18425
rect 32427 18376 32428 18416
rect 32468 18376 32469 18416
rect 32427 18367 32469 18376
rect 32428 17837 32468 18367
rect 32716 18005 32756 18544
rect 32811 18248 32853 18257
rect 32811 18208 32812 18248
rect 32852 18208 32853 18248
rect 32811 18199 32853 18208
rect 32715 17996 32757 18005
rect 32715 17956 32716 17996
rect 32756 17956 32757 17996
rect 32715 17947 32757 17956
rect 32427 17828 32469 17837
rect 32427 17788 32428 17828
rect 32468 17788 32469 17828
rect 32427 17779 32469 17788
rect 32331 17744 32373 17753
rect 32331 17704 32332 17744
rect 32372 17704 32373 17744
rect 32331 17695 32373 17704
rect 32139 17660 32181 17669
rect 32139 17620 32140 17660
rect 32180 17620 32181 17660
rect 32139 17611 32181 17620
rect 32332 16232 32372 17695
rect 32716 17576 32756 17585
rect 32716 17333 32756 17536
rect 32715 17324 32757 17333
rect 32715 17284 32716 17324
rect 32756 17284 32757 17324
rect 32715 17275 32757 17284
rect 32812 17324 32852 18199
rect 32907 17324 32949 17333
rect 32812 17284 32908 17324
rect 32948 17284 32949 17324
rect 32332 16183 32372 16192
rect 32139 15644 32181 15653
rect 32139 15604 32140 15644
rect 32180 15604 32181 15644
rect 32139 15595 32181 15604
rect 31755 14972 31797 14981
rect 31755 14932 31756 14972
rect 31796 14932 31797 14972
rect 31755 14923 31797 14932
rect 31755 14468 31797 14477
rect 31755 14428 31756 14468
rect 31796 14428 31797 14468
rect 31755 14419 31797 14428
rect 31563 14048 31605 14057
rect 31563 14008 31564 14048
rect 31604 14008 31605 14048
rect 31563 13999 31605 14008
rect 31660 14048 31700 14057
rect 30700 13880 30740 13889
rect 30604 13840 30700 13880
rect 30700 13831 30740 13840
rect 31660 13217 31700 14008
rect 31756 14048 31796 14419
rect 31852 14225 31892 15268
rect 32044 14813 32084 15520
rect 32140 15510 32180 15595
rect 32236 15560 32276 15569
rect 32043 14804 32085 14813
rect 32043 14764 32044 14804
rect 32084 14764 32085 14804
rect 32043 14755 32085 14764
rect 32236 14561 32276 15520
rect 32427 15560 32469 15569
rect 32427 15520 32428 15560
rect 32468 15520 32469 15560
rect 32427 15511 32469 15520
rect 32235 14552 32277 14561
rect 32235 14512 32236 14552
rect 32276 14512 32277 14552
rect 32235 14503 32277 14512
rect 32428 14477 32468 15511
rect 32715 14972 32757 14981
rect 32715 14932 32716 14972
rect 32756 14932 32757 14972
rect 32715 14923 32757 14932
rect 32619 14552 32661 14561
rect 32524 14512 32620 14552
rect 32660 14512 32661 14552
rect 32427 14468 32469 14477
rect 32427 14428 32428 14468
rect 32468 14428 32469 14468
rect 32427 14419 32469 14428
rect 31851 14216 31893 14225
rect 31851 14176 31852 14216
rect 31892 14176 31893 14216
rect 31851 14167 31893 14176
rect 31756 13999 31796 14008
rect 31852 14048 31892 14167
rect 32235 14132 32277 14141
rect 32235 14092 32236 14132
rect 32276 14092 32277 14132
rect 32235 14083 32277 14092
rect 31852 13999 31892 14008
rect 31948 14048 31988 14059
rect 31948 13973 31988 14008
rect 32236 14048 32276 14083
rect 32236 13997 32276 14008
rect 32524 14048 32564 14512
rect 32619 14503 32661 14512
rect 32620 14418 32660 14503
rect 32524 13999 32564 14008
rect 32620 14048 32660 14057
rect 32620 13973 32660 14008
rect 31947 13964 31989 13973
rect 31947 13924 31948 13964
rect 31988 13924 31989 13964
rect 31947 13915 31989 13924
rect 32619 13964 32661 13973
rect 32619 13924 32620 13964
rect 32660 13924 32661 13964
rect 32619 13915 32661 13924
rect 32620 13301 32660 13915
rect 32619 13292 32661 13301
rect 32619 13252 32620 13292
rect 32660 13252 32661 13292
rect 32619 13243 32661 13252
rect 31659 13208 31701 13217
rect 31659 13168 31660 13208
rect 31700 13168 31701 13208
rect 31659 13159 31701 13168
rect 32716 12980 32756 14923
rect 32812 14720 32852 17284
rect 32907 17275 32949 17284
rect 33004 16325 33044 18619
rect 33196 17753 33236 18619
rect 33292 18584 33332 18593
rect 33388 18584 33428 19510
rect 33580 19424 33620 19433
rect 33620 19384 33812 19424
rect 33580 19375 33620 19384
rect 33772 19256 33812 19384
rect 33772 19207 33812 19216
rect 33964 19256 34004 19265
rect 33868 19172 33908 19181
rect 33868 18761 33908 19132
rect 33867 18752 33909 18761
rect 33867 18712 33868 18752
rect 33908 18712 33909 18752
rect 33867 18703 33909 18712
rect 33332 18544 33428 18584
rect 33292 18535 33332 18544
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 33387 17996 33429 18005
rect 33387 17956 33388 17996
rect 33428 17956 33429 17996
rect 33387 17947 33429 17956
rect 33388 17862 33428 17947
rect 33195 17744 33237 17753
rect 33195 17704 33196 17744
rect 33236 17704 33237 17744
rect 33195 17695 33237 17704
rect 33292 17744 33332 17753
rect 33292 17072 33332 17704
rect 33483 17744 33525 17753
rect 33483 17704 33484 17744
rect 33524 17704 33525 17744
rect 33483 17695 33525 17704
rect 33484 17610 33524 17695
rect 33964 17333 34004 19216
rect 34156 18584 34196 20728
rect 34252 18593 34292 24592
rect 35116 23969 35156 25012
rect 35596 24977 35636 25255
rect 35692 25061 35732 25264
rect 35691 25052 35733 25061
rect 35691 25012 35692 25052
rect 35732 25012 35733 25052
rect 35691 25003 35733 25012
rect 35595 24968 35637 24977
rect 35595 24928 35596 24968
rect 35636 24928 35637 24968
rect 35595 24919 35637 24928
rect 35308 24632 35348 24641
rect 35211 24296 35253 24305
rect 35211 24256 35212 24296
rect 35252 24256 35253 24296
rect 35211 24247 35253 24256
rect 35115 23960 35157 23969
rect 35115 23920 35116 23960
rect 35156 23920 35157 23960
rect 35115 23911 35157 23920
rect 35212 23624 35252 24247
rect 35308 23960 35348 24592
rect 35500 23960 35540 23969
rect 35308 23920 35500 23960
rect 35500 23911 35540 23920
rect 35308 23624 35348 23633
rect 35212 23584 35308 23624
rect 35308 23575 35348 23584
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 35596 23060 35636 24919
rect 35692 24137 35732 25003
rect 35691 24128 35733 24137
rect 35691 24088 35692 24128
rect 35732 24088 35733 24128
rect 35691 24079 35733 24088
rect 35788 23213 35828 25936
rect 35884 25481 35924 26104
rect 35980 25901 36020 26104
rect 36076 26144 36116 26272
rect 36364 26228 36404 26272
rect 36364 26179 36404 26188
rect 36076 26095 36116 26104
rect 36267 26144 36309 26153
rect 36267 26104 36268 26144
rect 36308 26104 36309 26144
rect 36267 26095 36309 26104
rect 36459 26144 36501 26153
rect 36459 26104 36460 26144
rect 36500 26104 36501 26144
rect 36459 26095 36501 26104
rect 35979 25892 36021 25901
rect 35979 25852 35980 25892
rect 36020 25852 36021 25892
rect 35979 25843 36021 25852
rect 36171 25892 36213 25901
rect 36171 25852 36172 25892
rect 36212 25852 36213 25892
rect 36171 25843 36213 25852
rect 35883 25472 35925 25481
rect 35883 25432 35884 25472
rect 35924 25432 35925 25472
rect 35883 25423 35925 25432
rect 35884 25304 35924 25313
rect 35884 24809 35924 25264
rect 35980 25304 36020 25313
rect 35883 24800 35925 24809
rect 35883 24760 35884 24800
rect 35924 24760 35925 24800
rect 35883 24751 35925 24760
rect 35980 23792 36020 25264
rect 36075 25220 36117 25229
rect 36075 25180 36076 25220
rect 36116 25180 36117 25220
rect 36075 25171 36117 25180
rect 36076 24380 36116 25171
rect 36172 24641 36212 25843
rect 36268 24809 36308 26095
rect 36460 25985 36500 26095
rect 36459 25976 36501 25985
rect 36459 25936 36460 25976
rect 36500 25936 36501 25976
rect 36459 25927 36501 25936
rect 36555 24884 36597 24893
rect 36555 24844 36556 24884
rect 36596 24844 36597 24884
rect 36555 24835 36597 24844
rect 36267 24800 36309 24809
rect 36267 24760 36268 24800
rect 36308 24760 36309 24800
rect 36267 24751 36309 24760
rect 36171 24632 36213 24641
rect 36171 24592 36172 24632
rect 36212 24592 36213 24632
rect 36171 24583 36213 24592
rect 36172 24498 36212 24583
rect 36076 24340 36308 24380
rect 36171 23960 36213 23969
rect 36171 23920 36172 23960
rect 36212 23920 36213 23960
rect 36171 23911 36213 23920
rect 36075 23792 36117 23801
rect 35980 23752 36076 23792
rect 36116 23752 36117 23792
rect 36075 23743 36117 23752
rect 36172 23792 36212 23911
rect 36076 23658 36116 23743
rect 35787 23204 35829 23213
rect 35787 23164 35788 23204
rect 35828 23164 35829 23204
rect 35787 23155 35829 23164
rect 35596 23020 35828 23060
rect 35211 22532 35253 22541
rect 35211 22492 35212 22532
rect 35252 22492 35253 22532
rect 35211 22483 35253 22492
rect 35212 22398 35252 22483
rect 35691 22196 35733 22205
rect 35691 22156 35692 22196
rect 35732 22156 35733 22196
rect 35691 22147 35733 22156
rect 35212 22112 35252 22121
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 35212 21701 35252 22072
rect 35692 22062 35732 22147
rect 35211 21692 35253 21701
rect 35211 21652 35212 21692
rect 35252 21652 35253 21692
rect 35211 21643 35253 21652
rect 35788 21617 35828 23020
rect 35980 22952 36020 22961
rect 36020 22912 36116 22952
rect 35980 22903 36020 22912
rect 36076 22280 36116 22912
rect 36076 22231 36116 22240
rect 36172 21953 36212 23752
rect 36268 23792 36308 24340
rect 36556 24044 36596 24835
rect 36939 24632 36981 24641
rect 36939 24592 36940 24632
rect 36980 24592 36981 24632
rect 36939 24583 36981 24592
rect 36556 23995 36596 24004
rect 36268 23633 36308 23752
rect 36364 23792 36404 23801
rect 36556 23792 36596 23801
rect 36404 23752 36556 23792
rect 36364 23743 36404 23752
rect 36556 23743 36596 23752
rect 36651 23792 36693 23801
rect 36651 23752 36652 23792
rect 36692 23752 36693 23792
rect 36651 23743 36693 23752
rect 36748 23792 36788 23801
rect 36267 23624 36309 23633
rect 36267 23584 36268 23624
rect 36308 23584 36309 23624
rect 36267 23575 36309 23584
rect 36267 23372 36309 23381
rect 36267 23332 36268 23372
rect 36308 23332 36309 23372
rect 36267 23323 36309 23332
rect 36268 23120 36308 23323
rect 36652 23204 36692 23743
rect 36652 23155 36692 23164
rect 36268 23071 36308 23080
rect 36556 23120 36596 23129
rect 36459 22616 36501 22625
rect 36459 22576 36460 22616
rect 36500 22576 36501 22616
rect 36459 22567 36501 22576
rect 36267 22196 36309 22205
rect 36267 22156 36268 22196
rect 36308 22156 36309 22196
rect 36267 22147 36309 22156
rect 36171 21944 36213 21953
rect 36171 21904 36172 21944
rect 36212 21904 36213 21944
rect 36171 21895 36213 21904
rect 36172 21776 36212 21785
rect 36268 21776 36308 22147
rect 36212 21736 36308 21776
rect 36172 21727 36212 21736
rect 36076 21617 36116 21702
rect 36460 21617 36500 22567
rect 36556 21785 36596 23080
rect 36748 22625 36788 23752
rect 36844 23792 36884 23801
rect 36844 23297 36884 23752
rect 36843 23288 36885 23297
rect 36843 23248 36844 23288
rect 36884 23248 36885 23288
rect 36843 23239 36885 23248
rect 36940 23060 36980 24583
rect 37036 24473 37076 26347
rect 37228 25901 37268 26776
rect 38380 26648 38420 26657
rect 38380 26153 38420 26608
rect 38379 26144 38421 26153
rect 38379 26104 38380 26144
rect 38420 26104 38421 26144
rect 38379 26095 38421 26104
rect 38091 26060 38133 26069
rect 38091 26020 38092 26060
rect 38132 26020 38133 26060
rect 38091 26011 38133 26020
rect 37227 25892 37269 25901
rect 37227 25852 37228 25892
rect 37268 25852 37269 25892
rect 37227 25843 37269 25852
rect 38092 25481 38132 26011
rect 38091 25472 38133 25481
rect 38091 25432 38092 25472
rect 38132 25432 38133 25472
rect 38091 25423 38133 25432
rect 37227 25304 37269 25313
rect 37227 25264 37228 25304
rect 37268 25264 37269 25304
rect 37227 25255 37269 25264
rect 37612 25304 37652 25313
rect 37228 25170 37268 25255
rect 37035 24464 37077 24473
rect 37035 24424 37036 24464
rect 37076 24424 37077 24464
rect 37612 24464 37652 25264
rect 38380 25145 38420 26095
rect 38475 25892 38517 25901
rect 38475 25852 38476 25892
rect 38516 25852 38517 25892
rect 38475 25843 38517 25852
rect 38476 25304 38516 25843
rect 38476 25229 38516 25264
rect 38475 25220 38517 25229
rect 38475 25180 38476 25220
rect 38516 25180 38517 25220
rect 38475 25171 38517 25180
rect 38379 25136 38421 25145
rect 38476 25140 38516 25171
rect 38379 25096 38380 25136
rect 38420 25096 38421 25136
rect 38379 25087 38421 25096
rect 38572 24968 38612 26860
rect 38668 26851 38708 26860
rect 38859 26900 38901 26909
rect 38859 26860 38860 26900
rect 38900 26860 38901 26900
rect 38859 26851 38901 26860
rect 38956 26312 38996 27616
rect 39532 28288 39860 28328
rect 40204 28328 40244 28337
rect 39532 27152 39572 28288
rect 39820 28160 39860 28169
rect 39724 28120 39820 28160
rect 39627 27236 39669 27245
rect 39627 27196 39628 27236
rect 39668 27196 39669 27236
rect 39627 27187 39669 27196
rect 39148 27112 39572 27152
rect 39051 26900 39093 26909
rect 39051 26860 39052 26900
rect 39092 26860 39093 26900
rect 39051 26851 39093 26860
rect 39052 26766 39092 26851
rect 38860 26272 38996 26312
rect 39148 26312 39188 27112
rect 39436 26900 39476 26909
rect 39628 26900 39668 27187
rect 39476 26860 39668 26900
rect 39436 26851 39476 26860
rect 39724 26741 39764 28120
rect 39820 28111 39860 28120
rect 39819 27656 39861 27665
rect 39819 27616 39820 27656
rect 39860 27616 39861 27656
rect 39819 27607 39861 27616
rect 39820 26816 39860 27607
rect 40108 27404 40148 27413
rect 39820 26767 39860 26776
rect 39916 26816 39956 26827
rect 40108 26825 40148 27364
rect 40204 26900 40244 28288
rect 40395 28328 40437 28337
rect 40395 28288 40396 28328
rect 40436 28288 40437 28328
rect 40395 28279 40437 28288
rect 40492 28328 40532 28337
rect 40780 28328 40820 28876
rect 40532 28288 40820 28328
rect 40876 28328 40916 29632
rect 41068 29168 41108 31051
rect 41643 30764 41685 30773
rect 41643 30724 41644 30764
rect 41684 30724 41685 30764
rect 41643 30715 41685 30724
rect 41452 30680 41492 30691
rect 41452 30605 41492 30640
rect 41644 30680 41684 30715
rect 41644 30629 41684 30640
rect 41739 30680 41781 30689
rect 41739 30640 41740 30680
rect 41780 30640 41781 30680
rect 41739 30631 41781 30640
rect 41451 30596 41493 30605
rect 41451 30556 41452 30596
rect 41492 30556 41493 30596
rect 41451 30547 41493 30556
rect 41740 30546 41780 30631
rect 42124 30605 42164 32647
rect 42123 30596 42165 30605
rect 42123 30556 42124 30596
rect 42164 30556 42165 30596
rect 42123 30547 42165 30556
rect 41643 30512 41685 30521
rect 41643 30472 41644 30512
rect 41684 30472 41685 30512
rect 41643 30463 41685 30472
rect 41452 30428 41492 30437
rect 40972 29128 41068 29168
rect 40972 28421 41012 29128
rect 41068 29119 41108 29128
rect 41164 30388 41452 30428
rect 41067 29000 41109 29009
rect 41067 28960 41068 29000
rect 41108 28960 41109 29000
rect 41067 28951 41109 28960
rect 40971 28412 41013 28421
rect 40971 28372 40972 28412
rect 41012 28372 41013 28412
rect 40971 28363 41013 28372
rect 40492 28279 40532 28288
rect 40876 28279 40916 28288
rect 41068 28328 41108 28951
rect 41068 28279 41108 28288
rect 41164 28328 41204 30388
rect 41452 30379 41492 30388
rect 41356 29840 41396 29851
rect 41356 29765 41396 29800
rect 41548 29840 41588 29849
rect 41355 29756 41397 29765
rect 41355 29716 41356 29756
rect 41396 29716 41397 29756
rect 41355 29707 41397 29716
rect 41452 29756 41492 29765
rect 41452 29336 41492 29716
rect 41548 29681 41588 29800
rect 41547 29672 41589 29681
rect 41547 29632 41548 29672
rect 41588 29632 41589 29672
rect 41547 29623 41589 29632
rect 41260 29296 41492 29336
rect 41260 29009 41300 29296
rect 41356 29168 41396 29177
rect 41259 29000 41301 29009
rect 41259 28960 41260 29000
rect 41300 28960 41301 29000
rect 41259 28951 41301 28960
rect 41259 28412 41301 28421
rect 41259 28372 41260 28412
rect 41300 28372 41301 28412
rect 41259 28363 41301 28372
rect 41164 28279 41204 28288
rect 40971 28244 41013 28253
rect 40971 28204 40972 28244
rect 41012 28204 41013 28244
rect 40971 28195 41013 28204
rect 40300 28160 40340 28169
rect 40340 28120 40628 28160
rect 40300 28111 40340 28120
rect 40395 27740 40437 27749
rect 40395 27700 40396 27740
rect 40436 27700 40437 27740
rect 40395 27691 40437 27700
rect 40299 27656 40341 27665
rect 40299 27616 40300 27656
rect 40340 27616 40341 27656
rect 40299 27607 40341 27616
rect 40300 27522 40340 27607
rect 40396 27606 40436 27691
rect 40492 27656 40532 27665
rect 40492 27413 40532 27616
rect 40588 27656 40628 28120
rect 40972 28110 41012 28195
rect 40588 27607 40628 27616
rect 40971 27656 41013 27665
rect 40971 27616 40972 27656
rect 41012 27616 41013 27656
rect 40971 27607 41013 27616
rect 41164 27656 41204 27665
rect 40972 27522 41012 27607
rect 40491 27404 40533 27413
rect 40491 27364 40492 27404
rect 40532 27364 40533 27404
rect 40491 27355 40533 27364
rect 41067 27404 41109 27413
rect 41067 27364 41068 27404
rect 41108 27364 41109 27404
rect 41067 27355 41109 27364
rect 41068 27270 41108 27355
rect 40491 27152 40533 27161
rect 40491 27112 40492 27152
rect 40532 27112 40533 27152
rect 40491 27103 40533 27112
rect 40204 26860 40340 26900
rect 39916 26741 39956 26776
rect 40012 26816 40052 26825
rect 39723 26732 39765 26741
rect 39723 26692 39724 26732
rect 39764 26692 39765 26732
rect 39723 26683 39765 26692
rect 39915 26732 39957 26741
rect 39915 26692 39916 26732
rect 39956 26692 39957 26732
rect 39915 26683 39957 26692
rect 38860 25901 38900 26272
rect 39148 26263 39188 26272
rect 39244 26648 39284 26657
rect 39244 26237 39284 26608
rect 39627 26648 39669 26657
rect 39627 26608 39628 26648
rect 39668 26608 39669 26648
rect 39627 26599 39669 26608
rect 39628 26514 39668 26599
rect 39820 26237 39860 26281
rect 39243 26228 39285 26237
rect 39243 26188 39244 26228
rect 39284 26188 39285 26228
rect 39243 26179 39285 26188
rect 39819 26228 39861 26237
rect 40012 26228 40052 26776
rect 40107 26816 40149 26825
rect 40107 26776 40108 26816
rect 40148 26776 40149 26816
rect 40107 26767 40149 26776
rect 39819 26188 39820 26228
rect 39860 26188 39861 26228
rect 39819 26186 39861 26188
rect 39819 26179 39820 26186
rect 39340 26144 39380 26153
rect 39532 26144 39572 26153
rect 39380 26104 39476 26144
rect 39340 26095 39380 26104
rect 38955 26060 38997 26069
rect 38955 26020 38956 26060
rect 38996 26020 38997 26060
rect 38955 26011 38997 26020
rect 38956 25926 38996 26011
rect 38859 25892 38901 25901
rect 38859 25852 38860 25892
rect 38900 25852 38901 25892
rect 38859 25843 38901 25852
rect 39148 25892 39188 25901
rect 39148 25649 39188 25852
rect 39340 25892 39380 25901
rect 39147 25640 39189 25649
rect 39147 25600 39148 25640
rect 39188 25600 39189 25640
rect 39147 25591 39189 25600
rect 39148 25220 39188 25591
rect 39340 25313 39380 25852
rect 39436 25397 39476 26104
rect 39532 25733 39572 26104
rect 39628 26144 39668 26153
rect 39860 26179 39861 26186
rect 39916 26188 40052 26228
rect 39820 26137 39860 26146
rect 39628 26060 39668 26104
rect 39628 26020 39860 26060
rect 39820 25976 39860 26020
rect 39820 25927 39860 25936
rect 39531 25724 39573 25733
rect 39531 25684 39532 25724
rect 39572 25684 39573 25724
rect 39531 25675 39573 25684
rect 39531 25556 39573 25565
rect 39531 25516 39532 25556
rect 39572 25516 39573 25556
rect 39531 25507 39573 25516
rect 39435 25388 39477 25397
rect 39435 25348 39436 25388
rect 39476 25348 39477 25388
rect 39435 25339 39477 25348
rect 39339 25304 39381 25313
rect 39339 25264 39340 25304
rect 39380 25264 39381 25304
rect 39339 25255 39381 25264
rect 39532 25220 39572 25507
rect 39627 25304 39669 25313
rect 39627 25264 39628 25304
rect 39668 25264 39669 25304
rect 39627 25255 39669 25264
rect 39819 25304 39861 25313
rect 39819 25264 39820 25304
rect 39860 25264 39861 25304
rect 39819 25255 39861 25264
rect 39916 25304 39956 26188
rect 40108 26144 40148 26767
rect 40203 26732 40245 26741
rect 40203 26692 40204 26732
rect 40244 26692 40245 26732
rect 40203 26683 40245 26692
rect 40012 26130 40052 26139
rect 40108 26095 40148 26104
rect 40012 25565 40052 26090
rect 40011 25556 40053 25565
rect 40011 25516 40012 25556
rect 40052 25516 40053 25556
rect 40011 25507 40053 25516
rect 40107 25388 40149 25397
rect 40107 25348 40108 25388
rect 40148 25348 40149 25388
rect 40107 25339 40149 25348
rect 39148 25180 39284 25220
rect 39147 25052 39189 25061
rect 39147 25012 39148 25052
rect 39188 25012 39189 25052
rect 39147 25003 39189 25012
rect 38380 24928 38612 24968
rect 37995 24800 38037 24809
rect 37995 24760 37996 24800
rect 38036 24760 38037 24800
rect 37995 24751 38037 24760
rect 37708 24464 37748 24473
rect 37612 24424 37708 24464
rect 37035 24415 37077 24424
rect 37708 24415 37748 24424
rect 37036 23381 37076 24415
rect 37324 24380 37364 24389
rect 37324 23801 37364 24340
rect 37515 24128 37557 24137
rect 37515 24088 37516 24128
rect 37556 24088 37557 24128
rect 37515 24079 37557 24088
rect 37323 23792 37365 23801
rect 37323 23752 37324 23792
rect 37364 23752 37365 23792
rect 37323 23743 37365 23752
rect 37035 23372 37077 23381
rect 37035 23332 37036 23372
rect 37076 23332 37077 23372
rect 37035 23323 37077 23332
rect 37323 23204 37365 23213
rect 37323 23164 37324 23204
rect 37364 23164 37365 23204
rect 37323 23155 37365 23164
rect 37516 23204 37556 24079
rect 37899 23288 37941 23297
rect 37899 23248 37900 23288
rect 37940 23248 37941 23288
rect 37899 23239 37941 23248
rect 37516 23164 37844 23204
rect 37132 23120 37172 23129
rect 37132 23060 37172 23080
rect 36844 23020 36980 23060
rect 37036 23020 37172 23060
rect 37228 23120 37268 23129
rect 36747 22616 36789 22625
rect 36747 22576 36748 22616
rect 36788 22576 36789 22616
rect 36747 22567 36789 22576
rect 36844 22280 36884 23020
rect 36940 22952 36980 22961
rect 37036 22952 37076 23020
rect 36980 22912 37076 22952
rect 37131 22952 37173 22961
rect 37131 22912 37132 22952
rect 37172 22912 37173 22952
rect 36940 22903 36980 22912
rect 37131 22903 37173 22912
rect 36940 22280 36980 22289
rect 36844 22240 36940 22280
rect 36940 22231 36980 22240
rect 37132 22112 37172 22903
rect 37228 22625 37268 23080
rect 37324 23120 37364 23155
rect 37324 23069 37364 23080
rect 37227 22616 37269 22625
rect 37227 22576 37228 22616
rect 37268 22576 37269 22616
rect 37227 22567 37269 22576
rect 36652 22072 37172 22112
rect 36555 21776 36597 21785
rect 36555 21736 36556 21776
rect 36596 21736 36597 21776
rect 36555 21727 36597 21736
rect 35787 21608 35829 21617
rect 35787 21568 35788 21608
rect 35828 21568 35829 21608
rect 35787 21559 35829 21568
rect 36075 21608 36117 21617
rect 36075 21568 36076 21608
rect 36116 21568 36117 21608
rect 36075 21559 36117 21568
rect 36267 21608 36309 21617
rect 36267 21568 36268 21608
rect 36308 21568 36309 21608
rect 36267 21559 36309 21568
rect 36364 21608 36404 21617
rect 36171 21524 36213 21533
rect 36171 21484 36172 21524
rect 36212 21484 36213 21524
rect 36171 21475 36213 21484
rect 35692 21440 35732 21449
rect 35692 20768 35732 21400
rect 35692 20719 35732 20728
rect 35308 20684 35348 20693
rect 34636 20600 34676 20609
rect 34444 20560 34636 20600
rect 34444 19937 34484 20560
rect 34636 20551 34676 20560
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 35308 20264 35348 20644
rect 36075 20516 36117 20525
rect 36075 20476 36076 20516
rect 36116 20476 36117 20516
rect 36075 20467 36117 20476
rect 35692 20264 35732 20273
rect 35308 20224 35692 20264
rect 35692 20215 35732 20224
rect 34828 20096 34868 20105
rect 34828 19937 34868 20056
rect 34924 20096 34964 20105
rect 35116 20096 35156 20105
rect 34443 19928 34485 19937
rect 34443 19888 34444 19928
rect 34484 19888 34485 19928
rect 34443 19879 34485 19888
rect 34827 19928 34869 19937
rect 34827 19888 34828 19928
rect 34868 19888 34869 19928
rect 34827 19879 34869 19888
rect 34924 19685 34964 20056
rect 35020 20056 35116 20096
rect 35020 19853 35060 20056
rect 35116 20047 35156 20056
rect 35500 20096 35540 20105
rect 35116 19928 35156 19937
rect 35500 19928 35540 20056
rect 35156 19888 35540 19928
rect 35596 20096 35636 20105
rect 35116 19879 35156 19888
rect 35019 19844 35061 19853
rect 35019 19804 35020 19844
rect 35060 19804 35061 19844
rect 35019 19795 35061 19804
rect 34923 19676 34965 19685
rect 34923 19636 34924 19676
rect 34964 19636 34965 19676
rect 34923 19627 34965 19636
rect 35596 19508 35636 20056
rect 35788 20096 35828 20105
rect 35980 20096 36020 20105
rect 35828 20056 35980 20096
rect 35788 20047 35828 20056
rect 35980 20047 36020 20056
rect 36076 20096 36116 20467
rect 36076 20047 36116 20056
rect 36172 20096 36212 21475
rect 36268 21474 36308 21559
rect 36364 21440 36404 21568
rect 36459 21608 36501 21617
rect 36459 21568 36460 21608
rect 36500 21568 36501 21608
rect 36459 21559 36501 21568
rect 36556 21608 36596 21617
rect 36652 21608 36692 22072
rect 36747 21692 36789 21701
rect 36747 21652 36748 21692
rect 36788 21652 36789 21692
rect 36747 21643 36789 21652
rect 36596 21568 36692 21608
rect 36748 21608 36788 21643
rect 36556 21559 36596 21568
rect 36748 21557 36788 21568
rect 36652 21440 36692 21449
rect 36364 21400 36652 21440
rect 36652 21391 36692 21400
rect 36556 20768 36596 20777
rect 36172 20047 36212 20056
rect 36268 20096 36308 20105
rect 36268 19937 36308 20056
rect 36267 19928 36309 19937
rect 36267 19888 36268 19928
rect 36308 19888 36309 19928
rect 36267 19879 36309 19888
rect 35788 19508 35828 19517
rect 35596 19468 35788 19508
rect 35692 19256 35732 19265
rect 35596 19216 35692 19256
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 35307 18668 35349 18677
rect 35307 18628 35308 18668
rect 35348 18628 35349 18668
rect 35307 18619 35349 18628
rect 34156 18509 34196 18544
rect 34251 18584 34293 18593
rect 34251 18544 34252 18584
rect 34292 18544 34293 18584
rect 34251 18535 34293 18544
rect 34155 18500 34197 18509
rect 34155 18460 34156 18500
rect 34196 18460 34197 18500
rect 34155 18451 34197 18460
rect 35308 18500 35348 18619
rect 35308 18451 35348 18460
rect 35499 18500 35541 18509
rect 35499 18460 35500 18500
rect 35540 18460 35541 18500
rect 35499 18451 35541 18460
rect 34156 18420 34196 18451
rect 34828 17912 34868 17921
rect 34868 17872 35060 17912
rect 34828 17863 34868 17872
rect 34347 17828 34389 17837
rect 34347 17788 34348 17828
rect 34388 17788 34389 17828
rect 34347 17779 34389 17788
rect 34348 17694 34388 17779
rect 34156 17576 34196 17585
rect 34060 17536 34156 17576
rect 33963 17324 34005 17333
rect 33963 17284 33964 17324
rect 34004 17284 34005 17324
rect 33963 17275 34005 17284
rect 33580 17081 33620 17166
rect 34060 17165 34100 17536
rect 34156 17527 34196 17536
rect 34347 17576 34389 17585
rect 34347 17536 34348 17576
rect 34388 17536 34389 17576
rect 34347 17527 34389 17536
rect 34059 17156 34101 17165
rect 34059 17116 34060 17156
rect 34100 17116 34101 17156
rect 34059 17107 34101 17116
rect 33388 17072 33428 17081
rect 33196 17032 33388 17072
rect 33003 16316 33045 16325
rect 33003 16276 33004 16316
rect 33044 16276 33045 16316
rect 33003 16267 33045 16276
rect 33196 15737 33236 17032
rect 33388 17023 33428 17032
rect 33579 17072 33621 17081
rect 33579 17032 33580 17072
rect 33620 17032 33621 17072
rect 33579 17023 33621 17032
rect 33772 17072 33812 17081
rect 33484 16904 33524 16913
rect 33772 16904 33812 17032
rect 33524 16864 33812 16904
rect 33868 17072 33908 17081
rect 33484 16855 33524 16864
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 33868 16493 33908 17032
rect 34060 17072 34100 17107
rect 34060 17021 34100 17032
rect 34252 17072 34292 17081
rect 34060 16904 34100 16913
rect 34252 16904 34292 17032
rect 34100 16864 34292 16904
rect 34060 16855 34100 16864
rect 34059 16736 34101 16745
rect 34059 16696 34060 16736
rect 34100 16696 34101 16736
rect 34059 16687 34101 16696
rect 33867 16484 33909 16493
rect 33867 16444 33868 16484
rect 33908 16444 33909 16484
rect 33867 16435 33909 16444
rect 33771 16316 33813 16325
rect 33771 16276 33772 16316
rect 33812 16276 33813 16316
rect 33771 16267 33813 16276
rect 33772 16232 33812 16267
rect 33772 16181 33812 16192
rect 34060 16232 34100 16687
rect 34251 16484 34293 16493
rect 34251 16444 34252 16484
rect 34292 16444 34293 16484
rect 34251 16435 34293 16444
rect 34060 16183 34100 16192
rect 34156 16148 34196 16157
rect 33484 16064 33524 16073
rect 34156 16064 34196 16108
rect 33484 15980 33524 16024
rect 33868 16024 34196 16064
rect 33868 15980 33908 16024
rect 34252 15980 34292 16435
rect 33388 15940 33908 15980
rect 34060 15940 34292 15980
rect 33195 15728 33237 15737
rect 33195 15688 33196 15728
rect 33236 15688 33237 15728
rect 33195 15679 33237 15688
rect 33388 15560 33428 15940
rect 33963 15896 34005 15905
rect 33963 15856 33964 15896
rect 34004 15856 34005 15896
rect 33963 15847 34005 15856
rect 33483 15812 33525 15821
rect 33483 15772 33484 15812
rect 33524 15772 33525 15812
rect 33483 15763 33525 15772
rect 33196 15520 33388 15560
rect 32907 14972 32949 14981
rect 32907 14932 32908 14972
rect 32948 14932 32949 14972
rect 33196 14972 33236 15520
rect 33388 15511 33428 15520
rect 33484 15560 33524 15763
rect 33964 15728 34004 15847
rect 33964 15679 34004 15688
rect 33484 15308 33524 15520
rect 33580 15560 33620 15571
rect 33580 15485 33620 15520
rect 33676 15560 33716 15569
rect 33868 15560 33908 15569
rect 33716 15520 33868 15560
rect 33676 15511 33716 15520
rect 33868 15511 33908 15520
rect 34060 15560 34100 15940
rect 34348 15569 34388 17527
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 34636 17072 34676 17081
rect 35020 17072 35060 17872
rect 35115 17324 35157 17333
rect 35115 17284 35116 17324
rect 35156 17284 35157 17324
rect 35115 17275 35157 17284
rect 34676 17032 35060 17072
rect 34636 17023 34676 17032
rect 35116 16988 35156 17275
rect 35500 17072 35540 18451
rect 35596 17333 35636 19216
rect 35692 19207 35732 19216
rect 35788 19004 35828 19468
rect 36076 19424 36116 19433
rect 35884 19256 35924 19265
rect 36076 19256 36116 19384
rect 35924 19216 36116 19256
rect 36268 19256 36308 19879
rect 36364 19256 36404 19265
rect 36268 19216 36364 19256
rect 35884 19207 35924 19216
rect 36364 19207 36404 19216
rect 36460 19256 36500 19265
rect 36460 19088 36500 19216
rect 36364 19048 36500 19088
rect 35788 18964 35924 19004
rect 35787 18668 35829 18677
rect 35787 18628 35788 18668
rect 35828 18628 35829 18668
rect 35787 18619 35829 18628
rect 35691 18584 35733 18593
rect 35691 18544 35692 18584
rect 35732 18544 35733 18584
rect 35691 18535 35733 18544
rect 35692 18425 35732 18535
rect 35788 18534 35828 18619
rect 35884 18584 35924 18964
rect 36171 18668 36213 18677
rect 36171 18628 36172 18668
rect 36212 18628 36213 18668
rect 36171 18619 36213 18628
rect 35884 18535 35924 18544
rect 35980 18584 36020 18593
rect 36020 18544 36116 18584
rect 35980 18535 36020 18544
rect 35691 18416 35733 18425
rect 35691 18376 35692 18416
rect 35732 18376 35733 18416
rect 35691 18367 35733 18376
rect 36076 18080 36116 18544
rect 36172 18534 36212 18619
rect 36364 18257 36404 19048
rect 36556 19004 36596 20728
rect 37516 19853 37556 23164
rect 37804 23120 37844 23164
rect 37900 23154 37940 23239
rect 37804 23071 37844 23080
rect 37996 23120 38036 24751
rect 38091 23792 38133 23801
rect 38091 23752 38092 23792
rect 38132 23752 38133 23792
rect 38091 23743 38133 23752
rect 37611 23060 37653 23069
rect 37611 23020 37612 23060
rect 37652 23020 37653 23060
rect 37611 23011 37653 23020
rect 37612 20273 37652 23011
rect 37996 22961 38036 23080
rect 38092 23120 38132 23743
rect 38092 23071 38132 23080
rect 37995 22952 38037 22961
rect 37995 22912 37996 22952
rect 38036 22912 38037 22952
rect 37995 22903 38037 22912
rect 38091 22196 38133 22205
rect 38091 22156 38092 22196
rect 38132 22156 38133 22196
rect 38091 22147 38133 22156
rect 38092 22112 38132 22147
rect 38092 21701 38132 22072
rect 38091 21692 38133 21701
rect 38091 21652 38092 21692
rect 38132 21652 38133 21692
rect 38091 21643 38133 21652
rect 38380 21113 38420 24928
rect 39148 24800 39188 25003
rect 39148 24751 39188 24760
rect 39244 24548 39284 25180
rect 39436 25180 39572 25220
rect 39340 24548 39380 24557
rect 39244 24508 39340 24548
rect 39340 24499 39380 24508
rect 39243 24128 39285 24137
rect 39243 24088 39244 24128
rect 39284 24088 39285 24128
rect 39243 24079 39285 24088
rect 38859 23960 38901 23969
rect 38859 23920 38860 23960
rect 38900 23920 38901 23960
rect 38859 23911 38901 23920
rect 38763 23792 38805 23801
rect 38763 23752 38764 23792
rect 38804 23752 38805 23792
rect 38763 23743 38805 23752
rect 38860 23792 38900 23911
rect 38860 23743 38900 23752
rect 38956 23792 38996 23801
rect 38764 23658 38804 23743
rect 38956 23633 38996 23752
rect 39244 23792 39284 24079
rect 39244 23743 39284 23752
rect 39436 23792 39476 25180
rect 39628 25136 39668 25255
rect 39723 25220 39765 25229
rect 39723 25180 39724 25220
rect 39764 25180 39765 25220
rect 39723 25171 39765 25180
rect 39052 23708 39092 23717
rect 38955 23624 38997 23633
rect 38955 23584 38956 23624
rect 38996 23584 38997 23624
rect 38955 23575 38997 23584
rect 38476 23129 38516 23214
rect 38475 23120 38517 23129
rect 38475 23080 38476 23120
rect 38516 23080 38517 23120
rect 38475 23071 38517 23080
rect 38860 23120 38900 23129
rect 38860 22448 38900 23080
rect 39052 22700 39092 23668
rect 39340 23624 39380 23633
rect 39147 23120 39189 23129
rect 39147 23080 39148 23120
rect 39188 23080 39189 23120
rect 39147 23071 39189 23080
rect 38860 22399 38900 22408
rect 38956 22660 39092 22700
rect 38956 22280 38996 22660
rect 39052 22532 39092 22541
rect 39148 22532 39188 23071
rect 39092 22492 39188 22532
rect 39052 22483 39092 22492
rect 39052 22280 39092 22289
rect 38956 22240 39052 22280
rect 39052 22231 39092 22240
rect 39243 22280 39285 22289
rect 39243 22240 39244 22280
rect 39284 22240 39285 22280
rect 39243 22231 39285 22240
rect 39340 22280 39380 23584
rect 39436 23060 39476 23752
rect 39532 25096 39628 25136
rect 39532 23792 39572 25096
rect 39628 25087 39668 25096
rect 39628 24632 39668 24641
rect 39628 24473 39668 24592
rect 39627 24464 39669 24473
rect 39627 24424 39628 24464
rect 39668 24424 39669 24464
rect 39627 24415 39669 24424
rect 39532 23743 39572 23752
rect 39724 23120 39764 25171
rect 39820 24800 39860 25255
rect 39916 25061 39956 25264
rect 40012 25304 40052 25315
rect 40012 25229 40052 25264
rect 40108 25304 40148 25339
rect 40108 25253 40148 25264
rect 40204 25229 40244 26683
rect 40300 26237 40340 26860
rect 40396 26816 40436 26827
rect 40396 26741 40436 26776
rect 40395 26732 40437 26741
rect 40395 26692 40396 26732
rect 40436 26692 40437 26732
rect 40395 26683 40437 26692
rect 40299 26228 40341 26237
rect 40299 26188 40300 26228
rect 40340 26188 40341 26228
rect 40299 26179 40341 26188
rect 40011 25220 40053 25229
rect 40011 25180 40012 25220
rect 40052 25180 40053 25220
rect 40011 25171 40053 25180
rect 40203 25220 40245 25229
rect 40203 25180 40204 25220
rect 40244 25180 40245 25220
rect 40203 25171 40245 25180
rect 39915 25052 39957 25061
rect 40300 25052 40340 26179
rect 40492 26060 40532 27103
rect 40875 27068 40917 27077
rect 40875 27028 40876 27068
rect 40916 27028 40917 27068
rect 40875 27019 40917 27028
rect 41068 27068 41108 27077
rect 41164 27068 41204 27616
rect 41260 27488 41300 28363
rect 41356 28328 41396 29128
rect 41451 29168 41493 29177
rect 41451 29128 41452 29168
rect 41492 29128 41493 29168
rect 41451 29119 41493 29128
rect 41452 29034 41492 29119
rect 41547 28664 41589 28673
rect 41547 28624 41548 28664
rect 41588 28624 41589 28664
rect 41547 28615 41589 28624
rect 41451 28580 41493 28589
rect 41451 28540 41452 28580
rect 41492 28540 41493 28580
rect 41451 28531 41493 28540
rect 41452 28446 41492 28531
rect 41356 27833 41396 28288
rect 41451 28328 41493 28337
rect 41451 28288 41452 28328
rect 41492 28288 41493 28328
rect 41451 28279 41493 28288
rect 41548 28328 41588 28615
rect 41355 27824 41397 27833
rect 41355 27784 41356 27824
rect 41396 27784 41397 27824
rect 41355 27775 41397 27784
rect 41356 27488 41396 27497
rect 41260 27448 41356 27488
rect 41260 27245 41300 27448
rect 41356 27439 41396 27448
rect 41259 27236 41301 27245
rect 41259 27196 41260 27236
rect 41300 27196 41301 27236
rect 41259 27187 41301 27196
rect 41108 27028 41204 27068
rect 41068 27019 41108 27028
rect 40684 26816 40724 26825
rect 40684 26405 40724 26776
rect 40779 26816 40821 26825
rect 40779 26776 40780 26816
rect 40820 26776 40821 26816
rect 40779 26767 40821 26776
rect 40780 26682 40820 26767
rect 40683 26396 40725 26405
rect 40683 26356 40684 26396
rect 40724 26356 40725 26396
rect 40683 26347 40725 26356
rect 40492 26011 40532 26020
rect 40684 25976 40724 25985
rect 40876 25976 40916 27019
rect 41452 26993 41492 28279
rect 41548 28253 41588 28288
rect 41547 28244 41589 28253
rect 41547 28204 41548 28244
rect 41588 28204 41589 28244
rect 41547 28195 41589 28204
rect 41548 27572 41588 27581
rect 41548 27413 41588 27532
rect 41547 27404 41589 27413
rect 41547 27364 41548 27404
rect 41588 27364 41589 27404
rect 41547 27355 41589 27364
rect 41451 26984 41493 26993
rect 41260 26944 41452 26984
rect 41492 26944 41493 26984
rect 41260 26816 41300 26944
rect 41451 26935 41493 26944
rect 41644 26909 41684 30463
rect 42220 30353 42260 32899
rect 42700 32814 42740 32899
rect 42891 32696 42933 32705
rect 42891 32656 42892 32696
rect 42932 32656 42933 32696
rect 42891 32647 42933 32656
rect 42892 32562 42932 32647
rect 42411 32528 42453 32537
rect 42411 32488 42412 32528
rect 42452 32488 42453 32528
rect 42411 32479 42453 32488
rect 42316 32192 42356 32201
rect 42316 31193 42356 32152
rect 42412 32192 42452 32479
rect 42315 31184 42357 31193
rect 42315 31144 42316 31184
rect 42356 31144 42357 31184
rect 42315 31135 42357 31144
rect 42315 30596 42357 30605
rect 42315 30556 42316 30596
rect 42356 30556 42357 30596
rect 42315 30547 42357 30556
rect 42219 30344 42261 30353
rect 42219 30304 42220 30344
rect 42260 30304 42261 30344
rect 42219 30295 42261 30304
rect 42123 30008 42165 30017
rect 42123 29968 42124 30008
rect 42164 29968 42165 30008
rect 42123 29959 42165 29968
rect 41835 29756 41877 29765
rect 41835 29716 41836 29756
rect 41876 29716 41877 29756
rect 41835 29707 41877 29716
rect 41739 29672 41781 29681
rect 41739 29632 41740 29672
rect 41780 29632 41781 29672
rect 41739 29623 41781 29632
rect 41740 29000 41780 29623
rect 41740 28951 41780 28960
rect 41739 28832 41781 28841
rect 41739 28792 41740 28832
rect 41780 28792 41781 28832
rect 41739 28783 41781 28792
rect 41740 28328 41780 28783
rect 41740 28279 41780 28288
rect 41836 28160 41876 29707
rect 41932 29168 41972 29177
rect 41932 28589 41972 29128
rect 42028 29168 42068 29177
rect 42028 29009 42068 29128
rect 42124 29168 42164 29959
rect 42220 29168 42260 29177
rect 42124 29128 42220 29168
rect 42027 29000 42069 29009
rect 42027 28960 42028 29000
rect 42068 28960 42069 29000
rect 42027 28951 42069 28960
rect 41931 28580 41973 28589
rect 41931 28540 41932 28580
rect 41972 28540 41973 28580
rect 41931 28531 41973 28540
rect 42124 28496 42164 29128
rect 42220 29119 42260 29128
rect 42219 28916 42261 28925
rect 42219 28876 42220 28916
rect 42260 28876 42261 28916
rect 42219 28867 42261 28876
rect 42220 28782 42260 28867
rect 42316 28757 42356 30547
rect 42412 29849 42452 32152
rect 42508 32192 42548 32201
rect 42508 31025 42548 32152
rect 42604 32192 42644 32201
rect 42892 32192 42932 32201
rect 42644 32152 42740 32192
rect 42604 32143 42644 32152
rect 42603 31184 42645 31193
rect 42603 31144 42604 31184
rect 42644 31144 42645 31184
rect 42603 31135 42645 31144
rect 42507 31016 42549 31025
rect 42507 30976 42508 31016
rect 42548 30976 42549 31016
rect 42507 30967 42549 30976
rect 42508 30848 42548 30967
rect 42508 30799 42548 30808
rect 42604 30689 42644 31135
rect 42603 30680 42645 30689
rect 42603 30640 42604 30680
rect 42644 30640 42645 30680
rect 42603 30631 42645 30640
rect 42700 30680 42740 32152
rect 42796 32152 42892 32192
rect 42796 31604 42836 32152
rect 42892 32143 42932 32152
rect 43084 32192 43124 32201
rect 42988 31940 43028 31949
rect 42796 31555 42836 31564
rect 42892 31900 42988 31940
rect 42892 31277 42932 31900
rect 42988 31891 43028 31900
rect 43084 31436 43124 32152
rect 43372 32192 43412 32201
rect 43756 32192 43796 32201
rect 43852 32192 43892 32992
rect 46252 32957 46292 34336
rect 46444 34376 46484 34385
rect 46636 34376 46676 34504
rect 46484 34336 46580 34376
rect 46444 34327 46484 34336
rect 46540 33872 46580 34336
rect 46636 34327 46676 34336
rect 47020 34376 47060 34385
rect 47116 34376 47156 35008
rect 48556 34964 48596 34973
rect 48596 34924 48980 34964
rect 48556 34915 48596 34924
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 48940 34385 48980 34924
rect 49228 34553 49268 34638
rect 49227 34544 49269 34553
rect 49227 34504 49228 34544
rect 49268 34504 49269 34544
rect 49227 34495 49269 34504
rect 47060 34336 47156 34376
rect 47884 34376 47924 34385
rect 48939 34376 48981 34385
rect 47924 34336 48020 34376
rect 47020 34327 47060 34336
rect 47884 34327 47924 34336
rect 47019 34208 47061 34217
rect 47019 34168 47020 34208
rect 47060 34168 47061 34208
rect 47019 34159 47061 34168
rect 46732 33872 46772 33881
rect 46540 33832 46732 33872
rect 46732 33823 46772 33832
rect 46828 33704 46868 33713
rect 46636 33664 46828 33704
rect 46636 33140 46676 33664
rect 46828 33655 46868 33664
rect 46924 33704 46964 33713
rect 46827 33200 46869 33209
rect 46827 33160 46828 33200
rect 46868 33160 46869 33200
rect 46827 33151 46869 33160
rect 46348 33100 46676 33140
rect 46059 32948 46101 32957
rect 46059 32908 46060 32948
rect 46100 32908 46101 32948
rect 46059 32899 46101 32908
rect 46251 32948 46293 32957
rect 46251 32908 46252 32948
rect 46292 32908 46293 32948
rect 46251 32899 46293 32908
rect 45868 32864 45908 32873
rect 44715 32528 44757 32537
rect 44715 32488 44716 32528
rect 44756 32488 44757 32528
rect 44715 32479 44757 32488
rect 43412 32152 43700 32192
rect 43372 32143 43412 32152
rect 43660 31688 43700 32152
rect 43796 32152 43892 32192
rect 44619 32192 44661 32201
rect 44619 32152 44620 32192
rect 44660 32152 44661 32192
rect 43756 32143 43796 32152
rect 44619 32143 44661 32152
rect 44620 32058 44660 32143
rect 43660 31648 44084 31688
rect 44044 31604 44084 31648
rect 44044 31555 44084 31564
rect 42988 31396 43124 31436
rect 42891 31268 42933 31277
rect 42891 31228 42892 31268
rect 42932 31228 42933 31268
rect 42891 31219 42933 31228
rect 42795 30848 42837 30857
rect 42795 30808 42796 30848
rect 42836 30808 42837 30848
rect 42795 30799 42837 30808
rect 42796 30714 42836 30799
rect 42700 30631 42740 30640
rect 42892 30680 42932 31219
rect 42988 30848 43028 31396
rect 43468 31352 43508 31363
rect 43756 31352 43796 31361
rect 43180 31325 43220 31334
rect 43084 31268 43124 31279
rect 43084 31193 43124 31228
rect 43083 31184 43125 31193
rect 43083 31144 43084 31184
rect 43124 31144 43125 31184
rect 43083 31135 43125 31144
rect 43180 31100 43220 31285
rect 43468 31277 43508 31312
rect 43564 31312 43756 31352
rect 43467 31268 43509 31277
rect 43467 31228 43468 31268
rect 43508 31228 43509 31268
rect 43467 31219 43509 31228
rect 43468 31109 43508 31219
rect 43179 30941 43220 31100
rect 43467 31100 43509 31109
rect 43467 31060 43468 31100
rect 43508 31060 43509 31100
rect 43467 31051 43509 31060
rect 43179 30932 43221 30941
rect 43564 30932 43604 31312
rect 43756 31303 43796 31312
rect 43852 31352 43892 31361
rect 44044 31352 44084 31361
rect 43852 31193 43892 31312
rect 43948 31312 44044 31352
rect 43851 31184 43893 31193
rect 43851 31144 43852 31184
rect 43892 31144 43893 31184
rect 43851 31135 43893 31144
rect 43179 30892 43180 30932
rect 43220 30892 43221 30932
rect 43179 30883 43221 30892
rect 43276 30892 43604 30932
rect 42988 30808 43124 30848
rect 42892 30631 42932 30640
rect 42988 30680 43028 30689
rect 42988 30521 43028 30640
rect 42987 30512 43029 30521
rect 42987 30472 42988 30512
rect 43028 30472 43029 30512
rect 42987 30463 43029 30472
rect 42507 30428 42549 30437
rect 42507 30388 42508 30428
rect 42548 30388 42549 30428
rect 42507 30379 42549 30388
rect 42508 30294 42548 30379
rect 42795 30344 42837 30353
rect 42795 30304 42796 30344
rect 42836 30304 42837 30344
rect 42795 30295 42837 30304
rect 42411 29840 42453 29849
rect 42411 29800 42412 29840
rect 42452 29800 42453 29840
rect 42411 29791 42453 29800
rect 42412 29000 42452 29009
rect 42315 28748 42357 28757
rect 42315 28708 42316 28748
rect 42356 28708 42357 28748
rect 42315 28699 42357 28708
rect 41740 28120 41876 28160
rect 42028 28456 42164 28496
rect 41740 27077 41780 28120
rect 41739 27068 41781 27077
rect 41739 27028 41740 27068
rect 41780 27028 41781 27068
rect 41739 27019 41781 27028
rect 42028 26984 42068 28456
rect 42124 28328 42164 28337
rect 42412 28328 42452 28960
rect 42164 28288 42452 28328
rect 42124 28279 42164 28288
rect 42603 28244 42645 28253
rect 42603 28204 42604 28244
rect 42644 28204 42645 28244
rect 42603 28195 42645 28204
rect 42028 26944 42260 26984
rect 41643 26900 41685 26909
rect 41643 26860 41644 26900
rect 41684 26860 41685 26900
rect 41643 26851 41685 26860
rect 41068 26776 41260 26816
rect 41068 25976 41108 26776
rect 41260 26767 41300 26776
rect 41356 26816 41396 26825
rect 41356 26396 41396 26776
rect 41452 26816 41492 26825
rect 41452 26405 41492 26776
rect 42028 26816 42068 26825
rect 42068 26776 42164 26816
rect 42028 26767 42068 26776
rect 41644 26732 41684 26741
rect 41164 26356 41396 26396
rect 41451 26396 41493 26405
rect 41451 26356 41452 26396
rect 41492 26356 41493 26396
rect 41164 26144 41204 26356
rect 41451 26347 41493 26356
rect 41164 26095 41204 26104
rect 41259 26144 41301 26153
rect 41452 26144 41492 26153
rect 41259 26104 41260 26144
rect 41300 26104 41301 26144
rect 41259 26095 41301 26104
rect 41356 26104 41452 26144
rect 41260 26010 41300 26095
rect 40724 25936 40916 25976
rect 40972 25936 41108 25976
rect 40684 25808 40724 25936
rect 40588 25768 40724 25808
rect 40588 25640 40628 25768
rect 40779 25724 40821 25733
rect 40684 25684 40780 25724
rect 40820 25684 40821 25724
rect 40588 25600 40632 25640
rect 40395 25556 40437 25565
rect 40592 25556 40632 25600
rect 40395 25516 40396 25556
rect 40436 25516 40437 25556
rect 40395 25507 40437 25516
rect 40588 25516 40632 25556
rect 40396 25422 40436 25507
rect 40588 25387 40628 25516
rect 40588 25338 40628 25347
rect 39915 25012 39916 25052
rect 39956 25012 39957 25052
rect 39915 25003 39957 25012
rect 40108 25012 40340 25052
rect 39820 24760 40052 24800
rect 40012 24716 40052 24760
rect 40012 24667 40052 24676
rect 39915 24632 39957 24641
rect 39915 24592 39916 24632
rect 39956 24592 39957 24632
rect 39915 24583 39957 24592
rect 39916 24498 39956 24583
rect 40011 24464 40053 24473
rect 40011 24424 40012 24464
rect 40052 24424 40053 24464
rect 40011 24415 40053 24424
rect 39436 23020 39572 23060
rect 39340 22231 39380 22240
rect 39244 22146 39284 22231
rect 38956 21608 38996 21617
rect 38379 21104 38421 21113
rect 38379 21064 38380 21104
rect 38420 21064 38421 21104
rect 38379 21055 38421 21064
rect 38380 20945 38420 21055
rect 38379 20936 38421 20945
rect 38379 20896 38380 20936
rect 38420 20896 38421 20936
rect 38379 20887 38421 20896
rect 38476 20936 38516 20945
rect 38516 20896 38708 20936
rect 38476 20887 38516 20896
rect 38188 20768 38228 20777
rect 37708 20600 37748 20609
rect 37611 20264 37653 20273
rect 37611 20224 37612 20264
rect 37652 20224 37653 20264
rect 37611 20215 37653 20224
rect 37708 20096 37748 20560
rect 37996 20264 38036 20273
rect 38188 20264 38228 20728
rect 38284 20768 38324 20777
rect 38475 20768 38517 20777
rect 38324 20728 38420 20768
rect 38284 20719 38324 20728
rect 38036 20224 38228 20264
rect 38283 20264 38325 20273
rect 38283 20224 38284 20264
rect 38324 20224 38325 20264
rect 37996 20215 38036 20224
rect 38283 20215 38325 20224
rect 37804 20096 37844 20105
rect 37708 20056 37804 20096
rect 37708 19937 37748 20056
rect 37804 20047 37844 20056
rect 37900 20096 37940 20105
rect 37707 19928 37749 19937
rect 37707 19888 37708 19928
rect 37748 19888 37749 19928
rect 37707 19879 37749 19888
rect 37515 19844 37557 19853
rect 37515 19804 37516 19844
rect 37556 19804 37557 19844
rect 37515 19795 37557 19804
rect 37900 19685 37940 20056
rect 38092 20096 38132 20105
rect 38284 20096 38324 20215
rect 38092 19937 38132 20056
rect 38188 20056 38284 20096
rect 38091 19928 38133 19937
rect 38091 19888 38092 19928
rect 38132 19888 38133 19928
rect 38091 19879 38133 19888
rect 37899 19676 37941 19685
rect 37899 19636 37900 19676
rect 37940 19636 37941 19676
rect 37899 19627 37941 19636
rect 37036 19424 37076 19433
rect 36460 18964 36596 19004
rect 36652 19384 37036 19424
rect 36460 18509 36500 18964
rect 36556 18584 36596 18593
rect 36652 18584 36692 19384
rect 37036 19375 37076 19384
rect 36596 18544 36692 18584
rect 36748 19256 36788 19265
rect 36556 18535 36596 18544
rect 36459 18500 36501 18509
rect 36459 18460 36460 18500
rect 36500 18460 36501 18500
rect 36459 18451 36501 18460
rect 36363 18248 36405 18257
rect 36363 18208 36364 18248
rect 36404 18208 36405 18248
rect 36363 18199 36405 18208
rect 36651 18248 36693 18257
rect 36651 18208 36652 18248
rect 36692 18208 36693 18248
rect 36651 18199 36693 18208
rect 36076 18040 36596 18080
rect 36556 17996 36596 18040
rect 36556 17947 36596 17956
rect 36459 17912 36501 17921
rect 36459 17872 36460 17912
rect 36500 17872 36501 17912
rect 36459 17863 36501 17872
rect 36460 17744 36500 17863
rect 36460 17695 36500 17704
rect 36652 17744 36692 18199
rect 36652 17695 36692 17704
rect 35595 17324 35637 17333
rect 35595 17284 35596 17324
rect 35636 17284 35637 17324
rect 35595 17275 35637 17284
rect 35500 17023 35540 17032
rect 34828 16948 35156 16988
rect 34731 16484 34773 16493
rect 34731 16444 34732 16484
rect 34772 16444 34773 16484
rect 34731 16435 34773 16444
rect 34444 16400 34484 16409
rect 34484 16360 34676 16400
rect 34444 16351 34484 16360
rect 34636 16232 34676 16360
rect 34732 16350 34772 16435
rect 34636 16183 34676 16192
rect 34828 16232 34868 16948
rect 36651 16820 36693 16829
rect 36651 16780 36652 16820
rect 36692 16780 36693 16820
rect 36651 16771 36693 16780
rect 36652 16686 36692 16771
rect 36748 16316 36788 19216
rect 37420 18584 37460 18595
rect 37420 18509 37460 18544
rect 37419 18500 37461 18509
rect 37419 18460 37420 18500
rect 37460 18460 37461 18500
rect 37419 18451 37461 18460
rect 37035 17996 37077 18005
rect 37035 17956 37036 17996
rect 37076 17956 37077 17996
rect 37035 17947 37077 17956
rect 37036 17862 37076 17947
rect 37900 17912 37940 17921
rect 36843 17828 36885 17837
rect 36843 17788 36844 17828
rect 36884 17788 36885 17828
rect 36843 17779 36885 17788
rect 36844 17501 36884 17779
rect 37036 17576 37076 17585
rect 36843 17492 36885 17501
rect 36843 17452 36844 17492
rect 36884 17452 36885 17492
rect 36843 17443 36885 17452
rect 36940 17072 36980 17081
rect 37036 17072 37076 17536
rect 36980 17032 37076 17072
rect 37132 17072 37172 17081
rect 36844 16325 36884 16344
rect 36843 16316 36885 16325
rect 36748 16276 36844 16316
rect 36884 16276 36885 16316
rect 36843 16267 36885 16276
rect 36844 16249 36884 16267
rect 36844 16200 36884 16209
rect 34828 16183 34868 16192
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 35595 15812 35637 15821
rect 35595 15772 35596 15812
rect 35636 15772 35637 15812
rect 35595 15763 35637 15772
rect 36363 15812 36405 15821
rect 36940 15812 36980 17032
rect 37132 16913 37172 17032
rect 37324 17072 37364 17081
rect 37131 16904 37173 16913
rect 37131 16864 37132 16904
rect 37172 16864 37173 16904
rect 37131 16855 37173 16864
rect 37036 16820 37076 16829
rect 37036 16241 37076 16780
rect 37035 16232 37077 16241
rect 37035 16192 37036 16232
rect 37076 16192 37077 16232
rect 37035 16183 37077 16192
rect 37132 16232 37172 16855
rect 37324 16493 37364 17032
rect 37708 17072 37748 17081
rect 37900 17072 37940 17872
rect 38091 17156 38133 17165
rect 38091 17116 38092 17156
rect 38132 17116 38133 17156
rect 38091 17107 38133 17116
rect 37748 17032 37940 17072
rect 37708 17023 37748 17032
rect 37323 16484 37365 16493
rect 37323 16444 37324 16484
rect 37364 16444 37365 16484
rect 37323 16435 37365 16444
rect 37995 16484 38037 16493
rect 37995 16444 37996 16484
rect 38036 16444 38037 16484
rect 37995 16435 38037 16444
rect 37515 16400 37557 16409
rect 37515 16360 37516 16400
rect 37556 16360 37557 16400
rect 37515 16351 37557 16360
rect 37516 16266 37556 16351
rect 37996 16350 38036 16435
rect 37132 16183 37172 16192
rect 37707 16232 37749 16241
rect 37707 16192 37708 16232
rect 37748 16192 37749 16232
rect 37707 16183 37749 16192
rect 37804 16232 37844 16241
rect 36363 15772 36364 15812
rect 36404 15772 36405 15812
rect 36363 15763 36405 15772
rect 36844 15772 36980 15812
rect 37228 16148 37268 16157
rect 34827 15728 34869 15737
rect 34827 15688 34828 15728
rect 34868 15688 34869 15728
rect 34827 15679 34869 15688
rect 35211 15728 35253 15737
rect 35211 15688 35212 15728
rect 35252 15688 35253 15728
rect 34060 15511 34100 15520
rect 34156 15560 34196 15569
rect 33579 15476 33621 15485
rect 33579 15436 33580 15476
rect 33620 15436 33621 15476
rect 33579 15427 33621 15436
rect 34156 15401 34196 15520
rect 34347 15560 34389 15569
rect 34347 15520 34348 15560
rect 34388 15520 34389 15560
rect 34347 15511 34389 15520
rect 34155 15392 34197 15401
rect 34155 15352 34156 15392
rect 34196 15352 34197 15392
rect 34155 15343 34197 15352
rect 33484 15268 33812 15308
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 33196 14932 33524 14972
rect 32907 14923 32949 14932
rect 32908 14838 32948 14923
rect 33099 14888 33141 14897
rect 33099 14848 33100 14888
rect 33140 14848 33236 14888
rect 33099 14839 33141 14848
rect 33100 14820 33140 14839
rect 32812 14671 32852 14680
rect 33004 14720 33044 14729
rect 32908 13880 32948 13889
rect 33004 13880 33044 14680
rect 33196 14720 33236 14848
rect 33387 14804 33429 14813
rect 33387 14764 33388 14804
rect 33428 14764 33429 14804
rect 33387 14755 33429 14764
rect 33196 14671 33236 14680
rect 33388 14720 33428 14755
rect 33388 14669 33428 14680
rect 33484 14720 33524 14932
rect 33484 14671 33524 14680
rect 33292 14552 33332 14561
rect 33196 14512 33292 14552
rect 32948 13840 33044 13880
rect 33100 14006 33140 14015
rect 32908 13831 32948 13840
rect 33100 13553 33140 13966
rect 32811 13544 32853 13553
rect 32811 13504 32812 13544
rect 32852 13504 32853 13544
rect 32811 13495 32853 13504
rect 33099 13544 33141 13553
rect 33099 13504 33100 13544
rect 33140 13504 33141 13544
rect 33099 13495 33141 13504
rect 32812 13460 32852 13495
rect 32812 13409 32852 13420
rect 33196 13292 33236 14512
rect 33292 14503 33332 14512
rect 33772 14225 33812 15268
rect 34348 14897 34388 15511
rect 34828 14972 34868 15679
rect 34924 15569 34964 15654
rect 35116 15653 35156 15684
rect 35211 15679 35253 15688
rect 35115 15644 35157 15653
rect 35115 15604 35116 15644
rect 35156 15604 35157 15644
rect 35115 15595 35157 15604
rect 34923 15560 34965 15569
rect 34923 15520 34924 15560
rect 34964 15520 34965 15560
rect 34923 15511 34965 15520
rect 35116 15560 35156 15595
rect 34923 15392 34965 15401
rect 34923 15352 34924 15392
rect 34964 15352 34965 15392
rect 34923 15343 34965 15352
rect 34924 15258 34964 15343
rect 34828 14923 34868 14932
rect 34347 14888 34389 14897
rect 34347 14848 34348 14888
rect 34388 14848 34389 14888
rect 34347 14839 34389 14848
rect 35116 14813 35156 15520
rect 35212 15560 35252 15679
rect 35212 15511 35252 15520
rect 35403 15476 35445 15485
rect 35403 15436 35404 15476
rect 35444 15436 35445 15476
rect 35403 15427 35445 15436
rect 35211 14888 35253 14897
rect 35211 14848 35212 14888
rect 35252 14848 35253 14888
rect 35211 14839 35253 14848
rect 35115 14804 35157 14813
rect 35115 14764 35116 14804
rect 35156 14764 35157 14804
rect 35115 14755 35157 14764
rect 34347 14720 34389 14729
rect 34347 14680 34348 14720
rect 34388 14680 34389 14720
rect 34347 14671 34389 14680
rect 33771 14216 33813 14225
rect 33771 14176 33772 14216
rect 33812 14176 33813 14216
rect 33771 14167 33813 14176
rect 33484 14048 33524 14057
rect 34348 14048 34388 14671
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 33524 14008 33812 14048
rect 33484 13999 33524 14008
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 33772 13460 33812 14008
rect 34348 13999 34388 14008
rect 33580 13420 33812 13460
rect 33580 13376 33620 13420
rect 33580 13327 33620 13336
rect 33118 13252 33236 13292
rect 34923 13292 34965 13301
rect 34923 13252 34924 13292
rect 34964 13252 34965 13292
rect 33118 13219 33158 13252
rect 34923 13243 34965 13252
rect 32811 13208 32853 13217
rect 32811 13168 32812 13208
rect 32852 13168 32853 13208
rect 32811 13159 32853 13168
rect 33004 13208 33044 13217
rect 33118 13170 33158 13179
rect 34924 13208 34964 13243
rect 35020 13217 35060 13302
rect 32812 13074 32852 13159
rect 33004 12980 33044 13168
rect 34924 13157 34964 13168
rect 35019 13208 35061 13217
rect 35116 13208 35156 14755
rect 35019 13168 35020 13208
rect 35060 13168 35156 13208
rect 35212 13208 35252 14839
rect 35307 14720 35349 14729
rect 35307 14680 35308 14720
rect 35348 14680 35349 14720
rect 35307 14671 35349 14680
rect 35019 13159 35061 13168
rect 35212 13133 35252 13168
rect 35211 13124 35253 13133
rect 35211 13084 35212 13124
rect 35252 13084 35253 13124
rect 35211 13075 35253 13084
rect 35116 13040 35156 13049
rect 35212 13044 35252 13075
rect 35116 12980 35156 13000
rect 32716 12940 33044 12980
rect 35020 12940 35156 12980
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 29931 12496 29932 12536
rect 29972 12496 30260 12536
rect 31371 12536 31413 12545
rect 31371 12496 31372 12536
rect 31412 12496 31413 12536
rect 29931 12487 29973 12496
rect 31371 12487 31413 12496
rect 33868 12536 33908 12545
rect 29932 12402 29972 12487
rect 31372 12402 31412 12487
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 33868 11957 33908 12496
rect 34252 12536 34292 12545
rect 33867 11948 33909 11957
rect 33867 11908 33868 11948
rect 33908 11908 33909 11948
rect 33867 11899 33909 11908
rect 34252 11864 34292 12496
rect 35020 12368 35060 12940
rect 35116 12536 35156 12545
rect 35308 12536 35348 14671
rect 35156 12496 35348 12536
rect 35116 12487 35156 12496
rect 35020 12328 35156 12368
rect 34827 11948 34869 11957
rect 34827 11908 34828 11948
rect 34868 11908 34869 11948
rect 34827 11899 34869 11908
rect 34348 11864 34388 11873
rect 34252 11824 34348 11864
rect 34348 11815 34388 11824
rect 34828 11814 34868 11899
rect 35019 11864 35061 11873
rect 35019 11824 35020 11864
rect 35060 11824 35061 11864
rect 35019 11815 35061 11824
rect 34827 11696 34869 11705
rect 34827 11656 34828 11696
rect 34868 11656 34869 11696
rect 34827 11647 34869 11656
rect 35020 11696 35060 11815
rect 35020 11647 35060 11656
rect 35116 11696 35156 12328
rect 35116 11647 35156 11656
rect 35307 11696 35349 11705
rect 35307 11656 35308 11696
rect 35348 11656 35349 11696
rect 35307 11647 35349 11656
rect 35404 11696 35444 15427
rect 35500 13796 35540 13805
rect 35500 13301 35540 13756
rect 35499 13292 35541 13301
rect 35499 13252 35500 13292
rect 35540 13252 35541 13292
rect 35499 13243 35541 13252
rect 35596 12980 35636 15763
rect 36267 15728 36309 15737
rect 36267 15688 36268 15728
rect 36308 15688 36309 15728
rect 36267 15679 36309 15688
rect 35979 15560 36021 15569
rect 35979 15520 35980 15560
rect 36020 15520 36021 15560
rect 35979 15511 36021 15520
rect 36268 15560 36308 15679
rect 36268 15511 36308 15520
rect 36364 15560 36404 15763
rect 36364 15511 36404 15520
rect 36460 15560 36500 15571
rect 35692 15392 35732 15401
rect 35692 15149 35732 15352
rect 35691 15140 35733 15149
rect 35691 15100 35692 15140
rect 35732 15100 35733 15140
rect 35691 15091 35733 15100
rect 35980 14729 36020 15511
rect 36460 15485 36500 15520
rect 36556 15560 36596 15569
rect 36748 15560 36788 15569
rect 36596 15520 36748 15560
rect 36556 15511 36596 15520
rect 36748 15511 36788 15520
rect 36459 15476 36501 15485
rect 36459 15436 36460 15476
rect 36500 15436 36501 15476
rect 36459 15427 36501 15436
rect 36844 15401 36884 15772
rect 37228 15737 37268 16108
rect 37708 16098 37748 16183
rect 37227 15728 37269 15737
rect 37227 15688 37228 15728
rect 37268 15688 37269 15728
rect 37227 15679 37269 15688
rect 37804 15653 37844 16192
rect 37996 16232 38036 16241
rect 38092 16232 38132 17107
rect 38036 16192 38132 16232
rect 36939 15644 36981 15653
rect 36939 15604 36940 15644
rect 36980 15604 36981 15644
rect 36939 15595 36981 15604
rect 37803 15644 37845 15653
rect 37803 15604 37804 15644
rect 37844 15604 37845 15644
rect 37803 15595 37845 15604
rect 36940 15560 36980 15595
rect 36940 15509 36980 15520
rect 37036 15560 37076 15569
rect 37515 15560 37557 15569
rect 37076 15520 37364 15560
rect 37036 15511 37076 15520
rect 36555 15392 36597 15401
rect 36555 15352 36556 15392
rect 36596 15352 36597 15392
rect 36555 15343 36597 15352
rect 36843 15392 36885 15401
rect 36843 15352 36844 15392
rect 36884 15352 36885 15392
rect 36843 15343 36885 15352
rect 35979 14720 36021 14729
rect 35979 14680 35980 14720
rect 36020 14680 36021 14720
rect 35979 14671 36021 14680
rect 35980 14586 36020 14671
rect 36556 13208 36596 15343
rect 36748 15308 36788 15317
rect 36748 14729 36788 15268
rect 36843 15140 36885 15149
rect 36843 15100 36844 15140
rect 36884 15100 36885 15140
rect 36843 15091 36885 15100
rect 36747 14720 36789 14729
rect 36747 14680 36748 14720
rect 36788 14680 36789 14720
rect 36747 14671 36789 14680
rect 36844 14720 36884 15091
rect 36844 14671 36884 14680
rect 37227 14720 37269 14729
rect 37227 14680 37228 14720
rect 37268 14680 37269 14720
rect 37227 14671 37269 14680
rect 37228 14586 37268 14671
rect 37324 14477 37364 15520
rect 37515 15520 37516 15560
rect 37556 15520 37557 15560
rect 37515 15511 37557 15520
rect 37516 15426 37556 15511
rect 37420 14552 37460 14561
rect 37323 14468 37365 14477
rect 37323 14428 37324 14468
rect 37364 14428 37365 14468
rect 37323 14419 37365 14428
rect 37420 14393 37460 14512
rect 37419 14384 37461 14393
rect 37419 14344 37420 14384
rect 37460 14344 37461 14384
rect 37419 14335 37461 14344
rect 37131 14132 37173 14141
rect 37131 14092 37132 14132
rect 37172 14092 37173 14132
rect 37131 14083 37173 14092
rect 36747 13376 36789 13385
rect 36747 13336 36748 13376
rect 36788 13336 36789 13376
rect 36747 13327 36789 13336
rect 35979 13124 36021 13133
rect 35979 13084 35980 13124
rect 36020 13084 36021 13124
rect 35979 13075 36021 13084
rect 34828 11562 34868 11647
rect 35308 11562 35348 11647
rect 35404 11537 35444 11656
rect 35500 12940 35636 12980
rect 35500 11696 35540 12940
rect 35595 12368 35637 12377
rect 35595 12328 35596 12368
rect 35636 12328 35637 12368
rect 35595 12319 35637 12328
rect 35500 11621 35540 11656
rect 35596 11696 35636 12319
rect 35596 11647 35636 11656
rect 35499 11612 35541 11621
rect 35499 11572 35500 11612
rect 35540 11572 35541 11612
rect 35499 11563 35541 11572
rect 35403 11528 35445 11537
rect 35403 11488 35404 11528
rect 35444 11488 35445 11528
rect 35403 11479 35445 11488
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 35980 11033 36020 13075
rect 36556 12713 36596 13168
rect 36748 13208 36788 13327
rect 36652 13124 36692 13133
rect 36555 12704 36597 12713
rect 36555 12664 36556 12704
rect 36596 12664 36597 12704
rect 36555 12655 36597 12664
rect 36267 12368 36309 12377
rect 36652 12368 36692 13084
rect 36748 12980 36788 13168
rect 36940 13124 36980 13133
rect 36748 12940 36884 12980
rect 36748 12536 36788 12545
rect 36748 12377 36788 12496
rect 36844 12536 36884 12940
rect 36844 12487 36884 12496
rect 36267 12328 36268 12368
rect 36308 12328 36309 12368
rect 36267 12319 36309 12328
rect 36556 12328 36692 12368
rect 36747 12368 36789 12377
rect 36747 12328 36748 12368
rect 36788 12328 36789 12368
rect 36268 12234 36308 12319
rect 36460 12284 36500 12293
rect 36171 11948 36213 11957
rect 36171 11908 36172 11948
rect 36212 11908 36213 11948
rect 36171 11899 36213 11908
rect 36172 11696 36212 11899
rect 36267 11864 36309 11873
rect 36267 11824 36268 11864
rect 36308 11824 36309 11864
rect 36267 11815 36309 11824
rect 36268 11730 36308 11815
rect 36172 11647 36212 11656
rect 36364 11696 36404 11705
rect 36460 11696 36500 12244
rect 36404 11656 36500 11696
rect 36556 11696 36596 12328
rect 36747 12319 36789 12328
rect 36651 11864 36693 11873
rect 36651 11824 36652 11864
rect 36692 11824 36693 11864
rect 36651 11815 36693 11824
rect 36364 11647 36404 11656
rect 36556 11647 36596 11656
rect 36652 11696 36692 11815
rect 36652 11647 36692 11656
rect 36748 11528 36788 12319
rect 36844 11948 36884 11957
rect 36940 11948 36980 13084
rect 37132 12536 37172 14083
rect 37323 14048 37365 14057
rect 37323 14008 37324 14048
rect 37364 14008 37365 14048
rect 37323 13999 37365 14008
rect 37324 13914 37364 13999
rect 37324 13208 37364 13217
rect 37324 12980 37364 13168
rect 37324 12940 37460 12980
rect 37132 12487 37172 12496
rect 37420 12368 37460 12940
rect 37420 12319 37460 12328
rect 36884 11908 36980 11948
rect 36844 11899 36884 11908
rect 37036 11864 37076 11873
rect 37076 11824 37172 11864
rect 37036 11815 37076 11824
rect 36843 11696 36885 11705
rect 36843 11656 36844 11696
rect 36884 11656 36885 11696
rect 36843 11647 36885 11656
rect 36844 11562 36884 11647
rect 36460 11488 36788 11528
rect 35979 11024 36021 11033
rect 35979 10984 35980 11024
rect 36020 10984 36021 11024
rect 35979 10975 36021 10984
rect 36460 11024 36500 11488
rect 36555 11108 36597 11117
rect 36555 11068 36556 11108
rect 36596 11068 36597 11108
rect 36555 11059 36597 11068
rect 36460 10975 36500 10984
rect 36556 11024 36596 11059
rect 36748 11033 36788 11118
rect 37036 11033 37076 11118
rect 36556 10973 36596 10984
rect 36747 11024 36789 11033
rect 36747 10984 36748 11024
rect 36788 10984 36789 11024
rect 36747 10975 36789 10984
rect 36940 11024 36980 11033
rect 36748 10856 36788 10865
rect 36940 10856 36980 10984
rect 37035 11024 37077 11033
rect 37035 10984 37036 11024
rect 37076 10984 37077 11024
rect 37035 10975 37077 10984
rect 37132 10856 37172 11824
rect 37996 11705 38036 16192
rect 38092 15392 38132 15401
rect 38092 14729 38132 15352
rect 38091 14720 38133 14729
rect 38091 14680 38092 14720
rect 38132 14680 38133 14720
rect 38091 14671 38133 14680
rect 38188 14552 38228 20056
rect 38284 20047 38324 20056
rect 38283 19928 38325 19937
rect 38283 19888 38284 19928
rect 38324 19888 38325 19928
rect 38283 19879 38325 19888
rect 38284 18005 38324 19879
rect 38380 19844 38420 20728
rect 38475 20728 38476 20768
rect 38516 20728 38517 20768
rect 38475 20719 38517 20728
rect 38668 20768 38708 20896
rect 38956 20777 38996 21568
rect 39052 21608 39092 21617
rect 39052 20945 39092 21568
rect 39147 21608 39189 21617
rect 39147 21568 39148 21608
rect 39188 21568 39189 21608
rect 39147 21559 39189 21568
rect 39244 21608 39284 21617
rect 39284 21568 39380 21608
rect 39244 21559 39284 21568
rect 39148 21474 39188 21559
rect 39051 20936 39093 20945
rect 39051 20896 39052 20936
rect 39092 20896 39093 20936
rect 39051 20887 39093 20896
rect 38668 20719 38708 20728
rect 38955 20768 38997 20777
rect 38955 20728 38956 20768
rect 38996 20728 38997 20768
rect 38955 20719 38997 20728
rect 39052 20768 39092 20777
rect 39147 20768 39189 20777
rect 39092 20728 39148 20768
rect 39188 20728 39189 20768
rect 39052 20719 39092 20728
rect 39147 20719 39189 20728
rect 38476 20634 38516 20719
rect 39340 20189 39380 21568
rect 39436 21440 39476 21449
rect 39436 20777 39476 21400
rect 39435 20768 39477 20777
rect 39435 20728 39436 20768
rect 39476 20728 39477 20768
rect 39435 20719 39477 20728
rect 39435 20600 39477 20609
rect 39435 20560 39436 20600
rect 39476 20560 39477 20600
rect 39435 20551 39477 20560
rect 39339 20180 39381 20189
rect 39339 20140 39340 20180
rect 39380 20140 39381 20180
rect 39339 20131 39381 20140
rect 38476 20096 38516 20105
rect 38476 19853 38516 20056
rect 38668 20096 38708 20105
rect 38668 19937 38708 20056
rect 38860 20096 38900 20105
rect 39147 20096 39189 20105
rect 38900 20056 38996 20096
rect 38860 20047 38900 20056
rect 38667 19928 38709 19937
rect 38667 19888 38668 19928
rect 38708 19888 38709 19928
rect 38667 19879 38709 19888
rect 38380 19676 38420 19804
rect 38475 19844 38517 19853
rect 38475 19804 38476 19844
rect 38516 19804 38517 19844
rect 38475 19795 38517 19804
rect 38764 19844 38804 19853
rect 38804 19804 38900 19844
rect 38764 19795 38804 19804
rect 38380 19636 38708 19676
rect 38380 19424 38420 19433
rect 38380 18677 38420 19384
rect 38572 19256 38612 19265
rect 38668 19256 38708 19636
rect 38764 19256 38804 19265
rect 38668 19216 38764 19256
rect 38379 18668 38421 18677
rect 38379 18628 38380 18668
rect 38420 18628 38421 18668
rect 38379 18619 38421 18628
rect 38572 18509 38612 19216
rect 38764 19207 38804 19216
rect 38860 19256 38900 19804
rect 38956 19265 38996 20056
rect 39147 20056 39148 20096
rect 39188 20056 39189 20096
rect 39147 20047 39189 20056
rect 39148 19962 39188 20047
rect 39051 19844 39093 19853
rect 39051 19804 39052 19844
rect 39092 19804 39093 19844
rect 39051 19795 39093 19804
rect 39052 19508 39092 19795
rect 39052 19459 39092 19468
rect 38860 19207 38900 19216
rect 38955 19256 38997 19265
rect 38955 19216 38956 19256
rect 38996 19216 38997 19256
rect 38955 19207 38997 19216
rect 39340 19256 39380 20131
rect 39436 19433 39476 20551
rect 39532 19685 39572 23020
rect 39724 20768 39764 23080
rect 39916 20768 39956 20777
rect 39724 20728 39916 20768
rect 39916 20719 39956 20728
rect 40012 20180 40052 24415
rect 40108 24389 40148 25012
rect 40491 24968 40533 24977
rect 40491 24928 40492 24968
rect 40532 24928 40533 24968
rect 40491 24919 40533 24928
rect 40492 24632 40532 24919
rect 40587 24884 40629 24893
rect 40587 24844 40588 24884
rect 40628 24844 40629 24884
rect 40587 24835 40629 24844
rect 40588 24800 40628 24835
rect 40588 24749 40628 24760
rect 40492 24583 40532 24592
rect 40684 24632 40724 25684
rect 40779 25675 40821 25684
rect 40876 25220 40916 25229
rect 40876 24977 40916 25180
rect 40875 24968 40917 24977
rect 40875 24928 40876 24968
rect 40916 24928 40917 24968
rect 40875 24919 40917 24928
rect 40684 24557 40724 24592
rect 40780 24632 40820 24641
rect 40203 24548 40245 24557
rect 40203 24508 40204 24548
rect 40244 24508 40245 24548
rect 40203 24499 40245 24508
rect 40683 24548 40725 24557
rect 40683 24508 40684 24548
rect 40724 24508 40725 24548
rect 40780 24548 40820 24592
rect 40972 24632 41012 25936
rect 41260 25304 41300 25313
rect 41163 24884 41205 24893
rect 41163 24844 41164 24884
rect 41204 24844 41205 24884
rect 41163 24835 41205 24844
rect 40875 24548 40917 24557
rect 40780 24508 40876 24548
rect 40916 24508 40917 24548
rect 40683 24499 40725 24508
rect 40875 24499 40917 24508
rect 40107 24380 40149 24389
rect 40107 24340 40108 24380
rect 40148 24340 40149 24380
rect 40107 24331 40149 24340
rect 40204 24044 40244 24499
rect 40684 24468 40724 24499
rect 40204 23995 40244 24004
rect 40300 24380 40340 24389
rect 40972 24380 41012 24592
rect 41068 24557 41108 24642
rect 41164 24641 41204 24835
rect 41163 24632 41205 24641
rect 41163 24592 41164 24632
rect 41204 24592 41205 24632
rect 41163 24583 41205 24592
rect 41067 24548 41109 24557
rect 41067 24508 41068 24548
rect 41108 24508 41109 24548
rect 41067 24499 41109 24508
rect 41164 24498 41204 24583
rect 41260 24464 41300 25264
rect 41356 24632 41396 26104
rect 41452 26095 41492 26104
rect 41452 25976 41492 25985
rect 41644 25976 41684 26692
rect 41739 26732 41781 26741
rect 41739 26692 41740 26732
rect 41780 26692 41781 26732
rect 41739 26683 41781 26692
rect 41492 25936 41684 25976
rect 41452 25927 41492 25936
rect 41356 24592 41492 24632
rect 41356 24464 41396 24473
rect 41260 24424 41356 24464
rect 41356 24415 41396 24424
rect 40972 24340 41204 24380
rect 40108 23792 40148 23801
rect 40108 23465 40148 23752
rect 40300 23792 40340 24340
rect 40684 23960 40724 23971
rect 40684 23885 40724 23920
rect 40875 23960 40917 23969
rect 40875 23920 40876 23960
rect 40916 23920 40917 23960
rect 40875 23911 40917 23920
rect 40491 23876 40533 23885
rect 40491 23836 40492 23876
rect 40532 23836 40533 23876
rect 40491 23827 40533 23836
rect 40683 23876 40725 23885
rect 40683 23836 40684 23876
rect 40724 23836 40725 23876
rect 40683 23827 40725 23836
rect 40300 23743 40340 23752
rect 40107 23456 40149 23465
rect 40107 23416 40108 23456
rect 40148 23416 40149 23456
rect 40107 23407 40149 23416
rect 40203 22112 40245 22121
rect 40203 22072 40204 22112
rect 40244 22072 40245 22112
rect 40203 22063 40245 22072
rect 39724 20140 40052 20180
rect 39531 19676 39573 19685
rect 39531 19636 39532 19676
rect 39572 19636 39573 19676
rect 39531 19627 39573 19636
rect 39435 19424 39477 19433
rect 39435 19384 39436 19424
rect 39476 19384 39477 19424
rect 39435 19375 39477 19384
rect 39340 19207 39380 19216
rect 39435 19256 39477 19265
rect 39724 19256 39764 20140
rect 40204 19340 40244 22063
rect 40492 21029 40532 23827
rect 40779 23792 40821 23801
rect 40779 23752 40780 23792
rect 40820 23752 40821 23792
rect 40779 23743 40821 23752
rect 40876 23792 40916 23911
rect 40876 23743 40916 23752
rect 41068 23792 41108 23801
rect 40780 23330 40820 23743
rect 40972 23708 41012 23717
rect 40876 23330 40916 23382
rect 40780 23290 40917 23330
rect 40875 23288 40917 23290
rect 40875 23248 40876 23288
rect 40916 23248 40917 23288
rect 40875 23239 40917 23248
rect 40972 23060 41012 23668
rect 41068 23330 41108 23752
rect 41068 23281 41108 23290
rect 40780 23020 41012 23060
rect 40780 22289 40820 23020
rect 41164 22616 41204 24340
rect 41452 24044 41492 24592
rect 41643 24380 41685 24389
rect 41643 24340 41644 24380
rect 41684 24340 41685 24380
rect 41643 24331 41685 24340
rect 41452 23969 41492 24004
rect 41451 23960 41493 23969
rect 41451 23920 41452 23960
rect 41492 23920 41493 23960
rect 41451 23911 41493 23920
rect 41259 23876 41301 23885
rect 41452 23880 41492 23911
rect 41259 23836 41260 23876
rect 41300 23836 41301 23876
rect 41259 23827 41301 23836
rect 41260 23742 41300 23827
rect 41452 23624 41492 23633
rect 40876 22576 41204 22616
rect 41260 23584 41452 23624
rect 40684 22280 40724 22289
rect 40684 21701 40724 22240
rect 40779 22280 40821 22289
rect 40779 22240 40780 22280
rect 40820 22240 40821 22280
rect 40779 22231 40821 22240
rect 40780 22146 40820 22231
rect 40683 21692 40725 21701
rect 40683 21652 40684 21692
rect 40724 21652 40725 21692
rect 40683 21643 40725 21652
rect 40876 21608 40916 22576
rect 40972 22448 41012 22457
rect 41012 22408 41204 22448
rect 40972 22399 41012 22408
rect 40972 22280 41012 22289
rect 40972 22112 41012 22240
rect 41164 22280 41204 22408
rect 41164 22231 41204 22240
rect 41260 22112 41300 23584
rect 41452 23575 41492 23584
rect 41355 23288 41397 23297
rect 41355 23248 41356 23288
rect 41396 23248 41397 23288
rect 41355 23239 41397 23248
rect 41356 23204 41396 23239
rect 41644 23213 41684 24331
rect 41740 23717 41780 26683
rect 42124 25976 42164 26776
rect 42124 25927 42164 25936
rect 42123 25304 42165 25313
rect 42123 25264 42124 25304
rect 42164 25264 42165 25304
rect 42123 25255 42165 25264
rect 42124 25170 42164 25255
rect 42220 23885 42260 26944
rect 42315 24632 42357 24641
rect 42315 24592 42316 24632
rect 42356 24592 42357 24632
rect 42315 24583 42357 24592
rect 42316 24498 42356 24583
rect 42219 23876 42261 23885
rect 42219 23836 42220 23876
rect 42260 23836 42261 23876
rect 42219 23827 42261 23836
rect 41739 23708 41781 23717
rect 41739 23668 41740 23708
rect 41780 23668 41781 23708
rect 41739 23659 41781 23668
rect 41356 23153 41396 23164
rect 41643 23204 41685 23213
rect 41643 23164 41644 23204
rect 41684 23164 41685 23204
rect 41643 23155 41685 23164
rect 40972 22072 41300 22112
rect 41452 23120 41492 23129
rect 41355 21944 41397 21953
rect 41452 21944 41492 23080
rect 41547 22952 41589 22961
rect 41547 22912 41548 22952
rect 41588 22912 41589 22952
rect 41547 22903 41589 22912
rect 41548 22280 41588 22903
rect 41548 22231 41588 22240
rect 41355 21904 41356 21944
rect 41396 21904 41492 21944
rect 41355 21895 41397 21904
rect 41259 21692 41301 21701
rect 41259 21652 41260 21692
rect 41300 21652 41301 21692
rect 41259 21643 41301 21652
rect 41164 21608 41204 21617
rect 40876 21568 41164 21608
rect 40491 21020 40533 21029
rect 40491 20980 40492 21020
rect 40532 20980 40533 21020
rect 40491 20971 40533 20980
rect 41068 20600 41108 20609
rect 40972 20560 41068 20600
rect 40972 20189 41012 20560
rect 41068 20551 41108 20560
rect 40971 20180 41013 20189
rect 40971 20140 40972 20180
rect 41012 20140 41013 20180
rect 40971 20131 41013 20140
rect 40779 19928 40821 19937
rect 40779 19888 40780 19928
rect 40820 19888 40821 19928
rect 40779 19879 40821 19888
rect 40780 19794 40820 19879
rect 40395 19676 40437 19685
rect 40395 19636 40396 19676
rect 40436 19636 40437 19676
rect 40395 19627 40437 19636
rect 40396 19550 40436 19627
rect 40779 19592 40821 19601
rect 40779 19552 40780 19592
rect 40820 19552 40821 19592
rect 40396 19510 40628 19550
rect 40779 19543 40821 19552
rect 40588 19508 40628 19510
rect 40588 19459 40628 19468
rect 40396 19424 40436 19435
rect 40396 19349 40436 19384
rect 40780 19351 40820 19543
rect 40204 19291 40244 19300
rect 40395 19340 40437 19349
rect 40395 19300 40396 19340
rect 40436 19300 40437 19340
rect 40780 19302 40820 19311
rect 40395 19291 40437 19300
rect 39435 19216 39436 19256
rect 39476 19216 39477 19256
rect 39435 19207 39477 19216
rect 39628 19216 39724 19256
rect 38668 19088 38708 19097
rect 38708 19048 38804 19088
rect 38668 19039 38708 19048
rect 38764 18668 38804 19048
rect 39436 18761 39476 19207
rect 39435 18752 39477 18761
rect 39435 18712 39436 18752
rect 39476 18712 39477 18752
rect 39435 18703 39477 18712
rect 38764 18619 38804 18628
rect 38667 18584 38709 18593
rect 38667 18544 38668 18584
rect 38708 18544 38709 18584
rect 38667 18535 38709 18544
rect 39148 18584 39188 18593
rect 39188 18544 39476 18584
rect 39148 18535 39188 18544
rect 38571 18500 38613 18509
rect 38571 18460 38572 18500
rect 38612 18460 38613 18500
rect 38571 18451 38613 18460
rect 38572 18332 38612 18343
rect 38572 18257 38612 18292
rect 38571 18248 38613 18257
rect 38571 18208 38572 18248
rect 38612 18208 38613 18248
rect 38571 18199 38613 18208
rect 38283 17996 38325 18005
rect 38283 17956 38284 17996
rect 38324 17956 38325 17996
rect 38283 17947 38325 17956
rect 38283 17324 38325 17333
rect 38283 17284 38284 17324
rect 38324 17284 38325 17324
rect 38283 17275 38325 17284
rect 38284 15560 38324 17275
rect 38572 17072 38612 17081
rect 38668 17072 38708 18535
rect 39436 17912 39476 18544
rect 39436 17863 39476 17872
rect 38955 17828 38997 17837
rect 38955 17788 38956 17828
rect 38996 17788 38997 17828
rect 38955 17779 38997 17788
rect 38612 17032 38708 17072
rect 38475 16400 38517 16409
rect 38475 16360 38476 16400
rect 38516 16360 38517 16400
rect 38475 16351 38517 16360
rect 38379 15644 38421 15653
rect 38379 15604 38380 15644
rect 38420 15604 38421 15644
rect 38379 15595 38421 15604
rect 38284 15511 38324 15520
rect 38380 15510 38420 15595
rect 38476 15560 38516 16351
rect 38572 15569 38612 17032
rect 38476 15511 38516 15520
rect 38571 15560 38613 15569
rect 38571 15520 38572 15560
rect 38612 15520 38613 15560
rect 38571 15511 38613 15520
rect 38572 14720 38612 15511
rect 38092 14512 38228 14552
rect 38380 14680 38572 14720
rect 38092 11957 38132 14512
rect 38284 14048 38324 14057
rect 38380 14048 38420 14680
rect 38572 14671 38612 14680
rect 38571 14468 38613 14477
rect 38571 14428 38572 14468
rect 38612 14428 38613 14468
rect 38571 14419 38613 14428
rect 38572 14216 38612 14419
rect 38572 14167 38612 14176
rect 38324 14008 38420 14048
rect 38476 14048 38516 14057
rect 38188 13208 38228 13217
rect 38284 13208 38324 14008
rect 38228 13168 38324 13208
rect 38091 11948 38133 11957
rect 38091 11908 38092 11948
rect 38132 11908 38133 11948
rect 38091 11899 38133 11908
rect 37995 11696 38037 11705
rect 37995 11656 37996 11696
rect 38036 11656 38037 11696
rect 37995 11647 38037 11656
rect 38092 11621 38132 11899
rect 37611 11612 37653 11621
rect 37611 11572 37612 11612
rect 37652 11572 37653 11612
rect 37611 11563 37653 11572
rect 38091 11612 38133 11621
rect 38091 11572 38092 11612
rect 38132 11572 38133 11612
rect 38091 11563 38133 11572
rect 37515 11528 37557 11537
rect 37515 11488 37516 11528
rect 37556 11488 37557 11528
rect 37515 11479 37557 11488
rect 37228 11024 37268 11033
rect 37420 11024 37460 11033
rect 37268 10984 37420 11024
rect 37228 10975 37268 10984
rect 37420 10975 37460 10984
rect 37516 11024 37556 11479
rect 37516 10975 37556 10984
rect 37612 11024 37652 11563
rect 37612 10975 37652 10984
rect 37707 11024 37749 11033
rect 37707 10984 37708 11024
rect 37748 10984 37749 11024
rect 37707 10975 37749 10984
rect 37708 10890 37748 10975
rect 36788 10816 36980 10856
rect 37036 10816 37172 10856
rect 36748 10807 36788 10816
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 36459 10184 36501 10193
rect 36459 10144 36460 10184
rect 36500 10144 36501 10184
rect 36459 10135 36501 10144
rect 36844 10184 36884 10193
rect 37036 10184 37076 10816
rect 37228 10772 37268 10781
rect 37228 10193 37268 10732
rect 36884 10144 37076 10184
rect 37227 10184 37269 10193
rect 37227 10144 37228 10184
rect 37268 10144 37269 10184
rect 36844 10135 36884 10144
rect 37227 10135 37269 10144
rect 37708 10184 37748 10193
rect 38188 10184 38228 13168
rect 38476 13133 38516 14008
rect 38571 14048 38613 14057
rect 38571 14008 38572 14048
rect 38612 14008 38613 14048
rect 38571 13999 38613 14008
rect 38668 14048 38708 14057
rect 38475 13124 38517 13133
rect 38475 13084 38476 13124
rect 38516 13084 38517 13124
rect 38475 13075 38517 13084
rect 38572 11024 38612 13999
rect 38668 13217 38708 14008
rect 38763 14048 38805 14057
rect 38763 14008 38764 14048
rect 38804 14008 38805 14048
rect 38763 13999 38805 14008
rect 38764 13914 38804 13999
rect 38667 13208 38709 13217
rect 38667 13168 38668 13208
rect 38708 13168 38709 13208
rect 38667 13159 38709 13168
rect 38859 12032 38901 12041
rect 38859 11992 38860 12032
rect 38900 11992 38901 12032
rect 38859 11983 38901 11992
rect 38860 11948 38900 11983
rect 38860 11897 38900 11908
rect 38859 11696 38901 11705
rect 38859 11656 38860 11696
rect 38900 11656 38901 11696
rect 38859 11647 38901 11656
rect 38860 11562 38900 11647
rect 38859 11360 38901 11369
rect 38859 11320 38860 11360
rect 38900 11320 38901 11360
rect 38859 11311 38901 11320
rect 38572 10975 38612 10984
rect 38860 11024 38900 11311
rect 38956 11276 38996 17779
rect 39243 16484 39285 16493
rect 39243 16444 39244 16484
rect 39284 16444 39285 16484
rect 39243 16435 39285 16444
rect 39052 15560 39092 15569
rect 39052 15308 39092 15520
rect 39147 15560 39189 15569
rect 39147 15520 39148 15560
rect 39188 15520 39189 15560
rect 39147 15511 39189 15520
rect 39244 15560 39284 16435
rect 39244 15511 39284 15520
rect 39148 15426 39188 15511
rect 39436 15308 39476 15317
rect 39052 15268 39436 15308
rect 39436 15259 39476 15268
rect 39435 14720 39477 14729
rect 39435 14680 39436 14720
rect 39476 14680 39477 14720
rect 39435 14671 39477 14680
rect 39339 14636 39381 14645
rect 39339 14596 39340 14636
rect 39380 14596 39381 14636
rect 39339 14587 39381 14596
rect 39340 14468 39380 14587
rect 39436 14586 39476 14671
rect 39340 14428 39476 14468
rect 39147 14384 39189 14393
rect 39147 14344 39148 14384
rect 39188 14344 39189 14384
rect 39147 14335 39189 14344
rect 39148 14057 39188 14335
rect 39339 14300 39381 14309
rect 39339 14260 39340 14300
rect 39380 14260 39381 14300
rect 39339 14251 39381 14260
rect 39147 14048 39189 14057
rect 39147 14008 39148 14048
rect 39188 14008 39189 14048
rect 39147 13999 39189 14008
rect 39244 14048 39284 14059
rect 39148 13914 39188 13999
rect 39244 13973 39284 14008
rect 39340 14048 39380 14251
rect 39436 14216 39476 14428
rect 39436 14167 39476 14176
rect 39628 14141 39668 19216
rect 39724 19207 39764 19216
rect 40972 19256 41012 20131
rect 40972 19207 41012 19216
rect 41068 19256 41108 19265
rect 41164 19256 41204 21568
rect 41260 21558 41300 21643
rect 41356 21608 41396 21895
rect 41356 21559 41396 21568
rect 41644 21188 41684 23155
rect 41740 23120 41780 23659
rect 41740 23071 41780 23080
rect 42604 23060 42644 28195
rect 42796 26648 42836 30295
rect 43084 29765 43124 30808
rect 43179 30701 43219 30883
rect 43276 30764 43316 30892
rect 43948 30848 43988 31312
rect 44044 31303 44084 31312
rect 43852 30808 43988 30848
rect 43276 30715 43316 30724
rect 43371 30764 43413 30773
rect 43371 30724 43372 30764
rect 43412 30724 43413 30764
rect 43371 30715 43413 30724
rect 43179 30652 43219 30661
rect 43372 30680 43412 30715
rect 43756 30689 43796 30774
rect 43372 30629 43412 30640
rect 43755 30680 43797 30689
rect 43755 30640 43756 30680
rect 43796 30640 43797 30680
rect 43755 30631 43797 30640
rect 43755 30512 43797 30521
rect 43755 30472 43756 30512
rect 43796 30472 43797 30512
rect 43755 30463 43797 30472
rect 43756 30378 43796 30463
rect 43852 30017 43892 30808
rect 43947 30680 43989 30689
rect 43947 30640 43948 30680
rect 43988 30640 43989 30680
rect 43947 30631 43989 30640
rect 44044 30680 44084 30689
rect 44620 30680 44660 30689
rect 44084 30640 44620 30680
rect 44044 30631 44084 30640
rect 43948 30546 43988 30631
rect 44236 30512 44276 30521
rect 43851 30008 43893 30017
rect 43851 29968 43852 30008
rect 43892 29968 43893 30008
rect 43851 29959 43893 29968
rect 43852 29840 43892 29849
rect 44236 29840 44276 30472
rect 44620 30101 44660 30640
rect 44716 30680 44756 32479
rect 45003 32192 45045 32201
rect 45003 32152 45004 32192
rect 45044 32152 45045 32192
rect 45003 32143 45045 32152
rect 44811 31688 44853 31697
rect 44811 31648 44812 31688
rect 44852 31648 44853 31688
rect 44811 31639 44853 31648
rect 44812 31025 44852 31639
rect 45004 31361 45044 32143
rect 45772 31940 45812 31949
rect 45003 31352 45045 31361
rect 45003 31312 45004 31352
rect 45044 31312 45045 31352
rect 45003 31303 45045 31312
rect 44811 31016 44853 31025
rect 44811 30976 44812 31016
rect 44852 30976 44853 31016
rect 44811 30967 44853 30976
rect 44716 30631 44756 30640
rect 44812 30680 44852 30967
rect 44812 30631 44852 30640
rect 44908 30680 44948 30689
rect 44715 30260 44757 30269
rect 44715 30220 44716 30260
rect 44756 30220 44757 30260
rect 44715 30211 44757 30220
rect 44619 30092 44661 30101
rect 44619 30052 44620 30092
rect 44660 30052 44661 30092
rect 44619 30043 44661 30052
rect 43892 29800 44276 29840
rect 44716 29840 44756 30211
rect 43852 29791 43892 29800
rect 44716 29791 44756 29800
rect 43083 29756 43125 29765
rect 43083 29716 43084 29756
rect 43124 29716 43125 29756
rect 43083 29707 43125 29716
rect 43468 29756 43508 29765
rect 43468 29345 43508 29716
rect 43467 29336 43509 29345
rect 43467 29296 43468 29336
rect 43508 29296 43509 29336
rect 43467 29287 43509 29296
rect 44908 29168 44948 30640
rect 45004 30269 45044 31303
rect 45772 30941 45812 31900
rect 45771 30932 45813 30941
rect 45771 30892 45772 30932
rect 45812 30892 45813 30932
rect 45771 30883 45813 30892
rect 45868 30680 45908 32824
rect 46060 32864 46100 32899
rect 46060 32813 46100 32824
rect 46156 32864 46196 32873
rect 45964 32696 46004 32705
rect 45964 32276 46004 32656
rect 46060 32276 46100 32285
rect 45964 32236 46060 32276
rect 46060 32227 46100 32236
rect 46156 31613 46196 32824
rect 46348 31781 46388 33100
rect 46444 32864 46484 32873
rect 46732 32864 46772 32873
rect 46484 32824 46580 32864
rect 46444 32815 46484 32824
rect 46443 32612 46485 32621
rect 46443 32572 46444 32612
rect 46484 32572 46485 32612
rect 46443 32563 46485 32572
rect 46444 32192 46484 32563
rect 46444 32143 46484 32152
rect 46347 31772 46389 31781
rect 46347 31732 46348 31772
rect 46388 31732 46389 31772
rect 46347 31723 46389 31732
rect 46155 31604 46197 31613
rect 46155 31564 46156 31604
rect 46196 31564 46197 31604
rect 46155 31555 46197 31564
rect 46060 30680 46100 30689
rect 45868 30640 46060 30680
rect 45964 30269 46004 30640
rect 46060 30631 46100 30640
rect 46252 30680 46292 30689
rect 46252 30512 46292 30640
rect 46156 30472 46292 30512
rect 46348 30680 46388 30689
rect 46060 30428 46100 30437
rect 45003 30260 45045 30269
rect 45003 30220 45004 30260
rect 45044 30220 45045 30260
rect 45003 30211 45045 30220
rect 45963 30260 46005 30269
rect 45963 30220 45964 30260
rect 46004 30220 46005 30260
rect 45963 30211 46005 30220
rect 46060 30185 46100 30388
rect 46059 30176 46101 30185
rect 46059 30136 46060 30176
rect 46100 30136 46101 30176
rect 46059 30127 46101 30136
rect 45867 30092 45909 30101
rect 45867 30052 45868 30092
rect 45908 30052 45909 30092
rect 45867 30043 45909 30052
rect 45868 29958 45908 30043
rect 46060 30008 46100 30017
rect 45964 29968 46060 30008
rect 45003 29336 45045 29345
rect 45003 29296 45004 29336
rect 45044 29296 45045 29336
rect 45003 29287 45045 29296
rect 45004 29202 45044 29287
rect 44908 29119 44948 29128
rect 45099 29168 45141 29177
rect 45099 29128 45100 29168
rect 45140 29128 45141 29168
rect 45099 29119 45141 29128
rect 45196 29168 45236 29177
rect 45100 29034 45140 29119
rect 45196 28580 45236 29128
rect 45964 29168 46004 29968
rect 46060 29959 46100 29968
rect 46156 29588 46196 30472
rect 46348 30353 46388 30640
rect 46347 30344 46389 30353
rect 46347 30304 46348 30344
rect 46388 30304 46389 30344
rect 46347 30295 46389 30304
rect 46251 30176 46293 30185
rect 46251 30136 46252 30176
rect 46292 30136 46293 30176
rect 46251 30127 46293 30136
rect 46060 29548 46196 29588
rect 46060 29252 46100 29548
rect 46060 29177 46100 29212
rect 46155 29252 46197 29261
rect 46155 29212 46156 29252
rect 46196 29212 46197 29252
rect 46252 29252 46292 30127
rect 46347 30092 46389 30101
rect 46347 30052 46348 30092
rect 46388 30052 46389 30092
rect 46347 30043 46389 30052
rect 46348 29840 46388 30043
rect 46348 29791 46388 29800
rect 46444 29840 46484 29851
rect 46540 29840 46580 32824
rect 46732 32108 46772 32824
rect 46828 32864 46868 33151
rect 46828 32815 46868 32824
rect 46924 32537 46964 33664
rect 47020 33704 47060 34159
rect 47020 33209 47060 33664
rect 47019 33200 47061 33209
rect 47019 33160 47020 33200
rect 47060 33160 47061 33200
rect 47019 33151 47061 33160
rect 47116 33032 47156 33041
rect 47116 32873 47156 32992
rect 47308 33032 47348 33041
rect 47115 32864 47157 32873
rect 47115 32824 47116 32864
rect 47156 32824 47157 32864
rect 47115 32815 47157 32824
rect 47308 32621 47348 32992
rect 47787 32948 47829 32957
rect 47787 32908 47788 32948
rect 47828 32908 47829 32948
rect 47787 32899 47829 32908
rect 47692 32864 47732 32873
rect 47307 32612 47349 32621
rect 47307 32572 47308 32612
rect 47348 32572 47349 32612
rect 47307 32563 47349 32572
rect 46923 32528 46965 32537
rect 46923 32488 46924 32528
rect 46964 32488 46965 32528
rect 46923 32479 46965 32488
rect 47307 32192 47349 32201
rect 47307 32152 47308 32192
rect 47348 32152 47349 32192
rect 47307 32143 47349 32152
rect 46732 32068 46868 32108
rect 46828 31949 46868 32068
rect 47308 32058 47348 32143
rect 46827 31940 46869 31949
rect 46827 31900 46828 31940
rect 46868 31900 46869 31940
rect 46827 31891 46869 31900
rect 46731 31604 46773 31613
rect 46731 31564 46732 31604
rect 46772 31564 46773 31604
rect 46731 31555 46773 31564
rect 46732 31470 46772 31555
rect 46635 31352 46677 31361
rect 46635 31312 46636 31352
rect 46676 31312 46677 31352
rect 46635 31303 46677 31312
rect 46828 31352 46868 31891
rect 46828 31303 46868 31312
rect 47211 31352 47253 31361
rect 47211 31312 47212 31352
rect 47252 31312 47253 31352
rect 47211 31303 47253 31312
rect 46636 31218 46676 31303
rect 47212 30689 47252 31303
rect 47211 30680 47253 30689
rect 47211 30640 47212 30680
rect 47252 30640 47253 30680
rect 47211 30631 47253 30640
rect 46828 30512 46868 30521
rect 46732 29840 46772 29849
rect 46540 29800 46732 29840
rect 46444 29765 46484 29800
rect 46443 29756 46485 29765
rect 46443 29716 46444 29756
rect 46484 29716 46485 29756
rect 46443 29707 46485 29716
rect 46348 29252 46388 29261
rect 46252 29212 46348 29252
rect 46155 29203 46197 29212
rect 46348 29203 46388 29212
rect 45964 29119 46004 29128
rect 46059 29168 46101 29177
rect 46059 29128 46060 29168
rect 46100 29128 46101 29168
rect 46059 29119 46101 29128
rect 46156 29168 46196 29203
rect 46060 29088 46100 29119
rect 46156 29117 46196 29128
rect 45292 28580 45332 28589
rect 45196 28540 45292 28580
rect 45292 28531 45332 28540
rect 44332 28496 44372 28505
rect 42988 28328 43028 28337
rect 42892 26816 42932 26825
rect 42988 26816 43028 28288
rect 44140 28160 44180 28169
rect 44140 27833 44180 28120
rect 44139 27824 44181 27833
rect 44139 27784 44140 27824
rect 44180 27784 44181 27824
rect 44139 27775 44181 27784
rect 43563 27740 43605 27749
rect 43563 27700 43564 27740
rect 43604 27700 43605 27740
rect 43563 27691 43605 27700
rect 43275 27656 43317 27665
rect 43275 27616 43276 27656
rect 43316 27616 43317 27656
rect 43275 27607 43317 27616
rect 43083 27404 43125 27413
rect 43083 27364 43084 27404
rect 43124 27364 43125 27404
rect 43083 27355 43125 27364
rect 42932 26776 43028 26816
rect 42892 26767 42932 26776
rect 42796 26608 42932 26648
rect 42700 24632 42740 24641
rect 42740 24592 42836 24632
rect 42700 24583 42740 24592
rect 42796 23960 42836 24592
rect 42796 23911 42836 23920
rect 42892 23060 42932 26608
rect 42988 25313 43028 26776
rect 43084 26228 43124 27355
rect 43276 26825 43316 27607
rect 43564 27606 43604 27691
rect 43948 27656 43988 27665
rect 44332 27656 44372 28456
rect 45004 28328 45044 28337
rect 45004 27833 45044 28288
rect 45100 28328 45140 28337
rect 45003 27824 45045 27833
rect 45003 27784 45004 27824
rect 45044 27784 45045 27824
rect 45003 27775 45045 27784
rect 43988 27616 44372 27656
rect 44812 27656 44852 27665
rect 43948 27607 43988 27616
rect 43371 27152 43413 27161
rect 43371 27112 43372 27152
rect 43412 27112 43413 27152
rect 43371 27103 43413 27112
rect 43275 26816 43317 26825
rect 43275 26776 43276 26816
rect 43316 26776 43317 26816
rect 43275 26767 43317 26776
rect 43179 26228 43221 26237
rect 43084 26188 43180 26228
rect 43220 26188 43221 26228
rect 42987 25304 43029 25313
rect 42987 25264 42988 25304
rect 43028 25264 43029 25304
rect 42987 25255 43029 25264
rect 43084 23060 43124 26188
rect 43179 26179 43221 26188
rect 43180 26160 43220 26179
rect 43276 25136 43316 25145
rect 43276 24809 43316 25096
rect 43275 24800 43317 24809
rect 43275 24760 43276 24800
rect 43316 24760 43317 24800
rect 43275 24751 43317 24760
rect 43372 23549 43412 27103
rect 44715 26900 44757 26909
rect 44715 26860 44716 26900
rect 44756 26860 44757 26900
rect 44715 26851 44757 26860
rect 44044 26648 44084 26657
rect 44044 26405 44084 26608
rect 44043 26396 44085 26405
rect 44043 26356 44044 26396
rect 44084 26356 44085 26396
rect 44043 26347 44085 26356
rect 43659 26144 43701 26153
rect 43659 26104 43660 26144
rect 43700 26104 43701 26144
rect 43659 26095 43701 26104
rect 44044 26144 44084 26153
rect 43660 26010 43700 26095
rect 43659 25892 43701 25901
rect 43659 25852 43660 25892
rect 43700 25852 43701 25892
rect 43659 25843 43701 25852
rect 43660 25313 43700 25843
rect 44044 25472 44084 26104
rect 44140 25472 44180 25481
rect 44044 25432 44140 25472
rect 44140 25423 44180 25432
rect 43659 25304 43701 25313
rect 43659 25264 43660 25304
rect 43700 25264 43701 25304
rect 43659 25255 43701 25264
rect 43564 24632 43604 24660
rect 43660 24632 43700 25255
rect 44043 25220 44085 25229
rect 44043 25180 44044 25220
rect 44084 25180 44085 25220
rect 44043 25171 44085 25180
rect 43604 24592 43700 24632
rect 43564 24583 43604 24592
rect 43371 23540 43413 23549
rect 43371 23500 43372 23540
rect 43412 23500 43413 23540
rect 43371 23491 43413 23500
rect 42604 23020 42740 23060
rect 42892 23020 43028 23060
rect 43084 23020 43220 23060
rect 42027 22952 42069 22961
rect 42027 22912 42028 22952
rect 42068 22912 42069 22952
rect 42027 22903 42069 22912
rect 42028 22818 42068 22903
rect 42411 22280 42453 22289
rect 42411 22240 42412 22280
rect 42452 22240 42453 22280
rect 42411 22231 42453 22240
rect 42412 22146 42452 22231
rect 42411 21692 42453 21701
rect 42411 21652 42412 21692
rect 42452 21652 42453 21692
rect 42411 21643 42453 21652
rect 42412 21558 42452 21643
rect 42507 21608 42549 21617
rect 42507 21568 42508 21608
rect 42548 21568 42549 21608
rect 42507 21559 42549 21568
rect 41356 21148 41684 21188
rect 41260 19433 41300 19518
rect 41259 19424 41301 19433
rect 41259 19384 41260 19424
rect 41300 19384 41301 19424
rect 41259 19375 41301 19384
rect 41108 19216 41204 19256
rect 41260 19256 41300 19265
rect 41356 19256 41396 21148
rect 41547 21020 41589 21029
rect 41547 20980 41548 21020
rect 41588 20980 41589 21020
rect 41547 20971 41589 20980
rect 41300 19216 41396 19256
rect 41452 20096 41492 20105
rect 41068 19207 41108 19216
rect 41260 19207 41300 19216
rect 41452 19181 41492 20056
rect 41548 19340 41588 20971
rect 41932 20936 41972 20945
rect 41836 20096 41876 20105
rect 41932 20096 41972 20896
rect 42411 20936 42453 20945
rect 42411 20896 42412 20936
rect 42452 20896 42453 20936
rect 42411 20887 42453 20896
rect 42412 20768 42452 20887
rect 42508 20777 42548 21559
rect 42700 20852 42740 23020
rect 42892 22952 42932 22961
rect 42796 21608 42836 21617
rect 42892 21608 42932 22912
rect 42836 21568 42932 21608
rect 42796 21559 42836 21568
rect 42892 20852 42932 20861
rect 42700 20812 42892 20852
rect 42892 20803 42932 20812
rect 42412 20719 42452 20728
rect 42507 20768 42549 20777
rect 42507 20728 42508 20768
rect 42548 20728 42549 20768
rect 42507 20719 42549 20728
rect 42604 20768 42644 20777
rect 42508 20634 42548 20719
rect 42316 20600 42356 20609
rect 41876 20056 41972 20096
rect 42220 20560 42316 20600
rect 41836 20047 41876 20056
rect 41643 19592 41685 19601
rect 41643 19552 41644 19592
rect 41684 19552 41685 19592
rect 41643 19543 41685 19552
rect 41548 19291 41588 19300
rect 41451 19172 41493 19181
rect 41451 19132 41452 19172
rect 41492 19132 41493 19172
rect 41451 19123 41493 19132
rect 40971 19088 41013 19097
rect 40971 19048 40972 19088
rect 41012 19048 41013 19088
rect 40971 19039 41013 19048
rect 40203 18668 40245 18677
rect 40203 18628 40204 18668
rect 40244 18628 40245 18668
rect 40203 18619 40245 18628
rect 40011 18584 40053 18593
rect 40011 18544 40012 18584
rect 40052 18544 40053 18584
rect 40011 18535 40053 18544
rect 40012 18450 40052 18535
rect 39819 17744 39861 17753
rect 39819 17704 39820 17744
rect 39860 17704 39861 17744
rect 39819 17695 39861 17704
rect 40204 17744 40244 18619
rect 40395 18500 40437 18509
rect 40395 18460 40396 18500
rect 40436 18460 40437 18500
rect 40395 18451 40437 18460
rect 40204 17695 40244 17704
rect 39820 17610 39860 17695
rect 39723 16904 39765 16913
rect 39723 16864 39724 16904
rect 39764 16864 39765 16904
rect 39723 16855 39765 16864
rect 39724 16770 39764 16855
rect 40107 16316 40149 16325
rect 40107 16276 40108 16316
rect 40148 16276 40149 16316
rect 40107 16267 40149 16276
rect 39820 16232 39860 16241
rect 39820 16073 39860 16192
rect 40012 16232 40052 16241
rect 39916 16148 39956 16157
rect 39819 16064 39861 16073
rect 39819 16024 39820 16064
rect 39860 16024 39861 16064
rect 39819 16015 39861 16024
rect 39724 15560 39764 15569
rect 39724 14561 39764 15520
rect 39820 15560 39860 16015
rect 39916 15905 39956 16108
rect 39915 15896 39957 15905
rect 39915 15856 39916 15896
rect 39956 15856 39957 15896
rect 39915 15847 39957 15856
rect 39820 15511 39860 15520
rect 40012 15485 40052 16192
rect 40108 15560 40148 16267
rect 40204 16148 40244 16157
rect 40204 15989 40244 16108
rect 40203 15980 40245 15989
rect 40203 15940 40204 15980
rect 40244 15940 40245 15980
rect 40203 15931 40245 15940
rect 40299 15896 40341 15905
rect 40299 15856 40300 15896
rect 40340 15856 40341 15896
rect 40299 15847 40341 15856
rect 40108 15511 40148 15520
rect 40203 15560 40245 15569
rect 40203 15520 40204 15560
rect 40244 15520 40245 15560
rect 40203 15511 40245 15520
rect 40011 15476 40053 15485
rect 40011 15436 40012 15476
rect 40052 15436 40053 15476
rect 40011 15427 40053 15436
rect 40012 15056 40052 15427
rect 40012 15016 40148 15056
rect 40012 14888 40052 14897
rect 39820 14848 40012 14888
rect 39820 14720 39860 14848
rect 40012 14839 40052 14848
rect 39820 14671 39860 14680
rect 40011 14720 40053 14729
rect 40011 14680 40012 14720
rect 40052 14680 40053 14720
rect 40011 14671 40053 14680
rect 40012 14586 40052 14671
rect 39723 14552 39765 14561
rect 39723 14512 39724 14552
rect 39764 14512 39765 14552
rect 39723 14503 39765 14512
rect 40108 14468 40148 15016
rect 40204 14720 40244 15511
rect 40300 15392 40340 15847
rect 40396 15560 40436 18451
rect 40876 16988 40916 16997
rect 40972 16988 41012 19039
rect 41163 18752 41205 18761
rect 41163 18712 41164 18752
rect 41204 18712 41205 18752
rect 41163 18703 41205 18712
rect 41164 18618 41204 18703
rect 41067 18584 41109 18593
rect 41067 18544 41068 18584
rect 41108 18544 41109 18584
rect 41067 18535 41109 18544
rect 41068 17744 41108 18535
rect 41547 18416 41589 18425
rect 41547 18376 41548 18416
rect 41588 18376 41589 18416
rect 41547 18367 41589 18376
rect 41068 17695 41108 17704
rect 41164 18332 41204 18341
rect 41164 17333 41204 18292
rect 41548 18282 41588 18367
rect 41644 18173 41684 19543
rect 41931 19424 41973 19433
rect 41931 19384 41932 19424
rect 41972 19384 41973 19424
rect 41931 19375 41973 19384
rect 41932 19256 41972 19375
rect 41932 19207 41972 19216
rect 42028 19256 42068 19265
rect 41740 19088 41780 19097
rect 41740 18500 41780 19048
rect 42028 18761 42068 19216
rect 42220 19256 42260 20560
rect 42316 20551 42356 20560
rect 42604 20021 42644 20728
rect 42891 20600 42933 20609
rect 42891 20560 42892 20600
rect 42932 20560 42933 20600
rect 42891 20551 42933 20560
rect 42795 20516 42837 20525
rect 42795 20476 42796 20516
rect 42836 20476 42837 20516
rect 42795 20467 42837 20476
rect 42700 20096 42740 20105
rect 42603 20012 42645 20021
rect 42603 19972 42604 20012
rect 42644 19972 42645 20012
rect 42603 19963 42645 19972
rect 42507 19676 42549 19685
rect 42507 19636 42508 19676
rect 42548 19636 42549 19676
rect 42507 19627 42549 19636
rect 42220 19207 42260 19216
rect 42315 19256 42357 19265
rect 42315 19216 42316 19256
rect 42356 19216 42357 19256
rect 42315 19207 42357 19216
rect 42123 19172 42165 19181
rect 42123 19132 42124 19172
rect 42164 19132 42165 19172
rect 42123 19123 42165 19132
rect 42124 19038 42164 19123
rect 42027 18752 42069 18761
rect 42027 18712 42028 18752
rect 42068 18712 42069 18752
rect 42027 18703 42069 18712
rect 41932 18584 41972 18593
rect 41643 18164 41685 18173
rect 41643 18124 41644 18164
rect 41684 18124 41685 18164
rect 41643 18115 41685 18124
rect 41740 18005 41780 18460
rect 41836 18544 41932 18584
rect 41739 17996 41781 18005
rect 41739 17956 41740 17996
rect 41780 17956 41781 17996
rect 41739 17947 41781 17956
rect 41836 17828 41876 18544
rect 41932 18535 41972 18544
rect 42123 18584 42165 18593
rect 42123 18544 42124 18584
rect 42164 18544 42165 18584
rect 42123 18535 42165 18544
rect 42220 18584 42260 18593
rect 42124 18450 42164 18535
rect 42027 18416 42069 18425
rect 42027 18376 42028 18416
rect 42068 18376 42069 18416
rect 42027 18367 42069 18376
rect 41644 17788 41876 17828
rect 41932 18332 41972 18341
rect 41163 17324 41205 17333
rect 41163 17284 41164 17324
rect 41204 17284 41205 17324
rect 41163 17275 41205 17284
rect 41644 17240 41684 17788
rect 41932 17753 41972 18292
rect 41931 17744 41973 17753
rect 41931 17704 41932 17744
rect 41972 17704 41973 17744
rect 41931 17695 41973 17704
rect 41644 17191 41684 17200
rect 41932 17165 41972 17196
rect 41931 17156 41973 17165
rect 41931 17116 41932 17156
rect 41972 17116 41973 17156
rect 41931 17107 41973 17116
rect 41067 17072 41109 17081
rect 41067 17032 41068 17072
rect 41108 17032 41109 17072
rect 41067 17023 41109 17032
rect 41740 17072 41780 17081
rect 40916 16948 41012 16988
rect 40876 16939 40916 16948
rect 41068 16904 41108 17023
rect 41451 16988 41493 16997
rect 41451 16948 41452 16988
rect 41492 16948 41493 16988
rect 41451 16939 41493 16948
rect 40588 16232 40628 16241
rect 40491 15980 40533 15989
rect 40491 15940 40492 15980
rect 40532 15940 40533 15980
rect 40491 15931 40533 15940
rect 40492 15728 40532 15931
rect 40588 15737 40628 16192
rect 41068 15896 41108 16864
rect 41452 16854 41492 16939
rect 41260 16820 41300 16829
rect 41300 16780 41396 16820
rect 41260 16771 41300 16780
rect 41356 16736 41396 16780
rect 41740 16736 41780 17032
rect 41835 17072 41877 17081
rect 41835 17032 41836 17072
rect 41876 17032 41877 17072
rect 41835 17023 41877 17032
rect 41932 17072 41972 17107
rect 41836 16938 41876 17023
rect 41356 16696 41780 16736
rect 41068 15856 41300 15896
rect 40492 15679 40532 15688
rect 40587 15728 40629 15737
rect 40587 15688 40588 15728
rect 40628 15688 40629 15728
rect 40587 15679 40629 15688
rect 40396 15511 40436 15520
rect 40491 15560 40533 15569
rect 40588 15560 40628 15569
rect 40491 15520 40492 15560
rect 40532 15520 40588 15560
rect 40491 15511 40533 15520
rect 40588 15511 40628 15520
rect 40684 15560 40724 15569
rect 40684 15392 40724 15520
rect 40875 15560 40917 15569
rect 40875 15520 40876 15560
rect 40916 15520 40917 15560
rect 40875 15511 40917 15520
rect 40300 15352 40724 15392
rect 40876 15392 40916 15511
rect 40876 15343 40916 15352
rect 40204 14671 40244 14680
rect 40300 14720 40340 14729
rect 39916 14428 40148 14468
rect 39819 14216 39861 14225
rect 39819 14176 39820 14216
rect 39860 14176 39861 14216
rect 39819 14167 39861 14176
rect 39627 14132 39669 14141
rect 39627 14092 39628 14132
rect 39668 14092 39669 14132
rect 39627 14083 39669 14092
rect 39340 13999 39380 14008
rect 39820 14048 39860 14167
rect 39820 13999 39860 14008
rect 39916 14048 39956 14428
rect 40012 14216 40052 14225
rect 40300 14216 40340 14680
rect 41164 14720 41204 14729
rect 41164 14225 41204 14680
rect 41260 14720 41300 15856
rect 40052 14176 40340 14216
rect 41163 14216 41205 14225
rect 41163 14176 41164 14216
rect 41204 14176 41205 14216
rect 40012 14167 40052 14176
rect 41163 14167 41205 14176
rect 39916 13999 39956 14008
rect 40108 14048 40148 14057
rect 39243 13964 39285 13973
rect 39243 13924 39244 13964
rect 39284 13924 39285 13964
rect 39243 13915 39285 13924
rect 40108 13889 40148 14008
rect 40300 14048 40340 14057
rect 40107 13880 40149 13889
rect 40107 13840 40108 13880
rect 40148 13840 40149 13880
rect 40107 13831 40149 13840
rect 39339 13376 39381 13385
rect 39339 13336 39340 13376
rect 39380 13336 39381 13376
rect 39339 13327 39381 13336
rect 39340 13242 39380 13327
rect 40300 13133 40340 14008
rect 40395 14048 40437 14057
rect 40395 14008 40396 14048
rect 40436 14008 40437 14048
rect 40395 13999 40437 14008
rect 40684 14048 40724 14057
rect 40724 14008 40820 14048
rect 40684 13999 40724 14008
rect 40299 13124 40341 13133
rect 40299 13084 40300 13124
rect 40340 13084 40341 13124
rect 40299 13075 40341 13084
rect 39148 12536 39188 12545
rect 39148 12041 39188 12496
rect 39532 12536 39572 12545
rect 40396 12536 40436 13999
rect 40780 13376 40820 14008
rect 41260 13973 41300 14680
rect 41356 14720 41396 16696
rect 41452 16232 41492 16241
rect 41492 16192 41588 16232
rect 41452 16183 41492 16192
rect 41356 14309 41396 14680
rect 41452 14552 41492 14561
rect 41355 14300 41397 14309
rect 41355 14260 41356 14300
rect 41396 14260 41397 14300
rect 41355 14251 41397 14260
rect 41259 13964 41301 13973
rect 41259 13924 41260 13964
rect 41300 13924 41301 13964
rect 41259 13915 41301 13924
rect 40780 13327 40820 13336
rect 39572 12496 39764 12536
rect 39532 12487 39572 12496
rect 39531 12368 39573 12377
rect 39531 12328 39532 12368
rect 39572 12328 39573 12368
rect 39531 12319 39573 12328
rect 39147 12032 39189 12041
rect 39147 11992 39148 12032
rect 39188 11992 39189 12032
rect 39147 11983 39189 11992
rect 39436 11864 39476 11873
rect 39148 11824 39436 11864
rect 39052 11696 39092 11705
rect 39052 11360 39092 11656
rect 39148 11696 39188 11824
rect 39436 11815 39476 11824
rect 39148 11647 39188 11656
rect 39340 11696 39380 11705
rect 39052 11320 39188 11360
rect 38956 11236 39092 11276
rect 38860 10975 38900 10984
rect 38955 11024 38997 11033
rect 38955 10984 38956 11024
rect 38996 10984 38997 11024
rect 38955 10975 38997 10984
rect 38860 10436 38900 10445
rect 38956 10436 38996 10975
rect 39052 10688 39092 11236
rect 39148 10949 39188 11320
rect 39340 11117 39380 11656
rect 39532 11696 39572 12319
rect 39724 11864 39764 12496
rect 40396 12487 40436 12496
rect 40683 12536 40725 12545
rect 40683 12496 40684 12536
rect 40724 12496 40725 12536
rect 40683 12487 40725 12496
rect 39724 11815 39764 11824
rect 39435 11612 39477 11621
rect 39435 11572 39436 11612
rect 39476 11572 39477 11612
rect 39435 11563 39477 11572
rect 39339 11108 39381 11117
rect 39339 11068 39340 11108
rect 39380 11068 39381 11108
rect 39339 11059 39381 11068
rect 39436 11024 39476 11563
rect 39532 11369 39572 11656
rect 39531 11360 39573 11369
rect 39531 11320 39532 11360
rect 39572 11320 39573 11360
rect 39531 11311 39573 11320
rect 39436 10975 39476 10984
rect 39628 11024 39668 11033
rect 39147 10940 39189 10949
rect 39147 10900 39148 10940
rect 39188 10900 39189 10940
rect 39147 10891 39189 10900
rect 39531 10940 39573 10949
rect 39531 10900 39532 10940
rect 39572 10900 39573 10940
rect 39531 10891 39573 10900
rect 39244 10856 39284 10865
rect 39244 10772 39284 10816
rect 39532 10806 39572 10891
rect 39244 10732 39476 10772
rect 39436 10688 39476 10732
rect 39628 10688 39668 10984
rect 40684 11024 40724 12487
rect 40684 10975 40724 10984
rect 39052 10648 39284 10688
rect 39436 10648 39668 10688
rect 40012 10856 40052 10865
rect 38900 10396 39188 10436
rect 38860 10387 38900 10396
rect 37748 10144 38228 10184
rect 37708 10135 37748 10144
rect 36460 10050 36500 10135
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 39148 9512 39188 10396
rect 39244 9848 39284 10648
rect 39820 10184 39860 10193
rect 40012 10184 40052 10816
rect 39860 10144 40052 10184
rect 40684 10184 40724 10193
rect 39820 10135 39860 10144
rect 39339 10100 39381 10109
rect 39339 10060 39340 10100
rect 39380 10060 39381 10100
rect 39339 10051 39381 10060
rect 39436 10100 39476 10109
rect 39476 10060 39764 10100
rect 39436 10051 39476 10060
rect 39340 9932 39380 10051
rect 39340 9892 39572 9932
rect 39244 9808 39380 9848
rect 39244 9512 39284 9521
rect 39148 9472 39244 9512
rect 39244 9463 39284 9472
rect 39340 9512 39380 9808
rect 39340 9463 39380 9472
rect 39532 9512 39572 9892
rect 39724 9764 39764 10060
rect 39724 9724 40244 9764
rect 40204 9680 40244 9724
rect 40684 9689 40724 10144
rect 40971 10100 41013 10109
rect 40971 10060 40972 10100
rect 41012 10060 41013 10100
rect 40971 10051 41013 10060
rect 40204 9631 40244 9640
rect 40683 9680 40725 9689
rect 40683 9640 40684 9680
rect 40724 9640 40725 9680
rect 40683 9631 40725 9640
rect 40875 9596 40917 9605
rect 40875 9556 40876 9596
rect 40916 9556 40917 9596
rect 40875 9547 40917 9556
rect 39532 9463 39572 9472
rect 40012 9512 40052 9521
rect 39532 9344 39572 9353
rect 40012 9344 40052 9472
rect 40107 9512 40149 9521
rect 40107 9472 40108 9512
rect 40148 9472 40149 9512
rect 40107 9463 40149 9472
rect 40300 9512 40340 9521
rect 40684 9512 40724 9521
rect 40340 9472 40684 9512
rect 40300 9463 40340 9472
rect 40684 9463 40724 9472
rect 40779 9512 40821 9521
rect 40779 9472 40780 9512
rect 40820 9472 40821 9512
rect 40779 9463 40821 9472
rect 40876 9512 40916 9547
rect 40108 9378 40148 9463
rect 40780 9378 40820 9463
rect 40876 9461 40916 9472
rect 40972 9512 41012 10051
rect 41260 9605 41300 13915
rect 41259 9596 41301 9605
rect 41259 9556 41260 9596
rect 41300 9556 41301 9596
rect 41259 9547 41301 9556
rect 41356 9521 41396 14251
rect 41452 13208 41492 14512
rect 41548 14057 41588 16192
rect 41835 15980 41877 15989
rect 41835 15940 41836 15980
rect 41876 15940 41877 15980
rect 41835 15931 41877 15940
rect 41836 15560 41876 15931
rect 41932 15896 41972 17032
rect 42028 15989 42068 18367
rect 42220 18341 42260 18544
rect 42219 18332 42261 18341
rect 42219 18292 42220 18332
rect 42260 18292 42261 18332
rect 42219 18283 42261 18292
rect 42123 18164 42165 18173
rect 42123 18124 42124 18164
rect 42164 18124 42165 18164
rect 42123 18115 42165 18124
rect 42124 16904 42164 18115
rect 42220 17576 42260 17585
rect 42220 17249 42260 17536
rect 42219 17240 42261 17249
rect 42219 17200 42220 17240
rect 42260 17200 42261 17240
rect 42219 17191 42261 17200
rect 42220 17072 42260 17081
rect 42316 17072 42356 19207
rect 42508 18668 42548 19627
rect 42604 19592 42644 19963
rect 42700 19853 42740 20056
rect 42699 19844 42741 19853
rect 42699 19804 42700 19844
rect 42740 19804 42741 19844
rect 42699 19795 42741 19804
rect 42604 19552 42740 19592
rect 42603 18668 42645 18677
rect 42508 18628 42604 18668
rect 42644 18628 42645 18668
rect 42603 18619 42645 18628
rect 42412 18584 42452 18593
rect 42604 18584 42644 18619
rect 42452 18544 42548 18584
rect 42412 18535 42452 18544
rect 42412 18341 42452 18426
rect 42508 18425 42548 18544
rect 42604 18534 42644 18544
rect 42700 18584 42740 19552
rect 42796 19265 42836 20467
rect 42795 19256 42837 19265
rect 42795 19216 42796 19256
rect 42836 19216 42837 19256
rect 42795 19207 42837 19216
rect 42796 19122 42836 19207
rect 42700 18535 42740 18544
rect 42795 18584 42837 18593
rect 42795 18544 42796 18584
rect 42836 18544 42837 18584
rect 42795 18535 42837 18544
rect 42507 18416 42549 18425
rect 42507 18376 42508 18416
rect 42548 18376 42549 18416
rect 42507 18367 42549 18376
rect 42411 18332 42453 18341
rect 42411 18292 42412 18332
rect 42452 18292 42453 18332
rect 42411 18283 42453 18292
rect 42604 17837 42644 17868
rect 42603 17828 42645 17837
rect 42603 17788 42604 17828
rect 42644 17788 42645 17828
rect 42603 17779 42645 17788
rect 42604 17744 42644 17779
rect 42796 17753 42836 18535
rect 42892 18509 42932 20551
rect 42988 20180 43028 23020
rect 43180 22952 43220 23020
rect 43084 22912 43220 22952
rect 43084 20861 43124 22912
rect 43563 22532 43605 22541
rect 43563 22492 43564 22532
rect 43604 22492 43605 22532
rect 43563 22483 43605 22492
rect 43564 22398 43604 22483
rect 43660 22289 43700 24592
rect 44044 23792 44084 25171
rect 44139 25052 44181 25061
rect 44139 25012 44140 25052
rect 44180 25012 44181 25052
rect 44139 25003 44181 25012
rect 43852 23752 44044 23792
rect 43852 23060 43892 23752
rect 44044 23743 44084 23752
rect 44140 23792 44180 25003
rect 44716 24716 44756 26851
rect 44812 26144 44852 27616
rect 44907 27068 44949 27077
rect 44907 27028 44908 27068
rect 44948 27028 44949 27068
rect 44907 27019 44949 27028
rect 44908 26934 44948 27019
rect 45004 26816 45044 27775
rect 45100 27077 45140 28288
rect 45292 28328 45332 28337
rect 45099 27068 45141 27077
rect 45099 27028 45100 27068
rect 45140 27028 45141 27068
rect 45099 27019 45141 27028
rect 45292 26993 45332 28288
rect 45484 28328 45524 28337
rect 45291 26984 45333 26993
rect 45291 26944 45292 26984
rect 45332 26944 45333 26984
rect 45291 26935 45333 26944
rect 45100 26816 45140 26825
rect 45004 26776 45100 26816
rect 45100 26767 45140 26776
rect 45196 26816 45236 26825
rect 44908 26648 44948 26657
rect 45003 26648 45045 26657
rect 44948 26608 45004 26648
rect 45044 26608 45045 26648
rect 44908 26599 44948 26608
rect 45003 26599 45045 26608
rect 44908 26144 44948 26153
rect 44812 26104 44908 26144
rect 44908 25985 44948 26104
rect 44907 25976 44949 25985
rect 44907 25936 44908 25976
rect 44948 25936 44949 25976
rect 44907 25927 44949 25936
rect 44907 25388 44949 25397
rect 44907 25348 44908 25388
rect 44948 25348 44949 25388
rect 44907 25339 44949 25348
rect 44812 25304 44852 25313
rect 44812 24800 44852 25264
rect 44908 25304 44948 25339
rect 44908 25253 44948 25264
rect 45004 25136 45044 26599
rect 45099 26144 45141 26153
rect 45099 26104 45100 26144
rect 45140 26104 45141 26144
rect 45099 26095 45141 26104
rect 45100 25556 45140 26095
rect 45100 25507 45140 25516
rect 45196 25481 45236 26776
rect 45292 26816 45332 26825
rect 45195 25472 45237 25481
rect 45195 25432 45196 25472
rect 45236 25432 45237 25472
rect 45292 25472 45332 26776
rect 45388 26816 45428 26825
rect 45484 26816 45524 28288
rect 45675 28328 45717 28337
rect 45675 28288 45676 28328
rect 45716 28288 45717 28328
rect 45675 28279 45717 28288
rect 45772 28328 45812 28337
rect 45676 28194 45716 28279
rect 45580 28160 45620 28169
rect 45580 27749 45620 28120
rect 45579 27740 45621 27749
rect 45579 27700 45580 27740
rect 45620 27700 45621 27740
rect 45579 27691 45621 27700
rect 45772 27068 45812 28288
rect 46347 28328 46389 28337
rect 46347 28288 46348 28328
rect 46388 28288 46389 28328
rect 46347 28279 46389 28288
rect 45963 27824 46005 27833
rect 45963 27784 45964 27824
rect 46004 27784 46005 27824
rect 45963 27775 46005 27784
rect 45964 27690 46004 27775
rect 46348 27581 46388 28279
rect 46443 27824 46485 27833
rect 46443 27784 46444 27824
rect 46484 27784 46485 27824
rect 46443 27775 46485 27784
rect 46444 27740 46484 27775
rect 46444 27689 46484 27700
rect 46539 27740 46581 27749
rect 46539 27700 46540 27740
rect 46580 27700 46581 27740
rect 46539 27691 46581 27700
rect 46636 27740 46676 29800
rect 46732 29791 46772 29800
rect 46732 29168 46772 29177
rect 46828 29168 46868 30472
rect 47115 30344 47157 30353
rect 47115 30304 47116 30344
rect 47156 30304 47157 30344
rect 47115 30295 47157 30304
rect 46923 30260 46965 30269
rect 46923 30220 46924 30260
rect 46964 30220 46965 30260
rect 46923 30211 46965 30220
rect 46772 29128 46868 29168
rect 46732 29119 46772 29128
rect 46636 27700 46868 27740
rect 46540 27656 46580 27691
rect 46540 27605 46580 27616
rect 46347 27572 46389 27581
rect 46347 27532 46348 27572
rect 46388 27532 46389 27572
rect 46347 27523 46389 27532
rect 46156 27404 46196 27413
rect 45868 27068 45908 27077
rect 45772 27028 45868 27068
rect 45868 27019 45908 27028
rect 45675 26984 45717 26993
rect 46059 26984 46101 26993
rect 45675 26944 45676 26984
rect 45716 26944 45812 26984
rect 45675 26935 45717 26944
rect 45428 26776 45524 26816
rect 45580 26816 45620 26825
rect 45388 26767 45428 26776
rect 45580 25901 45620 26776
rect 45676 26816 45716 26825
rect 45772 26816 45812 26944
rect 46059 26944 46060 26984
rect 46100 26944 46101 26984
rect 46059 26935 46101 26944
rect 45868 26816 45908 26825
rect 45772 26776 45868 26816
rect 45676 26657 45716 26776
rect 45675 26648 45717 26657
rect 45675 26608 45676 26648
rect 45716 26608 45717 26648
rect 45675 26599 45717 26608
rect 45771 25976 45813 25985
rect 45771 25936 45772 25976
rect 45812 25936 45813 25976
rect 45771 25927 45813 25936
rect 45579 25892 45621 25901
rect 45579 25852 45580 25892
rect 45620 25852 45621 25892
rect 45579 25843 45621 25852
rect 45483 25472 45525 25481
rect 45292 25432 45428 25472
rect 45195 25423 45237 25432
rect 45100 25304 45140 25313
rect 45292 25304 45332 25313
rect 45140 25264 45292 25304
rect 45100 25255 45140 25264
rect 45292 25255 45332 25264
rect 45388 25304 45428 25432
rect 45483 25432 45484 25472
rect 45524 25432 45525 25472
rect 45483 25423 45525 25432
rect 45388 25229 45428 25264
rect 45484 25304 45524 25423
rect 45580 25313 45620 25843
rect 45387 25220 45429 25229
rect 45387 25180 45388 25220
rect 45428 25180 45429 25220
rect 45387 25171 45429 25180
rect 45388 25140 45428 25171
rect 45004 25096 45140 25136
rect 45004 24800 45044 24809
rect 44812 24760 45004 24800
rect 45004 24751 45044 24760
rect 44716 24676 44852 24716
rect 44427 24632 44469 24641
rect 44427 24592 44428 24632
rect 44468 24592 44469 24632
rect 44427 24583 44469 24592
rect 44235 24296 44277 24305
rect 44235 24256 44236 24296
rect 44276 24256 44277 24296
rect 44235 24247 44277 24256
rect 43947 23624 43989 23633
rect 43947 23584 43948 23624
rect 43988 23584 43989 23624
rect 43947 23575 43989 23584
rect 43948 23490 43988 23575
rect 43852 23020 43988 23060
rect 43659 22280 43701 22289
rect 43659 22240 43660 22280
rect 43700 22240 43701 22280
rect 43659 22231 43701 22240
rect 43564 22112 43604 22121
rect 43564 21953 43604 22072
rect 43563 21944 43605 21953
rect 43563 21904 43564 21944
rect 43604 21904 43605 21944
rect 43563 21895 43605 21904
rect 43660 21608 43700 22231
rect 43660 21559 43700 21568
rect 43852 21020 43892 21029
rect 43468 20980 43852 21020
rect 43083 20852 43125 20861
rect 43468 20852 43508 20980
rect 43852 20971 43892 20980
rect 43948 20945 43988 23020
rect 44043 21608 44085 21617
rect 44043 21568 44044 21608
rect 44084 21568 44085 21608
rect 44043 21559 44085 21568
rect 43947 20936 43989 20945
rect 43947 20896 43948 20936
rect 43988 20896 43989 20936
rect 43947 20887 43989 20896
rect 43083 20812 43084 20852
rect 43124 20812 43125 20852
rect 43083 20803 43125 20812
rect 43372 20812 43468 20852
rect 43083 20600 43125 20609
rect 43083 20560 43084 20600
rect 43124 20560 43125 20600
rect 43083 20551 43125 20560
rect 43275 20600 43317 20609
rect 43275 20560 43276 20600
rect 43316 20560 43317 20600
rect 43275 20551 43317 20560
rect 43084 20466 43124 20551
rect 43276 20466 43316 20551
rect 43083 20180 43125 20189
rect 42988 20140 43084 20180
rect 43124 20140 43125 20180
rect 43083 20131 43125 20140
rect 43275 20180 43317 20189
rect 43275 20140 43276 20180
rect 43316 20140 43317 20180
rect 43275 20131 43317 20140
rect 43083 20012 43125 20021
rect 43083 19972 43084 20012
rect 43124 19972 43125 20012
rect 43083 19963 43125 19972
rect 42987 19844 43029 19853
rect 42987 19804 42988 19844
rect 43028 19804 43029 19844
rect 42987 19795 43029 19804
rect 42891 18500 42933 18509
rect 42891 18460 42892 18500
rect 42932 18460 42933 18500
rect 42891 18451 42933 18460
rect 42891 18332 42933 18341
rect 42891 18292 42892 18332
rect 42932 18292 42933 18332
rect 42891 18283 42933 18292
rect 42892 18173 42932 18283
rect 42891 18164 42933 18173
rect 42891 18124 42892 18164
rect 42932 18124 42933 18164
rect 42891 18115 42933 18124
rect 42604 17300 42644 17704
rect 42795 17744 42837 17753
rect 42795 17704 42796 17744
rect 42836 17704 42837 17744
rect 42795 17695 42837 17704
rect 42892 17744 42932 17753
rect 42699 17660 42741 17669
rect 42699 17620 42700 17660
rect 42740 17620 42741 17660
rect 42699 17611 42741 17620
rect 42700 17526 42740 17611
rect 42796 17610 42836 17695
rect 42604 17260 42740 17300
rect 42603 17156 42645 17165
rect 42603 17116 42604 17156
rect 42644 17116 42645 17156
rect 42603 17107 42645 17116
rect 42260 17032 42356 17072
rect 42220 17023 42260 17032
rect 42124 16864 42260 16904
rect 42027 15980 42069 15989
rect 42027 15940 42028 15980
rect 42068 15940 42069 15980
rect 42027 15931 42069 15940
rect 41932 15856 41973 15896
rect 41933 15812 41973 15856
rect 41933 15772 42164 15812
rect 42027 15560 42069 15569
rect 41876 15520 41972 15560
rect 41836 15511 41876 15520
rect 41836 15308 41876 15317
rect 41740 15268 41836 15308
rect 41547 14048 41589 14057
rect 41547 14008 41548 14048
rect 41588 14008 41589 14048
rect 41547 13999 41589 14008
rect 41548 13914 41588 13999
rect 41452 13159 41492 13168
rect 41643 13208 41685 13217
rect 41643 13168 41644 13208
rect 41684 13168 41685 13208
rect 41643 13159 41685 13168
rect 41740 13208 41780 15268
rect 41836 15259 41876 15268
rect 41932 13889 41972 15520
rect 42027 15520 42028 15560
rect 42068 15520 42069 15560
rect 42027 15511 42069 15520
rect 42124 15560 42164 15772
rect 42124 15511 42164 15520
rect 42028 15426 42068 15511
rect 42220 15392 42260 16864
rect 42124 15352 42260 15392
rect 41931 13880 41973 13889
rect 41931 13840 41932 13880
rect 41972 13840 41973 13880
rect 41931 13831 41973 13840
rect 41740 13159 41780 13168
rect 41547 13124 41589 13133
rect 41547 13084 41548 13124
rect 41588 13084 41589 13124
rect 41547 13075 41589 13084
rect 41548 12990 41588 13075
rect 41644 13074 41684 13159
rect 41932 13124 41972 13831
rect 41836 13084 41972 13124
rect 41836 12980 41876 13084
rect 41740 12940 41876 12980
rect 41547 12368 41589 12377
rect 41547 12328 41548 12368
rect 41588 12328 41589 12368
rect 41547 12319 41589 12328
rect 41548 12234 41588 12319
rect 41547 11696 41589 11705
rect 41547 11656 41548 11696
rect 41588 11656 41589 11696
rect 41547 11647 41589 11656
rect 41548 11562 41588 11647
rect 41740 10520 41780 12940
rect 42124 12704 42164 15352
rect 42219 14720 42261 14729
rect 42219 14680 42220 14720
rect 42260 14680 42261 14720
rect 42219 14671 42261 14680
rect 41836 12664 42164 12704
rect 41836 11864 41876 12664
rect 41931 12536 41973 12545
rect 41931 12496 41932 12536
rect 41972 12496 41973 12536
rect 41931 12487 41973 12496
rect 42028 12536 42068 12547
rect 42220 12536 42260 14671
rect 42316 12965 42356 17032
rect 42508 17072 42548 17081
rect 42411 16484 42453 16493
rect 42411 16444 42412 16484
rect 42452 16444 42453 16484
rect 42411 16435 42453 16444
rect 42412 13637 42452 16435
rect 42508 16325 42548 17032
rect 42604 17022 42644 17107
rect 42507 16316 42549 16325
rect 42507 16276 42508 16316
rect 42548 16276 42549 16316
rect 42507 16267 42549 16276
rect 42603 16064 42645 16073
rect 42603 16024 42604 16064
rect 42644 16024 42645 16064
rect 42603 16015 42645 16024
rect 42604 15930 42644 16015
rect 42507 15560 42549 15569
rect 42507 15520 42508 15560
rect 42548 15520 42549 15560
rect 42507 15511 42549 15520
rect 42411 13628 42453 13637
rect 42411 13588 42412 13628
rect 42452 13588 42453 13628
rect 42411 13579 42453 13588
rect 42508 13460 42548 15511
rect 42700 14729 42740 17260
rect 42892 17240 42932 17704
rect 42988 17249 43028 19795
rect 43084 19592 43124 19963
rect 43276 19769 43316 20131
rect 43275 19760 43317 19769
rect 43275 19720 43276 19760
rect 43316 19720 43317 19760
rect 43275 19711 43317 19720
rect 43084 19552 43220 19592
rect 43180 19298 43220 19552
rect 43084 19256 43124 19265
rect 43180 19249 43220 19258
rect 43084 18929 43124 19216
rect 43083 18920 43125 18929
rect 43083 18880 43084 18920
rect 43124 18880 43125 18920
rect 43083 18871 43125 18880
rect 43179 18668 43221 18677
rect 43179 18628 43180 18668
rect 43220 18628 43221 18668
rect 43179 18619 43221 18628
rect 43083 18500 43125 18509
rect 43083 18460 43084 18500
rect 43124 18460 43125 18500
rect 43083 18451 43125 18460
rect 43084 18089 43124 18451
rect 43083 18080 43125 18089
rect 43083 18040 43084 18080
rect 43124 18040 43125 18080
rect 43083 18031 43125 18040
rect 43083 17660 43125 17669
rect 43083 17620 43084 17660
rect 43124 17620 43125 17660
rect 43083 17611 43125 17620
rect 43084 17526 43124 17611
rect 42796 17200 42932 17240
rect 42987 17240 43029 17249
rect 42987 17200 42988 17240
rect 43028 17200 43029 17240
rect 42796 16409 42836 17200
rect 42987 17191 43029 17200
rect 42891 17072 42933 17081
rect 43180 17072 43220 18619
rect 42891 17032 42892 17072
rect 42932 17032 42933 17072
rect 42891 17023 42933 17032
rect 42988 17032 43220 17072
rect 42892 16904 42932 17023
rect 42892 16855 42932 16864
rect 42795 16400 42837 16409
rect 42795 16360 42796 16400
rect 42836 16360 42837 16400
rect 42795 16351 42837 16360
rect 42988 16232 43028 17032
rect 43276 16988 43316 19711
rect 43276 16939 43316 16948
rect 43083 16904 43125 16913
rect 43083 16864 43084 16904
rect 43124 16864 43125 16904
rect 43083 16855 43125 16864
rect 43084 16661 43124 16855
rect 43372 16745 43412 20812
rect 43468 20803 43508 20812
rect 43659 20852 43701 20861
rect 43659 20812 43660 20852
rect 43700 20812 43701 20852
rect 43659 20803 43701 20812
rect 44044 20852 44084 21559
rect 44044 20803 44084 20812
rect 43660 20718 43700 20803
rect 44140 20777 44180 23752
rect 44236 23792 44276 24247
rect 44428 24044 44468 24583
rect 44716 24380 44756 24391
rect 44716 24305 44756 24340
rect 44715 24296 44757 24305
rect 44715 24256 44716 24296
rect 44756 24256 44757 24296
rect 44715 24247 44757 24256
rect 44428 23995 44468 24004
rect 44236 23743 44276 23752
rect 44428 23792 44468 23801
rect 44428 23633 44468 23752
rect 44619 23792 44661 23801
rect 44619 23752 44620 23792
rect 44660 23752 44661 23792
rect 44619 23743 44661 23752
rect 44716 23792 44756 23801
rect 44620 23658 44660 23743
rect 44427 23624 44469 23633
rect 44427 23584 44428 23624
rect 44468 23584 44469 23624
rect 44427 23575 44469 23584
rect 44523 23540 44565 23549
rect 44523 23500 44524 23540
rect 44564 23500 44565 23540
rect 44523 23491 44565 23500
rect 44524 20852 44564 23491
rect 44716 23288 44756 23752
rect 44716 23239 44756 23248
rect 44619 23204 44661 23213
rect 44619 23164 44620 23204
rect 44660 23164 44661 23204
rect 44619 23155 44661 23164
rect 44620 23120 44660 23155
rect 44620 23069 44660 23080
rect 44812 23120 44852 24676
rect 44908 24632 44948 24641
rect 44908 24473 44948 24592
rect 45100 24632 45140 25096
rect 45484 25061 45524 25264
rect 45579 25304 45621 25313
rect 45579 25264 45580 25304
rect 45620 25264 45621 25304
rect 45579 25255 45621 25264
rect 45772 25304 45812 25927
rect 45772 25255 45812 25264
rect 45580 25170 45620 25255
rect 45483 25052 45525 25061
rect 45483 25012 45484 25052
rect 45524 25012 45525 25052
rect 45483 25003 45525 25012
rect 44907 24464 44949 24473
rect 44907 24424 44908 24464
rect 44948 24424 44949 24464
rect 44907 24415 44949 24424
rect 44908 23297 44948 24415
rect 45003 23960 45045 23969
rect 45003 23920 45004 23960
rect 45044 23920 45045 23960
rect 45003 23911 45045 23920
rect 45004 23792 45044 23911
rect 45004 23717 45044 23752
rect 45003 23708 45045 23717
rect 45003 23668 45004 23708
rect 45044 23668 45045 23708
rect 45003 23659 45045 23668
rect 45003 23456 45045 23465
rect 45003 23416 45004 23456
rect 45044 23416 45045 23456
rect 45003 23407 45045 23416
rect 44907 23288 44949 23297
rect 44907 23248 44908 23288
rect 44948 23248 44949 23288
rect 44907 23239 44949 23248
rect 44812 23071 44852 23080
rect 44908 23120 44948 23129
rect 44908 22784 44948 23080
rect 44716 22744 44948 22784
rect 44716 21776 44756 22744
rect 45004 22700 45044 23407
rect 45100 23045 45140 24592
rect 45196 24632 45236 24641
rect 45196 24305 45236 24592
rect 45868 24473 45908 26776
rect 46060 26564 46100 26935
rect 46156 26816 46196 27364
rect 46348 27068 46388 27523
rect 46348 27019 46388 27028
rect 46636 26993 46676 27700
rect 46828 27656 46868 27700
rect 46828 27607 46868 27616
rect 46924 27656 46964 30211
rect 47116 30092 47156 30295
rect 47116 30043 47156 30052
rect 47212 29924 47252 30631
rect 47020 29884 47252 29924
rect 47020 29840 47060 29884
rect 47595 29840 47637 29849
rect 47020 29791 47060 29800
rect 47212 29827 47252 29836
rect 47595 29800 47596 29840
rect 47636 29800 47637 29840
rect 47595 29791 47637 29800
rect 47212 29765 47252 29787
rect 47211 29756 47253 29765
rect 47211 29716 47212 29756
rect 47252 29716 47253 29756
rect 47211 29707 47253 29716
rect 47212 28925 47252 29707
rect 47596 29168 47636 29791
rect 47596 29119 47636 29128
rect 47211 28916 47253 28925
rect 47211 28876 47212 28916
rect 47252 28876 47253 28916
rect 47211 28867 47253 28876
rect 47500 28496 47540 28505
rect 47211 27824 47253 27833
rect 47211 27784 47212 27824
rect 47252 27784 47253 27824
rect 47211 27775 47253 27784
rect 47116 27656 47156 27665
rect 46924 27616 47116 27656
rect 46635 26984 46677 26993
rect 46635 26944 46636 26984
rect 46676 26944 46677 26984
rect 46635 26935 46677 26944
rect 46443 26816 46485 26825
rect 46156 26803 46283 26816
rect 46156 26776 46243 26803
rect 46443 26776 46444 26816
rect 46484 26776 46485 26816
rect 46443 26767 46485 26776
rect 46635 26816 46677 26825
rect 46635 26776 46636 26816
rect 46676 26776 46677 26816
rect 46635 26767 46677 26776
rect 46828 26816 46868 26825
rect 46243 26754 46283 26763
rect 46060 26524 46196 26564
rect 46059 25892 46101 25901
rect 46059 25852 46060 25892
rect 46100 25852 46101 25892
rect 46059 25843 46101 25852
rect 46060 25758 46100 25843
rect 46059 25472 46101 25481
rect 46059 25432 46060 25472
rect 46100 25432 46101 25472
rect 46059 25423 46101 25432
rect 45867 24464 45909 24473
rect 45867 24424 45868 24464
rect 45908 24424 45909 24464
rect 45867 24415 45909 24424
rect 45195 24296 45237 24305
rect 45195 24256 45196 24296
rect 45236 24256 45237 24296
rect 45195 24247 45237 24256
rect 45387 24296 45429 24305
rect 45387 24256 45388 24296
rect 45428 24256 45429 24296
rect 45387 24247 45429 24256
rect 45195 23960 45237 23969
rect 45195 23920 45196 23960
rect 45236 23920 45237 23960
rect 45195 23911 45237 23920
rect 45099 23036 45141 23045
rect 45099 22996 45100 23036
rect 45140 22996 45141 23036
rect 45099 22987 45141 22996
rect 44812 22660 45044 22700
rect 44812 22280 44852 22660
rect 45196 22532 45236 23911
rect 45292 23792 45332 23801
rect 45292 23129 45332 23752
rect 45388 23792 45428 24247
rect 45676 23960 45716 23969
rect 45716 23920 45908 23960
rect 45676 23911 45716 23920
rect 45388 23743 45428 23752
rect 45868 23792 45908 23920
rect 45868 23743 45908 23752
rect 45963 23792 46005 23801
rect 45963 23752 45964 23792
rect 46004 23752 46005 23792
rect 45963 23743 46005 23752
rect 46060 23792 46100 25423
rect 46156 25304 46196 26524
rect 46444 25481 46484 26767
rect 46636 26682 46676 26767
rect 46732 26732 46772 26741
rect 46635 25640 46677 25649
rect 46635 25600 46636 25640
rect 46676 25600 46677 25640
rect 46635 25591 46677 25600
rect 46443 25472 46485 25481
rect 46443 25432 46444 25472
rect 46484 25432 46485 25472
rect 46443 25423 46485 25432
rect 46156 23969 46196 25264
rect 46444 25304 46484 25313
rect 46444 25061 46484 25264
rect 46539 25304 46581 25313
rect 46539 25264 46540 25304
rect 46580 25264 46581 25304
rect 46539 25255 46581 25264
rect 46540 25170 46580 25255
rect 46443 25052 46485 25061
rect 46443 25012 46444 25052
rect 46484 25012 46485 25052
rect 46443 25003 46485 25012
rect 46636 24632 46676 25591
rect 46732 25397 46772 26692
rect 46828 25556 46868 26776
rect 46924 25649 46964 27616
rect 47116 27607 47156 27616
rect 47116 27404 47156 27413
rect 47020 26816 47060 26825
rect 47116 26816 47156 27364
rect 47212 26825 47252 27775
rect 47308 27656 47348 27667
rect 47308 27581 47348 27616
rect 47403 27656 47445 27665
rect 47403 27616 47404 27656
rect 47444 27616 47445 27656
rect 47403 27607 47445 27616
rect 47307 27572 47349 27581
rect 47307 27532 47308 27572
rect 47348 27532 47349 27572
rect 47307 27523 47349 27532
rect 47404 27522 47444 27607
rect 47060 26776 47156 26816
rect 47211 26816 47253 26825
rect 47211 26776 47212 26816
rect 47252 26776 47253 26816
rect 47020 26767 47060 26776
rect 47211 26767 47253 26776
rect 47404 26816 47444 26825
rect 47500 26816 47540 28456
rect 47692 27833 47732 32824
rect 47788 32814 47828 32899
rect 47883 32864 47925 32873
rect 47883 32824 47884 32864
rect 47924 32824 47925 32864
rect 47883 32815 47925 32824
rect 47884 32730 47924 32815
rect 47980 32201 48020 34336
rect 48939 34336 48940 34376
rect 48980 34336 48981 34376
rect 48939 34327 48981 34336
rect 49228 34376 49268 34387
rect 49420 34376 49460 34385
rect 49228 34301 49268 34336
rect 49324 34336 49420 34376
rect 49227 34292 49269 34301
rect 49227 34252 49228 34292
rect 49268 34252 49269 34292
rect 49227 34243 49269 34252
rect 49035 34208 49077 34217
rect 49035 34168 49036 34208
rect 49076 34168 49172 34208
rect 49035 34159 49077 34168
rect 49036 34074 49076 34159
rect 49035 33704 49077 33713
rect 49035 33664 49036 33704
rect 49076 33664 49077 33704
rect 49035 33655 49077 33664
rect 48844 33536 48884 33545
rect 48884 33496 48980 33536
rect 48844 33487 48884 33496
rect 48363 33452 48405 33461
rect 48363 33412 48364 33452
rect 48404 33412 48405 33452
rect 48363 33403 48405 33412
rect 48364 32864 48404 33403
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 48940 33140 48980 33496
rect 48844 33100 48980 33140
rect 48747 33032 48789 33041
rect 48747 32992 48748 33032
rect 48788 32992 48789 33032
rect 48747 32983 48789 32992
rect 48651 32948 48693 32957
rect 48651 32908 48652 32948
rect 48692 32908 48693 32948
rect 48651 32899 48693 32908
rect 48460 32864 48500 32873
rect 48364 32824 48460 32864
rect 48460 32815 48500 32824
rect 48652 32360 48692 32899
rect 48652 32311 48692 32320
rect 47979 32192 48021 32201
rect 47979 32152 47980 32192
rect 48020 32152 48021 32192
rect 47979 32143 48021 32152
rect 48363 32192 48405 32201
rect 48363 32152 48364 32192
rect 48404 32152 48405 32192
rect 48363 32143 48405 32152
rect 48748 32192 48788 32983
rect 48844 32864 48884 33100
rect 49036 32957 49076 33655
rect 49035 32948 49077 32957
rect 49035 32908 49036 32948
rect 49076 32908 49077 32948
rect 49035 32899 49077 32908
rect 48844 32815 48884 32824
rect 49132 32696 49172 34168
rect 49227 33704 49269 33713
rect 49227 33664 49228 33704
rect 49268 33664 49269 33704
rect 49227 33655 49269 33664
rect 49228 33570 49268 33655
rect 49227 33452 49269 33461
rect 49227 33412 49228 33452
rect 49268 33412 49269 33452
rect 49227 33403 49269 33412
rect 49228 33318 49268 33403
rect 49324 33140 49364 34336
rect 49420 34327 49460 34336
rect 49515 34376 49557 34385
rect 49515 34336 49516 34376
rect 49556 34336 49557 34376
rect 49515 34327 49557 34336
rect 49516 34242 49556 34327
rect 49036 32656 49172 32696
rect 49228 33100 49364 33140
rect 49420 33704 49460 33713
rect 48843 32612 48885 32621
rect 48843 32572 48844 32612
rect 48884 32572 48885 32612
rect 48843 32563 48885 32572
rect 48364 31352 48404 32143
rect 48460 31949 48500 32034
rect 48748 32033 48788 32152
rect 48844 32192 48884 32563
rect 48844 32143 48884 32152
rect 48940 32192 48980 32203
rect 48940 32117 48980 32152
rect 48939 32108 48981 32117
rect 48939 32068 48940 32108
rect 48980 32068 48981 32108
rect 48939 32059 48981 32068
rect 48747 32024 48789 32033
rect 48747 31984 48748 32024
rect 48788 31984 48789 32024
rect 48747 31975 48789 31984
rect 48459 31940 48501 31949
rect 49036 31940 49076 32656
rect 49228 32369 49268 33100
rect 49323 32612 49365 32621
rect 49323 32572 49324 32612
rect 49364 32572 49365 32612
rect 49323 32563 49365 32572
rect 49227 32360 49269 32369
rect 49227 32320 49228 32360
rect 49268 32320 49269 32360
rect 49227 32311 49269 32320
rect 49131 32192 49173 32201
rect 49131 32152 49132 32192
rect 49172 32152 49173 32192
rect 49131 32143 49173 32152
rect 49132 32058 49172 32143
rect 48459 31900 48460 31940
rect 48500 31900 48501 31940
rect 48459 31891 48501 31900
rect 48935 31900 49076 31940
rect 48935 31856 48975 31900
rect 49227 31856 49269 31865
rect 48935 31816 48980 31856
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 48556 31352 48596 31361
rect 48364 31312 48556 31352
rect 48268 30512 48308 30521
rect 48172 29840 48212 29849
rect 48268 29840 48308 30472
rect 48364 29849 48404 31312
rect 48556 31303 48596 31312
rect 48940 31352 48980 31816
rect 49227 31816 49228 31856
rect 49268 31816 49269 31856
rect 49227 31807 49269 31816
rect 49035 31604 49077 31613
rect 49035 31564 49036 31604
rect 49076 31564 49077 31604
rect 49035 31555 49077 31564
rect 49228 31604 49268 31807
rect 49228 31555 49268 31564
rect 49036 31361 49076 31555
rect 48940 31303 48980 31312
rect 49035 31352 49077 31361
rect 49227 31352 49269 31361
rect 49035 31312 49036 31352
rect 49076 31312 49077 31352
rect 49035 31303 49077 31312
rect 49132 31312 49228 31352
rect 49268 31312 49269 31352
rect 49036 31218 49076 31303
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 48212 29800 48308 29840
rect 48363 29840 48405 29849
rect 48363 29800 48364 29840
rect 48404 29800 48405 29840
rect 48172 29791 48212 29800
rect 48363 29791 48405 29800
rect 49035 29840 49077 29849
rect 49035 29800 49036 29840
rect 49076 29800 49077 29840
rect 49035 29791 49077 29800
rect 47788 29756 47828 29765
rect 47788 29009 47828 29716
rect 49036 29706 49076 29791
rect 49132 29681 49172 31312
rect 49227 31303 49269 31312
rect 49228 31218 49268 31303
rect 49228 30848 49268 30857
rect 49324 30848 49364 32563
rect 49420 32369 49460 33664
rect 49516 33704 49556 33713
rect 49419 32360 49461 32369
rect 49419 32320 49420 32360
rect 49460 32320 49461 32360
rect 49419 32311 49461 32320
rect 49516 31865 49556 33664
rect 49612 32864 49652 35176
rect 49707 35167 49749 35176
rect 49708 35082 49748 35167
rect 50283 34292 50325 34301
rect 50283 34252 50284 34292
rect 50324 34252 50325 34292
rect 50283 34243 50325 34252
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 49708 32864 49748 32873
rect 49612 32824 49708 32864
rect 49612 32360 49652 32824
rect 49708 32815 49748 32824
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 49612 32311 49652 32320
rect 50091 32192 50133 32201
rect 50091 32152 50092 32192
rect 50132 32152 50133 32192
rect 50091 32143 50133 32152
rect 49995 32108 50037 32117
rect 49995 32068 49996 32108
rect 50036 32068 50037 32108
rect 49995 32059 50037 32068
rect 49611 31940 49653 31949
rect 49611 31900 49612 31940
rect 49652 31900 49653 31940
rect 49611 31891 49653 31900
rect 49515 31856 49557 31865
rect 49515 31816 49516 31856
rect 49556 31816 49557 31856
rect 49515 31807 49557 31816
rect 49515 31184 49557 31193
rect 49515 31144 49516 31184
rect 49556 31144 49557 31184
rect 49515 31135 49557 31144
rect 49268 30808 49364 30848
rect 49228 30799 49268 30808
rect 49324 30689 49364 30808
rect 49323 30680 49365 30689
rect 49323 30640 49324 30680
rect 49364 30640 49365 30680
rect 49323 30631 49365 30640
rect 49420 30596 49460 30605
rect 49420 29840 49460 30556
rect 49324 29800 49460 29840
rect 49131 29672 49173 29681
rect 49131 29632 49132 29672
rect 49172 29632 49173 29672
rect 49131 29623 49173 29632
rect 47787 29000 47829 29009
rect 47787 28960 47788 29000
rect 47828 28960 47829 29000
rect 47787 28951 47829 28960
rect 48748 28925 48788 29010
rect 48747 28916 48789 28925
rect 48747 28876 48748 28916
rect 48788 28876 48789 28916
rect 48747 28867 48789 28876
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 49228 28496 49268 28505
rect 48843 28160 48885 28169
rect 48843 28120 48844 28160
rect 48884 28120 48885 28160
rect 48843 28111 48885 28120
rect 47691 27824 47733 27833
rect 47691 27784 47692 27824
rect 47732 27784 47733 27824
rect 47691 27775 47733 27784
rect 47788 27749 47828 27780
rect 47787 27740 47829 27749
rect 47787 27700 47788 27740
rect 47828 27700 47829 27740
rect 47787 27691 47829 27700
rect 48844 27740 48884 28111
rect 48844 27691 48884 27700
rect 47596 27656 47636 27665
rect 47596 26909 47636 27616
rect 47691 27656 47733 27665
rect 47691 27616 47692 27656
rect 47732 27616 47733 27656
rect 47691 27607 47733 27616
rect 47788 27656 47828 27691
rect 47692 27522 47732 27607
rect 47788 27581 47828 27616
rect 49228 27656 49268 28456
rect 49228 27607 49268 27616
rect 47787 27572 47829 27581
rect 47787 27532 47788 27572
rect 47828 27532 47829 27572
rect 47787 27523 47829 27532
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 47595 26900 47637 26909
rect 47595 26860 47596 26900
rect 47636 26860 47637 26900
rect 47595 26851 47637 26860
rect 47444 26776 47540 26816
rect 48267 26816 48309 26825
rect 48267 26776 48268 26816
rect 48308 26776 48309 26816
rect 47404 26767 47444 26776
rect 48267 26767 48309 26776
rect 47979 26648 48021 26657
rect 47979 26608 47980 26648
rect 48020 26608 48021 26648
rect 47979 26599 48021 26608
rect 47212 26144 47252 26153
rect 47115 26060 47157 26069
rect 47115 26020 47116 26060
rect 47156 26020 47157 26060
rect 47115 26011 47157 26020
rect 47019 25976 47061 25985
rect 47019 25936 47020 25976
rect 47060 25936 47061 25976
rect 47019 25927 47061 25936
rect 47020 25842 47060 25927
rect 46923 25640 46965 25649
rect 46923 25600 46924 25640
rect 46964 25600 46965 25640
rect 46923 25591 46965 25600
rect 46828 25507 46868 25516
rect 46731 25388 46773 25397
rect 46731 25348 46732 25388
rect 46772 25348 46964 25388
rect 46731 25339 46773 25348
rect 46732 25254 46772 25339
rect 46827 24884 46869 24893
rect 46827 24844 46828 24884
rect 46868 24844 46869 24884
rect 46827 24835 46869 24844
rect 46828 24800 46868 24835
rect 46828 24749 46868 24760
rect 46732 24632 46772 24641
rect 46636 24592 46732 24632
rect 46636 24053 46676 24592
rect 46732 24583 46772 24592
rect 46924 24632 46964 25348
rect 47020 25220 47060 25229
rect 47020 24893 47060 25180
rect 47019 24884 47061 24893
rect 47019 24844 47020 24884
rect 47060 24844 47061 24884
rect 47019 24835 47061 24844
rect 46924 24583 46964 24592
rect 47020 24632 47060 24641
rect 47116 24632 47156 26011
rect 47060 24592 47156 24632
rect 47020 24583 47060 24592
rect 46635 24044 46677 24053
rect 46635 24004 46636 24044
rect 46676 24004 46677 24044
rect 46635 23995 46677 24004
rect 46155 23960 46197 23969
rect 46155 23920 46156 23960
rect 46196 23920 46197 23960
rect 46155 23911 46197 23920
rect 45580 23248 45908 23288
rect 45484 23129 45524 23214
rect 45580 23204 45620 23248
rect 45580 23155 45620 23164
rect 45291 23120 45333 23129
rect 45291 23080 45292 23120
rect 45332 23080 45333 23120
rect 45291 23071 45333 23080
rect 45483 23120 45525 23129
rect 45483 23080 45484 23120
rect 45524 23080 45525 23120
rect 45483 23071 45525 23080
rect 45676 23120 45716 23129
rect 45580 23060 45620 23064
rect 45676 23060 45716 23080
rect 45868 23120 45908 23248
rect 45868 23071 45908 23080
rect 45964 23120 46004 23743
rect 46060 23465 46100 23752
rect 46059 23456 46101 23465
rect 46059 23416 46060 23456
rect 46100 23416 46101 23456
rect 46059 23407 46101 23416
rect 46636 23381 46676 23995
rect 46924 23960 46964 23969
rect 46732 23920 46924 23960
rect 46155 23372 46197 23381
rect 46155 23332 46156 23372
rect 46196 23332 46197 23372
rect 46155 23323 46197 23332
rect 46635 23372 46677 23381
rect 46635 23332 46636 23372
rect 46676 23332 46677 23372
rect 46635 23323 46677 23332
rect 45964 23071 46004 23080
rect 46156 23120 46196 23323
rect 46635 23204 46677 23213
rect 46635 23164 46636 23204
rect 46676 23164 46677 23204
rect 46635 23155 46677 23164
rect 46156 23060 46196 23080
rect 45580 23045 45812 23060
rect 45579 23036 45812 23045
rect 45579 22996 45580 23036
rect 45620 23020 45812 23036
rect 45620 22996 45621 23020
rect 45579 22987 45621 22996
rect 45196 22492 45620 22532
rect 44908 22448 44948 22457
rect 44948 22408 45428 22448
rect 44908 22399 44948 22408
rect 44812 22231 44852 22240
rect 45004 22280 45044 22289
rect 44812 21776 44852 21785
rect 44716 21736 44812 21776
rect 44812 21617 44852 21736
rect 44811 21608 44853 21617
rect 44811 21568 44812 21608
rect 44852 21568 44853 21608
rect 44811 21559 44853 21568
rect 44620 20852 44660 20861
rect 44524 20812 44620 20852
rect 44620 20803 44660 20812
rect 44139 20768 44181 20777
rect 44139 20728 44140 20768
rect 44180 20728 44181 20768
rect 44139 20719 44181 20728
rect 44812 20768 44852 21559
rect 45004 21440 45044 22240
rect 45004 21391 45044 21400
rect 45196 22280 45236 22289
rect 45003 20936 45045 20945
rect 45003 20896 45004 20936
rect 45044 20896 45045 20936
rect 45003 20887 45045 20896
rect 44812 20719 44852 20728
rect 44907 20768 44949 20777
rect 44907 20728 44908 20768
rect 44948 20728 44949 20768
rect 44907 20719 44949 20728
rect 45004 20768 45044 20887
rect 45004 20719 45044 20728
rect 45100 20768 45140 20777
rect 45196 20768 45236 22240
rect 45388 22280 45428 22408
rect 45292 22112 45332 22121
rect 45292 21785 45332 22072
rect 45291 21776 45333 21785
rect 45291 21736 45292 21776
rect 45332 21736 45333 21776
rect 45388 21776 45428 22240
rect 45483 22280 45525 22289
rect 45483 22240 45484 22280
rect 45524 22240 45525 22280
rect 45483 22231 45525 22240
rect 45484 22146 45524 22231
rect 45388 21736 45524 21776
rect 45291 21727 45333 21736
rect 45291 21608 45333 21617
rect 45291 21568 45292 21608
rect 45332 21568 45333 21608
rect 45291 21559 45333 21568
rect 45388 21608 45428 21617
rect 45292 21474 45332 21559
rect 45388 21533 45428 21568
rect 45387 21524 45429 21533
rect 45387 21484 45388 21524
rect 45428 21484 45429 21524
rect 45484 21524 45524 21736
rect 45580 21608 45620 22492
rect 45772 22364 45812 23020
rect 46060 23020 46196 23060
rect 46348 23120 46388 23129
rect 45772 22324 45908 22364
rect 45676 22280 45716 22289
rect 45676 21785 45716 22240
rect 45868 22280 45908 22324
rect 45772 22196 45812 22205
rect 45675 21776 45717 21785
rect 45675 21736 45676 21776
rect 45716 21736 45717 21776
rect 45675 21727 45717 21736
rect 45676 21608 45716 21617
rect 45580 21568 45676 21608
rect 45676 21559 45716 21568
rect 45484 21484 45620 21524
rect 45387 21475 45429 21484
rect 45388 21281 45428 21475
rect 45387 21272 45429 21281
rect 45387 21232 45388 21272
rect 45428 21232 45429 21272
rect 45387 21223 45429 21232
rect 45140 20728 45236 20768
rect 45483 20768 45525 20777
rect 45483 20728 45484 20768
rect 45524 20728 45525 20768
rect 45580 20768 45620 21484
rect 45676 20768 45716 20777
rect 45580 20728 45676 20768
rect 45100 20719 45140 20728
rect 45483 20719 45525 20728
rect 45676 20719 45716 20728
rect 45772 20768 45812 22156
rect 45868 21533 45908 22240
rect 45964 21608 46004 21617
rect 45867 21524 45909 21533
rect 45867 21484 45868 21524
rect 45908 21484 45909 21524
rect 45867 21475 45909 21484
rect 45772 20719 45812 20728
rect 44908 20634 44948 20719
rect 45484 20634 45524 20719
rect 44236 20600 44276 20609
rect 44236 20105 44276 20560
rect 44428 20600 44468 20609
rect 44235 20096 44277 20105
rect 44235 20056 44236 20096
rect 44276 20056 44277 20096
rect 44235 20047 44277 20056
rect 43851 20012 43893 20021
rect 43851 19972 43852 20012
rect 43892 19972 43893 20012
rect 43851 19963 43893 19972
rect 44331 20012 44373 20021
rect 44331 19972 44332 20012
rect 44372 19972 44373 20012
rect 44428 20012 44468 20560
rect 45003 20600 45045 20609
rect 45003 20560 45004 20600
rect 45044 20560 45045 20600
rect 45003 20551 45045 20560
rect 45580 20600 45620 20609
rect 45964 20600 46004 21568
rect 46060 20777 46100 23020
rect 46156 22952 46196 22961
rect 46348 22952 46388 23080
rect 46196 22912 46388 22952
rect 46156 22903 46196 22912
rect 46444 22448 46484 22457
rect 46251 22280 46293 22289
rect 46251 22240 46252 22280
rect 46292 22240 46293 22280
rect 46251 22231 46293 22240
rect 46252 21020 46292 22231
rect 46348 21608 46388 21617
rect 46444 21608 46484 22408
rect 46388 21568 46484 21608
rect 46348 21559 46388 21568
rect 46636 21524 46676 23155
rect 46732 23120 46772 23920
rect 46924 23911 46964 23920
rect 46732 23071 46772 23080
rect 47212 23060 47252 26104
rect 47980 26144 48020 26599
rect 47980 26095 48020 26104
rect 48172 26144 48212 26153
rect 48075 26060 48117 26069
rect 48075 26020 48076 26060
rect 48116 26020 48117 26060
rect 48075 26011 48117 26020
rect 47596 25976 47636 25985
rect 47500 25936 47596 25976
rect 47404 25304 47444 25313
rect 47500 25304 47540 25936
rect 47596 25927 47636 25936
rect 48076 25926 48116 26011
rect 47979 25640 48021 25649
rect 47979 25600 47980 25640
rect 48020 25600 48021 25640
rect 47979 25591 48021 25600
rect 47444 25264 47540 25304
rect 47404 25255 47444 25264
rect 47595 23792 47637 23801
rect 47595 23752 47596 23792
rect 47636 23752 47637 23792
rect 47595 23743 47637 23752
rect 47596 23120 47636 23743
rect 47596 23071 47636 23080
rect 46924 23020 47252 23060
rect 46731 22280 46773 22289
rect 46731 22240 46732 22280
rect 46772 22240 46773 22280
rect 46731 22231 46773 22240
rect 46444 21484 46676 21524
rect 46348 21020 46388 21029
rect 46252 20980 46348 21020
rect 46348 20971 46388 20980
rect 46059 20768 46101 20777
rect 46059 20728 46060 20768
rect 46100 20728 46101 20768
rect 46059 20719 46101 20728
rect 46348 20768 46388 20777
rect 46444 20768 46484 21484
rect 46539 21356 46581 21365
rect 46539 21316 46540 21356
rect 46580 21316 46581 21356
rect 46539 21307 46581 21316
rect 46388 20728 46484 20768
rect 46540 20768 46580 21307
rect 46348 20719 46388 20728
rect 46540 20719 46580 20728
rect 46636 20768 46676 20777
rect 46732 20768 46772 22231
rect 46676 20728 46772 20768
rect 46636 20719 46676 20728
rect 45620 20560 46004 20600
rect 45580 20551 45620 20560
rect 44907 20180 44949 20189
rect 44907 20140 44908 20180
rect 44948 20140 44949 20180
rect 44907 20131 44949 20140
rect 44524 20012 44564 20021
rect 44428 19972 44524 20012
rect 44331 19963 44373 19972
rect 43852 19878 43892 19963
rect 44043 19928 44085 19937
rect 44043 19888 44044 19928
rect 44084 19888 44085 19928
rect 44043 19879 44085 19888
rect 43468 19424 43508 19433
rect 43508 19384 43604 19424
rect 43468 19375 43508 19384
rect 43564 18584 43604 19384
rect 44044 19256 44084 19879
rect 44044 19207 44084 19216
rect 44332 19844 44372 19963
rect 43660 19172 43700 19181
rect 43700 19132 43988 19172
rect 43660 19123 43700 19132
rect 43851 18920 43893 18929
rect 43851 18880 43852 18920
rect 43892 18880 43893 18920
rect 43851 18871 43893 18880
rect 43659 18752 43701 18761
rect 43659 18712 43660 18752
rect 43700 18712 43701 18752
rect 43659 18703 43701 18712
rect 43660 18668 43700 18703
rect 43660 18617 43700 18628
rect 43564 18535 43604 18544
rect 43756 18584 43796 18593
rect 43468 17744 43508 17753
rect 43508 17704 43604 17744
rect 43468 17695 43508 17704
rect 43564 16904 43604 17704
rect 43756 16913 43796 18544
rect 43564 16855 43604 16864
rect 43755 16904 43797 16913
rect 43755 16864 43756 16904
rect 43796 16864 43797 16904
rect 43755 16855 43797 16864
rect 43852 16820 43892 18871
rect 43948 18752 43988 19132
rect 44332 18929 44372 19804
rect 44524 19601 44564 19972
rect 44715 19928 44757 19937
rect 44715 19888 44716 19928
rect 44756 19888 44757 19928
rect 44715 19879 44757 19888
rect 44716 19794 44756 19879
rect 44523 19592 44565 19601
rect 44523 19552 44524 19592
rect 44564 19552 44565 19592
rect 44523 19543 44565 19552
rect 44908 19256 44948 20131
rect 44908 19207 44948 19216
rect 44619 19088 44661 19097
rect 44619 19048 44620 19088
rect 44660 19048 44661 19088
rect 44619 19039 44661 19048
rect 44331 18920 44373 18929
rect 44331 18880 44332 18920
rect 44372 18880 44373 18920
rect 44331 18871 44373 18880
rect 44044 18752 44084 18761
rect 43948 18712 44044 18752
rect 44044 18703 44084 18712
rect 44139 18752 44181 18761
rect 44139 18712 44140 18752
rect 44180 18712 44181 18752
rect 44139 18703 44181 18712
rect 43947 18584 43989 18593
rect 43947 18544 43948 18584
rect 43988 18544 43989 18584
rect 43947 18535 43989 18544
rect 44140 18584 44180 18703
rect 44620 18677 44660 19039
rect 44427 18668 44469 18677
rect 44427 18628 44428 18668
rect 44468 18628 44469 18668
rect 44427 18619 44469 18628
rect 44619 18668 44661 18677
rect 44619 18628 44620 18668
rect 44660 18628 44661 18668
rect 44619 18619 44661 18628
rect 44140 18535 44180 18544
rect 44236 18584 44276 18593
rect 43948 17837 43988 18535
rect 44236 18416 44276 18544
rect 44428 18584 44468 18619
rect 44428 18533 44468 18544
rect 44620 18584 44660 18619
rect 44620 18533 44660 18544
rect 44524 18416 44564 18425
rect 44236 18376 44524 18416
rect 44524 18367 44564 18376
rect 43947 17828 43989 17837
rect 43947 17788 43948 17828
rect 43988 17788 43989 17828
rect 43947 17779 43989 17788
rect 44043 17744 44085 17753
rect 44043 17704 44044 17744
rect 44084 17704 44085 17744
rect 44043 17695 44085 17704
rect 44332 17744 44372 17753
rect 44044 17156 44084 17695
rect 44332 17249 44372 17704
rect 44907 17576 44949 17585
rect 44907 17536 44908 17576
rect 44948 17536 44949 17576
rect 44907 17527 44949 17536
rect 44331 17240 44373 17249
rect 44331 17200 44332 17240
rect 44372 17200 44373 17240
rect 44331 17191 44373 17200
rect 44044 17107 44084 17116
rect 43947 17072 43989 17081
rect 43947 17032 43948 17072
rect 43988 17032 43989 17072
rect 43947 17023 43989 17032
rect 44140 17072 44180 17081
rect 43948 16938 43988 17023
rect 44140 16913 44180 17032
rect 44715 17072 44757 17081
rect 44715 17032 44716 17072
rect 44756 17032 44757 17072
rect 44715 17023 44757 17032
rect 44524 16988 44564 16997
rect 44139 16904 44181 16913
rect 44139 16864 44140 16904
rect 44180 16864 44181 16904
rect 44139 16855 44181 16864
rect 43852 16780 43988 16820
rect 43371 16736 43413 16745
rect 43371 16696 43372 16736
rect 43412 16696 43413 16736
rect 43371 16687 43413 16696
rect 43083 16652 43125 16661
rect 43083 16612 43084 16652
rect 43124 16612 43125 16652
rect 43083 16603 43125 16612
rect 43083 16400 43125 16409
rect 43083 16360 43084 16400
rect 43124 16360 43125 16400
rect 43083 16351 43125 16360
rect 43084 16266 43124 16351
rect 43172 16316 43214 16325
rect 43172 16276 43173 16316
rect 43213 16276 43214 16316
rect 43172 16267 43214 16276
rect 42988 15569 43028 16192
rect 43173 16247 43213 16267
rect 43173 16181 43213 16207
rect 43756 16232 43796 16241
rect 43796 16192 43892 16232
rect 43756 16183 43796 16192
rect 43372 16148 43412 16157
rect 43372 15905 43412 16108
rect 43371 15896 43413 15905
rect 43371 15856 43372 15896
rect 43412 15856 43413 15896
rect 43371 15847 43413 15856
rect 42987 15560 43029 15569
rect 42987 15520 42988 15560
rect 43028 15520 43029 15560
rect 42987 15511 43029 15520
rect 43179 15560 43221 15569
rect 43179 15520 43180 15560
rect 43220 15520 43221 15560
rect 43179 15511 43221 15520
rect 42699 14720 42741 14729
rect 42699 14680 42700 14720
rect 42740 14680 42741 14720
rect 42699 14671 42741 14680
rect 42892 14720 42932 14729
rect 42700 14586 42740 14671
rect 42796 14552 42836 14561
rect 42699 14216 42741 14225
rect 42699 14176 42700 14216
rect 42740 14176 42741 14216
rect 42699 14167 42741 14176
rect 42603 14132 42645 14141
rect 42603 14092 42604 14132
rect 42644 14092 42645 14132
rect 42603 14083 42645 14092
rect 42604 13796 42644 14083
rect 42700 14082 42740 14167
rect 42796 13922 42836 14512
rect 42892 14141 42932 14680
rect 42987 14720 43029 14729
rect 42987 14680 42988 14720
rect 43028 14680 43029 14720
rect 42987 14671 43029 14680
rect 43180 14720 43220 15511
rect 43852 15392 43892 16192
rect 43852 15343 43892 15352
rect 43180 14671 43220 14680
rect 43275 14720 43317 14729
rect 43275 14680 43276 14720
rect 43316 14680 43317 14720
rect 43275 14671 43317 14680
rect 43372 14720 43412 14729
rect 42988 14586 43028 14671
rect 43276 14586 43316 14671
rect 42891 14132 42933 14141
rect 42891 14092 42892 14132
rect 42932 14092 42933 14132
rect 42891 14083 42933 14092
rect 43179 14132 43221 14141
rect 43179 14092 43180 14132
rect 43220 14092 43221 14132
rect 43179 14083 43221 14092
rect 43180 13998 43220 14083
rect 43276 14048 43316 14057
rect 43372 14048 43412 14680
rect 43316 14008 43412 14048
rect 43564 14048 43604 14057
rect 42796 13882 43124 13922
rect 42892 13796 42932 13805
rect 42604 13756 42836 13796
rect 42699 13628 42741 13637
rect 42699 13588 42700 13628
rect 42740 13588 42741 13628
rect 42699 13579 42741 13588
rect 42412 13420 42548 13460
rect 42315 12956 42357 12965
rect 42315 12916 42316 12956
rect 42356 12916 42357 12956
rect 42315 12907 42357 12916
rect 41932 12402 41972 12487
rect 42028 12461 42068 12496
rect 42124 12496 42220 12536
rect 42027 12452 42069 12461
rect 42027 12412 42028 12452
rect 42068 12412 42069 12452
rect 42027 12403 42069 12412
rect 41836 11824 42068 11864
rect 41835 11696 41877 11705
rect 41835 11656 41836 11696
rect 41876 11656 41877 11696
rect 41835 11647 41877 11656
rect 41836 11562 41876 11647
rect 41932 11612 41972 11621
rect 41644 10480 41780 10520
rect 41644 10277 41684 10480
rect 41836 10436 41876 10445
rect 41932 10436 41972 11572
rect 42028 10529 42068 11824
rect 42124 11696 42164 12496
rect 42220 12487 42260 12496
rect 42412 12536 42452 13420
rect 42700 13208 42740 13579
rect 42796 13460 42836 13756
rect 42796 13217 42836 13420
rect 42700 12980 42740 13168
rect 42795 13208 42837 13217
rect 42795 13168 42796 13208
rect 42836 13168 42837 13208
rect 42795 13159 42837 13168
rect 42892 13208 42932 13756
rect 42892 13159 42932 13168
rect 43084 13208 43124 13882
rect 43276 13553 43316 14008
rect 43467 13880 43509 13889
rect 43467 13840 43468 13880
rect 43508 13840 43509 13880
rect 43467 13831 43509 13840
rect 43275 13544 43317 13553
rect 43275 13504 43276 13544
rect 43316 13504 43317 13544
rect 43275 13495 43317 13504
rect 43084 13159 43124 13168
rect 43468 13208 43508 13831
rect 43468 13159 43508 13168
rect 42700 12940 43124 12980
rect 43564 12965 43604 14008
rect 43659 14048 43701 14057
rect 43659 14008 43660 14048
rect 43700 14008 43701 14048
rect 43659 13999 43701 14008
rect 43660 13301 43700 13999
rect 43851 13880 43893 13889
rect 43851 13840 43852 13880
rect 43892 13840 43893 13880
rect 43851 13831 43893 13840
rect 43852 13746 43892 13831
rect 43659 13292 43701 13301
rect 43659 13252 43660 13292
rect 43700 13252 43701 13292
rect 43659 13243 43701 13252
rect 42412 12487 42452 12496
rect 42507 12536 42549 12545
rect 42507 12496 42508 12536
rect 42548 12496 42549 12536
rect 42507 12487 42549 12496
rect 42604 12536 42644 12545
rect 42508 12402 42548 12487
rect 42220 12284 42260 12293
rect 42260 12244 42452 12284
rect 42220 12235 42260 12244
rect 42220 11864 42260 11873
rect 42260 11824 42356 11864
rect 42220 11815 42260 11824
rect 42124 11656 42260 11696
rect 42027 10520 42069 10529
rect 42027 10480 42028 10520
rect 42068 10480 42069 10520
rect 42027 10471 42069 10480
rect 41740 10396 41836 10436
rect 41876 10396 41972 10436
rect 41643 10268 41685 10277
rect 41643 10228 41644 10268
rect 41684 10228 41685 10268
rect 41643 10219 41685 10228
rect 41740 10109 41780 10396
rect 41836 10387 41876 10396
rect 41931 10268 41973 10277
rect 41931 10228 41932 10268
rect 41972 10228 41973 10268
rect 42028 10268 42068 10471
rect 42220 10277 42260 11656
rect 42316 11444 42356 11824
rect 42412 11696 42452 12244
rect 42604 12041 42644 12496
rect 42987 12452 43029 12461
rect 42987 12412 42988 12452
rect 43028 12412 43029 12452
rect 42987 12403 43029 12412
rect 42892 12368 42932 12377
rect 42603 12032 42645 12041
rect 42603 11992 42604 12032
rect 42644 11992 42645 12032
rect 42603 11983 42645 11992
rect 42604 11705 42644 11983
rect 42412 11647 42452 11656
rect 42603 11696 42645 11705
rect 42603 11656 42604 11696
rect 42644 11656 42645 11696
rect 42603 11647 42645 11656
rect 42796 11696 42836 11705
rect 42892 11696 42932 12328
rect 42836 11656 42932 11696
rect 42796 11647 42836 11656
rect 42316 11404 42932 11444
rect 42603 11192 42645 11201
rect 42603 11152 42604 11192
rect 42644 11152 42645 11192
rect 42603 11143 42645 11152
rect 42604 11058 42644 11143
rect 42892 11024 42932 11404
rect 42892 10975 42932 10984
rect 42315 10940 42357 10949
rect 42315 10900 42316 10940
rect 42356 10900 42357 10940
rect 42315 10891 42357 10900
rect 42316 10436 42356 10891
rect 42124 10268 42164 10277
rect 42028 10228 42124 10268
rect 41931 10219 41973 10228
rect 42124 10219 42164 10228
rect 42219 10268 42261 10277
rect 42219 10228 42220 10268
rect 42260 10228 42261 10268
rect 42219 10219 42261 10228
rect 41835 10184 41877 10193
rect 41835 10144 41836 10184
rect 41876 10144 41877 10184
rect 41835 10135 41877 10144
rect 41739 10100 41781 10109
rect 41739 10060 41740 10100
rect 41780 10060 41781 10100
rect 41739 10051 41781 10060
rect 40972 9463 41012 9472
rect 41355 9512 41397 9521
rect 41355 9472 41356 9512
rect 41396 9472 41397 9512
rect 41355 9463 41397 9472
rect 41740 9512 41780 10051
rect 41740 9463 41780 9472
rect 41836 9512 41876 10135
rect 41932 9512 41972 10219
rect 42316 10193 42356 10396
rect 42988 10772 43028 12403
rect 43084 11024 43124 12940
rect 43275 12956 43317 12965
rect 43275 12916 43276 12956
rect 43316 12916 43317 12956
rect 43275 12907 43317 12916
rect 43563 12956 43605 12965
rect 43563 12916 43564 12956
rect 43604 12916 43605 12956
rect 43563 12907 43605 12916
rect 43276 11621 43316 12907
rect 43660 11696 43700 13243
rect 43948 12980 43988 16780
rect 44140 16493 44180 16855
rect 44524 16745 44564 16948
rect 44716 16904 44756 17023
rect 44908 16988 44948 17527
rect 44908 16939 44948 16948
rect 44716 16855 44756 16864
rect 44523 16736 44565 16745
rect 44523 16696 44524 16736
rect 44564 16696 44565 16736
rect 44523 16687 44565 16696
rect 44139 16484 44181 16493
rect 44139 16444 44140 16484
rect 44180 16444 44181 16484
rect 44139 16435 44181 16444
rect 44620 16232 44660 16241
rect 44660 16192 44756 16232
rect 44620 16183 44660 16192
rect 44619 14048 44661 14057
rect 44619 14008 44620 14048
rect 44660 14008 44661 14048
rect 44619 13999 44661 14008
rect 44620 13914 44660 13999
rect 44716 13301 44756 16192
rect 45004 15317 45044 20551
rect 45676 20105 45716 20136
rect 45675 20096 45717 20105
rect 45675 20056 45676 20096
rect 45716 20056 45717 20096
rect 45675 20047 45717 20056
rect 45291 20012 45333 20021
rect 45291 19972 45292 20012
rect 45332 19972 45333 20012
rect 45291 19963 45333 19972
rect 45676 20012 45716 20047
rect 45100 19844 45140 19853
rect 45100 16997 45140 19804
rect 45292 19349 45332 19963
rect 45484 19844 45524 19853
rect 45291 19340 45333 19349
rect 45291 19300 45292 19340
rect 45332 19300 45333 19340
rect 45291 19291 45333 19300
rect 45195 18668 45237 18677
rect 45195 18628 45196 18668
rect 45236 18628 45237 18668
rect 45195 18619 45237 18628
rect 45099 16988 45141 16997
rect 45099 16948 45100 16988
rect 45140 16948 45141 16988
rect 45099 16939 45141 16948
rect 45100 16820 45140 16829
rect 45100 16409 45140 16780
rect 45099 16400 45141 16409
rect 45099 16360 45100 16400
rect 45140 16360 45141 16400
rect 45099 16351 45141 16360
rect 45003 15308 45045 15317
rect 45003 15268 45004 15308
rect 45044 15268 45045 15308
rect 45003 15259 45045 15268
rect 45100 14888 45140 14897
rect 45004 14848 45100 14888
rect 45004 14048 45044 14848
rect 45100 14839 45140 14848
rect 45004 13999 45044 14008
rect 45196 13805 45236 18619
rect 45484 18593 45524 19804
rect 45483 18584 45525 18593
rect 45483 18544 45484 18584
rect 45524 18544 45525 18584
rect 45483 18535 45525 18544
rect 45676 17828 45716 19972
rect 46732 19928 46772 19937
rect 46636 19888 46732 19928
rect 46636 19256 46676 19888
rect 46732 19879 46772 19888
rect 46636 19207 46676 19216
rect 46252 19172 46292 19181
rect 46060 19088 46100 19097
rect 46060 18677 46100 19048
rect 46059 18668 46101 18677
rect 46059 18628 46060 18668
rect 46100 18628 46101 18668
rect 46059 18619 46101 18628
rect 46252 18425 46292 19132
rect 46732 18584 46772 18593
rect 46444 18544 46732 18584
rect 46251 18416 46293 18425
rect 46251 18376 46252 18416
rect 46292 18376 46293 18416
rect 46251 18367 46293 18376
rect 46444 17996 46484 18544
rect 46732 18535 46772 18544
rect 46827 18584 46869 18593
rect 46827 18544 46828 18584
rect 46868 18544 46869 18584
rect 46827 18535 46869 18544
rect 46828 18450 46868 18535
rect 46827 18332 46869 18341
rect 46827 18292 46828 18332
rect 46868 18292 46869 18332
rect 46827 18283 46869 18292
rect 46828 18089 46868 18283
rect 46827 18080 46869 18089
rect 46827 18040 46828 18080
rect 46868 18040 46869 18080
rect 46827 18031 46869 18040
rect 46444 17947 46484 17956
rect 45580 17788 45716 17828
rect 46443 17828 46485 17837
rect 46443 17788 46444 17828
rect 46484 17788 46485 17828
rect 45580 17669 45620 17788
rect 46443 17779 46485 17788
rect 46828 17828 46868 18031
rect 46828 17779 46868 17788
rect 45772 17744 45812 17753
rect 45676 17704 45772 17744
rect 45579 17660 45621 17669
rect 45579 17620 45580 17660
rect 45620 17620 45621 17660
rect 45579 17611 45621 17620
rect 45484 17576 45524 17585
rect 45292 17536 45484 17576
rect 45292 16325 45332 17536
rect 45484 17527 45524 17536
rect 45579 17492 45621 17501
rect 45579 17452 45580 17492
rect 45620 17452 45621 17492
rect 45579 17443 45621 17452
rect 45483 17408 45525 17417
rect 45483 17368 45484 17408
rect 45524 17368 45525 17408
rect 45483 17359 45525 17368
rect 45388 17081 45428 17166
rect 45387 17072 45429 17081
rect 45387 17032 45388 17072
rect 45428 17032 45429 17072
rect 45387 17023 45429 17032
rect 45484 16904 45524 17359
rect 45388 16864 45524 16904
rect 45291 16316 45333 16325
rect 45291 16276 45292 16316
rect 45332 16276 45333 16316
rect 45291 16267 45333 16276
rect 45292 16157 45332 16267
rect 45291 16148 45333 16157
rect 45291 16108 45292 16148
rect 45332 16108 45333 16148
rect 45291 16099 45333 16108
rect 45388 15392 45428 16864
rect 45483 16064 45525 16073
rect 45483 16024 45484 16064
rect 45524 16024 45525 16064
rect 45580 16064 45620 17443
rect 45676 17072 45716 17704
rect 45772 17695 45812 17704
rect 45963 17744 46005 17753
rect 45963 17704 45964 17744
rect 46004 17704 46005 17744
rect 45963 17695 46005 17704
rect 46156 17744 46196 17753
rect 45868 17660 45908 17669
rect 45771 17156 45813 17165
rect 45771 17116 45772 17156
rect 45812 17116 45813 17156
rect 45771 17107 45813 17116
rect 45676 16997 45716 17032
rect 45675 16988 45717 16997
rect 45675 16948 45676 16988
rect 45716 16948 45717 16988
rect 45675 16939 45717 16948
rect 45772 16484 45812 17107
rect 45772 16435 45812 16444
rect 45868 16232 45908 17620
rect 45964 17610 46004 17695
rect 46156 17165 46196 17704
rect 46251 17744 46293 17753
rect 46251 17704 46252 17744
rect 46292 17704 46293 17744
rect 46251 17695 46293 17704
rect 46444 17744 46484 17779
rect 46252 17610 46292 17695
rect 46155 17156 46197 17165
rect 46155 17116 46156 17156
rect 46196 17116 46197 17156
rect 46155 17107 46197 17116
rect 46252 17072 46292 17081
rect 46059 16820 46101 16829
rect 46059 16780 46060 16820
rect 46100 16780 46101 16820
rect 46059 16771 46101 16780
rect 46060 16686 46100 16771
rect 46252 16484 46292 17032
rect 46252 16435 46292 16444
rect 46251 16316 46293 16325
rect 46251 16276 46252 16316
rect 46292 16276 46293 16316
rect 46251 16267 46293 16276
rect 45964 16232 46004 16241
rect 45868 16192 45964 16232
rect 45964 16183 46004 16192
rect 46059 16232 46101 16241
rect 46252 16232 46292 16267
rect 46059 16192 46060 16232
rect 46100 16192 46196 16232
rect 46059 16183 46101 16192
rect 46060 16098 46100 16183
rect 45771 16064 45813 16073
rect 45580 16024 45716 16064
rect 45483 16015 45525 16024
rect 45484 15560 45524 16015
rect 45484 15511 45524 15520
rect 45580 15560 45620 15569
rect 45580 15392 45620 15520
rect 45388 15352 45620 15392
rect 45676 15560 45716 16024
rect 45771 16024 45772 16064
rect 45812 16024 45813 16064
rect 45771 16015 45813 16024
rect 45772 15930 45812 16015
rect 46059 15896 46101 15905
rect 46059 15856 46060 15896
rect 46100 15856 46101 15896
rect 46059 15847 46101 15856
rect 46060 15728 46100 15847
rect 46060 15679 46100 15688
rect 45676 15392 45716 15520
rect 45772 15560 45812 15569
rect 45964 15560 46004 15569
rect 45812 15520 45964 15560
rect 45772 15511 45812 15520
rect 45964 15511 46004 15520
rect 46156 15560 46196 16192
rect 46252 16181 46292 16192
rect 46156 15511 46196 15520
rect 46252 15560 46292 15569
rect 45676 15352 45812 15392
rect 45195 13796 45237 13805
rect 45195 13756 45196 13796
rect 45236 13756 45237 13796
rect 45195 13747 45237 13756
rect 44331 13292 44373 13301
rect 44331 13252 44332 13292
rect 44372 13252 44373 13292
rect 44331 13243 44373 13252
rect 44715 13292 44757 13301
rect 44715 13252 44716 13292
rect 44756 13252 44757 13292
rect 44715 13243 44757 13252
rect 44332 13208 44372 13243
rect 44332 13157 44372 13168
rect 43660 11647 43700 11656
rect 43852 12940 43988 12980
rect 45388 12965 45428 15352
rect 45483 13544 45525 13553
rect 45483 13504 45484 13544
rect 45524 13504 45525 13544
rect 45483 13495 45525 13504
rect 45484 13460 45524 13495
rect 45484 13409 45524 13420
rect 45579 13292 45621 13301
rect 45579 13252 45580 13292
rect 45620 13252 45621 13292
rect 45579 13243 45621 13252
rect 45387 12956 45429 12965
rect 43275 11612 43317 11621
rect 43275 11572 43276 11612
rect 43316 11572 43317 11612
rect 43275 11563 43317 11572
rect 43084 10975 43124 10984
rect 42315 10184 42357 10193
rect 42315 10144 42316 10184
rect 42356 10144 42357 10184
rect 42315 10135 42357 10144
rect 42508 9808 42836 9848
rect 42028 9640 42452 9680
rect 42028 9512 42068 9640
rect 41932 9472 42028 9512
rect 41836 9463 41876 9472
rect 42028 9463 42068 9472
rect 42220 9512 42260 9521
rect 39572 9304 40052 9344
rect 41547 9344 41589 9353
rect 41547 9304 41548 9344
rect 41588 9304 41589 9344
rect 39532 9295 39572 9304
rect 41547 9295 41589 9304
rect 41931 9344 41973 9353
rect 41931 9304 41932 9344
rect 41972 9304 41973 9344
rect 41931 9295 41973 9304
rect 42028 9344 42068 9353
rect 42220 9344 42260 9472
rect 42068 9304 42260 9344
rect 42316 9512 42356 9521
rect 42028 9295 42068 9304
rect 41548 9210 41588 9295
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 41547 8756 41589 8765
rect 41547 8716 41548 8756
rect 41588 8716 41589 8756
rect 41547 8707 41589 8716
rect 41548 8588 41588 8707
rect 41932 8672 41972 9295
rect 42316 9269 42356 9472
rect 42315 9260 42357 9269
rect 42315 9220 42316 9260
rect 42356 9220 42357 9260
rect 42315 9211 42357 9220
rect 41932 8623 41972 8632
rect 41548 8539 41588 8548
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 42412 8093 42452 9640
rect 42508 9512 42548 9808
rect 42699 9680 42741 9689
rect 42699 9640 42700 9680
rect 42740 9640 42741 9680
rect 42699 9631 42741 9640
rect 42796 9680 42836 9808
rect 42988 9773 43028 10732
rect 43564 10352 43604 10361
rect 43604 10312 43796 10352
rect 43564 10303 43604 10312
rect 42987 9764 43029 9773
rect 42987 9724 42988 9764
rect 43028 9724 43029 9764
rect 42987 9715 43029 9724
rect 42796 9631 42836 9640
rect 43083 9680 43125 9689
rect 43083 9640 43084 9680
rect 43124 9640 43125 9680
rect 43083 9631 43125 9640
rect 43659 9680 43701 9689
rect 43659 9640 43660 9680
rect 43700 9640 43701 9680
rect 43659 9631 43701 9640
rect 42508 9463 42548 9472
rect 42508 9260 42548 9269
rect 42508 8765 42548 9220
rect 42507 8756 42549 8765
rect 42507 8716 42508 8756
rect 42548 8716 42549 8756
rect 42507 8707 42549 8716
rect 42700 8672 42740 9631
rect 42987 9596 43029 9605
rect 42987 9556 42988 9596
rect 43028 9556 43029 9596
rect 42987 9547 43029 9556
rect 42891 9512 42933 9521
rect 42891 9472 42892 9512
rect 42932 9472 42933 9512
rect 42891 9463 42933 9472
rect 42988 9512 43028 9547
rect 42892 9378 42932 9463
rect 42988 9353 43028 9472
rect 43084 9512 43124 9631
rect 43084 9463 43124 9472
rect 42987 9344 43029 9353
rect 42987 9304 42988 9344
rect 43028 9304 43029 9344
rect 42987 9295 43029 9304
rect 43660 9092 43700 9631
rect 43756 9512 43796 10312
rect 43852 10277 43892 12940
rect 45387 12916 45388 12956
rect 45428 12916 45429 12956
rect 45387 12907 45429 12916
rect 45292 12536 45332 12545
rect 44811 12032 44853 12041
rect 44811 11992 44812 12032
rect 44852 11992 44853 12032
rect 44811 11983 44853 11992
rect 44812 11948 44852 11983
rect 45292 11957 45332 12496
rect 44812 11897 44852 11908
rect 45291 11948 45333 11957
rect 45291 11908 45292 11948
rect 45332 11908 45333 11948
rect 45291 11899 45333 11908
rect 45004 11864 45044 11873
rect 43947 11108 43989 11117
rect 43947 11068 43948 11108
rect 43988 11068 43989 11108
rect 43947 11059 43989 11068
rect 43948 11024 43988 11059
rect 43851 10268 43893 10277
rect 43851 10228 43852 10268
rect 43892 10228 43893 10268
rect 43851 10219 43893 10228
rect 43948 10184 43988 10984
rect 44140 11024 44180 11035
rect 44140 10949 44180 10984
rect 44332 11024 44372 11033
rect 44716 11024 44756 11033
rect 45004 11024 45044 11824
rect 44372 10984 44660 11024
rect 44332 10975 44372 10984
rect 44139 10940 44181 10949
rect 44139 10900 44140 10940
rect 44180 10900 44181 10940
rect 44139 10891 44181 10900
rect 44044 10772 44084 10781
rect 44084 10732 44564 10772
rect 44044 10723 44084 10732
rect 44331 10604 44373 10613
rect 44331 10564 44332 10604
rect 44372 10564 44373 10604
rect 44331 10555 44373 10564
rect 44139 10268 44181 10277
rect 44139 10228 44140 10268
rect 44180 10228 44181 10268
rect 44139 10219 44181 10228
rect 43948 10135 43988 10144
rect 43852 10100 43892 10109
rect 43852 9689 43892 10060
rect 43851 9680 43893 9689
rect 43851 9640 43852 9680
rect 43892 9640 43893 9680
rect 43851 9631 43893 9640
rect 43948 9512 43988 9521
rect 43756 9472 43948 9512
rect 43948 9463 43988 9472
rect 44140 9512 44180 10219
rect 44236 10184 44276 10193
rect 44236 9857 44276 10144
rect 44235 9848 44277 9857
rect 44235 9808 44236 9848
rect 44276 9808 44277 9848
rect 44235 9799 44277 9808
rect 44043 9260 44085 9269
rect 44043 9220 44044 9260
rect 44084 9220 44085 9260
rect 44043 9211 44085 9220
rect 44044 9126 44084 9211
rect 43660 9052 43988 9092
rect 43948 8924 43988 9052
rect 43948 8875 43988 8884
rect 44140 8765 44180 9472
rect 44236 9437 44276 9799
rect 44235 9428 44277 9437
rect 44235 9388 44236 9428
rect 44276 9388 44277 9428
rect 44235 9379 44277 9388
rect 44139 8756 44181 8765
rect 44139 8716 44140 8756
rect 44180 8716 44181 8756
rect 44139 8707 44181 8716
rect 42795 8672 42837 8681
rect 42700 8632 42796 8672
rect 42836 8632 42837 8672
rect 42795 8623 42837 8632
rect 42796 8538 42836 8623
rect 44140 8588 44180 8597
rect 43948 8504 43988 8513
rect 43988 8464 44084 8504
rect 43948 8455 43988 8464
rect 42411 8084 42453 8093
rect 42411 8044 42412 8084
rect 42452 8044 42453 8084
rect 42411 8035 42453 8044
rect 44044 8000 44084 8464
rect 44140 8177 44180 8548
rect 44139 8168 44181 8177
rect 44139 8128 44140 8168
rect 44180 8128 44181 8168
rect 44139 8119 44181 8128
rect 44140 8000 44180 8009
rect 44044 7960 44140 8000
rect 44140 7951 44180 7960
rect 44236 8000 44276 8009
rect 44332 8000 44372 10555
rect 44524 10184 44564 10732
rect 44620 10436 44660 10984
rect 44756 10984 45044 11024
rect 45580 11024 45620 13243
rect 45675 13208 45717 13217
rect 45675 13168 45676 13208
rect 45716 13168 45717 13208
rect 45675 13159 45717 13168
rect 45772 13208 45812 15352
rect 46252 14972 46292 15520
rect 46444 15485 46484 17704
rect 46539 17744 46581 17753
rect 46539 17704 46540 17744
rect 46580 17704 46581 17744
rect 46539 17695 46581 17704
rect 46540 17576 46580 17695
rect 46636 17576 46676 17585
rect 46540 17536 46636 17576
rect 46443 15476 46485 15485
rect 46443 15436 46444 15476
rect 46484 15436 46485 15476
rect 46443 15427 46485 15436
rect 46348 14972 46388 14981
rect 46252 14932 46348 14972
rect 46348 14923 46388 14932
rect 46060 14720 46100 14729
rect 45964 14680 46060 14720
rect 45964 14225 46004 14680
rect 46060 14671 46100 14680
rect 46155 14720 46197 14729
rect 46155 14680 46156 14720
rect 46196 14680 46197 14720
rect 46155 14671 46197 14680
rect 46348 14720 46388 14729
rect 46444 14720 46484 15427
rect 46540 14729 46580 17536
rect 46636 17527 46676 17536
rect 46636 17072 46676 17081
rect 46636 16400 46676 17032
rect 46732 16400 46772 16409
rect 46636 16360 46732 16400
rect 46732 16351 46772 16360
rect 46388 14680 46484 14720
rect 46539 14720 46581 14729
rect 46539 14680 46540 14720
rect 46580 14680 46581 14720
rect 46348 14671 46388 14680
rect 46539 14671 46581 14680
rect 46156 14586 46196 14671
rect 46924 14309 46964 23020
rect 47980 22541 48020 25591
rect 48172 25061 48212 26104
rect 48268 25985 48308 26767
rect 48747 26648 48789 26657
rect 48747 26608 48748 26648
rect 48788 26608 48789 26648
rect 48747 26599 48789 26608
rect 48748 26228 48788 26599
rect 48748 26179 48788 26188
rect 49132 26144 49172 26153
rect 48556 25985 48596 26070
rect 49132 25985 49172 26104
rect 48267 25976 48309 25985
rect 48267 25936 48268 25976
rect 48308 25936 48309 25976
rect 48267 25927 48309 25936
rect 48555 25976 48597 25985
rect 48555 25936 48556 25976
rect 48596 25936 48597 25976
rect 48555 25927 48597 25936
rect 49131 25976 49173 25985
rect 49131 25936 49132 25976
rect 49172 25936 49173 25976
rect 49131 25927 49173 25936
rect 48268 25304 48308 25927
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 49324 25565 49364 29800
rect 49419 29672 49461 29681
rect 49419 29632 49420 29672
rect 49460 29632 49461 29672
rect 49419 29623 49461 29632
rect 49420 28328 49460 29623
rect 49516 29345 49556 31135
rect 49612 30848 49652 31891
rect 49996 31781 50036 32059
rect 50092 32058 50132 32143
rect 49995 31772 50037 31781
rect 50284 31772 50324 34243
rect 50380 32705 50420 35923
rect 50572 35216 50612 36007
rect 50955 35972 50997 35981
rect 50955 35932 50956 35972
rect 50996 35932 50997 35972
rect 50955 35923 50997 35932
rect 50956 35838 50996 35923
rect 51340 35888 51380 35897
rect 51051 35804 51093 35813
rect 51051 35764 51052 35804
rect 51092 35764 51093 35804
rect 51051 35755 51093 35764
rect 50764 35720 50804 35729
rect 50572 35167 50612 35176
rect 50668 35680 50764 35720
rect 50475 34376 50517 34385
rect 50475 34336 50476 34376
rect 50516 34336 50517 34376
rect 50475 34327 50517 34336
rect 50572 34376 50612 34385
rect 50476 34242 50516 34327
rect 50475 33452 50517 33461
rect 50475 33412 50476 33452
rect 50516 33412 50517 33452
rect 50475 33403 50517 33412
rect 50379 32696 50421 32705
rect 50379 32656 50380 32696
rect 50420 32656 50421 32696
rect 50476 32696 50516 33403
rect 50572 32873 50612 34336
rect 50668 34376 50708 35680
rect 50764 35671 50804 35680
rect 50956 35216 50996 35225
rect 50956 34628 50996 35176
rect 50956 34579 50996 34588
rect 50668 33200 50708 34336
rect 50764 34376 50804 34385
rect 50956 34376 50996 34385
rect 50804 34336 50956 34376
rect 51052 34376 51092 35755
rect 51148 35048 51188 35057
rect 51340 35048 51380 35848
rect 51532 35888 51572 35897
rect 52396 35888 52436 35897
rect 52492 35888 52532 36520
rect 55660 35897 55700 37351
rect 55756 36476 55796 37360
rect 55947 37400 55989 37409
rect 55947 37360 55948 37400
rect 55988 37360 55989 37400
rect 55947 37351 55989 37360
rect 56044 37400 56084 37409
rect 55948 37266 55988 37351
rect 55852 37232 55892 37241
rect 55852 36821 55892 37192
rect 55851 36812 55893 36821
rect 55851 36772 55852 36812
rect 55892 36772 55893 36812
rect 55851 36763 55893 36772
rect 55947 36728 55989 36737
rect 55947 36688 55948 36728
rect 55988 36688 55989 36728
rect 55947 36679 55989 36688
rect 55948 36594 55988 36679
rect 56044 36569 56084 37360
rect 57388 37400 57428 37409
rect 56235 37232 56277 37241
rect 56235 37192 56236 37232
rect 56276 37192 56277 37232
rect 56235 37183 56277 37192
rect 56236 37098 56276 37183
rect 57388 36737 57428 37360
rect 58252 37400 58292 38023
rect 58252 37351 58292 37360
rect 57579 37232 57621 37241
rect 57579 37192 57580 37232
rect 57620 37192 57621 37232
rect 57579 37183 57621 37192
rect 57580 36821 57620 37183
rect 57579 36812 57621 36821
rect 57579 36772 57580 36812
rect 57620 36772 57621 36812
rect 57579 36763 57621 36772
rect 56427 36728 56469 36737
rect 57292 36728 57332 36737
rect 56427 36688 56428 36728
rect 56468 36688 56469 36728
rect 56427 36679 56469 36688
rect 57196 36688 57292 36728
rect 56043 36560 56085 36569
rect 56043 36520 56044 36560
rect 56084 36520 56085 36560
rect 56043 36511 56085 36520
rect 56331 36476 56373 36485
rect 55756 36436 55988 36476
rect 51572 35848 51764 35888
rect 51532 35839 51572 35848
rect 51435 35804 51477 35813
rect 51435 35764 51436 35804
rect 51476 35764 51477 35804
rect 51435 35755 51477 35764
rect 51436 35670 51476 35755
rect 51531 35300 51573 35309
rect 51531 35260 51532 35300
rect 51572 35260 51573 35300
rect 51531 35251 51573 35260
rect 51188 35008 51380 35048
rect 51436 35216 51476 35225
rect 51148 34999 51188 35008
rect 51243 34544 51285 34553
rect 51243 34504 51244 34544
rect 51284 34504 51285 34544
rect 51243 34495 51285 34504
rect 51148 34376 51188 34385
rect 51052 34336 51148 34376
rect 50764 34327 50804 34336
rect 50956 34327 50996 34336
rect 51148 34327 51188 34336
rect 51244 34376 51284 34495
rect 51436 34385 51476 35176
rect 51532 35216 51572 35251
rect 51532 35165 51572 35176
rect 51244 34327 51284 34336
rect 51435 34376 51477 34385
rect 51435 34336 51436 34376
rect 51476 34336 51477 34376
rect 51435 34327 51477 34336
rect 51627 33788 51669 33797
rect 51627 33748 51628 33788
rect 51668 33748 51669 33788
rect 51627 33739 51669 33748
rect 51628 33654 51668 33739
rect 51724 33461 51764 35848
rect 52436 35848 52532 35888
rect 53285 35888 53325 35897
rect 55564 35888 55604 35897
rect 52396 35839 52436 35848
rect 52012 35804 52052 35813
rect 52012 35384 52052 35764
rect 52299 35804 52341 35813
rect 52299 35764 52300 35804
rect 52340 35764 52341 35804
rect 52299 35755 52341 35764
rect 52204 35384 52244 35393
rect 52012 35344 52204 35384
rect 52204 35335 52244 35344
rect 51820 35216 51860 35227
rect 51820 35141 51860 35176
rect 52108 35216 52148 35225
rect 51819 35132 51861 35141
rect 51819 35092 51820 35132
rect 51860 35092 51861 35132
rect 51819 35083 51861 35092
rect 52108 35057 52148 35176
rect 52300 35216 52340 35755
rect 53285 35636 53325 35848
rect 54892 35848 55564 35888
rect 54412 35720 54452 35729
rect 54452 35680 54548 35720
rect 54412 35671 54452 35680
rect 53285 35596 53396 35636
rect 52300 35167 52340 35176
rect 52396 35344 52724 35384
rect 52396 35216 52436 35344
rect 52684 35300 52724 35344
rect 52684 35251 52724 35260
rect 52779 35300 52821 35309
rect 52779 35260 52780 35300
rect 52820 35260 52821 35300
rect 52779 35251 52821 35260
rect 52396 35167 52436 35176
rect 52588 35216 52628 35225
rect 52107 35048 52149 35057
rect 52107 35008 52108 35048
rect 52148 35008 52149 35048
rect 52107 34999 52149 35008
rect 52204 34553 52244 34638
rect 52012 34544 52052 34553
rect 52012 33704 52052 34504
rect 52203 34544 52245 34553
rect 52588 34544 52628 35176
rect 52780 35216 52820 35251
rect 53356 35225 53396 35596
rect 54508 35309 54548 35680
rect 54507 35300 54549 35309
rect 54507 35260 54508 35300
rect 54548 35260 54549 35300
rect 54507 35251 54549 35260
rect 54892 35300 54932 35848
rect 55564 35839 55604 35848
rect 55659 35888 55701 35897
rect 55659 35848 55660 35888
rect 55700 35848 55701 35888
rect 55659 35839 55701 35848
rect 55852 35888 55892 35897
rect 55948 35888 55988 36436
rect 56331 36436 56332 36476
rect 56372 36436 56373 36476
rect 56331 36427 56373 36436
rect 56044 35888 56084 35897
rect 55948 35848 56044 35888
rect 55852 35729 55892 35848
rect 56044 35839 56084 35848
rect 56140 35888 56180 35897
rect 55756 35720 55796 35729
rect 54892 35251 54932 35260
rect 55180 35680 55756 35720
rect 55180 35300 55220 35680
rect 55756 35671 55796 35680
rect 55851 35720 55893 35729
rect 55851 35680 55852 35720
rect 55892 35680 55893 35720
rect 55851 35671 55893 35680
rect 55467 35552 55509 35561
rect 55467 35512 55468 35552
rect 55508 35512 55509 35552
rect 55467 35503 55509 35512
rect 55180 35251 55220 35260
rect 52780 35165 52820 35176
rect 53355 35216 53397 35225
rect 53355 35176 53356 35216
rect 53396 35176 53397 35216
rect 53355 35167 53397 35176
rect 53739 35132 53781 35141
rect 53739 35092 53740 35132
rect 53780 35092 53781 35132
rect 53739 35083 53781 35092
rect 52203 34504 52204 34544
rect 52244 34504 52245 34544
rect 52203 34495 52245 34504
rect 52396 34504 52628 34544
rect 52203 34376 52245 34385
rect 52203 34336 52204 34376
rect 52244 34336 52245 34376
rect 52203 34327 52245 34336
rect 52396 34376 52436 34504
rect 52204 34242 52244 34327
rect 52012 33655 52052 33664
rect 51723 33452 51765 33461
rect 51723 33412 51724 33452
rect 51764 33412 51765 33452
rect 51723 33403 51765 33412
rect 50668 33160 50804 33200
rect 50764 33041 50804 33160
rect 50763 33032 50805 33041
rect 50763 32992 50764 33032
rect 50804 32992 50805 33032
rect 50763 32983 50805 32992
rect 50571 32864 50613 32873
rect 50571 32824 50572 32864
rect 50612 32824 50613 32864
rect 50571 32815 50613 32824
rect 51052 32864 51092 32873
rect 50763 32780 50805 32789
rect 50763 32740 50764 32780
rect 50804 32740 50805 32780
rect 50763 32731 50805 32740
rect 50476 32656 50612 32696
rect 50379 32647 50421 32656
rect 50475 32360 50517 32369
rect 50475 32320 50476 32360
rect 50516 32320 50517 32360
rect 50475 32311 50517 32320
rect 50476 32276 50516 32311
rect 50476 32225 50516 32236
rect 49995 31732 49996 31772
rect 50036 31732 50037 31772
rect 49995 31723 50037 31732
rect 50092 31732 50324 31772
rect 50380 32192 50420 32201
rect 49708 31361 49748 31446
rect 49707 31352 49749 31361
rect 49707 31312 49708 31352
rect 49748 31312 49749 31352
rect 49707 31303 49749 31312
rect 49900 31352 49940 31361
rect 49900 31193 49940 31312
rect 49996 31352 50036 31723
rect 50092 31361 50132 31732
rect 50188 31604 50228 31613
rect 50380 31604 50420 32152
rect 50572 32192 50612 32656
rect 50667 32612 50709 32621
rect 50667 32572 50668 32612
rect 50708 32572 50709 32612
rect 50667 32563 50709 32572
rect 50572 32143 50612 32152
rect 50475 31772 50517 31781
rect 50475 31732 50476 31772
rect 50516 31732 50517 31772
rect 50475 31723 50517 31732
rect 50228 31564 50420 31604
rect 50188 31555 50228 31564
rect 49996 31303 50036 31312
rect 50091 31352 50133 31361
rect 50091 31312 50092 31352
rect 50132 31312 50133 31352
rect 50091 31303 50133 31312
rect 50379 31352 50421 31361
rect 50379 31312 50380 31352
rect 50420 31312 50421 31352
rect 50379 31303 50421 31312
rect 50476 31352 50516 31723
rect 50476 31303 50516 31312
rect 50572 31352 50612 31361
rect 50668 31352 50708 32563
rect 50612 31312 50708 31352
rect 50572 31303 50612 31312
rect 50187 31268 50229 31277
rect 50187 31228 50188 31268
rect 50228 31228 50229 31268
rect 50187 31219 50229 31228
rect 49707 31184 49749 31193
rect 49804 31184 49844 31193
rect 49707 31144 49708 31184
rect 49748 31144 49804 31184
rect 49707 31135 49749 31144
rect 49804 31135 49844 31144
rect 49899 31184 49941 31193
rect 49899 31144 49900 31184
rect 49940 31144 49941 31184
rect 49899 31135 49941 31144
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 49612 30808 49748 30848
rect 49612 30680 49652 30689
rect 49515 29336 49557 29345
rect 49515 29296 49516 29336
rect 49556 29296 49557 29336
rect 49515 29287 49557 29296
rect 49516 29168 49556 29177
rect 49612 29168 49652 30640
rect 49708 30680 49748 30808
rect 49708 30631 49748 30640
rect 49803 30680 49845 30689
rect 49803 30640 49804 30680
rect 49844 30640 49845 30680
rect 49803 30631 49845 30640
rect 49900 30680 49940 30689
rect 49804 30546 49844 30631
rect 49900 30092 49940 30640
rect 50188 30596 50228 31219
rect 50380 30848 50420 31303
rect 50764 31193 50804 32731
rect 50860 32696 50900 32705
rect 50860 31781 50900 32656
rect 51052 32621 51092 32824
rect 51244 32864 51284 32875
rect 51244 32789 51284 32824
rect 51148 32780 51188 32789
rect 51051 32612 51093 32621
rect 51051 32572 51052 32612
rect 51092 32572 51093 32612
rect 51051 32563 51093 32572
rect 50955 32360 50997 32369
rect 51148 32360 51188 32740
rect 51243 32780 51285 32789
rect 51243 32740 51244 32780
rect 51284 32740 51285 32780
rect 51243 32731 51285 32740
rect 50955 32320 50956 32360
rect 50996 32320 50997 32360
rect 50955 32311 50997 32320
rect 51052 32320 51188 32360
rect 50859 31772 50901 31781
rect 50859 31732 50860 31772
rect 50900 31732 50901 31772
rect 50859 31723 50901 31732
rect 50859 31352 50901 31361
rect 50859 31312 50860 31352
rect 50900 31312 50901 31352
rect 50859 31303 50901 31312
rect 50860 31218 50900 31303
rect 50475 31184 50517 31193
rect 50475 31144 50476 31184
rect 50516 31144 50517 31184
rect 50475 31135 50517 31144
rect 50763 31184 50805 31193
rect 50763 31144 50764 31184
rect 50804 31144 50805 31184
rect 50956 31184 50996 32311
rect 51052 31352 51092 32320
rect 51148 32192 51188 32201
rect 51148 31604 51188 32152
rect 51532 32192 51572 32201
rect 51572 32152 51668 32192
rect 51532 32143 51572 32152
rect 51436 31604 51476 31613
rect 51148 31564 51436 31604
rect 51436 31555 51476 31564
rect 51628 31520 51668 32152
rect 51628 31471 51668 31480
rect 51148 31352 51188 31361
rect 51052 31312 51148 31352
rect 51148 31303 51188 31312
rect 51244 31352 51284 31361
rect 51244 31184 51284 31312
rect 50956 31144 51284 31184
rect 51436 31352 51476 31361
rect 51724 31352 51764 33403
rect 52396 33200 52436 34336
rect 52492 34376 52532 34385
rect 52492 33545 52532 34336
rect 52876 33704 52916 33713
rect 52491 33536 52533 33545
rect 52491 33496 52492 33536
rect 52532 33496 52533 33536
rect 52491 33487 52533 33496
rect 52204 33160 52436 33200
rect 52204 32789 52244 33160
rect 52300 33032 52340 33041
rect 52876 33032 52916 33664
rect 53451 33536 53493 33545
rect 53451 33496 53452 33536
rect 53492 33496 53493 33536
rect 53451 33487 53493 33496
rect 52340 32992 52916 33032
rect 52300 32983 52340 32992
rect 52203 32780 52245 32789
rect 52203 32740 52204 32780
rect 52244 32740 52245 32780
rect 52203 32731 52245 32740
rect 51819 32192 51861 32201
rect 51819 32152 51820 32192
rect 51860 32152 51861 32192
rect 51819 32143 51861 32152
rect 52396 32192 52436 32992
rect 52588 32864 52628 32873
rect 53452 32864 53492 33487
rect 53740 33377 53780 35083
rect 53836 34376 53876 34385
rect 53739 33368 53781 33377
rect 53739 33328 53740 33368
rect 53780 33328 53781 33368
rect 53739 33319 53781 33328
rect 53643 33032 53685 33041
rect 53643 32992 53644 33032
rect 53684 32992 53685 33032
rect 53643 32983 53685 32992
rect 52628 32824 52724 32864
rect 52588 32815 52628 32824
rect 50763 31135 50805 31144
rect 50380 30799 50420 30808
rect 50476 30689 50516 31135
rect 50571 30848 50613 30857
rect 50571 30808 50572 30848
rect 50612 30808 50613 30848
rect 51436 30848 51476 31312
rect 51532 31312 51764 31352
rect 51532 30857 51572 31312
rect 51531 30848 51573 30857
rect 51436 30808 51477 30848
rect 50571 30799 50613 30808
rect 50475 30680 50517 30689
rect 50475 30640 50476 30680
rect 50516 30640 50517 30680
rect 50475 30631 50517 30640
rect 50572 30680 50612 30799
rect 51437 30764 51477 30808
rect 51531 30808 51532 30848
rect 51572 30808 51573 30848
rect 51531 30799 51573 30808
rect 51436 30724 51477 30764
rect 51159 30701 51199 30710
rect 50572 30631 50612 30640
rect 50764 30680 50804 30689
rect 50188 30353 50228 30556
rect 50379 30428 50421 30437
rect 50284 30388 50380 30428
rect 50420 30388 50421 30428
rect 50187 30344 50229 30353
rect 50187 30304 50188 30344
rect 50228 30304 50229 30344
rect 50187 30295 50229 30304
rect 50188 30092 50228 30101
rect 49900 30052 50188 30092
rect 50188 30043 50228 30052
rect 50188 29672 50228 29681
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 49803 29336 49845 29345
rect 49803 29296 49804 29336
rect 49844 29296 49845 29336
rect 49803 29287 49845 29296
rect 50091 29336 50133 29345
rect 50091 29296 50092 29336
rect 50132 29296 50133 29336
rect 50091 29287 50133 29296
rect 50188 29336 50228 29632
rect 50284 29513 50324 30388
rect 50379 30379 50421 30388
rect 50380 30294 50420 30379
rect 50379 29924 50421 29933
rect 50379 29884 50380 29924
rect 50420 29884 50421 29924
rect 50379 29875 50421 29884
rect 50380 29790 50420 29875
rect 50283 29504 50325 29513
rect 50283 29464 50284 29504
rect 50324 29464 50325 29504
rect 50476 29504 50516 30631
rect 50668 30428 50708 30437
rect 50668 30269 50708 30388
rect 50667 30260 50709 30269
rect 50667 30220 50668 30260
rect 50708 30220 50709 30260
rect 50667 30211 50709 30220
rect 50764 30008 50804 30640
rect 50956 30680 50996 30689
rect 51199 30689 51284 30701
rect 51199 30680 51285 30689
rect 51199 30661 51244 30680
rect 51159 30652 51199 30661
rect 50956 30596 50996 30640
rect 51243 30640 51244 30661
rect 51284 30640 51285 30680
rect 51243 30631 51285 30640
rect 51340 30596 51380 30605
rect 50956 30556 51188 30596
rect 51052 30428 51092 30437
rect 50668 29968 50804 30008
rect 50860 30388 51052 30428
rect 50572 29681 50612 29766
rect 50571 29672 50613 29681
rect 50571 29632 50572 29672
rect 50612 29632 50613 29672
rect 50571 29623 50613 29632
rect 50476 29464 50612 29504
rect 50283 29455 50325 29464
rect 50188 29296 50516 29336
rect 49556 29128 49652 29168
rect 49707 29168 49749 29177
rect 49707 29128 49708 29168
rect 49748 29128 49749 29168
rect 49516 29119 49556 29128
rect 49707 29119 49749 29128
rect 49804 29168 49844 29287
rect 49804 29119 49844 29128
rect 50092 29168 50132 29287
rect 50092 29119 50132 29128
rect 49708 29034 49748 29119
rect 49515 29000 49557 29009
rect 50188 29000 50228 29296
rect 50476 29252 50516 29296
rect 50476 29203 50516 29212
rect 50380 29168 50420 29179
rect 50380 29093 50420 29128
rect 50379 29084 50421 29093
rect 50379 29044 50380 29084
rect 50420 29044 50421 29084
rect 50379 29035 50421 29044
rect 49515 28960 49516 29000
rect 49556 28960 49557 29000
rect 49515 28951 49557 28960
rect 49804 28960 50228 29000
rect 50283 29000 50325 29009
rect 50283 28960 50284 29000
rect 50324 28960 50325 29000
rect 49516 28866 49556 28951
rect 49611 28832 49653 28841
rect 49611 28792 49612 28832
rect 49652 28792 49653 28832
rect 49611 28783 49653 28792
rect 49420 28279 49460 28288
rect 49612 28328 49652 28783
rect 49612 28279 49652 28288
rect 49708 28328 49748 28337
rect 49804 28328 49844 28960
rect 50283 28951 50325 28960
rect 49748 28288 49844 28328
rect 49900 28328 49940 28337
rect 49708 28279 49748 28288
rect 49516 28160 49556 28169
rect 49900 28160 49940 28288
rect 49995 28328 50037 28337
rect 49995 28288 49996 28328
rect 50036 28288 50037 28328
rect 49995 28279 50037 28288
rect 50188 28328 50228 28337
rect 49996 28194 50036 28279
rect 50092 28169 50132 28254
rect 49556 28120 49940 28160
rect 50091 28160 50133 28169
rect 50091 28120 50092 28160
rect 50132 28120 50133 28160
rect 49516 28111 49556 28120
rect 50091 28111 50133 28120
rect 50188 28085 50228 28288
rect 50187 28076 50229 28085
rect 50187 28036 50188 28076
rect 50228 28036 50229 28076
rect 50187 28027 50229 28036
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 50092 27656 50132 27665
rect 49419 27572 49461 27581
rect 49419 27532 49420 27572
rect 49460 27532 49461 27572
rect 49419 27523 49461 27532
rect 49420 27068 49460 27523
rect 50092 27245 50132 27616
rect 49611 27236 49653 27245
rect 49611 27196 49612 27236
rect 49652 27196 49653 27236
rect 49611 27187 49653 27196
rect 50091 27236 50133 27245
rect 50091 27196 50092 27236
rect 50132 27196 50133 27236
rect 50091 27187 50133 27196
rect 49420 27019 49460 27028
rect 49612 26825 49652 27187
rect 50284 26993 50324 28951
rect 50572 28841 50612 29464
rect 50668 29000 50708 29968
rect 50860 29924 50900 30388
rect 51052 30379 51092 30388
rect 50955 30260 50997 30269
rect 51148 30260 51188 30556
rect 51340 30260 51380 30556
rect 50955 30220 50956 30260
rect 50996 30220 50997 30260
rect 50955 30211 50997 30220
rect 51052 30220 51188 30260
rect 51244 30220 51380 30260
rect 50764 29884 50900 29924
rect 50764 29840 50804 29884
rect 50956 29840 50996 30211
rect 51052 30017 51092 30220
rect 51244 30092 51284 30220
rect 51436 30101 51476 30724
rect 51532 30714 51572 30799
rect 51724 30512 51764 30521
rect 51628 30472 51724 30512
rect 51531 30176 51573 30185
rect 51531 30136 51532 30176
rect 51572 30136 51573 30176
rect 51531 30127 51573 30136
rect 51148 30052 51284 30092
rect 51435 30092 51477 30101
rect 51435 30052 51436 30092
rect 51476 30052 51477 30092
rect 51051 30008 51093 30017
rect 51051 29968 51052 30008
rect 51092 29968 51093 30008
rect 51051 29959 51093 29968
rect 50764 29791 50804 29800
rect 50860 29800 50996 29840
rect 51052 29840 51092 29851
rect 50860 29798 50900 29800
rect 51052 29765 51092 29800
rect 50860 29177 50900 29758
rect 51051 29756 51093 29765
rect 51051 29716 51052 29756
rect 51092 29716 51093 29756
rect 51051 29707 51093 29716
rect 50956 29672 50996 29681
rect 50956 29513 50996 29632
rect 51148 29588 51188 30052
rect 51435 30043 51477 30052
rect 51339 30008 51381 30017
rect 51339 29968 51340 30008
rect 51380 29968 51381 30008
rect 51339 29959 51381 29968
rect 51052 29548 51188 29588
rect 51244 29756 51284 29765
rect 50955 29504 50997 29513
rect 50955 29464 50956 29504
rect 50996 29464 50997 29504
rect 50955 29455 50997 29464
rect 51052 29261 51092 29548
rect 51244 29513 51284 29716
rect 51243 29504 51285 29513
rect 51243 29464 51244 29504
rect 51284 29464 51285 29504
rect 51243 29455 51285 29464
rect 51051 29252 51093 29261
rect 51051 29212 51052 29252
rect 51092 29212 51093 29252
rect 51051 29203 51093 29212
rect 50859 29168 50901 29177
rect 50859 29128 50860 29168
rect 50900 29128 50901 29168
rect 50859 29119 50901 29128
rect 50764 29000 50804 29009
rect 50668 28960 50764 29000
rect 50764 28951 50804 28960
rect 50956 28916 50996 28927
rect 51052 28916 51092 29203
rect 51340 29093 51380 29959
rect 51436 29765 51476 30043
rect 51435 29756 51477 29765
rect 51435 29716 51436 29756
rect 51476 29716 51477 29756
rect 51435 29707 51477 29716
rect 51148 29084 51188 29093
rect 51339 29084 51381 29093
rect 51188 29044 51284 29084
rect 51148 29035 51188 29044
rect 51052 28876 51188 28916
rect 50956 28841 50996 28876
rect 50571 28832 50613 28841
rect 50571 28792 50572 28832
rect 50612 28792 50613 28832
rect 50571 28783 50613 28792
rect 50955 28832 50997 28841
rect 50955 28792 50956 28832
rect 50996 28792 50997 28832
rect 50955 28783 50997 28792
rect 50475 28748 50517 28757
rect 50475 28708 50476 28748
rect 50516 28708 50517 28748
rect 50475 28699 50517 28708
rect 50476 28328 50516 28699
rect 50955 28664 50997 28673
rect 50955 28624 50956 28664
rect 50996 28624 50997 28664
rect 50955 28615 50997 28624
rect 50476 28279 50516 28288
rect 50572 28328 50612 28337
rect 50380 28160 50420 28171
rect 50572 28169 50612 28288
rect 50668 28328 50708 28337
rect 50380 28085 50420 28120
rect 50571 28160 50613 28169
rect 50571 28120 50572 28160
rect 50612 28120 50613 28160
rect 50571 28111 50613 28120
rect 50379 28076 50421 28085
rect 50379 28036 50380 28076
rect 50420 28036 50421 28076
rect 50379 28027 50421 28036
rect 50379 27908 50421 27917
rect 50379 27868 50380 27908
rect 50420 27868 50421 27908
rect 50379 27859 50421 27868
rect 50283 26984 50325 26993
rect 50092 26944 50284 26984
rect 50324 26944 50325 26984
rect 49611 26816 49653 26825
rect 49611 26776 49612 26816
rect 49652 26776 49653 26816
rect 49611 26767 49653 26776
rect 50092 26816 50132 26944
rect 50283 26935 50325 26944
rect 50092 26767 50132 26776
rect 50283 26816 50325 26825
rect 50283 26776 50284 26816
rect 50324 26776 50325 26816
rect 50283 26767 50325 26776
rect 50380 26816 50420 27859
rect 50572 26984 50612 28111
rect 50668 27917 50708 28288
rect 50667 27908 50709 27917
rect 50667 27868 50668 27908
rect 50708 27868 50709 27908
rect 50667 27859 50709 27868
rect 50380 26767 50420 26776
rect 50476 26944 50612 26984
rect 49515 26732 49557 26741
rect 49515 26692 49516 26732
rect 49556 26692 49557 26732
rect 49515 26683 49557 26692
rect 49420 26648 49460 26657
rect 49420 26321 49460 26608
rect 49419 26312 49461 26321
rect 49419 26272 49420 26312
rect 49460 26272 49461 26312
rect 49419 26263 49461 26272
rect 49323 25556 49365 25565
rect 49323 25516 49324 25556
rect 49364 25516 49365 25556
rect 49323 25507 49365 25516
rect 48171 25052 48213 25061
rect 48171 25012 48172 25052
rect 48212 25012 48213 25052
rect 48171 25003 48213 25012
rect 48268 23801 48308 25264
rect 49420 25136 49460 25147
rect 49420 25061 49460 25096
rect 49419 25052 49461 25061
rect 49419 25012 49420 25052
rect 49460 25012 49461 25052
rect 49419 25003 49461 25012
rect 48556 24464 48596 24473
rect 48556 24380 48596 24424
rect 48364 24340 48596 24380
rect 48267 23792 48309 23801
rect 48267 23752 48268 23792
rect 48308 23752 48309 23792
rect 48364 23792 48404 24340
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 48747 24044 48789 24053
rect 48747 24004 48748 24044
rect 48788 24004 48789 24044
rect 48747 23995 48789 24004
rect 48460 23792 48500 23801
rect 48364 23752 48460 23792
rect 48267 23743 48309 23752
rect 48460 23743 48500 23752
rect 48075 23708 48117 23717
rect 48075 23668 48076 23708
rect 48116 23668 48117 23708
rect 48075 23659 48117 23668
rect 48076 23574 48116 23659
rect 48748 23288 48788 23995
rect 49323 23792 49365 23801
rect 49323 23752 49324 23792
rect 49364 23752 49365 23792
rect 49323 23743 49365 23752
rect 49324 23658 49364 23743
rect 48748 23129 48788 23248
rect 49035 23288 49077 23297
rect 49035 23248 49036 23288
rect 49076 23248 49077 23288
rect 49035 23239 49077 23248
rect 48747 23120 48789 23129
rect 48747 23080 48748 23120
rect 48788 23080 48789 23120
rect 48747 23071 48789 23080
rect 48939 23120 48981 23129
rect 48939 23080 48940 23120
rect 48980 23080 48981 23120
rect 48939 23071 48981 23080
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 47979 22532 48021 22541
rect 48940 22532 48980 23071
rect 47979 22492 47980 22532
rect 48020 22492 48021 22532
rect 47979 22483 48021 22492
rect 48652 22492 48980 22532
rect 48172 22448 48212 22457
rect 48076 22408 48172 22448
rect 47212 21608 47252 21617
rect 47212 20189 47252 21568
rect 47691 21356 47733 21365
rect 47691 21316 47692 21356
rect 47732 21316 47733 21356
rect 47691 21307 47733 21316
rect 47692 20768 47732 21307
rect 47692 20719 47732 20728
rect 48076 20768 48116 22408
rect 48172 22399 48212 22408
rect 48555 22280 48597 22289
rect 48555 22240 48556 22280
rect 48596 22240 48597 22280
rect 48555 22231 48597 22240
rect 48652 22280 48692 22492
rect 49036 22448 49076 23239
rect 49516 23060 49556 26683
rect 49612 26153 49652 26767
rect 50187 26732 50229 26741
rect 50187 26692 50188 26732
rect 50228 26692 50229 26732
rect 50187 26683 50229 26692
rect 50188 26598 50228 26683
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 50187 26480 50229 26489
rect 50187 26440 50188 26480
rect 50228 26440 50229 26480
rect 50187 26431 50229 26440
rect 50188 26321 50228 26431
rect 50187 26312 50229 26321
rect 50187 26272 50188 26312
rect 50228 26272 50229 26312
rect 50187 26263 50229 26272
rect 49611 26144 49653 26153
rect 49611 26104 49612 26144
rect 49652 26104 49653 26144
rect 49611 26095 49653 26104
rect 49995 26144 50037 26153
rect 49995 26104 49996 26144
rect 50036 26104 50037 26144
rect 49995 26095 50037 26104
rect 49996 26010 50036 26095
rect 50284 25976 50324 26767
rect 50476 26312 50516 26944
rect 50572 26816 50612 26827
rect 50572 26741 50612 26776
rect 50668 26816 50708 26825
rect 50571 26732 50613 26741
rect 50571 26692 50572 26732
rect 50612 26692 50613 26732
rect 50571 26683 50613 26692
rect 50668 26321 50708 26776
rect 50860 26816 50900 26825
rect 50763 26648 50805 26657
rect 50763 26608 50764 26648
rect 50804 26608 50805 26648
rect 50763 26599 50805 26608
rect 50764 26514 50804 26599
rect 50667 26312 50709 26321
rect 50476 26272 50612 26312
rect 50284 25936 50420 25976
rect 49611 25556 49653 25565
rect 49611 25516 49612 25556
rect 49652 25516 49653 25556
rect 49611 25507 49653 25516
rect 49612 24557 49652 25507
rect 49995 25304 50037 25313
rect 49995 25264 49996 25304
rect 50036 25264 50037 25304
rect 49995 25255 50037 25264
rect 49996 25136 50036 25255
rect 49996 25096 50228 25136
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 50188 24800 50228 25096
rect 50380 24977 50420 25936
rect 50572 25472 50612 26272
rect 50667 26272 50668 26312
rect 50708 26272 50709 26312
rect 50667 26263 50709 26272
rect 50572 25432 50708 25472
rect 50668 25313 50708 25432
rect 50572 25304 50612 25313
rect 50572 25136 50612 25264
rect 50667 25304 50709 25313
rect 50667 25264 50668 25304
rect 50708 25264 50709 25304
rect 50667 25255 50709 25264
rect 50764 25304 50804 25313
rect 50764 25136 50804 25264
rect 50860 25304 50900 26776
rect 50860 25255 50900 25264
rect 50572 25096 50708 25136
rect 50764 25096 50805 25136
rect 50379 24968 50421 24977
rect 50379 24928 50380 24968
rect 50420 24928 50421 24968
rect 50379 24919 50421 24928
rect 50571 24968 50613 24977
rect 50571 24928 50572 24968
rect 50612 24928 50613 24968
rect 50571 24919 50613 24928
rect 50188 24751 50228 24760
rect 49707 24632 49749 24641
rect 49707 24592 49708 24632
rect 49748 24592 49749 24632
rect 49707 24583 49749 24592
rect 50379 24632 50421 24641
rect 50379 24592 50380 24632
rect 50420 24592 50421 24632
rect 50379 24583 50421 24592
rect 50572 24632 50612 24919
rect 50668 24893 50708 25096
rect 50765 25052 50805 25096
rect 50956 25052 50996 28615
rect 51052 28412 51092 28421
rect 51052 28253 51092 28372
rect 51051 28244 51093 28253
rect 51051 28204 51052 28244
rect 51092 28204 51093 28244
rect 51051 28195 51093 28204
rect 51148 26060 51188 28876
rect 51244 28580 51284 29044
rect 51339 29044 51340 29084
rect 51380 29044 51381 29084
rect 51339 29035 51381 29044
rect 51340 28916 51380 28925
rect 51436 28916 51476 29707
rect 51532 29084 51572 30127
rect 51628 29840 51668 30472
rect 51724 30463 51764 30472
rect 51723 29924 51765 29933
rect 51723 29884 51724 29924
rect 51764 29884 51765 29924
rect 51723 29875 51765 29884
rect 51628 29791 51668 29800
rect 51572 29044 51668 29084
rect 51532 29035 51572 29044
rect 51380 28876 51476 28916
rect 51340 28867 51380 28876
rect 51435 28664 51477 28673
rect 51435 28624 51436 28664
rect 51476 28624 51477 28664
rect 51435 28615 51477 28624
rect 51244 28531 51284 28540
rect 51243 28160 51285 28169
rect 51243 28120 51244 28160
rect 51284 28120 51285 28160
rect 51243 28111 51285 28120
rect 51244 28026 51284 28111
rect 51243 27908 51285 27917
rect 51243 27868 51244 27908
rect 51284 27868 51285 27908
rect 51243 27859 51285 27868
rect 51244 27824 51284 27859
rect 51244 27773 51284 27784
rect 51244 27404 51284 27413
rect 51244 26993 51284 27364
rect 51243 26984 51285 26993
rect 51243 26944 51244 26984
rect 51284 26944 51285 26984
rect 51243 26935 51285 26944
rect 51244 26816 51284 26825
rect 51244 26144 51284 26776
rect 51436 26564 51476 28615
rect 51628 27656 51668 29044
rect 51724 29009 51764 29875
rect 51820 29177 51860 32143
rect 52396 31361 52436 32152
rect 52395 31352 52437 31361
rect 52395 31312 52396 31352
rect 52436 31312 52437 31352
rect 52395 31303 52437 31312
rect 52491 29840 52533 29849
rect 52491 29800 52492 29840
rect 52532 29800 52533 29840
rect 52491 29791 52533 29800
rect 51819 29168 51861 29177
rect 51819 29128 51820 29168
rect 51860 29128 51861 29168
rect 51819 29119 51861 29128
rect 51820 29034 51860 29119
rect 52492 29093 52532 29791
rect 52491 29084 52533 29093
rect 52491 29044 52492 29084
rect 52532 29044 52533 29084
rect 52491 29035 52533 29044
rect 51723 29000 51765 29009
rect 51723 28960 51724 29000
rect 51764 28960 51765 29000
rect 51723 28951 51765 28960
rect 52492 28496 52532 28505
rect 51724 28421 51764 28452
rect 51723 28412 51765 28421
rect 51723 28372 51724 28412
rect 51764 28372 51765 28412
rect 51723 28363 51765 28372
rect 51724 28328 51764 28363
rect 51724 27917 51764 28288
rect 51819 28328 51861 28337
rect 51819 28288 51820 28328
rect 51860 28288 51861 28328
rect 51819 28279 51861 28288
rect 51916 28328 51956 28337
rect 52107 28328 52149 28337
rect 51956 28288 52052 28328
rect 51916 28279 51956 28288
rect 51723 27908 51765 27917
rect 51723 27868 51724 27908
rect 51764 27868 51765 27908
rect 51723 27859 51765 27868
rect 51723 27740 51765 27749
rect 51723 27700 51724 27740
rect 51764 27700 51765 27740
rect 51723 27691 51765 27700
rect 51628 27607 51668 27616
rect 51724 27606 51764 27691
rect 51820 27656 51860 28279
rect 51820 27607 51860 27616
rect 51915 27656 51957 27665
rect 51915 27616 51916 27656
rect 51956 27616 51957 27656
rect 51915 27607 51957 27616
rect 51916 27522 51956 27607
rect 51819 27404 51861 27413
rect 51819 27364 51820 27404
rect 51860 27364 51861 27404
rect 51819 27355 51861 27364
rect 51627 26984 51669 26993
rect 51627 26944 51628 26984
rect 51668 26944 51669 26984
rect 51627 26935 51669 26944
rect 51531 26816 51573 26825
rect 51531 26776 51532 26816
rect 51572 26776 51573 26816
rect 51531 26767 51573 26776
rect 51628 26816 51668 26935
rect 51628 26767 51668 26776
rect 51532 26682 51572 26767
rect 51436 26524 51572 26564
rect 51435 26144 51477 26153
rect 51244 26104 51436 26144
rect 51476 26104 51477 26144
rect 51435 26095 51477 26104
rect 51148 26020 51284 26060
rect 50764 25012 50996 25052
rect 51148 25892 51188 25901
rect 50667 24884 50709 24893
rect 50667 24844 50668 24884
rect 50708 24844 50709 24884
rect 50667 24835 50709 24844
rect 49611 24548 49653 24557
rect 49611 24508 49612 24548
rect 49652 24508 49653 24548
rect 49611 24499 49653 24508
rect 49708 24380 49748 24583
rect 49995 24548 50037 24557
rect 49995 24508 49996 24548
rect 50036 24508 50037 24548
rect 49995 24499 50037 24508
rect 49996 24414 50036 24499
rect 50380 24498 50420 24583
rect 50475 24464 50517 24473
rect 50475 24424 50476 24464
rect 50516 24424 50517 24464
rect 50475 24415 50517 24424
rect 49612 24340 49748 24380
rect 50188 24380 50228 24389
rect 50380 24380 50420 24389
rect 50228 24340 50324 24380
rect 49612 23288 49652 24340
rect 50188 24331 50228 24340
rect 50091 24044 50133 24053
rect 50091 24004 50092 24044
rect 50132 24004 50133 24044
rect 50091 23995 50133 24004
rect 50092 23633 50132 23995
rect 50187 23876 50229 23885
rect 50187 23836 50188 23876
rect 50228 23836 50229 23876
rect 50187 23827 50229 23836
rect 50091 23624 50133 23633
rect 50091 23584 50092 23624
rect 50132 23584 50133 23624
rect 50091 23575 50133 23584
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 49612 23239 49652 23248
rect 49995 23288 50037 23297
rect 49995 23248 49996 23288
rect 50036 23248 50037 23288
rect 49995 23239 50037 23248
rect 50092 23288 50141 23297
rect 50140 23248 50141 23288
rect 50092 23239 50141 23248
rect 49900 23129 49940 23214
rect 49899 23120 49941 23129
rect 49420 23036 49556 23060
rect 49804 23075 49844 23084
rect 49460 23020 49556 23036
rect 49420 22987 49460 22996
rect 49803 22996 49804 23045
rect 49899 23080 49900 23120
rect 49940 23080 49941 23120
rect 49899 23071 49941 23080
rect 49996 23120 50036 23239
rect 50100 23161 50140 23239
rect 49996 23071 50036 23080
rect 49844 22996 49845 23045
rect 49803 22987 49845 22996
rect 49612 22868 49652 22877
rect 48652 22231 48692 22240
rect 48748 22408 49076 22448
rect 49420 22828 49612 22868
rect 48748 22280 48788 22408
rect 48748 22231 48788 22240
rect 49420 22280 49460 22828
rect 49612 22819 49652 22828
rect 49420 22231 49460 22240
rect 49612 22280 49652 22289
rect 48556 22146 48596 22231
rect 48844 22112 48884 22121
rect 49516 22112 49556 22121
rect 48844 21608 48884 22072
rect 49132 22072 49516 22112
rect 48844 21559 48884 21568
rect 49035 21608 49077 21617
rect 49035 21568 49036 21608
rect 49076 21568 49077 21608
rect 49035 21559 49077 21568
rect 49132 21608 49172 22072
rect 49516 22063 49556 22072
rect 49612 21776 49652 22240
rect 49708 22280 49748 22289
rect 49804 22280 49844 22987
rect 50188 22364 50228 23827
rect 50284 23129 50324 24340
rect 50380 23885 50420 24340
rect 50379 23876 50421 23885
rect 50379 23836 50380 23876
rect 50420 23836 50421 23876
rect 50379 23827 50421 23836
rect 50476 23792 50516 24415
rect 50572 23969 50612 24592
rect 50668 24632 50708 24835
rect 50668 24583 50708 24592
rect 50764 24053 50804 25012
rect 51148 24893 51188 25852
rect 51147 24884 51189 24893
rect 51147 24844 51148 24884
rect 51188 24844 51189 24884
rect 51147 24835 51189 24844
rect 50860 24632 50900 24643
rect 50860 24557 50900 24592
rect 51052 24632 51092 24641
rect 50859 24548 50901 24557
rect 50859 24508 50860 24548
rect 50900 24508 50901 24548
rect 50859 24499 50901 24508
rect 50956 24380 50996 24389
rect 50860 24340 50956 24380
rect 50763 24044 50805 24053
rect 50763 24004 50764 24044
rect 50804 24004 50805 24044
rect 50763 23995 50805 24004
rect 50860 23969 50900 24340
rect 50956 24331 50996 24340
rect 50571 23960 50613 23969
rect 50571 23920 50572 23960
rect 50612 23920 50613 23960
rect 50571 23911 50613 23920
rect 50859 23960 50901 23969
rect 50859 23920 50860 23960
rect 50900 23920 50901 23960
rect 50859 23911 50901 23920
rect 50668 23792 50708 23801
rect 50476 23752 50612 23792
rect 50476 23624 50516 23633
rect 50476 23213 50516 23584
rect 50475 23204 50517 23213
rect 50475 23164 50476 23204
rect 50516 23164 50517 23204
rect 50475 23155 50517 23164
rect 50283 23120 50325 23129
rect 50283 23080 50284 23120
rect 50324 23080 50325 23120
rect 50283 23071 50325 23080
rect 50380 23120 50420 23129
rect 50380 23060 50420 23080
rect 50572 23060 50612 23752
rect 50668 23381 50708 23752
rect 50860 23792 50900 23911
rect 50955 23876 50997 23885
rect 50955 23836 50956 23876
rect 50996 23836 50997 23876
rect 50955 23827 50997 23836
rect 50860 23743 50900 23752
rect 50956 23792 50996 23827
rect 50956 23741 50996 23752
rect 50763 23708 50805 23717
rect 50763 23668 50764 23708
rect 50804 23668 50805 23708
rect 50763 23659 50805 23668
rect 50764 23574 50804 23659
rect 50667 23372 50709 23381
rect 50667 23332 50668 23372
rect 50708 23332 50709 23372
rect 50667 23323 50709 23332
rect 50859 23372 50901 23381
rect 50859 23332 50860 23372
rect 50900 23332 50901 23372
rect 50859 23323 50901 23332
rect 51052 23330 51092 24592
rect 51244 24548 51284 26020
rect 51436 25304 51476 26095
rect 51532 26060 51572 26524
rect 51723 26144 51765 26153
rect 51723 26104 51724 26144
rect 51764 26104 51765 26144
rect 51820 26144 51860 27355
rect 51916 27068 51956 27077
rect 52012 27068 52052 28288
rect 52107 28288 52108 28328
rect 52148 28288 52149 28328
rect 52107 28279 52149 28288
rect 52300 28328 52340 28337
rect 52108 28194 52148 28279
rect 52204 28244 52244 28253
rect 52107 27740 52149 27749
rect 52107 27700 52108 27740
rect 52148 27700 52149 27740
rect 52107 27691 52149 27700
rect 52108 27606 52148 27691
rect 52204 27665 52244 28204
rect 52300 28001 52340 28288
rect 52395 28160 52437 28169
rect 52395 28120 52396 28160
rect 52436 28120 52437 28160
rect 52395 28111 52437 28120
rect 52299 27992 52341 28001
rect 52299 27952 52300 27992
rect 52340 27952 52341 27992
rect 52299 27943 52341 27952
rect 52203 27656 52245 27665
rect 52203 27616 52204 27656
rect 52244 27616 52245 27656
rect 52203 27607 52245 27616
rect 52107 27404 52149 27413
rect 52107 27364 52108 27404
rect 52148 27364 52149 27404
rect 52107 27355 52149 27364
rect 51956 27028 52052 27068
rect 51916 27019 51956 27028
rect 52108 26900 52148 27355
rect 52108 26851 52148 26860
rect 52300 26825 52340 27943
rect 52396 27581 52436 28111
rect 52492 27656 52532 28456
rect 52587 28328 52629 28337
rect 52587 28288 52588 28328
rect 52628 28288 52629 28328
rect 52587 28279 52629 28288
rect 52492 27607 52532 27616
rect 52395 27572 52437 27581
rect 52395 27532 52396 27572
rect 52436 27532 52437 27572
rect 52395 27523 52437 27532
rect 52299 26816 52341 26825
rect 52299 26776 52300 26816
rect 52340 26776 52341 26816
rect 52299 26767 52341 26776
rect 52299 26648 52341 26657
rect 52299 26608 52300 26648
rect 52340 26608 52341 26648
rect 52299 26599 52341 26608
rect 52300 26321 52340 26599
rect 52588 26321 52628 28279
rect 52107 26312 52149 26321
rect 52107 26272 52108 26312
rect 52148 26272 52149 26312
rect 52107 26263 52149 26272
rect 52299 26312 52341 26321
rect 52299 26272 52300 26312
rect 52340 26272 52341 26312
rect 52299 26263 52341 26272
rect 52587 26312 52629 26321
rect 52587 26272 52588 26312
rect 52628 26272 52629 26312
rect 52587 26263 52629 26272
rect 52108 26228 52148 26263
rect 52012 26144 52052 26153
rect 51820 26104 52012 26144
rect 51723 26095 51765 26104
rect 51532 26011 51572 26020
rect 51724 25976 51764 26095
rect 51724 25927 51764 25936
rect 51819 25892 51861 25901
rect 51819 25852 51820 25892
rect 51860 25852 51861 25892
rect 51819 25843 51861 25852
rect 51820 25724 51860 25843
rect 51724 25684 51860 25724
rect 51724 25304 51764 25684
rect 51476 25264 51572 25304
rect 51436 25255 51476 25264
rect 51436 24800 51476 24809
rect 51339 24632 51381 24641
rect 51339 24592 51340 24632
rect 51380 24592 51381 24632
rect 51339 24583 51381 24592
rect 51244 24499 51284 24508
rect 51243 23960 51285 23969
rect 51243 23920 51244 23960
rect 51284 23920 51285 23960
rect 51243 23911 51285 23920
rect 51244 23806 51284 23911
rect 51147 23792 51189 23801
rect 51147 23752 51148 23792
rect 51188 23752 51189 23792
rect 51244 23757 51284 23766
rect 51340 23792 51380 24583
rect 51436 24557 51476 24760
rect 51435 24548 51477 24557
rect 51435 24508 51436 24548
rect 51476 24508 51477 24548
rect 51435 24499 51477 24508
rect 51532 24473 51572 25264
rect 51724 25255 51764 25264
rect 51820 25220 51860 25229
rect 51820 25136 51860 25180
rect 51724 25096 51860 25136
rect 51724 24893 51764 25096
rect 51916 25052 51956 26104
rect 52012 26095 52052 26104
rect 52108 25724 52148 26188
rect 51820 25012 51956 25052
rect 52012 25684 52148 25724
rect 52204 26144 52244 26153
rect 52300 26144 52340 26263
rect 52396 26144 52436 26153
rect 52300 26104 52396 26144
rect 51723 24884 51765 24893
rect 51723 24844 51724 24884
rect 51764 24844 51765 24884
rect 51723 24835 51765 24844
rect 51820 24557 51860 25012
rect 51915 24884 51957 24893
rect 51915 24844 51916 24884
rect 51956 24844 51957 24884
rect 51915 24835 51957 24844
rect 51819 24548 51861 24557
rect 51819 24508 51820 24548
rect 51860 24508 51861 24548
rect 51819 24499 51861 24508
rect 51531 24464 51573 24473
rect 51531 24424 51532 24464
rect 51572 24424 51573 24464
rect 51531 24415 51573 24424
rect 51819 24212 51861 24221
rect 51819 24172 51820 24212
rect 51860 24172 51861 24212
rect 51819 24163 51861 24172
rect 51436 23960 51476 23969
rect 51476 23920 51764 23960
rect 51436 23911 51476 23920
rect 51436 23792 51476 23801
rect 51147 23743 51189 23752
rect 51340 23752 51436 23792
rect 51148 23658 51188 23743
rect 51340 23624 51380 23752
rect 51436 23743 51476 23752
rect 51531 23792 51573 23801
rect 51531 23752 51532 23792
rect 51572 23752 51573 23792
rect 51531 23743 51573 23752
rect 51724 23792 51764 23920
rect 51724 23743 51764 23752
rect 51244 23584 51380 23624
rect 51435 23624 51477 23633
rect 51435 23584 51436 23624
rect 51476 23584 51477 23624
rect 51244 23540 51284 23584
rect 51435 23575 51477 23584
rect 50763 23204 50805 23213
rect 50763 23164 50764 23204
rect 50804 23164 50805 23204
rect 50763 23155 50805 23164
rect 50667 23120 50709 23129
rect 50667 23080 50668 23120
rect 50708 23080 50709 23120
rect 50667 23071 50709 23080
rect 50380 23020 50612 23060
rect 50379 22532 50421 22541
rect 50379 22492 50380 22532
rect 50420 22492 50421 22532
rect 50379 22483 50421 22492
rect 50380 22398 50420 22483
rect 50188 22315 50228 22324
rect 49748 22240 49844 22280
rect 50091 22280 50133 22289
rect 50091 22240 50092 22280
rect 50132 22240 50133 22280
rect 49708 22231 49748 22240
rect 50091 22231 50133 22240
rect 50092 22112 50132 22231
rect 50092 22072 50228 22112
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 49132 21559 49172 21568
rect 49420 21736 49652 21776
rect 49036 21474 49076 21559
rect 49420 21533 49460 21736
rect 49516 21608 49556 21617
rect 49419 21524 49461 21533
rect 49419 21484 49420 21524
rect 49460 21484 49461 21524
rect 49419 21475 49461 21484
rect 48364 21356 48404 21367
rect 48844 21365 48884 21450
rect 49516 21449 49556 21568
rect 49611 21608 49653 21617
rect 49611 21568 49612 21608
rect 49652 21568 49653 21608
rect 49611 21559 49653 21568
rect 49708 21608 49748 21617
rect 49612 21474 49652 21559
rect 49515 21440 49557 21449
rect 49515 21400 49516 21440
rect 49556 21400 49557 21440
rect 49708 21440 49748 21568
rect 50188 21608 50228 22072
rect 50379 21860 50421 21869
rect 49900 21440 49940 21449
rect 49708 21400 49900 21440
rect 49515 21391 49557 21400
rect 49900 21391 49940 21400
rect 48364 21281 48404 21316
rect 48843 21356 48885 21365
rect 48843 21316 48844 21356
rect 48884 21316 48885 21356
rect 48843 21307 48885 21316
rect 48363 21272 48405 21281
rect 48363 21232 48364 21272
rect 48404 21232 48405 21272
rect 48363 21223 48405 21232
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 50092 21020 50132 21029
rect 50188 21020 50228 21568
rect 50284 21820 50380 21860
rect 50420 21820 50421 21860
rect 50284 21608 50324 21820
rect 50379 21811 50421 21820
rect 50379 21692 50421 21701
rect 50379 21652 50380 21692
rect 50420 21652 50421 21692
rect 50379 21643 50421 21652
rect 50284 21029 50324 21568
rect 50132 20980 50228 21020
rect 50283 21020 50325 21029
rect 50283 20980 50284 21020
rect 50324 20980 50325 21020
rect 50092 20971 50132 20980
rect 50283 20971 50325 20980
rect 48076 20719 48116 20728
rect 48940 20768 48980 20777
rect 48940 20189 48980 20728
rect 50284 20768 50324 20777
rect 50380 20768 50420 21643
rect 50476 21608 50516 23020
rect 50668 22986 50708 23071
rect 50764 23070 50804 23155
rect 50763 22952 50805 22961
rect 50763 22912 50764 22952
rect 50804 22912 50805 22952
rect 50763 22903 50805 22912
rect 50572 22280 50612 22289
rect 50572 21869 50612 22240
rect 50764 22280 50804 22903
rect 50764 22231 50804 22240
rect 50668 22196 50708 22205
rect 50571 21860 50613 21869
rect 50571 21820 50572 21860
rect 50612 21820 50613 21860
rect 50571 21811 50613 21820
rect 50572 21608 50612 21617
rect 50476 21568 50572 21608
rect 50572 21559 50612 21568
rect 50668 21533 50708 22156
rect 50860 21776 50900 23323
rect 51052 23281 51092 23290
rect 51148 23500 51284 23540
rect 51148 22541 51188 23500
rect 51339 23204 51381 23213
rect 51339 23164 51340 23204
rect 51380 23164 51381 23204
rect 51244 23141 51284 23160
rect 51339 23155 51381 23164
rect 51244 23045 51284 23101
rect 51340 23070 51380 23155
rect 51436 23129 51476 23575
rect 51435 23120 51477 23129
rect 51435 23080 51436 23120
rect 51476 23080 51477 23120
rect 51435 23071 51477 23080
rect 51243 23036 51285 23045
rect 51243 22996 51244 23036
rect 51284 22996 51285 23036
rect 51243 22987 51285 22996
rect 51244 22956 51284 22987
rect 51436 22986 51476 23071
rect 51147 22532 51189 22541
rect 51147 22492 51148 22532
rect 51188 22492 51189 22532
rect 51147 22483 51189 22492
rect 50764 21736 50900 21776
rect 50667 21524 50709 21533
rect 50667 21484 50668 21524
rect 50708 21484 50709 21524
rect 50667 21475 50709 21484
rect 50764 21113 50804 21736
rect 51051 21692 51093 21701
rect 51051 21652 51052 21692
rect 51092 21652 51093 21692
rect 51051 21643 51093 21652
rect 50860 21608 50900 21619
rect 50860 21533 50900 21568
rect 50955 21608 50997 21617
rect 50955 21568 50956 21608
rect 50996 21568 50997 21608
rect 50955 21559 50997 21568
rect 50859 21524 50901 21533
rect 50859 21484 50860 21524
rect 50900 21484 50901 21524
rect 50859 21475 50901 21484
rect 50956 21474 50996 21559
rect 51052 21558 51092 21643
rect 51148 21608 51188 22483
rect 51148 21559 51188 21568
rect 51340 21440 51380 21449
rect 50763 21104 50805 21113
rect 50763 21064 50764 21104
rect 50804 21064 50805 21104
rect 50763 21055 50805 21064
rect 50324 20728 50420 20768
rect 50668 20768 50708 20777
rect 51340 20768 51380 21400
rect 51532 21281 51572 23743
rect 51820 23624 51860 24163
rect 51916 23708 51956 24835
rect 52012 24464 52052 25684
rect 52108 25556 52148 25565
rect 52204 25556 52244 26104
rect 52396 26095 52436 26104
rect 52588 26144 52628 26153
rect 52491 26060 52533 26069
rect 52588 26060 52628 26104
rect 52491 26020 52492 26060
rect 52532 26020 52628 26060
rect 52491 26011 52533 26020
rect 52684 25976 52724 32824
rect 53452 32815 53492 32824
rect 53547 32864 53589 32873
rect 53547 32824 53548 32864
rect 53588 32824 53589 32864
rect 53547 32815 53589 32824
rect 53644 32864 53684 32983
rect 53644 32815 53684 32824
rect 53740 32864 53780 32873
rect 53836 32864 53876 34336
rect 54028 34376 54068 34385
rect 53932 34208 53972 34217
rect 53932 33797 53972 34168
rect 54028 33881 54068 34336
rect 54124 34376 54164 34385
rect 54027 33872 54069 33881
rect 54027 33832 54028 33872
rect 54068 33832 54069 33872
rect 54027 33823 54069 33832
rect 53931 33788 53973 33797
rect 53931 33748 53932 33788
rect 53972 33748 53973 33788
rect 53931 33739 53973 33748
rect 54027 33704 54069 33713
rect 54027 33664 54028 33704
rect 54068 33664 54069 33704
rect 54027 33655 54069 33664
rect 54028 33620 54068 33655
rect 54028 33545 54068 33580
rect 54027 33536 54069 33545
rect 54027 33496 54028 33536
rect 54068 33496 54069 33536
rect 54027 33487 54069 33496
rect 54028 33456 54068 33487
rect 54027 33368 54069 33377
rect 54027 33328 54028 33368
rect 54068 33328 54069 33368
rect 54027 33319 54069 33328
rect 53780 32824 53876 32864
rect 53740 32815 53780 32824
rect 53548 32730 53588 32815
rect 53547 32612 53589 32621
rect 53547 32572 53548 32612
rect 53588 32572 53589 32612
rect 53547 32563 53589 32572
rect 53548 32360 53588 32563
rect 53548 32311 53588 32320
rect 53931 32192 53973 32201
rect 53931 32152 53932 32192
rect 53972 32152 53973 32192
rect 53931 32143 53973 32152
rect 53548 31940 53588 31951
rect 53548 31865 53588 31900
rect 53547 31856 53589 31865
rect 53547 31816 53548 31856
rect 53588 31816 53589 31856
rect 53547 31807 53589 31816
rect 53260 31339 53300 31348
rect 52876 31268 52916 31277
rect 52876 30521 52916 31228
rect 53260 31016 53300 31299
rect 53260 30976 53396 31016
rect 52875 30512 52917 30521
rect 52875 30472 52876 30512
rect 52916 30472 52917 30512
rect 52875 30463 52917 30472
rect 53356 30512 53396 30976
rect 53356 30463 53396 30472
rect 53644 29672 53684 29681
rect 53644 29261 53684 29632
rect 53643 29252 53685 29261
rect 53643 29212 53644 29252
rect 53684 29212 53685 29252
rect 53643 29203 53685 29212
rect 52972 29168 53012 29177
rect 52972 28505 53012 29128
rect 53356 29168 53396 29177
rect 53396 29128 53492 29168
rect 53356 29119 53396 29128
rect 52971 28496 53013 28505
rect 52971 28456 52972 28496
rect 53012 28456 53013 28496
rect 52971 28447 53013 28456
rect 53068 28328 53108 28337
rect 52588 25936 52724 25976
rect 52780 25976 52820 25985
rect 52492 25892 52532 25901
rect 52148 25516 52244 25556
rect 52396 25852 52492 25892
rect 52108 25507 52148 25516
rect 52107 25304 52149 25313
rect 52107 25264 52108 25304
rect 52148 25264 52149 25304
rect 52107 25255 52149 25264
rect 52108 24641 52148 25255
rect 52300 25220 52340 25229
rect 52204 24800 52244 24809
rect 52300 24800 52340 25180
rect 52244 24760 52340 24800
rect 52204 24751 52244 24760
rect 52107 24632 52149 24641
rect 52300 24632 52340 24641
rect 52107 24592 52108 24632
rect 52148 24592 52149 24632
rect 52107 24583 52149 24592
rect 52204 24592 52300 24632
rect 52204 24464 52244 24592
rect 52300 24583 52340 24592
rect 52396 24632 52436 25852
rect 52492 25843 52532 25852
rect 52588 25724 52628 25936
rect 52396 24583 52436 24592
rect 52492 25684 52628 25724
rect 52012 24424 52244 24464
rect 52107 23792 52149 23801
rect 52107 23752 52108 23792
rect 52148 23752 52149 23792
rect 52107 23743 52149 23752
rect 51916 23668 52052 23708
rect 51820 23584 51956 23624
rect 51819 23456 51861 23465
rect 51819 23416 51820 23456
rect 51860 23416 51861 23456
rect 51819 23407 51861 23416
rect 51724 23036 51764 23045
rect 51628 22280 51668 22289
rect 51724 22280 51764 22996
rect 51820 22625 51860 23407
rect 51819 22616 51861 22625
rect 51819 22576 51820 22616
rect 51860 22576 51861 22616
rect 51819 22567 51861 22576
rect 51668 22240 51764 22280
rect 51531 21272 51573 21281
rect 51531 21232 51532 21272
rect 51572 21232 51573 21272
rect 51531 21223 51573 21232
rect 50708 20728 51380 20768
rect 51532 20768 51572 20777
rect 51628 20768 51668 22240
rect 51916 21029 51956 23584
rect 52012 23540 52052 23668
rect 52108 23658 52148 23743
rect 52012 23500 52148 23540
rect 52011 23204 52053 23213
rect 52011 23164 52012 23204
rect 52052 23164 52053 23204
rect 52011 23155 52053 23164
rect 52012 22532 52052 23155
rect 52012 22483 52052 22492
rect 52108 22364 52148 23500
rect 52492 23129 52532 25684
rect 52684 25304 52724 25313
rect 52780 25304 52820 25936
rect 52724 25264 52820 25304
rect 52684 25255 52724 25264
rect 52587 25220 52629 25229
rect 52587 25180 52588 25220
rect 52628 25180 52629 25220
rect 52587 25171 52629 25180
rect 52588 24632 52628 25171
rect 52875 24632 52917 24641
rect 52588 24592 52724 24632
rect 52588 24464 52628 24473
rect 52588 23801 52628 24424
rect 52684 24053 52724 24592
rect 52875 24592 52876 24632
rect 52916 24592 52917 24632
rect 53068 24632 53108 28288
rect 53356 27656 53396 27665
rect 53356 27245 53396 27616
rect 53355 27236 53397 27245
rect 53355 27196 53356 27236
rect 53396 27196 53397 27236
rect 53355 27187 53397 27196
rect 53452 26984 53492 29128
rect 53932 29009 53972 32143
rect 54028 30437 54068 33319
rect 54124 32024 54164 34336
rect 54411 33872 54453 33881
rect 54411 33832 54412 33872
rect 54452 33832 54453 33872
rect 54411 33823 54453 33832
rect 54316 33704 54356 33713
rect 54316 33377 54356 33664
rect 54315 33368 54357 33377
rect 54315 33328 54316 33368
rect 54356 33328 54357 33368
rect 54315 33319 54357 33328
rect 54412 33140 54452 33823
rect 54508 33377 54548 35251
rect 54796 35216 54836 35225
rect 54796 35141 54836 35176
rect 54988 35216 55028 35225
rect 54795 35132 54837 35141
rect 54795 35092 54796 35132
rect 54836 35092 54837 35132
rect 54795 35083 54837 35092
rect 54604 33704 54644 33713
rect 54507 33368 54549 33377
rect 54507 33328 54508 33368
rect 54548 33328 54549 33368
rect 54507 33319 54549 33328
rect 54316 33100 54452 33140
rect 54220 32201 54260 32286
rect 54219 32192 54261 32201
rect 54219 32152 54220 32192
rect 54260 32152 54261 32192
rect 54219 32143 54261 32152
rect 54220 32024 54260 32033
rect 54124 31984 54220 32024
rect 54220 31975 54260 31984
rect 54123 31352 54165 31361
rect 54123 31312 54124 31352
rect 54164 31312 54165 31352
rect 54123 31303 54165 31312
rect 54124 31218 54164 31303
rect 54027 30428 54069 30437
rect 54027 30388 54028 30428
rect 54068 30388 54069 30428
rect 54027 30379 54069 30388
rect 54316 29261 54356 33100
rect 54412 32864 54452 32873
rect 54412 32789 54452 32824
rect 54507 32864 54549 32873
rect 54507 32824 54508 32864
rect 54548 32824 54549 32864
rect 54507 32815 54549 32824
rect 54604 32864 54644 33664
rect 54699 33704 54741 33713
rect 54699 33664 54700 33704
rect 54740 33664 54741 33704
rect 54699 33655 54741 33664
rect 54700 33570 54740 33655
rect 54796 33140 54836 35083
rect 54988 34889 55028 35176
rect 54987 34880 55029 34889
rect 54987 34840 54988 34880
rect 55028 34840 55029 34880
rect 54987 34831 55029 34840
rect 55084 33832 55412 33872
rect 54891 33788 54933 33797
rect 54891 33748 54892 33788
rect 54932 33748 54933 33788
rect 54891 33739 54933 33748
rect 54411 32780 54453 32789
rect 54411 32740 54412 32780
rect 54452 32740 54453 32780
rect 54411 32731 54453 32740
rect 54412 32360 54452 32731
rect 54508 32730 54548 32815
rect 54604 32705 54644 32824
rect 54700 33100 54836 33140
rect 54603 32696 54645 32705
rect 54603 32656 54604 32696
rect 54644 32656 54645 32696
rect 54603 32647 54645 32656
rect 54700 32369 54740 33100
rect 54795 32864 54837 32873
rect 54795 32824 54796 32864
rect 54836 32824 54837 32864
rect 54795 32815 54837 32824
rect 54892 32864 54932 33739
rect 54988 33536 55028 33545
rect 55084 33536 55124 33832
rect 55028 33496 55124 33536
rect 55180 33704 55220 33713
rect 54988 33487 55028 33496
rect 55180 33461 55220 33664
rect 55275 33704 55317 33713
rect 55275 33664 55276 33704
rect 55316 33664 55317 33704
rect 55275 33655 55317 33664
rect 55372 33704 55412 33832
rect 55372 33655 55412 33664
rect 55276 33570 55316 33655
rect 55468 33536 55508 35503
rect 55564 35216 55604 35225
rect 55564 34544 55604 35176
rect 55852 35057 55892 35671
rect 56140 35561 56180 35848
rect 56236 35888 56276 35897
rect 56139 35552 56181 35561
rect 56139 35512 56140 35552
rect 56180 35512 56181 35552
rect 56139 35503 56181 35512
rect 56043 35216 56085 35225
rect 56043 35176 56044 35216
rect 56084 35176 56085 35216
rect 56043 35167 56085 35176
rect 55851 35048 55893 35057
rect 55851 35008 55852 35048
rect 55892 35008 55893 35048
rect 55851 34999 55893 35008
rect 55852 34628 55892 34999
rect 55564 34495 55604 34504
rect 55660 34588 55892 34628
rect 55372 33496 55508 33536
rect 55179 33452 55221 33461
rect 55179 33412 55180 33452
rect 55220 33412 55221 33452
rect 55179 33403 55221 33412
rect 55372 33140 55412 33496
rect 55660 33140 55700 34588
rect 56044 34385 56084 35167
rect 56139 34880 56181 34889
rect 56139 34840 56140 34880
rect 56180 34840 56181 34880
rect 56139 34831 56181 34840
rect 55852 34376 55892 34385
rect 56043 34376 56085 34385
rect 55892 34336 55988 34376
rect 55852 34327 55892 34336
rect 54892 32815 54932 32824
rect 54988 33100 55412 33140
rect 55564 33100 55700 33140
rect 55852 33536 55892 33545
rect 54796 32730 54836 32815
rect 54988 32612 55028 33100
rect 55084 33032 55124 33041
rect 55124 32992 55316 33032
rect 55084 32983 55124 32992
rect 54796 32572 55028 32612
rect 55084 32864 55124 32873
rect 54699 32360 54741 32369
rect 54412 32320 54644 32360
rect 54412 32192 54452 32201
rect 54412 32117 54452 32152
rect 54507 32192 54549 32201
rect 54507 32152 54508 32192
rect 54548 32152 54549 32192
rect 54507 32143 54549 32152
rect 54411 32108 54453 32117
rect 54411 32068 54412 32108
rect 54452 32068 54453 32108
rect 54411 32059 54453 32068
rect 54412 31949 54452 32059
rect 54508 32058 54548 32143
rect 54411 31940 54453 31949
rect 54411 31900 54412 31940
rect 54452 31900 54453 31940
rect 54411 31891 54453 31900
rect 54604 31856 54644 32320
rect 54699 32320 54700 32360
rect 54740 32320 54741 32360
rect 54699 32311 54741 32320
rect 54508 31816 54644 31856
rect 54700 32192 54740 32201
rect 54508 29924 54548 31816
rect 54604 30680 54644 30689
rect 54700 30680 54740 32152
rect 54796 32192 54836 32572
rect 54891 32276 54933 32285
rect 54891 32236 54892 32276
rect 54932 32236 54933 32276
rect 54891 32227 54933 32236
rect 54796 30857 54836 32152
rect 54892 32192 54932 32227
rect 54892 32141 54932 32152
rect 54987 32192 55029 32201
rect 54987 32152 54988 32192
rect 55028 32152 55029 32192
rect 54987 32143 55029 32152
rect 54988 32058 55028 32143
rect 54987 31940 55029 31949
rect 54987 31900 54988 31940
rect 55028 31900 55029 31940
rect 54987 31891 55029 31900
rect 54795 30848 54837 30857
rect 54795 30808 54796 30848
rect 54836 30808 54837 30848
rect 54795 30799 54837 30808
rect 54644 30640 54740 30680
rect 54795 30680 54837 30689
rect 54795 30640 54796 30680
rect 54836 30640 54837 30680
rect 54604 30631 54644 30640
rect 54795 30631 54837 30640
rect 54892 30680 54932 30689
rect 54796 30546 54836 30631
rect 54603 30512 54645 30521
rect 54603 30472 54604 30512
rect 54644 30472 54645 30512
rect 54603 30463 54645 30472
rect 54604 30378 54644 30463
rect 54699 30260 54741 30269
rect 54699 30220 54700 30260
rect 54740 30220 54741 30260
rect 54699 30211 54741 30220
rect 54508 29875 54548 29884
rect 54700 30008 54740 30211
rect 54892 30092 54932 30640
rect 54988 30269 55028 31891
rect 54987 30260 55029 30269
rect 54987 30220 54988 30260
rect 55028 30220 55029 30260
rect 54987 30211 55029 30220
rect 55084 30185 55124 32824
rect 55276 32864 55316 32992
rect 55276 32815 55316 32824
rect 55371 32276 55413 32285
rect 55371 32236 55372 32276
rect 55412 32236 55413 32276
rect 55371 32227 55413 32236
rect 55275 32192 55317 32201
rect 55275 32152 55276 32192
rect 55316 32152 55317 32192
rect 55275 32143 55317 32152
rect 55276 31604 55316 32143
rect 55276 31555 55316 31564
rect 55372 31436 55412 32227
rect 55180 31396 55412 31436
rect 55180 30848 55220 31396
rect 55564 31352 55604 33100
rect 55660 32864 55700 32873
rect 55852 32864 55892 33496
rect 55700 32824 55892 32864
rect 55660 32815 55700 32824
rect 55659 32192 55701 32201
rect 55659 32152 55660 32192
rect 55700 32152 55701 32192
rect 55659 32143 55701 32152
rect 55852 32192 55892 32201
rect 55660 32058 55700 32143
rect 55756 31940 55796 31949
rect 55660 31352 55700 31361
rect 55564 31312 55660 31352
rect 55756 31352 55796 31900
rect 55852 31520 55892 32152
rect 55948 31781 55988 34336
rect 56043 34336 56044 34376
rect 56084 34336 56085 34376
rect 56043 34327 56085 34336
rect 56140 34376 56180 34831
rect 56236 34460 56276 35848
rect 56332 35888 56372 36427
rect 56332 34637 56372 35848
rect 56428 35216 56468 36679
rect 57099 36476 57141 36485
rect 57099 36436 57100 36476
rect 57140 36436 57141 36476
rect 57099 36427 57141 36436
rect 57100 36342 57140 36427
rect 56524 36016 56852 36056
rect 56524 35888 56564 36016
rect 56524 35839 56564 35848
rect 56619 35888 56661 35897
rect 56619 35848 56620 35888
rect 56660 35848 56661 35888
rect 56619 35839 56661 35848
rect 56716 35888 56756 35897
rect 56620 35754 56660 35839
rect 56716 35216 56756 35848
rect 56331 34628 56373 34637
rect 56331 34588 56332 34628
rect 56372 34588 56373 34628
rect 56331 34579 56373 34588
rect 56236 34420 56372 34460
rect 56140 34327 56180 34336
rect 56235 34292 56277 34301
rect 56235 34252 56236 34292
rect 56276 34252 56277 34292
rect 56235 34243 56277 34252
rect 56236 34158 56276 34243
rect 56332 32285 56372 34420
rect 56428 33140 56468 35176
rect 56524 35176 56756 35216
rect 56524 34628 56564 35176
rect 56524 34579 56564 34588
rect 56428 33100 56564 33140
rect 56524 32864 56564 33100
rect 56564 32824 56660 32864
rect 56524 32815 56564 32824
rect 56331 32276 56373 32285
rect 56331 32236 56332 32276
rect 56372 32236 56373 32276
rect 56331 32227 56373 32236
rect 55947 31772 55989 31781
rect 55947 31732 55948 31772
rect 55988 31732 55989 31772
rect 55947 31723 55989 31732
rect 55852 31480 56084 31520
rect 55852 31352 55892 31361
rect 55756 31312 55852 31352
rect 55275 31184 55317 31193
rect 55275 31144 55276 31184
rect 55316 31144 55317 31184
rect 55275 31135 55317 31144
rect 55563 31184 55605 31193
rect 55563 31144 55564 31184
rect 55604 31144 55605 31184
rect 55563 31135 55605 31144
rect 55276 31050 55316 31135
rect 55180 30808 55316 30848
rect 55180 30680 55220 30689
rect 55180 30437 55220 30640
rect 55179 30428 55221 30437
rect 55179 30388 55180 30428
rect 55220 30388 55221 30428
rect 55179 30379 55221 30388
rect 55083 30176 55125 30185
rect 55083 30136 55084 30176
rect 55124 30136 55125 30176
rect 55083 30127 55125 30136
rect 55276 30092 55316 30808
rect 55564 30764 55604 31135
rect 55564 30715 55604 30724
rect 55468 30680 55508 30689
rect 55468 30353 55508 30640
rect 55467 30344 55509 30353
rect 55467 30304 55468 30344
rect 55508 30304 55509 30344
rect 55660 30344 55700 31312
rect 55755 31184 55797 31193
rect 55755 31144 55756 31184
rect 55796 31144 55797 31184
rect 55755 31135 55797 31144
rect 55756 31050 55796 31135
rect 55852 30689 55892 31312
rect 55948 31352 55988 31361
rect 55948 31025 55988 31312
rect 55947 31016 55989 31025
rect 55947 30976 55948 31016
rect 55988 30976 55989 31016
rect 55947 30967 55989 30976
rect 56044 30848 56084 31480
rect 56620 31361 56660 32824
rect 56812 32201 56852 36016
rect 57099 35972 57141 35981
rect 57099 35932 57100 35972
rect 57140 35932 57141 35972
rect 57099 35923 57141 35932
rect 57100 35838 57140 35923
rect 56908 35720 56948 35729
rect 56908 35561 56948 35680
rect 56907 35552 56949 35561
rect 56907 35512 56908 35552
rect 56948 35512 56949 35552
rect 56907 35503 56949 35512
rect 57196 35225 57236 36688
rect 57292 36679 57332 36688
rect 57387 36728 57429 36737
rect 57387 36688 57388 36728
rect 57428 36688 57429 36728
rect 57387 36679 57429 36688
rect 57484 36728 57524 36737
rect 57291 36560 57333 36569
rect 57291 36520 57292 36560
rect 57332 36520 57333 36560
rect 57291 36511 57333 36520
rect 57292 36426 57332 36511
rect 57195 35216 57237 35225
rect 57195 35176 57196 35216
rect 57236 35176 57237 35216
rect 57195 35167 57237 35176
rect 57484 35141 57524 36688
rect 57580 36728 57620 36763
rect 57580 36678 57620 36688
rect 58348 36644 58388 38116
rect 58539 38156 58581 38165
rect 58539 38116 58540 38156
rect 58580 38116 58581 38156
rect 58539 38107 58581 38116
rect 58924 38156 58964 38165
rect 58540 38072 58580 38107
rect 58540 38021 58580 38032
rect 58924 37997 58964 38116
rect 59307 38156 59349 38165
rect 63340 38156 63380 38189
rect 59307 38116 59308 38156
rect 59348 38116 59349 38156
rect 59307 38107 59349 38116
rect 62668 38116 63380 38156
rect 59308 38022 59348 38107
rect 61612 38072 61652 38081
rect 61516 38032 61612 38072
rect 58732 37988 58772 37997
rect 58923 37988 58965 37997
rect 58772 37948 58868 37988
rect 58732 37939 58772 37948
rect 58828 37568 58868 37948
rect 58923 37948 58924 37988
rect 58964 37948 58965 37988
rect 58923 37939 58965 37948
rect 59115 37988 59157 37997
rect 59115 37948 59116 37988
rect 59156 37948 59157 37988
rect 59115 37939 59157 37948
rect 59116 37854 59156 37939
rect 59788 37568 59828 37577
rect 58828 37528 59060 37568
rect 58828 37400 58868 37409
rect 58635 37316 58677 37325
rect 58635 37276 58636 37316
rect 58676 37276 58677 37316
rect 58635 37267 58677 37276
rect 58636 37182 58676 37267
rect 58828 36905 58868 37360
rect 58924 37400 58964 37409
rect 58924 36989 58964 37360
rect 59020 37400 59060 37528
rect 58923 36980 58965 36989
rect 58923 36940 58924 36980
rect 58964 36940 58965 36980
rect 58923 36931 58965 36940
rect 58827 36896 58869 36905
rect 58827 36856 58828 36896
rect 58868 36856 58869 36896
rect 58827 36847 58869 36856
rect 58443 36812 58485 36821
rect 58443 36772 58444 36812
rect 58484 36772 58485 36812
rect 58443 36763 58485 36772
rect 58444 36678 58484 36763
rect 58540 36728 58580 36737
rect 58827 36728 58869 36737
rect 58580 36688 58676 36728
rect 58540 36679 58580 36688
rect 58060 36604 58388 36644
rect 58060 35636 58100 36604
rect 58156 36476 58196 36485
rect 58196 36436 58580 36476
rect 58156 36427 58196 36436
rect 58540 35888 58580 36436
rect 58636 36065 58676 36688
rect 58827 36688 58828 36728
rect 58868 36688 58869 36728
rect 58827 36679 58869 36688
rect 58828 36594 58868 36679
rect 59020 36233 59060 37360
rect 59116 37400 59156 37409
rect 59308 37400 59348 37409
rect 59156 37360 59308 37400
rect 59116 37351 59156 37360
rect 59308 37351 59348 37360
rect 59499 37400 59541 37409
rect 59499 37360 59500 37400
rect 59540 37360 59541 37400
rect 59499 37351 59541 37360
rect 59596 37400 59636 37411
rect 59403 37316 59445 37325
rect 59403 37276 59404 37316
rect 59444 37276 59445 37316
rect 59403 37267 59445 37276
rect 59307 37232 59349 37241
rect 59307 37192 59308 37232
rect 59348 37192 59349 37232
rect 59307 37183 59349 37192
rect 59116 36728 59156 36737
rect 59019 36224 59061 36233
rect 59019 36184 59020 36224
rect 59060 36184 59061 36224
rect 59019 36175 59061 36184
rect 58635 36056 58677 36065
rect 59116 36056 59156 36688
rect 58635 36016 58636 36056
rect 58676 36016 58677 36056
rect 58635 36007 58677 36016
rect 59020 36016 59156 36056
rect 58540 35839 58580 35848
rect 58635 35888 58677 35897
rect 58635 35848 58636 35888
rect 58676 35848 58677 35888
rect 58635 35839 58677 35848
rect 58732 35888 58772 35897
rect 58636 35754 58676 35839
rect 58251 35720 58293 35729
rect 58251 35680 58252 35720
rect 58292 35680 58293 35720
rect 58251 35671 58293 35680
rect 58060 35596 58196 35636
rect 57771 35216 57813 35225
rect 57771 35176 57772 35216
rect 57812 35176 57813 35216
rect 57771 35167 57813 35176
rect 57964 35216 58004 35227
rect 57483 35132 57525 35141
rect 57483 35092 57484 35132
rect 57524 35092 57525 35132
rect 57483 35083 57525 35092
rect 57772 35082 57812 35167
rect 57964 35141 58004 35176
rect 58060 35216 58100 35225
rect 57963 35132 58005 35141
rect 57963 35092 57964 35132
rect 58004 35092 58005 35132
rect 57963 35083 58005 35092
rect 57580 34964 57620 34975
rect 57772 34964 57812 34973
rect 57580 34889 57620 34924
rect 57676 34924 57772 34964
rect 57579 34880 57621 34889
rect 57579 34840 57580 34880
rect 57620 34840 57621 34880
rect 57579 34831 57621 34840
rect 57676 34628 57716 34924
rect 57772 34915 57812 34924
rect 57484 34588 57716 34628
rect 57484 34376 57524 34588
rect 58060 34553 58100 35176
rect 57772 34544 57812 34553
rect 58059 34544 58101 34553
rect 57812 34504 58004 34544
rect 57772 34495 57812 34504
rect 57484 34327 57524 34336
rect 57580 34376 57620 34385
rect 57580 32873 57620 34336
rect 57772 34376 57812 34385
rect 57772 34049 57812 34336
rect 57964 34376 58004 34504
rect 58059 34504 58060 34544
rect 58100 34504 58101 34544
rect 58059 34495 58101 34504
rect 57964 34327 58004 34336
rect 58059 34376 58101 34385
rect 58059 34336 58060 34376
rect 58100 34336 58101 34376
rect 58059 34327 58101 34336
rect 57771 34040 57813 34049
rect 57771 34000 57772 34040
rect 57812 34000 57813 34040
rect 57771 33991 57813 34000
rect 57579 32864 57621 32873
rect 57579 32824 57580 32864
rect 57620 32824 57621 32864
rect 57579 32815 57621 32824
rect 58060 32864 58100 34327
rect 58156 33125 58196 35596
rect 58252 34385 58292 35671
rect 58444 35048 58484 35057
rect 58251 34376 58293 34385
rect 58251 34336 58252 34376
rect 58292 34336 58293 34376
rect 58251 34327 58293 34336
rect 58348 34376 58388 34385
rect 58444 34376 58484 35008
rect 58732 34637 58772 35848
rect 58924 35888 58964 35897
rect 58924 35729 58964 35848
rect 59020 35804 59060 36016
rect 59115 35888 59157 35897
rect 59115 35848 59116 35888
rect 59156 35848 59157 35888
rect 59115 35839 59157 35848
rect 59212 35888 59252 35899
rect 59308 35897 59348 37183
rect 59404 37182 59444 37267
rect 59500 37266 59540 37351
rect 59596 37325 59636 37360
rect 59595 37316 59637 37325
rect 59595 37276 59596 37316
rect 59636 37276 59637 37316
rect 59595 37267 59637 37276
rect 59788 37148 59828 37528
rect 59500 37108 59828 37148
rect 60172 37400 60212 37409
rect 59500 36728 59540 37108
rect 59500 36679 59540 36688
rect 59499 36224 59541 36233
rect 59499 36184 59500 36224
rect 59540 36184 59541 36224
rect 59499 36175 59541 36184
rect 59500 35981 59540 36175
rect 59595 36056 59637 36065
rect 59595 36016 59596 36056
rect 59636 36016 59637 36056
rect 59595 36007 59637 36016
rect 59499 35972 59541 35981
rect 59499 35932 59500 35972
rect 59540 35932 59541 35972
rect 59499 35923 59541 35932
rect 59020 35755 59060 35764
rect 59116 35754 59156 35839
rect 59212 35813 59252 35848
rect 59307 35888 59349 35897
rect 59307 35848 59308 35888
rect 59348 35848 59349 35888
rect 59307 35839 59349 35848
rect 59404 35888 59444 35897
rect 59211 35804 59253 35813
rect 59211 35764 59212 35804
rect 59252 35764 59253 35804
rect 59211 35755 59253 35764
rect 58923 35720 58965 35729
rect 58923 35680 58924 35720
rect 58964 35680 58965 35720
rect 58923 35671 58965 35680
rect 58827 35132 58869 35141
rect 58827 35092 58828 35132
rect 58868 35092 58869 35132
rect 58827 35083 58869 35092
rect 58731 34628 58773 34637
rect 58731 34588 58732 34628
rect 58772 34588 58773 34628
rect 58731 34579 58773 34588
rect 58388 34336 58484 34376
rect 58348 34327 58388 34336
rect 58635 34208 58677 34217
rect 58635 34168 58636 34208
rect 58676 34168 58677 34208
rect 58635 34159 58677 34168
rect 58347 34040 58389 34049
rect 58347 34000 58348 34040
rect 58388 34000 58389 34040
rect 58347 33991 58389 34000
rect 58348 33872 58388 33991
rect 58443 33956 58485 33965
rect 58443 33916 58444 33956
rect 58484 33916 58485 33956
rect 58443 33907 58485 33916
rect 58348 33823 58388 33832
rect 58444 33704 58484 33907
rect 58539 33788 58581 33797
rect 58539 33748 58540 33788
rect 58580 33748 58581 33788
rect 58539 33739 58581 33748
rect 58444 33655 58484 33664
rect 58540 33704 58580 33739
rect 58540 33653 58580 33664
rect 58636 33704 58676 34159
rect 58347 33452 58389 33461
rect 58347 33412 58348 33452
rect 58388 33412 58389 33452
rect 58347 33403 58389 33412
rect 58155 33116 58197 33125
rect 58155 33076 58156 33116
rect 58196 33076 58197 33116
rect 58155 33067 58197 33076
rect 58252 32873 58292 32958
rect 58060 32815 58100 32824
rect 58251 32864 58293 32873
rect 58251 32824 58252 32864
rect 58292 32824 58293 32864
rect 58251 32815 58293 32824
rect 58348 32864 58388 33403
rect 58636 33140 58676 33664
rect 58828 33704 58868 35083
rect 59404 34796 59444 35848
rect 59596 35888 59636 36007
rect 59499 35804 59541 35813
rect 59499 35764 59500 35804
rect 59540 35764 59541 35804
rect 59499 35755 59541 35764
rect 59500 35670 59540 35755
rect 59596 35729 59636 35848
rect 59595 35720 59637 35729
rect 59595 35680 59596 35720
rect 59636 35680 59637 35720
rect 59595 35671 59637 35680
rect 59884 35216 59924 35225
rect 59788 35176 59884 35216
rect 59404 34756 59540 34796
rect 59403 34628 59445 34637
rect 59403 34588 59404 34628
rect 59444 34588 59445 34628
rect 59403 34579 59445 34588
rect 59212 34376 59252 34385
rect 59252 34336 59348 34376
rect 59212 34327 59252 34336
rect 58828 33655 58868 33664
rect 59020 33704 59060 33713
rect 58924 33461 58964 33546
rect 58923 33452 58965 33461
rect 58923 33412 58924 33452
rect 58964 33412 58965 33452
rect 58923 33403 58965 33412
rect 58923 33284 58965 33293
rect 58923 33244 58924 33284
rect 58964 33244 58965 33284
rect 58923 33235 58965 33244
rect 58636 33100 58772 33140
rect 58635 33032 58677 33041
rect 58635 32992 58636 33032
rect 58676 32992 58677 33032
rect 58635 32983 58677 32992
rect 58348 32815 58388 32824
rect 58155 32780 58197 32789
rect 58155 32740 58156 32780
rect 58196 32740 58197 32780
rect 58155 32731 58197 32740
rect 57675 32696 57717 32705
rect 57675 32656 57676 32696
rect 57716 32656 57717 32696
rect 57675 32647 57717 32656
rect 56811 32192 56853 32201
rect 56811 32152 56812 32192
rect 56852 32152 56853 32192
rect 56811 32143 56853 32152
rect 57195 31604 57237 31613
rect 57195 31564 57196 31604
rect 57236 31564 57237 31604
rect 57195 31555 57237 31564
rect 56524 31352 56564 31361
rect 56140 31268 56180 31279
rect 56140 31193 56180 31228
rect 56139 31184 56181 31193
rect 56139 31144 56140 31184
rect 56180 31144 56181 31184
rect 56139 31135 56181 31144
rect 56139 31016 56181 31025
rect 56139 30976 56140 31016
rect 56180 30976 56181 31016
rect 56139 30967 56181 30976
rect 55948 30808 56084 30848
rect 55851 30680 55893 30689
rect 55851 30640 55852 30680
rect 55892 30640 55893 30680
rect 55851 30631 55893 30640
rect 55852 30512 55892 30521
rect 55948 30512 55988 30808
rect 56140 30764 56180 30967
rect 56140 30715 56180 30724
rect 56236 30680 56276 30689
rect 55892 30472 55988 30512
rect 56044 30657 56084 30666
rect 55852 30463 55892 30472
rect 55660 30304 55892 30344
rect 55467 30295 55509 30304
rect 55468 30136 55796 30176
rect 55468 30092 55508 30136
rect 55276 30052 55508 30092
rect 54892 30043 54932 30052
rect 55563 30008 55605 30017
rect 54700 29849 54740 29968
rect 54988 29968 55564 30008
rect 55604 29968 55605 30008
rect 54795 29924 54837 29933
rect 54795 29884 54796 29924
rect 54836 29884 54932 29924
rect 54795 29875 54837 29884
rect 54699 29840 54741 29849
rect 54699 29800 54700 29840
rect 54740 29800 54741 29840
rect 54699 29791 54741 29800
rect 54892 29840 54932 29884
rect 54892 29791 54932 29800
rect 54988 29672 55028 29968
rect 55563 29959 55605 29968
rect 55564 29874 55604 29959
rect 55083 29840 55125 29849
rect 55083 29800 55084 29840
rect 55124 29800 55125 29840
rect 55083 29791 55125 29800
rect 55180 29840 55220 29849
rect 55468 29840 55508 29849
rect 55220 29800 55412 29840
rect 55180 29791 55220 29800
rect 55084 29706 55124 29791
rect 54892 29632 55028 29672
rect 54027 29252 54069 29261
rect 54027 29212 54028 29252
rect 54068 29212 54069 29252
rect 54027 29203 54069 29212
rect 54315 29252 54357 29261
rect 54315 29212 54316 29252
rect 54356 29212 54357 29252
rect 54315 29203 54357 29212
rect 53931 29000 53973 29009
rect 53931 28960 53932 29000
rect 53972 28960 53973 29000
rect 53931 28951 53973 28960
rect 53452 26935 53492 26944
rect 53259 26900 53301 26909
rect 53259 26860 53260 26900
rect 53300 26860 53301 26900
rect 53259 26851 53301 26860
rect 53260 26741 53300 26851
rect 53259 26732 53301 26741
rect 53259 26692 53260 26732
rect 53300 26692 53301 26732
rect 53259 26683 53301 26692
rect 53548 25304 53588 25313
rect 53548 24641 53588 25264
rect 53547 24632 53589 24641
rect 53068 24592 53204 24632
rect 52875 24583 52917 24592
rect 52683 24044 52725 24053
rect 52683 24004 52684 24044
rect 52724 24004 52725 24044
rect 52683 23995 52725 24004
rect 52587 23792 52629 23801
rect 52587 23752 52588 23792
rect 52628 23752 52629 23792
rect 52876 23792 52916 24583
rect 52972 23792 53012 23801
rect 52876 23752 52972 23792
rect 52587 23743 52629 23752
rect 52779 23288 52821 23297
rect 52779 23248 52780 23288
rect 52820 23248 52821 23288
rect 52779 23239 52821 23248
rect 52491 23120 52533 23129
rect 52683 23120 52725 23129
rect 52491 23080 52492 23120
rect 52532 23080 52533 23120
rect 52491 23071 52533 23080
rect 52588 23080 52684 23120
rect 52724 23080 52725 23120
rect 52203 23036 52245 23045
rect 52203 22996 52204 23036
rect 52244 22996 52245 23036
rect 52203 22987 52245 22996
rect 52012 22324 52148 22364
rect 52012 22028 52052 22324
rect 52204 22280 52244 22987
rect 52299 22952 52341 22961
rect 52299 22912 52300 22952
rect 52340 22912 52341 22952
rect 52299 22903 52341 22912
rect 52300 22818 52340 22903
rect 52395 22784 52437 22793
rect 52395 22744 52396 22784
rect 52436 22744 52437 22784
rect 52395 22735 52437 22744
rect 52396 22532 52436 22735
rect 52396 22483 52436 22492
rect 52588 22448 52628 23080
rect 52683 23071 52725 23080
rect 52683 22868 52725 22877
rect 52683 22828 52684 22868
rect 52724 22828 52725 22868
rect 52683 22819 52725 22828
rect 52492 22408 52628 22448
rect 52684 22532 52724 22819
rect 52300 22280 52340 22289
rect 52108 22269 52148 22278
rect 52204 22240 52300 22280
rect 52108 22205 52148 22229
rect 52107 22196 52149 22205
rect 52107 22156 52108 22196
rect 52148 22156 52149 22196
rect 52107 22147 52149 22156
rect 52108 22134 52148 22147
rect 52300 22037 52340 22240
rect 52299 22028 52341 22037
rect 52012 21988 52148 22028
rect 51915 21020 51957 21029
rect 51915 20980 51916 21020
rect 51956 20980 51957 21020
rect 51915 20971 51957 20980
rect 51572 20728 51668 20768
rect 50284 20719 50324 20728
rect 50668 20719 50708 20728
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 51532 20189 51572 20728
rect 51627 20516 51669 20525
rect 51627 20476 51628 20516
rect 51668 20476 51669 20516
rect 51627 20467 51669 20476
rect 47211 20180 47253 20189
rect 47211 20140 47212 20180
rect 47252 20140 47253 20180
rect 47211 20131 47253 20140
rect 47595 20180 47637 20189
rect 47595 20140 47596 20180
rect 47636 20140 47637 20180
rect 47595 20131 47637 20140
rect 48939 20180 48981 20189
rect 48939 20140 48940 20180
rect 48980 20140 48981 20180
rect 48939 20131 48981 20140
rect 50859 20180 50901 20189
rect 50859 20140 50860 20180
rect 50900 20140 50901 20180
rect 50859 20131 50901 20140
rect 51531 20180 51573 20189
rect 51531 20140 51532 20180
rect 51572 20140 51573 20180
rect 51531 20131 51573 20140
rect 47500 20012 47540 20021
rect 47308 19844 47348 19853
rect 47308 18752 47348 19804
rect 47500 19433 47540 19972
rect 47499 19424 47541 19433
rect 47499 19384 47500 19424
rect 47540 19384 47541 19424
rect 47499 19375 47541 19384
rect 47500 19256 47540 19265
rect 47596 19256 47636 20131
rect 49132 20096 49172 20105
rect 49036 20056 49132 20096
rect 47884 20012 47924 20021
rect 47692 19844 47732 19853
rect 47732 19804 47828 19844
rect 47692 19795 47732 19804
rect 47540 19216 47636 19256
rect 47500 19207 47540 19216
rect 47308 18712 47636 18752
rect 47020 18584 47060 18593
rect 47404 18584 47444 18593
rect 47060 18544 47404 18584
rect 47020 18535 47060 18544
rect 47404 18535 47444 18544
rect 47500 18584 47540 18595
rect 47500 18509 47540 18544
rect 47596 18584 47636 18712
rect 47499 18500 47541 18509
rect 47499 18460 47500 18500
rect 47540 18460 47541 18500
rect 47499 18451 47541 18460
rect 47019 18416 47061 18425
rect 47019 18376 47020 18416
rect 47060 18376 47061 18416
rect 47019 18367 47061 18376
rect 47020 18282 47060 18367
rect 47500 17501 47540 18451
rect 47499 17492 47541 17501
rect 47499 17452 47500 17492
rect 47540 17452 47541 17492
rect 47499 17443 47541 17452
rect 47596 17417 47636 18544
rect 47691 18584 47733 18593
rect 47691 18544 47692 18584
rect 47732 18544 47733 18584
rect 47691 18535 47733 18544
rect 47692 18450 47732 18535
rect 47788 18509 47828 19804
rect 47787 18500 47829 18509
rect 47787 18460 47788 18500
rect 47828 18460 47829 18500
rect 47787 18451 47829 18460
rect 47595 17408 47637 17417
rect 47595 17368 47596 17408
rect 47636 17368 47637 17408
rect 47595 17359 47637 17368
rect 47499 17240 47541 17249
rect 47499 17200 47500 17240
rect 47540 17200 47541 17240
rect 47499 17191 47541 17200
rect 47019 17072 47061 17081
rect 47019 17032 47020 17072
rect 47060 17032 47061 17072
rect 47019 17023 47061 17032
rect 47500 17072 47540 17191
rect 47020 14720 47060 17023
rect 47307 16904 47349 16913
rect 47307 16864 47308 16904
rect 47348 16864 47349 16904
rect 47307 16855 47349 16864
rect 47115 16820 47157 16829
rect 47115 16780 47116 16820
rect 47156 16780 47157 16820
rect 47115 16771 47157 16780
rect 47116 16232 47156 16771
rect 47116 16183 47156 16192
rect 47211 16232 47253 16241
rect 47211 16192 47212 16232
rect 47252 16192 47253 16232
rect 47211 16183 47253 16192
rect 47308 16232 47348 16855
rect 47403 16316 47445 16325
rect 47403 16276 47404 16316
rect 47444 16276 47445 16316
rect 47403 16267 47445 16276
rect 47212 16098 47252 16183
rect 47308 15905 47348 16192
rect 47307 15896 47349 15905
rect 47307 15856 47308 15896
rect 47348 15856 47349 15896
rect 47307 15847 47349 15856
rect 47404 15392 47444 16267
rect 47500 16241 47540 17032
rect 47884 16577 47924 19972
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 48939 19676 48981 19685
rect 48939 19636 48940 19676
rect 48980 19636 48981 19676
rect 48939 19627 48981 19636
rect 48940 19508 48980 19627
rect 48940 19459 48980 19468
rect 49036 19265 49076 20056
rect 49132 20047 49172 20056
rect 49324 20096 49364 20105
rect 49228 19844 49268 19853
rect 48940 19256 48980 19265
rect 48268 19216 48940 19256
rect 47883 16568 47925 16577
rect 47883 16528 47884 16568
rect 47924 16528 47925 16568
rect 47883 16519 47925 16528
rect 48268 16325 48308 19216
rect 48940 19207 48980 19216
rect 49035 19256 49077 19265
rect 49035 19216 49036 19256
rect 49076 19216 49077 19256
rect 49035 19207 49077 19216
rect 49132 19256 49172 19265
rect 48652 19088 48692 19097
rect 48692 19048 48884 19088
rect 48652 19039 48692 19048
rect 48651 18752 48693 18761
rect 48651 18712 48652 18752
rect 48692 18712 48693 18752
rect 48651 18703 48693 18712
rect 48364 18584 48404 18593
rect 48364 17081 48404 18544
rect 48652 18584 48692 18703
rect 48844 18593 48884 19048
rect 49035 18920 49077 18929
rect 49035 18880 49036 18920
rect 49076 18880 49077 18920
rect 49035 18871 49077 18880
rect 49036 18761 49076 18871
rect 49035 18752 49077 18761
rect 49035 18712 49036 18752
rect 49076 18712 49077 18752
rect 49035 18703 49077 18712
rect 49132 18677 49172 19216
rect 49228 19256 49268 19804
rect 49228 19207 49268 19216
rect 49227 18920 49269 18929
rect 49227 18880 49228 18920
rect 49268 18880 49269 18920
rect 49324 18920 49364 20056
rect 50092 19928 50132 19937
rect 49611 19676 49653 19685
rect 49611 19636 49612 19676
rect 49652 19636 49653 19676
rect 49611 19627 49653 19636
rect 49612 19256 49652 19627
rect 49612 19207 49652 19216
rect 49996 19256 50036 19265
rect 50092 19256 50132 19888
rect 50036 19216 50132 19256
rect 50860 19256 50900 20131
rect 51531 19592 51573 19601
rect 51531 19552 51532 19592
rect 51572 19552 51573 19592
rect 51531 19543 51573 19552
rect 49996 19207 50036 19216
rect 50860 19207 50900 19216
rect 49611 18920 49653 18929
rect 49324 18880 49556 18920
rect 49227 18871 49269 18880
rect 49131 18668 49173 18677
rect 49131 18628 49132 18668
rect 49172 18628 49173 18668
rect 49131 18619 49173 18628
rect 49228 18605 49268 18871
rect 49324 18677 49364 18762
rect 49323 18668 49365 18677
rect 49323 18628 49324 18668
rect 49364 18628 49365 18668
rect 49323 18619 49365 18628
rect 48652 18535 48692 18544
rect 48748 18584 48788 18593
rect 48843 18584 48885 18593
rect 48788 18544 48844 18584
rect 48884 18544 48980 18584
rect 49228 18556 49268 18565
rect 49420 18584 49460 18593
rect 48748 18535 48788 18544
rect 48843 18535 48885 18544
rect 48844 18450 48884 18535
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 48940 17996 48980 18544
rect 49420 18500 49460 18544
rect 49261 18460 49460 18500
rect 49036 18416 49076 18425
rect 49261 18416 49301 18460
rect 49076 18376 49301 18416
rect 49036 18367 49076 18376
rect 49516 18089 49556 18880
rect 49611 18880 49612 18920
rect 49652 18880 49653 18920
rect 49611 18871 49653 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 49612 18500 49652 18871
rect 51532 18509 51572 19543
rect 49803 18500 49845 18509
rect 49612 18460 49804 18500
rect 49844 18460 49845 18500
rect 49803 18451 49845 18460
rect 50476 18500 50516 18509
rect 49804 18366 49844 18451
rect 50476 18341 50516 18460
rect 50571 18500 50613 18509
rect 51340 18500 51380 18509
rect 50571 18460 50572 18500
rect 50612 18460 50613 18500
rect 50571 18451 50613 18460
rect 51244 18460 51340 18500
rect 49996 18332 50036 18341
rect 49515 18080 49557 18089
rect 49515 18040 49516 18080
rect 49556 18040 49557 18080
rect 49515 18031 49557 18040
rect 48652 17956 48980 17996
rect 48652 17744 48692 17956
rect 48939 17828 48981 17837
rect 48939 17788 48940 17828
rect 48980 17788 48981 17828
rect 48939 17779 48981 17788
rect 49515 17828 49557 17837
rect 49515 17788 49516 17828
rect 49556 17788 49557 17828
rect 49515 17779 49557 17788
rect 48652 17695 48692 17704
rect 48747 17744 48789 17753
rect 48747 17704 48748 17744
rect 48788 17704 48789 17744
rect 48747 17695 48789 17704
rect 48940 17744 48980 17779
rect 48748 17610 48788 17695
rect 48940 17693 48980 17704
rect 49420 17744 49460 17753
rect 48844 17576 48884 17585
rect 48884 17536 48980 17576
rect 48844 17527 48884 17536
rect 48363 17072 48405 17081
rect 48363 17032 48364 17072
rect 48404 17032 48405 17072
rect 48940 17072 48980 17536
rect 49420 17333 49460 17704
rect 49516 17694 49556 17779
rect 49612 17753 49652 17838
rect 49803 17828 49845 17837
rect 49803 17788 49804 17828
rect 49844 17788 49845 17828
rect 49803 17779 49845 17788
rect 49611 17744 49653 17753
rect 49611 17704 49612 17744
rect 49652 17704 49653 17744
rect 49611 17695 49653 17704
rect 49804 17744 49844 17779
rect 49804 17693 49844 17704
rect 49900 17744 49940 17753
rect 49900 17576 49940 17704
rect 49612 17536 49940 17576
rect 49996 17576 50036 18292
rect 50284 18332 50324 18341
rect 50475 18332 50517 18341
rect 50324 18292 50420 18332
rect 50284 18283 50324 18292
rect 50092 17996 50132 18005
rect 50132 17956 50324 17996
rect 50092 17947 50132 17956
rect 50092 17753 50132 17838
rect 50091 17744 50133 17753
rect 50091 17704 50092 17744
rect 50132 17704 50133 17744
rect 50091 17695 50133 17704
rect 50284 17744 50324 17956
rect 50380 17753 50420 18292
rect 50475 18292 50476 18332
rect 50516 18292 50517 18332
rect 50475 18283 50517 18292
rect 50284 17695 50324 17704
rect 50379 17744 50421 17753
rect 50379 17704 50380 17744
rect 50420 17704 50421 17744
rect 50379 17695 50421 17704
rect 50476 17585 50516 18283
rect 50475 17576 50517 17585
rect 49996 17536 50228 17576
rect 49419 17324 49461 17333
rect 49419 17284 49420 17324
rect 49460 17284 49461 17324
rect 49419 17275 49461 17284
rect 49612 17249 49652 17536
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 49611 17240 49653 17249
rect 49611 17200 49612 17240
rect 49652 17200 49653 17240
rect 49611 17191 49653 17200
rect 49227 17156 49269 17165
rect 49227 17116 49228 17156
rect 49268 17116 49269 17156
rect 49227 17107 49269 17116
rect 49132 17072 49172 17081
rect 48940 17032 49132 17072
rect 48363 17023 48405 17032
rect 49132 17023 49172 17032
rect 49228 17072 49268 17107
rect 49228 17021 49268 17032
rect 49420 17072 49460 17081
rect 49708 17072 49748 17081
rect 49460 17032 49708 17072
rect 49420 17023 49460 17032
rect 49708 17023 49748 17032
rect 49804 17072 49844 17081
rect 48651 16988 48693 16997
rect 48651 16948 48652 16988
rect 48692 16948 48693 16988
rect 48651 16939 48693 16948
rect 48652 16854 48692 16939
rect 49420 16820 49460 16829
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 49420 16325 49460 16780
rect 49611 16568 49653 16577
rect 49611 16528 49612 16568
rect 49652 16528 49653 16568
rect 49611 16519 49653 16528
rect 48267 16316 48309 16325
rect 48267 16276 48268 16316
rect 48308 16276 48309 16316
rect 48267 16267 48309 16276
rect 48651 16316 48693 16325
rect 48651 16276 48652 16316
rect 48692 16276 48693 16316
rect 48651 16267 48693 16276
rect 49419 16316 49461 16325
rect 49419 16276 49420 16316
rect 49460 16276 49461 16316
rect 49419 16267 49461 16276
rect 47499 16232 47541 16241
rect 47499 16192 47500 16232
rect 47540 16192 47541 16232
rect 47499 16183 47541 16192
rect 48652 16232 48692 16267
rect 48652 16181 48692 16192
rect 49036 16232 49076 16241
rect 47499 15896 47541 15905
rect 47499 15856 47500 15896
rect 47540 15856 47541 15896
rect 47499 15847 47541 15856
rect 48267 15896 48309 15905
rect 48267 15856 48268 15896
rect 48308 15856 48309 15896
rect 48267 15847 48309 15856
rect 47500 15560 47540 15847
rect 47500 15511 47540 15520
rect 47692 15560 47732 15569
rect 47404 15352 47540 15392
rect 47307 15056 47349 15065
rect 47307 15016 47308 15056
rect 47348 15016 47349 15056
rect 47307 15007 47349 15016
rect 47020 14468 47060 14680
rect 47308 14720 47348 15007
rect 47308 14671 47348 14680
rect 47404 14636 47444 14645
rect 47020 14428 47156 14468
rect 46923 14300 46965 14309
rect 46923 14260 46924 14300
rect 46964 14260 46965 14300
rect 46923 14251 46965 14260
rect 45963 14216 46005 14225
rect 45963 14176 45964 14216
rect 46004 14176 46005 14216
rect 45963 14167 46005 14176
rect 45868 14048 45908 14057
rect 45868 13385 45908 14008
rect 45867 13376 45909 13385
rect 45867 13336 45868 13376
rect 45908 13336 45909 13376
rect 45867 13327 45909 13336
rect 45676 13074 45716 13159
rect 45772 13049 45812 13168
rect 45868 13208 45908 13217
rect 45771 13040 45813 13049
rect 45771 13000 45772 13040
rect 45812 13000 45813 13040
rect 45771 12991 45813 13000
rect 45868 12965 45908 13168
rect 45964 13208 46004 14167
rect 46155 14048 46197 14057
rect 46155 14008 46156 14048
rect 46196 14008 46197 14048
rect 46155 13999 46197 14008
rect 46347 14048 46389 14057
rect 46347 14008 46348 14048
rect 46388 14008 46389 14048
rect 46347 13999 46389 14008
rect 46156 13460 46196 13999
rect 46156 13411 46196 13420
rect 45964 13159 46004 13168
rect 46155 13208 46197 13217
rect 46155 13168 46156 13208
rect 46196 13168 46197 13208
rect 46155 13159 46197 13168
rect 46348 13208 46388 13999
rect 46539 13292 46581 13301
rect 46539 13252 46540 13292
rect 46580 13252 46581 13292
rect 46539 13243 46581 13252
rect 46348 13159 46388 13168
rect 46444 13208 46484 13219
rect 46156 13074 46196 13159
rect 46444 13133 46484 13168
rect 46443 13124 46485 13133
rect 46443 13084 46444 13124
rect 46484 13084 46485 13124
rect 46443 13075 46485 13084
rect 45867 12956 45909 12965
rect 45867 12916 45868 12956
rect 45908 12916 45909 12956
rect 45867 12907 45909 12916
rect 45676 12536 45716 12545
rect 45676 11864 45716 12496
rect 45772 11864 45812 11873
rect 45676 11824 45772 11864
rect 45772 11815 45812 11824
rect 45868 11705 45908 12907
rect 46540 12536 46580 13243
rect 46540 12487 46580 12496
rect 46828 13208 46868 13217
rect 46828 12980 46868 13168
rect 46924 12980 46964 14251
rect 47019 14216 47061 14225
rect 47019 14176 47020 14216
rect 47060 14176 47061 14216
rect 47019 14167 47061 14176
rect 47020 14082 47060 14167
rect 46828 12940 46964 12980
rect 47116 12980 47156 14428
rect 47404 14225 47444 14596
rect 47403 14216 47445 14225
rect 47403 14176 47404 14216
rect 47444 14176 47445 14216
rect 47403 14167 47445 14176
rect 47212 14048 47252 14057
rect 47500 14048 47540 15352
rect 47596 15308 47636 15317
rect 47596 14300 47636 15268
rect 47692 14972 47732 15520
rect 47883 15560 47925 15569
rect 47883 15520 47884 15560
rect 47924 15520 47925 15560
rect 47883 15511 47925 15520
rect 48076 15560 48116 15569
rect 47884 15426 47924 15511
rect 47980 15308 48020 15317
rect 47692 14923 47732 14932
rect 47884 15268 47980 15308
rect 47596 14260 47828 14300
rect 47692 14132 47732 14141
rect 47596 14048 47636 14057
rect 47500 14008 47596 14048
rect 47212 13460 47252 14008
rect 47596 13469 47636 14008
rect 47692 13922 47732 14092
rect 47788 14057 47828 14260
rect 47787 14048 47829 14057
rect 47787 14008 47788 14048
rect 47828 14008 47829 14048
rect 47787 13999 47829 14008
rect 47884 14048 47924 15268
rect 47980 15259 48020 15268
rect 48076 15065 48116 15520
rect 48171 15560 48213 15569
rect 48171 15520 48172 15560
rect 48212 15520 48213 15560
rect 48171 15511 48213 15520
rect 48075 15056 48117 15065
rect 48075 15016 48076 15056
rect 48116 15016 48117 15056
rect 48075 15007 48117 15016
rect 48172 14888 48212 15511
rect 48076 14848 48212 14888
rect 48076 14729 48116 14848
rect 48075 14720 48117 14729
rect 48075 14680 48076 14720
rect 48116 14680 48117 14720
rect 48075 14671 48117 14680
rect 47884 13999 47924 14008
rect 47980 14636 48020 14645
rect 47980 13922 48020 14596
rect 47692 13882 48020 13922
rect 47212 13411 47252 13420
rect 47595 13460 47637 13469
rect 47595 13420 47596 13460
rect 47636 13420 47637 13460
rect 47595 13411 47637 13420
rect 47404 13376 47444 13387
rect 47404 13301 47444 13336
rect 47403 13292 47445 13301
rect 47403 13252 47404 13292
rect 47444 13252 47445 13292
rect 47403 13243 47445 13252
rect 48076 13217 48116 14671
rect 47884 13208 47924 13217
rect 47788 13168 47884 13208
rect 47116 12940 47636 12980
rect 45867 11696 45909 11705
rect 45867 11656 45868 11696
rect 45908 11656 45909 11696
rect 45867 11647 45909 11656
rect 46732 11192 46772 11203
rect 46828 11201 46868 12940
rect 47499 12788 47541 12797
rect 47499 12748 47500 12788
rect 47540 12748 47541 12788
rect 47499 12739 47541 12748
rect 46732 11117 46772 11152
rect 46827 11192 46869 11201
rect 46827 11152 46828 11192
rect 46868 11152 46869 11192
rect 46827 11143 46869 11152
rect 46731 11108 46773 11117
rect 46731 11068 46732 11108
rect 46772 11068 46773 11108
rect 46731 11059 46773 11068
rect 44716 10975 44756 10984
rect 45580 10975 45620 10984
rect 46251 10940 46293 10949
rect 46251 10900 46252 10940
rect 46292 10900 46293 10940
rect 46251 10891 46293 10900
rect 44812 10436 44852 10445
rect 44620 10396 44812 10436
rect 44812 10387 44852 10396
rect 44524 10135 44564 10144
rect 44620 10184 44660 10193
rect 44620 9596 44660 10144
rect 44811 10184 44853 10193
rect 44811 10144 44812 10184
rect 44852 10144 44853 10184
rect 44811 10135 44853 10144
rect 44812 10050 44852 10135
rect 44524 9556 44660 9596
rect 44524 9269 44564 9556
rect 45483 9512 45525 9521
rect 45483 9472 45484 9512
rect 45524 9472 45525 9512
rect 45483 9463 45525 9472
rect 44620 9344 44660 9353
rect 44523 9260 44565 9269
rect 44523 9220 44524 9260
rect 44564 9220 44565 9260
rect 44523 9211 44565 9220
rect 44524 8672 44564 8681
rect 44620 8672 44660 9304
rect 44564 8632 44660 8672
rect 45387 8672 45429 8681
rect 45387 8632 45388 8672
rect 45428 8632 45429 8672
rect 44524 8623 44564 8632
rect 45387 8623 45429 8632
rect 44811 8588 44853 8597
rect 44811 8548 44812 8588
rect 44852 8548 44853 8588
rect 44811 8539 44853 8548
rect 44427 8084 44469 8093
rect 44427 8044 44428 8084
rect 44468 8044 44469 8084
rect 44427 8035 44469 8044
rect 44276 7960 44372 8000
rect 44428 8000 44468 8035
rect 44236 7951 44276 7960
rect 44428 7949 44468 7960
rect 44716 8000 44756 8009
rect 44428 7832 44468 7841
rect 44716 7832 44756 7960
rect 44812 8000 44852 8539
rect 45388 8538 45428 8623
rect 44907 8168 44949 8177
rect 44907 8128 44908 8168
rect 44948 8128 44949 8168
rect 44907 8119 44949 8128
rect 44908 8034 44948 8119
rect 44812 7951 44852 7960
rect 45004 8000 45044 8009
rect 45388 8000 45428 8009
rect 45044 7960 45388 8000
rect 45004 7951 45044 7960
rect 45388 7951 45428 7960
rect 45484 8000 45524 9463
rect 45579 9344 45621 9353
rect 45579 9304 45580 9344
rect 45620 9304 45621 9344
rect 45579 9295 45621 9304
rect 44468 7792 44756 7832
rect 44428 7783 44468 7792
rect 45387 7748 45429 7757
rect 45387 7708 45388 7748
rect 45428 7708 45429 7748
rect 45387 7699 45429 7708
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 45388 7160 45428 7699
rect 45388 7111 45428 7120
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 45484 6413 45524 7960
rect 45580 8000 45620 9295
rect 46252 8177 46292 10891
rect 46828 10697 46868 11143
rect 46924 11024 46964 11035
rect 46924 10949 46964 10984
rect 47116 11024 47156 11033
rect 46923 10940 46965 10949
rect 46923 10900 46924 10940
rect 46964 10900 46965 10940
rect 46923 10891 46965 10900
rect 47020 10772 47060 10781
rect 46827 10688 46869 10697
rect 46827 10648 46828 10688
rect 46868 10648 46869 10688
rect 46827 10639 46869 10648
rect 46444 10312 46868 10352
rect 46347 10184 46389 10193
rect 46347 10144 46348 10184
rect 46388 10144 46389 10184
rect 46347 10135 46389 10144
rect 46348 10050 46388 10135
rect 46444 10100 46484 10312
rect 46444 10051 46484 10060
rect 46540 10184 46580 10193
rect 46540 9680 46580 10144
rect 46636 10184 46676 10193
rect 46828 10184 46868 10312
rect 46676 10144 46772 10184
rect 46636 10135 46676 10144
rect 46732 10016 46772 10144
rect 46828 10135 46868 10144
rect 47020 10100 47060 10732
rect 47116 10529 47156 10984
rect 47115 10520 47157 10529
rect 47115 10480 47116 10520
rect 47156 10480 47157 10520
rect 47115 10471 47157 10480
rect 46924 10060 47060 10100
rect 46924 10016 46964 10060
rect 46732 9976 46964 10016
rect 46540 9640 46868 9680
rect 46636 9512 46676 9521
rect 46347 9260 46389 9269
rect 46347 9220 46348 9260
rect 46388 9220 46389 9260
rect 46347 9211 46389 9220
rect 46348 9126 46388 9211
rect 46540 8924 46580 8933
rect 46636 8924 46676 9472
rect 46731 9512 46773 9521
rect 46731 9472 46732 9512
rect 46772 9472 46773 9512
rect 46731 9463 46773 9472
rect 46732 9378 46772 9463
rect 46731 9260 46773 9269
rect 46731 9220 46732 9260
rect 46772 9220 46773 9260
rect 46731 9211 46773 9220
rect 46580 8884 46676 8924
rect 46540 8875 46580 8884
rect 46635 8672 46677 8681
rect 46635 8632 46636 8672
rect 46676 8632 46677 8672
rect 46635 8623 46677 8632
rect 46732 8672 46772 9211
rect 46732 8623 46772 8632
rect 46540 8504 46580 8513
rect 46251 8168 46293 8177
rect 46251 8128 46252 8168
rect 46292 8128 46293 8168
rect 46251 8119 46293 8128
rect 46540 8009 46580 8464
rect 45580 6497 45620 7960
rect 45675 8000 45717 8009
rect 45675 7960 45676 8000
rect 45716 7960 45717 8000
rect 45675 7951 45717 7960
rect 46539 8000 46581 8009
rect 46539 7960 46540 8000
rect 46580 7960 46581 8000
rect 46539 7951 46581 7960
rect 45676 7866 45716 7951
rect 45964 7832 46004 7841
rect 45772 7160 45812 7169
rect 45964 7160 46004 7792
rect 46636 7169 46676 8623
rect 46828 8597 46868 9640
rect 47020 9512 47060 9523
rect 47116 9521 47156 10471
rect 47212 10184 47252 10193
rect 47252 10144 47348 10184
rect 47212 10135 47252 10144
rect 47020 9437 47060 9472
rect 47115 9512 47157 9521
rect 47115 9472 47116 9512
rect 47156 9472 47157 9512
rect 47115 9463 47157 9472
rect 47019 9428 47061 9437
rect 47019 9388 47020 9428
rect 47060 9388 47061 9428
rect 47019 9379 47061 9388
rect 47308 9344 47348 10144
rect 47308 9295 47348 9304
rect 46923 8756 46965 8765
rect 46923 8716 46924 8756
rect 46964 8716 46965 8756
rect 46923 8707 46965 8716
rect 46924 8672 46964 8707
rect 46924 8621 46964 8632
rect 46827 8588 46869 8597
rect 46827 8548 46828 8588
rect 46868 8548 46869 8588
rect 46827 8539 46869 8548
rect 46828 8454 46868 8539
rect 47500 8177 47540 12739
rect 47596 12536 47636 12940
rect 47692 12713 47732 12798
rect 47788 12797 47828 13168
rect 47884 13159 47924 13168
rect 48075 13208 48117 13217
rect 48075 13168 48076 13208
rect 48116 13168 48117 13208
rect 48075 13159 48117 13168
rect 48172 13208 48212 13217
rect 48268 13208 48308 15847
rect 48460 15392 48500 15401
rect 48364 15352 48460 15392
rect 49036 15392 49076 16192
rect 49612 15476 49652 16519
rect 49804 16400 49844 17032
rect 49900 17072 49940 17081
rect 49900 16913 49940 17032
rect 49995 17072 50037 17081
rect 49995 17032 49996 17072
rect 50036 17032 50037 17072
rect 49995 17023 50037 17032
rect 49996 16938 50036 17023
rect 50188 16913 50228 17536
rect 50475 17536 50476 17576
rect 50516 17536 50517 17576
rect 50475 17527 50517 17536
rect 50379 17240 50421 17249
rect 50379 17200 50380 17240
rect 50420 17200 50421 17240
rect 50379 17191 50421 17200
rect 50380 17072 50420 17191
rect 50380 17023 50420 17032
rect 49899 16904 49941 16913
rect 49899 16864 49900 16904
rect 49940 16864 49941 16904
rect 49899 16855 49941 16864
rect 50187 16904 50229 16913
rect 50187 16864 50188 16904
rect 50228 16864 50229 16904
rect 50187 16855 50229 16864
rect 50475 16820 50517 16829
rect 50475 16780 50476 16820
rect 50516 16780 50517 16820
rect 50475 16771 50517 16780
rect 49804 16360 50228 16400
rect 49899 16232 49941 16241
rect 49899 16192 49900 16232
rect 49940 16192 49941 16232
rect 49899 16183 49941 16192
rect 49900 16098 49940 16183
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 50188 15728 50228 16360
rect 50188 15679 50228 15688
rect 49996 15476 50036 15485
rect 50379 15476 50421 15485
rect 49612 15436 49996 15476
rect 49996 15427 50036 15436
rect 50284 15436 50380 15476
rect 50420 15436 50421 15476
rect 49132 15392 49172 15401
rect 49036 15352 49132 15392
rect 48364 14720 48404 15352
rect 48460 15343 48500 15352
rect 49132 15343 49172 15352
rect 50188 15308 50228 15317
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 48364 14671 48404 14680
rect 49228 14720 49268 14729
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 48843 13460 48885 13469
rect 48843 13420 48844 13460
rect 48884 13420 48885 13460
rect 48843 13411 48885 13420
rect 48556 13208 48596 13217
rect 48268 13168 48556 13208
rect 47979 13124 48021 13133
rect 47979 13084 47980 13124
rect 48020 13084 48021 13124
rect 47979 13075 48021 13084
rect 47980 12990 48020 13075
rect 48075 13040 48117 13049
rect 48075 13000 48076 13040
rect 48116 13000 48117 13040
rect 48075 12991 48117 13000
rect 47787 12788 47829 12797
rect 47787 12748 47788 12788
rect 47828 12748 47829 12788
rect 47787 12739 47829 12748
rect 47691 12704 47733 12713
rect 47691 12664 47692 12704
rect 47732 12664 47733 12704
rect 47691 12655 47733 12664
rect 47980 12536 48020 12545
rect 47596 12496 47980 12536
rect 47980 12487 48020 12496
rect 48076 12368 48116 12991
rect 48172 12980 48212 13168
rect 48556 13159 48596 13168
rect 48748 13208 48788 13217
rect 48652 13124 48692 13133
rect 48172 12940 48404 12980
rect 48172 12713 48212 12940
rect 48171 12704 48213 12713
rect 48171 12664 48172 12704
rect 48212 12664 48213 12704
rect 48171 12655 48213 12664
rect 48267 12620 48309 12629
rect 48267 12580 48268 12620
rect 48308 12580 48309 12620
rect 48267 12571 48309 12580
rect 48364 12620 48404 12940
rect 48364 12571 48404 12580
rect 48268 12536 48308 12571
rect 48652 12545 48692 13084
rect 48268 12485 48308 12496
rect 48651 12536 48693 12545
rect 48651 12496 48652 12536
rect 48692 12496 48693 12536
rect 48651 12487 48693 12496
rect 47980 12328 48116 12368
rect 48652 12368 48692 12377
rect 48748 12368 48788 13168
rect 48844 12536 48884 13411
rect 49228 13301 49268 14680
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 49227 13292 49269 13301
rect 49227 13252 49228 13292
rect 49268 13252 49269 13292
rect 49227 13243 49269 13252
rect 49612 13208 49652 13217
rect 49516 13168 49612 13208
rect 49228 13124 49268 13133
rect 48940 12704 48980 12713
rect 49228 12704 49268 13084
rect 49323 13124 49365 13133
rect 49323 13084 49324 13124
rect 49364 13084 49365 13124
rect 49323 13075 49365 13084
rect 48980 12664 49268 12704
rect 48940 12655 48980 12664
rect 48844 12487 48884 12496
rect 49035 12536 49077 12545
rect 49035 12496 49036 12536
rect 49076 12496 49077 12536
rect 49035 12487 49077 12496
rect 49132 12536 49172 12547
rect 48692 12328 48788 12368
rect 47692 12284 47732 12293
rect 47692 11696 47732 12244
rect 47788 11696 47828 11705
rect 47692 11656 47788 11696
rect 47788 11647 47828 11656
rect 47883 11696 47925 11705
rect 47883 11656 47884 11696
rect 47924 11656 47925 11696
rect 47883 11647 47925 11656
rect 47980 11696 48020 12328
rect 48652 12319 48692 12328
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 48267 11948 48309 11957
rect 48267 11908 48268 11948
rect 48308 11908 48309 11948
rect 48267 11899 48309 11908
rect 48268 11814 48308 11899
rect 48555 11864 48597 11873
rect 48555 11824 48556 11864
rect 48596 11824 48597 11864
rect 48555 11815 48597 11824
rect 48940 11864 48980 11873
rect 47980 11647 48020 11656
rect 48076 11696 48116 11705
rect 48268 11696 48308 11705
rect 48116 11656 48268 11696
rect 48076 11647 48116 11656
rect 48268 11647 48308 11656
rect 48459 11696 48501 11705
rect 48459 11656 48460 11696
rect 48500 11656 48501 11696
rect 48459 11647 48501 11656
rect 48556 11696 48596 11815
rect 48556 11647 48596 11656
rect 47884 11562 47924 11647
rect 48363 11612 48405 11621
rect 48363 11572 48364 11612
rect 48404 11572 48405 11612
rect 48363 11563 48405 11572
rect 48172 11192 48212 11201
rect 48364 11192 48404 11563
rect 48460 11562 48500 11647
rect 48212 11152 48404 11192
rect 48172 11143 48212 11152
rect 48940 11033 48980 11824
rect 49036 11705 49076 12487
rect 49132 12461 49172 12496
rect 49324 12536 49364 13075
rect 49516 12713 49556 13168
rect 49612 13159 49652 13168
rect 49707 13208 49749 13217
rect 49707 13168 49708 13208
rect 49748 13168 49749 13208
rect 49707 13159 49749 13168
rect 49708 12980 49748 13159
rect 49612 12940 49748 12980
rect 49515 12704 49557 12713
rect 49515 12664 49516 12704
rect 49556 12664 49557 12704
rect 49515 12655 49557 12664
rect 49131 12452 49173 12461
rect 49131 12412 49132 12452
rect 49172 12412 49173 12452
rect 49131 12403 49173 12412
rect 49228 11873 49268 11958
rect 49227 11864 49269 11873
rect 49227 11824 49228 11864
rect 49268 11824 49269 11864
rect 49227 11815 49269 11824
rect 49035 11696 49077 11705
rect 49035 11656 49036 11696
rect 49076 11656 49077 11696
rect 49035 11647 49077 11656
rect 49227 11696 49269 11705
rect 49227 11656 49228 11696
rect 49268 11656 49269 11696
rect 49324 11696 49364 12496
rect 49515 12536 49557 12545
rect 49515 12496 49516 12536
rect 49556 12496 49557 12536
rect 49515 12487 49557 12496
rect 49419 12452 49461 12461
rect 49419 12412 49420 12452
rect 49460 12412 49461 12452
rect 49419 12403 49461 12412
rect 49420 12318 49460 12403
rect 49516 12402 49556 12487
rect 49420 11696 49460 11705
rect 49324 11656 49420 11696
rect 49227 11647 49269 11656
rect 49420 11647 49460 11656
rect 49516 11696 49556 11707
rect 49228 11562 49268 11647
rect 49516 11621 49556 11656
rect 49515 11612 49557 11621
rect 49515 11572 49516 11612
rect 49556 11572 49557 11612
rect 49515 11563 49557 11572
rect 48939 11024 48981 11033
rect 48939 10984 48940 11024
rect 48980 10984 48981 11024
rect 48939 10975 48981 10984
rect 49324 11024 49364 11033
rect 49612 11024 49652 12940
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 49707 12704 49749 12713
rect 49707 12664 49708 12704
rect 49748 12664 49749 12704
rect 49707 12655 49749 12664
rect 49708 12368 49748 12655
rect 49708 12319 49748 12328
rect 50092 12284 50132 12293
rect 50092 11705 50132 12244
rect 50091 11696 50133 11705
rect 50091 11656 50092 11696
rect 50132 11656 50133 11696
rect 50091 11647 50133 11656
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 50188 11201 50228 15268
rect 50284 12452 50324 15436
rect 50379 15427 50421 15436
rect 50380 15342 50420 15427
rect 50379 15056 50421 15065
rect 50379 15016 50380 15056
rect 50420 15016 50421 15056
rect 50379 15007 50421 15016
rect 50380 14972 50420 15007
rect 50380 14921 50420 14932
rect 50476 13637 50516 16771
rect 50572 16409 50612 18451
rect 50764 18416 50804 18425
rect 50668 17744 50708 17753
rect 50764 17744 50804 18376
rect 50708 17704 50804 17744
rect 51148 18332 51188 18341
rect 50668 17695 50708 17704
rect 51148 17669 51188 18292
rect 51244 18005 51284 18460
rect 51340 18451 51380 18460
rect 51531 18500 51573 18509
rect 51531 18460 51532 18500
rect 51572 18460 51573 18500
rect 51531 18451 51573 18460
rect 51532 18366 51572 18451
rect 51339 18332 51381 18341
rect 51339 18292 51340 18332
rect 51380 18292 51381 18332
rect 51339 18283 51381 18292
rect 51243 17996 51285 18005
rect 51243 17956 51244 17996
rect 51284 17956 51285 17996
rect 51243 17947 51285 17956
rect 51147 17660 51189 17669
rect 51147 17620 51148 17660
rect 51188 17620 51189 17660
rect 51147 17611 51189 17620
rect 50667 17324 50709 17333
rect 50667 17284 50668 17324
rect 50708 17284 50709 17324
rect 50667 17275 50709 17284
rect 50668 17072 50708 17275
rect 50668 17023 50708 17032
rect 50763 17072 50805 17081
rect 51051 17072 51093 17081
rect 50763 17032 50764 17072
rect 50804 17032 50996 17072
rect 50763 17023 50805 17032
rect 50764 16938 50804 17023
rect 50667 16904 50709 16913
rect 50667 16864 50668 16904
rect 50708 16864 50709 16904
rect 50667 16855 50709 16864
rect 50571 16400 50613 16409
rect 50571 16360 50572 16400
rect 50612 16360 50613 16400
rect 50571 16351 50613 16360
rect 50571 15560 50613 15569
rect 50571 15520 50572 15560
rect 50612 15520 50613 15560
rect 50571 15511 50613 15520
rect 50572 15308 50612 15511
rect 50572 14141 50612 15268
rect 50571 14132 50613 14141
rect 50571 14092 50572 14132
rect 50612 14092 50613 14132
rect 50571 14083 50613 14092
rect 50475 13628 50517 13637
rect 50475 13588 50476 13628
rect 50516 13588 50517 13628
rect 50475 13579 50517 13588
rect 50475 13208 50517 13217
rect 50475 13168 50476 13208
rect 50516 13168 50517 13208
rect 50475 13159 50517 13168
rect 50476 13074 50516 13159
rect 50284 12403 50324 12412
rect 50283 11696 50325 11705
rect 50283 11656 50284 11696
rect 50324 11656 50325 11696
rect 50283 11647 50325 11656
rect 50187 11192 50229 11201
rect 50187 11152 50188 11192
rect 50228 11152 50229 11192
rect 50187 11143 50229 11152
rect 49364 10984 49652 11024
rect 50187 11024 50229 11033
rect 50187 10984 50188 11024
rect 50228 10984 50229 11024
rect 49324 10975 49364 10984
rect 50187 10975 50229 10984
rect 50188 10890 50228 10975
rect 49419 10688 49461 10697
rect 49419 10648 49420 10688
rect 49460 10648 49461 10688
rect 49419 10639 49461 10648
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 49227 10520 49269 10529
rect 49227 10480 49228 10520
rect 49268 10480 49269 10520
rect 49227 10471 49269 10480
rect 49228 10436 49268 10471
rect 49228 10385 49268 10396
rect 48076 10184 48116 10193
rect 47979 9428 48021 9437
rect 47979 9388 47980 9428
rect 48020 9388 48021 9428
rect 47979 9379 48021 9388
rect 46827 8168 46869 8177
rect 46827 8128 46828 8168
rect 46868 8128 46869 8168
rect 46827 8119 46869 8128
rect 47019 8168 47061 8177
rect 47019 8128 47020 8168
rect 47060 8128 47061 8168
rect 47019 8119 47061 8128
rect 47499 8168 47541 8177
rect 47499 8128 47500 8168
rect 47540 8128 47541 8168
rect 47499 8119 47541 8128
rect 47691 8168 47733 8177
rect 47691 8128 47692 8168
rect 47732 8128 47733 8168
rect 47691 8119 47733 8128
rect 46731 8000 46773 8009
rect 46731 7960 46732 8000
rect 46772 7960 46773 8000
rect 46731 7951 46773 7960
rect 46828 8000 46868 8119
rect 46732 7866 46772 7951
rect 45812 7120 46004 7160
rect 46635 7160 46677 7169
rect 46635 7120 46636 7160
rect 46676 7120 46677 7160
rect 45772 7111 45812 7120
rect 46635 7111 46677 7120
rect 46636 7026 46676 7111
rect 46828 6581 46868 7960
rect 47020 8000 47060 8119
rect 47020 7951 47060 7960
rect 47212 8000 47252 8009
rect 47020 7832 47060 7841
rect 47212 7832 47252 7960
rect 47307 8000 47349 8009
rect 47500 8000 47540 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 47404 7960 47500 8000
rect 47308 7866 47348 7951
rect 47060 7792 47252 7832
rect 47020 7783 47060 7792
rect 47115 7160 47157 7169
rect 47115 7120 47116 7160
rect 47156 7120 47157 7160
rect 47115 7111 47157 7120
rect 46827 6572 46869 6581
rect 46827 6532 46828 6572
rect 46868 6532 46869 6572
rect 46827 6523 46869 6532
rect 45579 6488 45621 6497
rect 45579 6448 45580 6488
rect 45620 6448 45621 6488
rect 45579 6439 45621 6448
rect 45483 6404 45525 6413
rect 45483 6364 45484 6404
rect 45524 6364 45525 6404
rect 45483 6355 45525 6364
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 46348 5816 46388 5825
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 45867 5060 45909 5069
rect 45867 5020 45868 5060
rect 45908 5020 45909 5060
rect 45867 5011 45909 5020
rect 45868 4926 45908 5011
rect 46252 4976 46292 4985
rect 46348 4976 46388 5776
rect 46292 4936 46388 4976
rect 47116 4976 47156 7111
rect 47212 6656 47252 6665
rect 47404 6656 47444 7960
rect 47500 7951 47540 7960
rect 47499 7748 47541 7757
rect 47499 7708 47500 7748
rect 47540 7708 47541 7748
rect 47499 7699 47541 7708
rect 47500 7614 47540 7699
rect 47499 7412 47541 7421
rect 47499 7372 47500 7412
rect 47540 7372 47541 7412
rect 47499 7363 47541 7372
rect 47252 6616 47444 6656
rect 47212 6607 47252 6616
rect 47308 6488 47348 6499
rect 47308 6413 47348 6448
rect 47403 6488 47445 6497
rect 47403 6448 47404 6488
rect 47444 6448 47445 6488
rect 47403 6439 47445 6448
rect 47500 6488 47540 7363
rect 47500 6439 47540 6448
rect 47692 6488 47732 8119
rect 47980 8000 48020 9379
rect 48076 8681 48116 10144
rect 48939 10184 48981 10193
rect 48939 10144 48940 10184
rect 48980 10144 48981 10184
rect 48939 10135 48981 10144
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 48459 8756 48501 8765
rect 48459 8716 48460 8756
rect 48500 8716 48501 8756
rect 48459 8707 48501 8716
rect 48075 8672 48117 8681
rect 48075 8632 48076 8672
rect 48116 8632 48117 8672
rect 48075 8623 48117 8632
rect 48460 8672 48500 8707
rect 48267 8168 48309 8177
rect 48267 8128 48268 8168
rect 48308 8128 48309 8168
rect 48267 8119 48309 8128
rect 48268 8000 48308 8119
rect 48020 7960 48212 8000
rect 47980 7951 48020 7960
rect 47787 7412 47829 7421
rect 47787 7372 47788 7412
rect 47828 7372 47829 7412
rect 47787 7363 47829 7372
rect 47979 7412 48021 7421
rect 47979 7372 47980 7412
rect 48020 7372 48021 7412
rect 47979 7363 48021 7372
rect 47788 7278 47828 7363
rect 47692 6439 47732 6448
rect 47883 6488 47925 6497
rect 47883 6448 47884 6488
rect 47924 6448 47925 6488
rect 47883 6439 47925 6448
rect 47980 6488 48020 7363
rect 47980 6439 48020 6448
rect 47307 6404 47349 6413
rect 47307 6364 47308 6404
rect 47348 6364 47349 6404
rect 47307 6355 47349 6364
rect 47308 5657 47348 6355
rect 47404 5825 47444 6439
rect 47884 6354 47924 6439
rect 47692 6236 47732 6245
rect 47500 6196 47692 6236
rect 47403 5816 47445 5825
rect 47403 5776 47404 5816
rect 47444 5776 47445 5816
rect 47403 5767 47445 5776
rect 46252 4927 46292 4936
rect 47116 4927 47156 4936
rect 47212 5648 47252 5657
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 47212 4136 47252 5608
rect 47307 5648 47349 5657
rect 47307 5608 47308 5648
rect 47348 5608 47349 5648
rect 47307 5599 47349 5608
rect 47404 5648 47444 5657
rect 47308 5480 47348 5489
rect 47308 5069 47348 5440
rect 47307 5060 47349 5069
rect 47307 5020 47308 5060
rect 47348 5020 47349 5060
rect 47307 5011 47349 5020
rect 47404 4817 47444 5608
rect 47500 5648 47540 6196
rect 47692 6187 47732 6196
rect 47595 5816 47637 5825
rect 47595 5776 47596 5816
rect 47636 5776 47637 5816
rect 47595 5767 47637 5776
rect 47500 5599 47540 5608
rect 47499 5480 47541 5489
rect 47499 5440 47500 5480
rect 47540 5440 47541 5480
rect 47499 5431 47541 5440
rect 47403 4808 47445 4817
rect 47403 4768 47404 4808
rect 47444 4768 47445 4808
rect 47403 4759 47445 4768
rect 47404 4136 47444 4145
rect 47212 4096 47404 4136
rect 47404 4087 47444 4096
rect 47500 4136 47540 5431
rect 47500 4087 47540 4096
rect 47596 4136 47636 5767
rect 48172 5648 48212 7960
rect 48268 7951 48308 7960
rect 48364 8000 48404 8009
rect 48267 7748 48309 7757
rect 48267 7708 48268 7748
rect 48308 7708 48309 7748
rect 48267 7699 48309 7708
rect 48172 5599 48212 5608
rect 48268 5396 48308 7699
rect 48364 7421 48404 7960
rect 48460 7757 48500 8632
rect 48652 8672 48692 8681
rect 48844 8672 48884 8681
rect 48940 8672 48980 10135
rect 49324 8840 49364 8849
rect 48555 8588 48597 8597
rect 48555 8548 48556 8588
rect 48596 8548 48597 8588
rect 48555 8539 48597 8548
rect 48556 8009 48596 8539
rect 48555 8000 48597 8009
rect 48555 7960 48556 8000
rect 48596 7960 48597 8000
rect 48555 7951 48597 7960
rect 48652 7832 48692 8632
rect 48652 7783 48692 7792
rect 48748 8632 48844 8672
rect 48884 8632 48980 8672
rect 49036 8672 49076 8683
rect 48748 7757 48788 8632
rect 48844 8623 48884 8632
rect 49036 8597 49076 8632
rect 49132 8672 49172 8681
rect 49035 8588 49077 8597
rect 49035 8548 49036 8588
rect 49076 8548 49077 8588
rect 49035 8539 49077 8548
rect 48940 8504 48980 8513
rect 48843 8168 48885 8177
rect 48843 8128 48844 8168
rect 48884 8128 48885 8168
rect 48843 8119 48885 8128
rect 48844 8013 48884 8119
rect 48940 8009 48980 8464
rect 49035 8252 49077 8261
rect 49035 8212 49036 8252
rect 49076 8212 49077 8252
rect 49035 8203 49077 8212
rect 48844 7964 48884 7973
rect 48939 8000 48981 8009
rect 48939 7960 48940 8000
rect 48980 7960 48981 8000
rect 48939 7951 48981 7960
rect 49036 8000 49076 8203
rect 49036 7951 49076 7960
rect 48940 7832 48980 7841
rect 48459 7748 48501 7757
rect 48459 7708 48460 7748
rect 48500 7708 48501 7748
rect 48459 7699 48501 7708
rect 48747 7748 48789 7757
rect 48747 7708 48748 7748
rect 48788 7708 48789 7748
rect 48940 7748 48980 7792
rect 49132 7748 49172 8632
rect 48940 7708 49172 7748
rect 48747 7699 48789 7708
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 48363 7412 48405 7421
rect 48363 7372 48364 7412
rect 48404 7372 48405 7412
rect 48363 7363 48405 7372
rect 49035 7412 49077 7421
rect 49035 7372 49036 7412
rect 49076 7372 49077 7412
rect 49035 7363 49077 7372
rect 48747 7244 48789 7253
rect 48747 7204 48748 7244
rect 48788 7204 48789 7244
rect 48747 7195 48789 7204
rect 48363 7160 48405 7169
rect 48363 7120 48364 7160
rect 48404 7120 48405 7160
rect 48363 7111 48405 7120
rect 48748 7160 48788 7195
rect 48364 7026 48404 7111
rect 48748 7109 48788 7120
rect 49036 6992 49076 7363
rect 49132 7160 49172 7169
rect 49324 7160 49364 8800
rect 49420 8009 49460 10639
rect 49515 10436 49557 10445
rect 49515 10396 49516 10436
rect 49556 10396 49557 10436
rect 49515 10387 49557 10396
rect 49419 8000 49461 8009
rect 49419 7960 49420 8000
rect 49460 7960 49461 8000
rect 49419 7951 49461 7960
rect 49420 7866 49460 7951
rect 49172 7120 49364 7160
rect 49132 7111 49172 7120
rect 49516 6992 49556 10387
rect 49803 10184 49845 10193
rect 49803 10144 49804 10184
rect 49844 10144 49845 10184
rect 49803 10135 49845 10144
rect 50188 10184 50228 10193
rect 49804 10050 49844 10135
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 50188 9344 50228 10144
rect 50284 9521 50324 11647
rect 50668 11033 50708 16855
rect 50956 16484 50996 17032
rect 51051 17032 51052 17072
rect 51092 17032 51093 17072
rect 51051 17023 51093 17032
rect 51052 16904 51092 17023
rect 51052 16855 51092 16864
rect 51052 16484 51092 16493
rect 50764 16444 51052 16484
rect 50764 15560 50804 16444
rect 51052 16435 51092 16444
rect 51148 15728 51188 17611
rect 51244 16988 51284 16997
rect 51244 16829 51284 16948
rect 51243 16820 51285 16829
rect 51243 16780 51244 16820
rect 51284 16780 51285 16820
rect 51243 16771 51285 16780
rect 51243 16232 51285 16241
rect 51243 16192 51244 16232
rect 51284 16192 51285 16232
rect 51243 16183 51285 16192
rect 50956 15688 51188 15728
rect 50764 15511 50804 15520
rect 50860 15560 50900 15569
rect 50956 15560 50996 15688
rect 50900 15520 50996 15560
rect 51051 15560 51093 15569
rect 51051 15520 51052 15560
rect 51092 15520 51093 15560
rect 50764 14636 50804 14645
rect 50764 13721 50804 14596
rect 50763 13712 50805 13721
rect 50763 13672 50764 13712
rect 50804 13672 50805 13712
rect 50763 13663 50805 13672
rect 50860 13301 50900 15520
rect 51051 15511 51093 15520
rect 51244 15560 51284 16183
rect 51340 15905 51380 18283
rect 51532 17744 51572 17753
rect 51435 17240 51477 17249
rect 51435 17200 51436 17240
rect 51476 17200 51477 17240
rect 51435 17191 51477 17200
rect 51436 17106 51476 17191
rect 51436 16820 51476 16829
rect 51436 16325 51476 16780
rect 51435 16316 51477 16325
rect 51435 16276 51436 16316
rect 51476 16276 51477 16316
rect 51435 16267 51477 16276
rect 51532 16241 51572 17704
rect 51628 17249 51668 20467
rect 52011 19088 52053 19097
rect 52011 19048 52012 19088
rect 52052 19048 52053 19088
rect 52011 19039 52053 19048
rect 52012 18954 52052 19039
rect 52108 18500 52148 21988
rect 52299 21988 52300 22028
rect 52340 21988 52341 22028
rect 52299 21979 52341 21988
rect 52299 21608 52341 21617
rect 52299 21568 52300 21608
rect 52340 21568 52341 21608
rect 52299 21559 52341 21568
rect 52396 21608 52436 21617
rect 52492 21608 52532 22408
rect 52588 22280 52628 22291
rect 52684 22289 52724 22492
rect 52588 22205 52628 22240
rect 52683 22280 52725 22289
rect 52683 22240 52684 22280
rect 52724 22240 52725 22280
rect 52683 22231 52725 22240
rect 52587 22196 52629 22205
rect 52587 22156 52588 22196
rect 52628 22156 52629 22196
rect 52587 22147 52629 22156
rect 52436 21568 52532 21608
rect 52587 21608 52629 21617
rect 52587 21568 52588 21608
rect 52628 21568 52629 21608
rect 52396 21559 52436 21568
rect 52587 21559 52629 21568
rect 52684 21608 52724 21617
rect 52780 21608 52820 23239
rect 52972 22961 53012 23752
rect 52971 22952 53013 22961
rect 52971 22912 52972 22952
rect 53012 22912 53013 22952
rect 52971 22903 53013 22912
rect 53164 22784 53204 24592
rect 53547 24592 53548 24632
rect 53588 24592 53589 24632
rect 53547 24583 53589 24592
rect 54028 24305 54068 29203
rect 54219 29168 54261 29177
rect 54219 29128 54220 29168
rect 54260 29128 54261 29168
rect 54219 29119 54261 29128
rect 54220 29034 54260 29119
rect 54316 28412 54356 29203
rect 54699 28832 54741 28841
rect 54699 28792 54700 28832
rect 54740 28792 54741 28832
rect 54699 28783 54741 28792
rect 54412 28412 54452 28421
rect 54316 28372 54412 28412
rect 54412 28363 54452 28372
rect 54507 27992 54549 28001
rect 54507 27952 54508 27992
rect 54548 27952 54549 27992
rect 54507 27943 54549 27952
rect 54508 27824 54548 27943
rect 54508 27775 54548 27784
rect 54700 27656 54740 28783
rect 54795 28496 54837 28505
rect 54795 28456 54796 28496
rect 54836 28456 54837 28496
rect 54795 28447 54837 28456
rect 54796 27824 54836 28447
rect 54796 27775 54836 27784
rect 54700 27607 54740 27616
rect 54892 27656 54932 29632
rect 55372 29336 55412 29800
rect 55372 29177 55412 29296
rect 55179 29168 55221 29177
rect 55179 29128 55180 29168
rect 55220 29128 55221 29168
rect 55179 29119 55221 29128
rect 55371 29168 55413 29177
rect 55371 29128 55372 29168
rect 55412 29128 55413 29168
rect 55371 29119 55413 29128
rect 55083 29000 55125 29009
rect 55083 28960 55084 29000
rect 55124 28960 55125 29000
rect 55083 28951 55125 28960
rect 55084 27740 55124 28951
rect 55180 28328 55220 29119
rect 55275 28580 55317 28589
rect 55275 28540 55276 28580
rect 55316 28540 55317 28580
rect 55275 28531 55317 28540
rect 55276 28446 55316 28531
rect 55372 28328 55412 29119
rect 55468 28589 55508 29800
rect 55660 29840 55700 29849
rect 55660 29681 55700 29800
rect 55659 29672 55701 29681
rect 55659 29632 55660 29672
rect 55700 29632 55701 29672
rect 55659 29623 55701 29632
rect 55564 29168 55604 29177
rect 55564 28841 55604 29128
rect 55660 29168 55700 29177
rect 55660 28925 55700 29128
rect 55756 29168 55796 30136
rect 55852 29933 55892 30304
rect 56044 30176 56084 30617
rect 56236 30353 56276 30640
rect 56524 30512 56564 31312
rect 56619 31352 56661 31361
rect 56619 31312 56620 31352
rect 56660 31312 56661 31352
rect 56619 31303 56661 31312
rect 56620 30512 56660 30521
rect 56524 30472 56620 30512
rect 56620 30463 56660 30472
rect 56235 30344 56277 30353
rect 56235 30304 56236 30344
rect 56276 30304 56277 30344
rect 56235 30295 56277 30304
rect 56044 30136 56276 30176
rect 56043 30008 56085 30017
rect 56043 29968 56044 30008
rect 56084 29968 56085 30008
rect 56043 29959 56085 29968
rect 55851 29924 55893 29933
rect 55851 29884 55852 29924
rect 55892 29884 55893 29924
rect 55851 29875 55893 29884
rect 55852 29840 55892 29875
rect 55852 29789 55892 29800
rect 56044 29840 56084 29959
rect 56236 29849 56276 30136
rect 56044 29791 56084 29800
rect 56140 29840 56180 29849
rect 55948 29672 55988 29681
rect 55948 29261 55988 29632
rect 56043 29672 56085 29681
rect 56043 29632 56044 29672
rect 56084 29632 56085 29672
rect 56043 29623 56085 29632
rect 55947 29252 55989 29261
rect 55947 29212 55948 29252
rect 55988 29212 55989 29252
rect 55947 29203 55989 29212
rect 55659 28916 55701 28925
rect 55659 28876 55660 28916
rect 55700 28876 55701 28916
rect 55659 28867 55701 28876
rect 55563 28832 55605 28841
rect 55563 28792 55564 28832
rect 55604 28792 55605 28832
rect 55563 28783 55605 28792
rect 55467 28580 55509 28589
rect 55467 28540 55468 28580
rect 55508 28540 55509 28580
rect 55467 28531 55509 28540
rect 55564 28328 55604 28337
rect 55180 28288 55316 28328
rect 55372 28288 55564 28328
rect 55179 27740 55221 27749
rect 55084 27700 55180 27740
rect 55220 27700 55221 27740
rect 55179 27691 55221 27700
rect 54892 27607 54932 27616
rect 54988 27656 55028 27665
rect 54988 27488 55028 27616
rect 55180 27656 55220 27691
rect 55180 27605 55220 27616
rect 55180 27488 55220 27497
rect 54988 27448 55180 27488
rect 55180 27439 55220 27448
rect 54219 27068 54261 27077
rect 54219 27028 54220 27068
rect 54260 27028 54261 27068
rect 54219 27019 54261 27028
rect 54220 26934 54260 27019
rect 55276 26816 55316 28288
rect 55564 28279 55604 28288
rect 55659 28328 55701 28337
rect 55659 28288 55660 28328
rect 55700 28288 55701 28328
rect 55659 28279 55701 28288
rect 55660 28194 55700 28279
rect 55756 28169 55796 29128
rect 55851 29168 55893 29177
rect 55851 29128 55852 29168
rect 55892 29128 55893 29168
rect 55851 29119 55893 29128
rect 55852 29034 55892 29119
rect 55947 28748 55989 28757
rect 55947 28708 55948 28748
rect 55988 28708 55989 28748
rect 55947 28699 55989 28708
rect 55948 28580 55988 28699
rect 55852 28540 55988 28580
rect 55755 28160 55797 28169
rect 55755 28120 55756 28160
rect 55796 28120 55797 28160
rect 55755 28111 55797 28120
rect 55372 27656 55412 27665
rect 55372 27581 55412 27616
rect 55468 27656 55508 27665
rect 55660 27656 55700 27665
rect 55508 27616 55660 27656
rect 55468 27607 55508 27616
rect 55371 27572 55413 27581
rect 55371 27532 55372 27572
rect 55412 27532 55413 27572
rect 55371 27523 55413 27532
rect 55372 26984 55412 27523
rect 55660 27077 55700 27616
rect 55756 27656 55796 28111
rect 55756 27607 55796 27616
rect 55852 27656 55892 28540
rect 55948 28328 55988 28337
rect 56044 28328 56084 29623
rect 55988 28288 56084 28328
rect 55948 28279 55988 28288
rect 55852 27607 55892 27616
rect 55947 27656 55989 27665
rect 55947 27616 55948 27656
rect 55988 27616 55989 27656
rect 55947 27607 55989 27616
rect 55948 27522 55988 27607
rect 55659 27068 55701 27077
rect 55659 27028 55660 27068
rect 55700 27028 55892 27068
rect 55659 27019 55701 27028
rect 55372 26944 55508 26984
rect 55372 26816 55412 26825
rect 55276 26776 55372 26816
rect 55468 26816 55508 26944
rect 55660 26934 55700 27019
rect 55468 26776 55700 26816
rect 55372 26767 55412 26776
rect 55467 26648 55509 26657
rect 55467 26608 55468 26648
rect 55508 26608 55509 26648
rect 55467 26599 55509 26608
rect 55468 26153 55508 26599
rect 55467 26144 55509 26153
rect 55467 26104 55468 26144
rect 55508 26104 55509 26144
rect 55467 26095 55509 26104
rect 55468 26010 55508 26095
rect 54891 25976 54933 25985
rect 54891 25936 54892 25976
rect 54932 25936 54933 25976
rect 54891 25927 54933 25936
rect 54699 25892 54741 25901
rect 54699 25852 54700 25892
rect 54740 25852 54741 25892
rect 54699 25843 54741 25852
rect 54700 25397 54740 25843
rect 54892 25842 54932 25927
rect 54699 25388 54741 25397
rect 54699 25348 54700 25388
rect 54740 25348 54741 25388
rect 54699 25339 54741 25348
rect 54700 25254 54740 25339
rect 55468 25313 55508 25398
rect 55275 25304 55317 25313
rect 55275 25264 55276 25304
rect 55316 25264 55317 25304
rect 55275 25255 55317 25264
rect 55467 25304 55509 25313
rect 55467 25264 55468 25304
rect 55508 25264 55509 25304
rect 55467 25255 55509 25264
rect 55564 25304 55604 25313
rect 55276 25170 55316 25255
rect 54699 25136 54741 25145
rect 54699 25096 54700 25136
rect 54740 25096 54741 25136
rect 54699 25087 54741 25096
rect 55372 25136 55412 25145
rect 54027 24296 54069 24305
rect 54027 24256 54028 24296
rect 54068 24256 54069 24296
rect 54027 24247 54069 24256
rect 54700 23801 54740 25087
rect 55372 24884 55412 25096
rect 55467 25136 55509 25145
rect 55467 25096 55468 25136
rect 55508 25096 55509 25136
rect 55467 25087 55509 25096
rect 54892 24844 55412 24884
rect 54892 24716 54932 24844
rect 54892 24667 54932 24676
rect 55179 24716 55221 24725
rect 55179 24676 55180 24716
rect 55220 24676 55221 24716
rect 55179 24667 55221 24676
rect 54699 23792 54741 23801
rect 54699 23752 54700 23792
rect 54740 23752 54741 23792
rect 54699 23743 54741 23752
rect 54796 23792 54836 23801
rect 54123 23624 54165 23633
rect 54123 23584 54124 23624
rect 54164 23584 54165 23624
rect 54123 23575 54165 23584
rect 54124 23490 54164 23575
rect 54315 23288 54357 23297
rect 54315 23248 54316 23288
rect 54356 23248 54357 23288
rect 54315 23239 54357 23248
rect 53643 23204 53685 23213
rect 53643 23164 53644 23204
rect 53684 23164 53685 23204
rect 53643 23155 53685 23164
rect 53644 23060 53684 23155
rect 54316 23060 54356 23239
rect 54796 23213 54836 23752
rect 55180 23792 55220 24667
rect 55276 24632 55316 24641
rect 55468 24632 55508 25087
rect 55316 24592 55508 24632
rect 55276 24583 55316 24592
rect 55564 24053 55604 25264
rect 55563 24044 55605 24053
rect 55563 24004 55564 24044
rect 55604 24004 55605 24044
rect 55563 23995 55605 24004
rect 55660 23792 55700 26776
rect 55852 26228 55892 27028
rect 56044 26657 56084 28288
rect 56140 28160 56180 29800
rect 56235 29840 56277 29849
rect 56235 29800 56236 29840
rect 56276 29800 56277 29840
rect 56235 29791 56277 29800
rect 56236 28328 56276 29791
rect 56331 29252 56373 29261
rect 56331 29212 56332 29252
rect 56372 29212 56373 29252
rect 56331 29203 56373 29212
rect 56332 29118 56372 29203
rect 56716 29168 56756 29177
rect 56427 28664 56469 28673
rect 56427 28624 56428 28664
rect 56468 28624 56469 28664
rect 56427 28615 56469 28624
rect 56428 28337 56468 28615
rect 56716 28496 56756 29128
rect 56812 28496 56852 28505
rect 56716 28456 56812 28496
rect 56812 28447 56852 28456
rect 56236 28279 56276 28288
rect 56427 28328 56469 28337
rect 56427 28288 56428 28328
rect 56468 28288 56469 28328
rect 56427 28279 56469 28288
rect 56332 28244 56372 28253
rect 56332 28160 56372 28204
rect 56428 28194 56468 28279
rect 56140 28120 56372 28160
rect 57099 28160 57141 28169
rect 57099 28120 57100 28160
rect 57140 28120 57141 28160
rect 57099 28111 57141 28120
rect 56811 27740 56853 27749
rect 56811 27700 56812 27740
rect 56852 27700 56853 27740
rect 56811 27691 56853 27700
rect 57100 27740 57140 28111
rect 57100 27691 57140 27700
rect 56331 27656 56373 27665
rect 56331 27616 56332 27656
rect 56372 27616 56373 27656
rect 56331 27607 56373 27616
rect 56236 26816 56276 26825
rect 56043 26648 56085 26657
rect 56043 26608 56044 26648
rect 56084 26608 56085 26648
rect 56043 26599 56085 26608
rect 55852 26179 55892 26188
rect 55755 26144 55797 26153
rect 55755 26104 55756 26144
rect 55796 26104 55797 26144
rect 55755 26095 55797 26104
rect 55756 26010 55796 26095
rect 56236 25985 56276 26776
rect 56332 26144 56372 27607
rect 56620 26732 56660 26741
rect 56428 26312 56468 26321
rect 56620 26312 56660 26692
rect 56468 26272 56660 26312
rect 56428 26263 56468 26272
rect 56332 26095 56372 26104
rect 56524 26144 56564 26153
rect 56235 25976 56277 25985
rect 56235 25936 56236 25976
rect 56276 25936 56277 25976
rect 56235 25927 56277 25936
rect 56140 25892 56180 25901
rect 55756 25472 55796 25481
rect 55756 25145 55796 25432
rect 56140 25304 56180 25852
rect 56236 25556 56276 25565
rect 56524 25556 56564 26104
rect 56620 26144 56660 26153
rect 56620 25976 56660 26104
rect 56812 26144 56852 27691
rect 57003 26312 57045 26321
rect 57003 26272 57004 26312
rect 57044 26272 57045 26312
rect 57003 26263 57045 26272
rect 56812 26095 56852 26104
rect 57004 26144 57044 26263
rect 57004 26095 57044 26104
rect 57100 26144 57140 26153
rect 56812 25976 56852 25985
rect 56620 25936 56812 25976
rect 56812 25927 56852 25936
rect 56276 25516 56564 25556
rect 56236 25313 56276 25516
rect 56140 25255 56180 25264
rect 56235 25304 56277 25313
rect 56235 25264 56236 25304
rect 56276 25264 56277 25304
rect 56235 25255 56277 25264
rect 56332 25304 56372 25313
rect 55755 25136 55797 25145
rect 55755 25096 55756 25136
rect 55796 25096 55797 25136
rect 55755 25087 55797 25096
rect 56139 24632 56181 24641
rect 56139 24592 56140 24632
rect 56180 24592 56181 24632
rect 56139 24583 56181 24592
rect 56140 24498 56180 24583
rect 56332 24557 56372 25264
rect 57100 25145 57140 26104
rect 57099 25136 57141 25145
rect 57099 25096 57100 25136
rect 57140 25096 57141 25136
rect 57099 25087 57141 25096
rect 56331 24548 56373 24557
rect 56331 24508 56332 24548
rect 56372 24508 56373 24548
rect 56331 24499 56373 24508
rect 57196 24473 57236 31555
rect 57387 31352 57429 31361
rect 57387 31312 57388 31352
rect 57428 31312 57429 31352
rect 57387 31303 57429 31312
rect 57579 31352 57621 31361
rect 57579 31312 57580 31352
rect 57620 31312 57621 31352
rect 57579 31303 57621 31312
rect 57388 31218 57428 31303
rect 57580 29168 57620 31303
rect 57676 30773 57716 32647
rect 58156 32646 58196 32731
rect 58252 32033 58292 32815
rect 58539 32780 58581 32789
rect 58539 32740 58540 32780
rect 58580 32740 58581 32780
rect 58539 32731 58581 32740
rect 58540 32646 58580 32731
rect 58348 32192 58388 32201
rect 58251 32024 58293 32033
rect 58251 31984 58252 32024
rect 58292 31984 58293 32024
rect 58251 31975 58293 31984
rect 58348 31781 58388 32152
rect 58636 32192 58676 32983
rect 58732 32276 58772 33100
rect 58924 32864 58964 33235
rect 59020 33125 59060 33664
rect 59212 33536 59252 33545
rect 59212 33293 59252 33496
rect 59211 33284 59253 33293
rect 59211 33244 59212 33284
rect 59252 33244 59253 33284
rect 59211 33235 59253 33244
rect 59019 33116 59061 33125
rect 59019 33076 59020 33116
rect 59060 33076 59061 33116
rect 59019 33067 59061 33076
rect 58924 32815 58964 32824
rect 58732 32227 58772 32236
rect 59020 32320 59252 32360
rect 58636 32143 58676 32152
rect 59020 32024 59060 32320
rect 59115 32192 59157 32201
rect 59115 32152 59116 32192
rect 59156 32152 59157 32192
rect 59115 32143 59157 32152
rect 59212 32192 59252 32320
rect 59308 32201 59348 34336
rect 59212 32143 59252 32152
rect 59307 32192 59349 32201
rect 59307 32152 59308 32192
rect 59348 32152 59349 32192
rect 59307 32143 59349 32152
rect 59404 32192 59444 34579
rect 59500 34133 59540 34756
rect 59788 34553 59828 35176
rect 59884 35167 59924 35176
rect 60172 35048 60212 37360
rect 60364 37400 60404 37409
rect 60267 37316 60309 37325
rect 60267 37276 60268 37316
rect 60308 37276 60309 37316
rect 60267 37267 60309 37276
rect 60268 37182 60308 37267
rect 60364 37232 60404 37360
rect 60460 37402 60500 37411
rect 60460 37316 60500 37362
rect 61132 37325 61172 37410
rect 61516 37400 61556 38032
rect 61612 38023 61652 38032
rect 62571 37988 62613 37997
rect 62571 37948 62572 37988
rect 62612 37948 62613 37988
rect 62571 37939 62613 37948
rect 61516 37351 61556 37360
rect 62379 37400 62421 37409
rect 62379 37360 62380 37400
rect 62420 37360 62421 37400
rect 62379 37351 62421 37360
rect 61131 37316 61173 37325
rect 60460 37276 60596 37316
rect 60364 37192 60500 37232
rect 60363 36896 60405 36905
rect 60363 36856 60364 36896
rect 60404 36856 60405 36896
rect 60363 36847 60405 36856
rect 60364 36728 60404 36847
rect 60364 36679 60404 36688
rect 60364 36056 60404 36065
rect 60268 35216 60308 35225
rect 60364 35216 60404 36016
rect 60308 35176 60404 35216
rect 60268 35167 60308 35176
rect 59884 35008 60212 35048
rect 59787 34544 59829 34553
rect 59787 34504 59788 34544
rect 59828 34504 59829 34544
rect 59787 34495 59829 34504
rect 59595 34208 59637 34217
rect 59595 34168 59596 34208
rect 59636 34168 59637 34208
rect 59595 34159 59637 34168
rect 59499 34124 59541 34133
rect 59499 34084 59500 34124
rect 59540 34084 59541 34124
rect 59499 34075 59541 34084
rect 59020 31975 59060 31984
rect 58347 31772 58389 31781
rect 58347 31732 58348 31772
rect 58388 31732 58389 31772
rect 58347 31723 58389 31732
rect 59116 31361 59156 32143
rect 59307 32024 59349 32033
rect 59307 31984 59308 32024
rect 59348 31984 59349 32024
rect 59307 31975 59349 31984
rect 59308 31890 59348 31975
rect 59307 31772 59349 31781
rect 59307 31732 59308 31772
rect 59348 31732 59349 31772
rect 59307 31723 59349 31732
rect 59115 31352 59157 31361
rect 59115 31312 59116 31352
rect 59156 31312 59157 31352
rect 59115 31303 59157 31312
rect 58540 31184 58580 31193
rect 57963 30848 58005 30857
rect 57963 30808 57964 30848
rect 58004 30808 58005 30848
rect 57963 30799 58005 30808
rect 57675 30764 57717 30773
rect 57675 30724 57676 30764
rect 57716 30724 57717 30764
rect 57675 30715 57717 30724
rect 57964 30714 58004 30799
rect 58540 30353 58580 31144
rect 59019 30932 59061 30941
rect 59019 30892 59020 30932
rect 59060 30892 59061 30932
rect 59019 30883 59061 30892
rect 58635 30680 58677 30689
rect 58635 30640 58636 30680
rect 58676 30640 58677 30680
rect 58635 30631 58677 30640
rect 58539 30344 58581 30353
rect 58539 30304 58540 30344
rect 58580 30304 58581 30344
rect 58539 30295 58581 30304
rect 58636 30008 58676 30631
rect 59020 30092 59060 30883
rect 59116 30680 59156 31303
rect 59116 30631 59156 30640
rect 59020 30052 59156 30092
rect 58636 29959 58676 29968
rect 58828 30008 58868 30019
rect 58828 29933 58868 29968
rect 58827 29924 58869 29933
rect 59020 29924 59060 29933
rect 58827 29884 58828 29924
rect 58868 29884 58869 29924
rect 58827 29875 58869 29884
rect 58924 29884 59020 29924
rect 57580 29119 57620 29128
rect 58732 28916 58772 28925
rect 58732 28673 58772 28876
rect 58731 28664 58773 28673
rect 58731 28624 58732 28664
rect 58772 28624 58773 28664
rect 58731 28615 58773 28624
rect 58636 28496 58676 28505
rect 58540 28456 58636 28496
rect 58676 28456 58868 28496
rect 58444 28412 58484 28421
rect 58444 27833 58484 28372
rect 58540 28085 58580 28456
rect 58636 28447 58676 28456
rect 58828 28412 58868 28456
rect 58828 28363 58868 28372
rect 58539 28076 58581 28085
rect 58539 28036 58540 28076
rect 58580 28036 58581 28076
rect 58539 28027 58581 28036
rect 58443 27824 58485 27833
rect 58443 27784 58444 27824
rect 58484 27784 58485 27824
rect 58443 27775 58485 27784
rect 57484 27656 57524 27665
rect 57484 26984 57524 27616
rect 58348 27656 58388 27665
rect 57963 27320 58005 27329
rect 57963 27280 57964 27320
rect 58004 27280 58005 27320
rect 57963 27271 58005 27280
rect 57580 26984 57620 26993
rect 57484 26944 57580 26984
rect 57580 26935 57620 26944
rect 57675 26984 57717 26993
rect 57675 26944 57676 26984
rect 57716 26944 57717 26984
rect 57675 26935 57717 26944
rect 57483 26816 57525 26825
rect 57483 26776 57484 26816
rect 57524 26776 57525 26816
rect 57483 26767 57525 26776
rect 57291 26144 57333 26153
rect 57291 26104 57292 26144
rect 57332 26104 57333 26144
rect 57291 26095 57333 26104
rect 57292 24548 57332 26095
rect 57484 26060 57524 26767
rect 57676 26312 57716 26935
rect 57676 26069 57716 26272
rect 57484 26011 57524 26020
rect 57675 26060 57717 26069
rect 57675 26020 57676 26060
rect 57716 26020 57717 26060
rect 57675 26011 57717 26020
rect 57387 25976 57429 25985
rect 57868 25976 57908 25985
rect 57387 25936 57388 25976
rect 57428 25936 57429 25976
rect 57387 25927 57429 25936
rect 57772 25936 57868 25976
rect 57388 25304 57428 25927
rect 57388 25255 57428 25264
rect 57772 25304 57812 25936
rect 57868 25927 57908 25936
rect 57772 25255 57812 25264
rect 57195 24464 57237 24473
rect 57195 24424 57196 24464
rect 57236 24424 57237 24464
rect 57195 24415 57237 24424
rect 55755 24044 55797 24053
rect 55755 24004 55756 24044
rect 55796 24004 55797 24044
rect 55755 23995 55797 24004
rect 55756 23910 55796 23995
rect 57292 23969 57332 24508
rect 57675 24380 57717 24389
rect 57675 24340 57676 24380
rect 57716 24340 57717 24380
rect 57675 24331 57717 24340
rect 55851 23960 55893 23969
rect 55851 23920 55852 23960
rect 55892 23920 55893 23960
rect 55851 23911 55893 23920
rect 57291 23960 57333 23969
rect 57291 23920 57292 23960
rect 57332 23920 57333 23960
rect 57291 23911 57333 23920
rect 55220 23752 55604 23792
rect 55180 23743 55220 23752
rect 54892 23624 54932 23633
rect 54795 23204 54837 23213
rect 54795 23164 54796 23204
rect 54836 23164 54837 23204
rect 54795 23155 54837 23164
rect 54603 23120 54645 23129
rect 54603 23080 54604 23120
rect 54644 23080 54740 23120
rect 54603 23071 54645 23080
rect 54700 23060 54740 23080
rect 54892 23060 54932 23584
rect 55276 23624 55316 23633
rect 55316 23584 55508 23624
rect 55276 23575 55316 23584
rect 55275 23204 55317 23213
rect 55275 23164 55276 23204
rect 55316 23164 55317 23204
rect 55275 23155 55317 23164
rect 55276 23060 55316 23155
rect 53644 23020 53695 23060
rect 53544 22868 53586 22877
rect 53544 22828 53545 22868
rect 53585 22828 53586 22868
rect 53544 22819 53586 22828
rect 53068 22744 53204 22784
rect 52875 22196 52917 22205
rect 52875 22156 52876 22196
rect 52916 22156 52917 22196
rect 52875 22147 52917 22156
rect 52724 21568 52820 21608
rect 52684 21559 52724 21568
rect 52300 20609 52340 21559
rect 52299 20600 52341 20609
rect 52299 20560 52300 20600
rect 52340 20560 52341 20600
rect 52299 20551 52341 20560
rect 52588 20525 52628 21559
rect 52683 21020 52725 21029
rect 52683 20980 52684 21020
rect 52724 20980 52725 21020
rect 52683 20971 52725 20980
rect 52684 20886 52724 20971
rect 52587 20516 52629 20525
rect 52587 20476 52588 20516
rect 52628 20476 52629 20516
rect 52587 20467 52629 20476
rect 52012 18460 52148 18500
rect 52300 18584 52340 18593
rect 51724 18332 51764 18341
rect 51764 18292 51860 18332
rect 51724 18283 51764 18292
rect 51627 17240 51669 17249
rect 51627 17200 51628 17240
rect 51668 17200 51669 17240
rect 51627 17191 51669 17200
rect 51723 17156 51765 17165
rect 51723 17116 51724 17156
rect 51764 17116 51765 17156
rect 51723 17107 51765 17116
rect 51627 17072 51669 17081
rect 51627 17032 51628 17072
rect 51668 17032 51669 17072
rect 51627 17023 51669 17032
rect 51628 16938 51668 17023
rect 51724 17022 51764 17107
rect 51820 17072 51860 18292
rect 51915 17744 51957 17753
rect 51915 17704 51916 17744
rect 51956 17704 51957 17744
rect 51915 17695 51957 17704
rect 51627 16568 51669 16577
rect 51627 16528 51628 16568
rect 51668 16528 51669 16568
rect 51627 16519 51669 16528
rect 51531 16232 51573 16241
rect 51531 16192 51532 16232
rect 51572 16192 51573 16232
rect 51531 16183 51573 16192
rect 51628 16232 51668 16519
rect 51723 16400 51765 16409
rect 51723 16360 51724 16400
rect 51764 16360 51765 16400
rect 51820 16400 51860 17032
rect 51916 16745 51956 17695
rect 51915 16736 51957 16745
rect 51915 16696 51916 16736
rect 51956 16696 51957 16736
rect 51915 16687 51957 16696
rect 51820 16360 51956 16400
rect 51723 16351 51765 16360
rect 51628 16183 51668 16192
rect 51724 16232 51764 16351
rect 51724 16183 51764 16192
rect 51819 16232 51861 16241
rect 51819 16192 51820 16232
rect 51860 16192 51861 16232
rect 51819 16183 51861 16192
rect 51820 16098 51860 16183
rect 51532 16064 51572 16073
rect 51436 16024 51532 16064
rect 51339 15896 51381 15905
rect 51339 15856 51340 15896
rect 51380 15856 51381 15896
rect 51339 15847 51381 15856
rect 51052 15426 51092 15511
rect 51244 15401 51284 15520
rect 51243 15392 51285 15401
rect 51243 15352 51244 15392
rect 51284 15352 51285 15392
rect 51243 15343 51285 15352
rect 51052 15308 51092 15317
rect 51052 14048 51092 15268
rect 51148 14720 51188 14729
rect 51188 14680 51380 14720
rect 51148 14671 51188 14680
rect 51243 14216 51285 14225
rect 51243 14176 51244 14216
rect 51284 14176 51285 14216
rect 51243 14167 51285 14176
rect 51148 14048 51188 14057
rect 51052 14008 51148 14048
rect 51148 13999 51188 14008
rect 51244 14048 51284 14167
rect 51244 13999 51284 14008
rect 51340 13922 51380 14680
rect 51436 14048 51476 16024
rect 51532 16015 51572 16024
rect 51819 15896 51861 15905
rect 51819 15856 51820 15896
rect 51860 15856 51861 15896
rect 51819 15847 51861 15856
rect 51724 15560 51764 15569
rect 51724 14309 51764 15520
rect 51723 14300 51765 14309
rect 51723 14260 51724 14300
rect 51764 14260 51765 14300
rect 51723 14251 51765 14260
rect 51436 13999 51476 14008
rect 51340 13882 51668 13922
rect 51628 13880 51668 13882
rect 51628 13831 51668 13840
rect 51436 13796 51476 13807
rect 51436 13721 51476 13756
rect 51435 13712 51477 13721
rect 51435 13672 51436 13712
rect 51476 13672 51477 13712
rect 51435 13663 51477 13672
rect 50955 13628 50997 13637
rect 50955 13588 50956 13628
rect 50996 13588 50997 13628
rect 50955 13579 50997 13588
rect 50859 13292 50901 13301
rect 50859 13252 50860 13292
rect 50900 13252 50901 13292
rect 50859 13243 50901 13252
rect 50956 12980 50996 13579
rect 51627 13460 51669 13469
rect 51627 13420 51628 13460
rect 51668 13420 51669 13460
rect 51627 13411 51669 13420
rect 51628 13326 51668 13411
rect 51628 13040 51668 13049
rect 50956 12940 51188 12980
rect 51148 12452 51188 12940
rect 51243 12956 51285 12965
rect 51243 12916 51244 12956
rect 51284 12916 51285 12956
rect 51243 12907 51285 12916
rect 51148 12403 51188 12412
rect 50956 12284 50996 12293
rect 51244 12284 51284 12907
rect 51628 12629 51668 13000
rect 51627 12620 51669 12629
rect 51627 12580 51628 12620
rect 51668 12580 51669 12620
rect 51627 12571 51669 12580
rect 51628 12452 51668 12461
rect 51820 12452 51860 15847
rect 51916 14552 51956 16360
rect 52012 16247 52052 18460
rect 52300 17501 52340 18544
rect 52684 18584 52724 18593
rect 52724 18544 52820 18584
rect 52684 18535 52724 18544
rect 52396 18332 52436 18341
rect 52299 17492 52341 17501
rect 52299 17452 52300 17492
rect 52340 17452 52341 17492
rect 52299 17443 52341 17452
rect 52299 17156 52341 17165
rect 52299 17116 52300 17156
rect 52340 17116 52341 17156
rect 52299 17107 52341 17116
rect 52300 17072 52340 17107
rect 52396 17081 52436 18292
rect 52588 18332 52628 18341
rect 52491 17408 52533 17417
rect 52491 17368 52492 17408
rect 52532 17368 52533 17408
rect 52491 17359 52533 17368
rect 52300 17021 52340 17032
rect 52395 17072 52437 17081
rect 52395 17032 52396 17072
rect 52436 17032 52437 17072
rect 52395 17023 52437 17032
rect 52492 16997 52532 17359
rect 52588 17333 52628 18292
rect 52684 17576 52724 17585
rect 52684 17417 52724 17536
rect 52683 17408 52725 17417
rect 52683 17368 52684 17408
rect 52724 17368 52725 17408
rect 52683 17359 52725 17368
rect 52587 17324 52629 17333
rect 52587 17284 52588 17324
rect 52628 17284 52629 17324
rect 52587 17275 52629 17284
rect 52780 17249 52820 18544
rect 52684 17240 52724 17249
rect 52779 17240 52821 17249
rect 52724 17200 52780 17240
rect 52820 17200 52821 17240
rect 52684 17191 52724 17200
rect 52779 17191 52821 17200
rect 52587 17156 52629 17165
rect 52587 17116 52588 17156
rect 52628 17116 52629 17156
rect 52587 17107 52629 17116
rect 52588 17072 52628 17107
rect 52780 17106 52820 17191
rect 52876 17165 52916 22147
rect 53068 17669 53108 22744
rect 53545 22596 53585 22819
rect 53655 22596 53695 23020
rect 54054 23036 54096 23045
rect 54054 22996 54055 23036
rect 54095 22996 54096 23036
rect 54316 23020 54385 23060
rect 54700 23020 54785 23060
rect 54892 23020 55185 23060
rect 54054 22987 54096 22996
rect 53944 22784 53986 22793
rect 53944 22744 53945 22784
rect 53985 22744 53986 22784
rect 53944 22735 53986 22744
rect 53945 22596 53985 22735
rect 54055 22596 54095 22987
rect 54345 22596 54385 23020
rect 54454 22952 54496 22961
rect 54454 22912 54455 22952
rect 54495 22912 54496 22952
rect 54454 22903 54496 22912
rect 54455 22596 54495 22903
rect 54745 22596 54785 23020
rect 54854 22784 54896 22793
rect 54854 22744 54855 22784
rect 54895 22744 54896 22784
rect 54854 22735 54896 22744
rect 54855 22596 54895 22735
rect 55145 22596 55185 23020
rect 55255 23020 55316 23060
rect 55255 22596 55295 23020
rect 55468 22784 55508 23584
rect 55564 23060 55604 23752
rect 55660 23743 55700 23752
rect 55852 23792 55892 23911
rect 55852 23743 55892 23752
rect 56140 23792 56180 23801
rect 56044 23624 56084 23633
rect 55948 23584 56044 23624
rect 55948 23060 55988 23584
rect 56044 23575 56084 23584
rect 56043 23372 56085 23381
rect 56140 23372 56180 23752
rect 56428 23792 56468 23801
rect 56043 23332 56044 23372
rect 56084 23332 56180 23372
rect 56332 23624 56372 23633
rect 56043 23323 56085 23332
rect 56044 23060 56084 23323
rect 55564 23020 55695 23060
rect 55468 22744 55585 22784
rect 55545 22596 55585 22744
rect 55655 22596 55695 23020
rect 55945 23020 55988 23060
rect 55945 22596 55985 23020
rect 56041 22996 56084 23060
rect 56332 23060 56372 23584
rect 56428 23297 56468 23752
rect 56620 23792 56660 23801
rect 56620 23465 56660 23752
rect 56908 23792 56948 23801
rect 56716 23624 56756 23633
rect 56619 23456 56661 23465
rect 56619 23416 56620 23456
rect 56660 23416 56661 23456
rect 56619 23407 56661 23416
rect 56427 23288 56469 23297
rect 56427 23248 56428 23288
rect 56468 23248 56469 23288
rect 56427 23239 56469 23248
rect 56428 23060 56468 23239
rect 56332 23020 56385 23060
rect 56428 23020 56495 23060
rect 56044 22784 56084 22996
rect 56044 22744 56095 22784
rect 56055 22596 56095 22744
rect 56345 22596 56385 23020
rect 56455 22596 56495 23020
rect 56716 22784 56756 23584
rect 56811 23456 56853 23465
rect 56811 23416 56812 23456
rect 56852 23416 56853 23456
rect 56811 23407 56853 23416
rect 56812 23060 56852 23407
rect 56908 23213 56948 23752
rect 57292 23792 57332 23801
rect 57004 23624 57044 23633
rect 56907 23204 56949 23213
rect 56907 23164 56908 23204
rect 56948 23164 56949 23204
rect 56907 23155 56949 23164
rect 57004 23060 57044 23584
rect 57292 23549 57332 23752
rect 57676 23792 57716 24331
rect 57388 23624 57428 23633
rect 57291 23540 57333 23549
rect 57291 23500 57292 23540
rect 57332 23500 57333 23540
rect 57291 23491 57333 23500
rect 57195 23204 57237 23213
rect 57195 23164 57196 23204
rect 57236 23164 57237 23204
rect 57195 23155 57237 23164
rect 57196 23060 57236 23155
rect 57388 23060 57428 23584
rect 57579 23540 57621 23549
rect 57579 23500 57580 23540
rect 57620 23500 57621 23540
rect 57579 23491 57621 23500
rect 57580 23204 57620 23491
rect 57676 23465 57716 23752
rect 57772 23624 57812 23633
rect 57675 23456 57717 23465
rect 57675 23416 57676 23456
rect 57716 23416 57717 23456
rect 57675 23407 57717 23416
rect 57580 23164 57716 23204
rect 57676 23060 57716 23164
rect 56812 23020 56895 23060
rect 57004 23020 57140 23060
rect 57196 23020 57295 23060
rect 57388 23020 57585 23060
rect 56716 22744 56785 22784
rect 56745 22596 56785 22744
rect 56855 22596 56895 23020
rect 57100 22784 57140 23020
rect 57100 22744 57185 22784
rect 57145 22596 57185 22744
rect 57255 22596 57295 23020
rect 57545 22596 57585 23020
rect 57655 23020 57716 23060
rect 57772 23060 57812 23584
rect 57964 23549 58004 27271
rect 58155 27068 58197 27077
rect 58155 27028 58156 27068
rect 58196 27028 58197 27068
rect 58155 27019 58197 27028
rect 58059 25136 58101 25145
rect 58059 25096 58060 25136
rect 58100 25096 58101 25136
rect 58059 25087 58101 25096
rect 58060 24725 58100 25087
rect 58059 24716 58101 24725
rect 58059 24676 58060 24716
rect 58100 24676 58101 24716
rect 58059 24667 58101 24676
rect 58060 24632 58100 24667
rect 58060 24582 58100 24592
rect 58156 24632 58196 27019
rect 58251 26984 58293 26993
rect 58251 26944 58252 26984
rect 58292 26944 58293 26984
rect 58251 26935 58293 26944
rect 58252 26900 58292 26935
rect 58252 26849 58292 26860
rect 58348 26312 58388 27616
rect 58443 27068 58485 27077
rect 58443 27028 58444 27068
rect 58484 27028 58485 27068
rect 58443 27019 58485 27028
rect 58444 26934 58484 27019
rect 58827 26816 58869 26825
rect 58827 26776 58828 26816
rect 58868 26776 58869 26816
rect 58827 26767 58869 26776
rect 58828 26648 58868 26767
rect 58348 26272 58484 26312
rect 58348 26144 58388 26153
rect 58252 26104 58348 26144
rect 58252 24800 58292 26104
rect 58348 26095 58388 26104
rect 58347 25976 58389 25985
rect 58347 25936 58348 25976
rect 58388 25936 58389 25976
rect 58347 25927 58389 25936
rect 58348 25842 58388 25927
rect 58444 25304 58484 26272
rect 58539 26144 58581 26153
rect 58539 26104 58540 26144
rect 58580 26104 58581 26144
rect 58539 26095 58581 26104
rect 58636 26144 58676 26153
rect 58540 26010 58580 26095
rect 58636 25976 58676 26104
rect 58828 26144 58868 26608
rect 58924 26489 58964 29884
rect 59020 29875 59060 29884
rect 59116 29756 59156 30052
rect 59020 29716 59156 29756
rect 59020 28748 59060 29716
rect 59212 29672 59252 29681
rect 59116 29632 59212 29672
rect 59116 29261 59156 29632
rect 59212 29623 59252 29632
rect 59308 29504 59348 31723
rect 59404 31613 59444 32152
rect 59596 32192 59636 34159
rect 59691 33704 59733 33713
rect 59691 33664 59692 33704
rect 59732 33664 59733 33704
rect 59691 33655 59733 33664
rect 59596 32143 59636 32152
rect 59692 32192 59732 33655
rect 59788 32864 59828 32873
rect 59788 32285 59828 32824
rect 59787 32276 59829 32285
rect 59787 32236 59788 32276
rect 59828 32236 59829 32276
rect 59787 32227 59829 32236
rect 59403 31604 59445 31613
rect 59403 31564 59404 31604
rect 59444 31564 59445 31604
rect 59403 31555 59445 31564
rect 59692 31520 59732 32152
rect 59884 32192 59924 35008
rect 60363 34208 60405 34217
rect 60363 34168 60364 34208
rect 60404 34168 60405 34208
rect 60363 34159 60405 34168
rect 59979 34124 60021 34133
rect 59979 34084 59980 34124
rect 60020 34084 60021 34124
rect 59979 34075 60021 34084
rect 59980 33545 60020 34075
rect 60364 34074 60404 34159
rect 60267 33788 60309 33797
rect 60267 33748 60268 33788
rect 60308 33748 60309 33788
rect 60267 33739 60309 33748
rect 59979 33536 60021 33545
rect 59979 33496 59980 33536
rect 60020 33496 60021 33536
rect 59979 33487 60021 33496
rect 59884 32108 59924 32152
rect 59813 32068 59924 32108
rect 59813 32024 59853 32068
rect 59788 31984 59853 32024
rect 59788 31781 59828 31984
rect 59883 31940 59925 31949
rect 59883 31900 59884 31940
rect 59924 31900 59925 31940
rect 59883 31891 59925 31900
rect 59884 31806 59924 31891
rect 59787 31772 59829 31781
rect 59787 31732 59788 31772
rect 59828 31732 59829 31772
rect 59787 31723 59829 31732
rect 59500 31480 59732 31520
rect 59500 30596 59540 31480
rect 59596 31352 59636 31361
rect 59596 30857 59636 31312
rect 59692 31352 59732 31361
rect 59692 31109 59732 31312
rect 59787 31352 59829 31361
rect 59787 31312 59788 31352
rect 59828 31312 59829 31352
rect 59787 31303 59829 31312
rect 59788 31218 59828 31303
rect 59883 31184 59925 31193
rect 59883 31144 59884 31184
rect 59924 31144 59925 31184
rect 59883 31135 59925 31144
rect 59691 31100 59733 31109
rect 59691 31060 59692 31100
rect 59732 31060 59733 31100
rect 59691 31051 59733 31060
rect 59884 31050 59924 31135
rect 59595 30848 59637 30857
rect 59980 30848 60020 33487
rect 60268 31604 60308 33739
rect 60460 33713 60500 37192
rect 60556 36737 60596 37276
rect 61131 37276 61132 37316
rect 61172 37276 61173 37316
rect 61131 37267 61173 37276
rect 62283 37316 62325 37325
rect 62283 37276 62284 37316
rect 62324 37276 62325 37316
rect 62283 37267 62325 37276
rect 61803 36980 61845 36989
rect 61803 36940 61804 36980
rect 61844 36940 61845 36980
rect 61803 36931 61845 36940
rect 61131 36896 61173 36905
rect 61131 36856 61132 36896
rect 61172 36856 61173 36896
rect 61131 36847 61173 36856
rect 60555 36728 60597 36737
rect 60555 36688 60556 36728
rect 60596 36688 60597 36728
rect 60555 36679 60597 36688
rect 61132 35216 61172 36847
rect 61707 36728 61749 36737
rect 61707 36688 61708 36728
rect 61748 36688 61749 36728
rect 61707 36679 61749 36688
rect 61804 36728 61844 36931
rect 62284 36896 62324 37267
rect 62380 36905 62420 37351
rect 62284 36847 62324 36856
rect 62379 36896 62421 36905
rect 62379 36856 62380 36896
rect 62420 36856 62421 36896
rect 62379 36847 62421 36856
rect 61708 36594 61748 36679
rect 61516 36476 61556 36485
rect 61516 35729 61556 36436
rect 61515 35720 61557 35729
rect 61515 35680 61516 35720
rect 61556 35680 61557 35720
rect 61515 35671 61557 35680
rect 61132 35167 61172 35176
rect 61804 35132 61844 36688
rect 61900 36728 61940 36737
rect 61900 35981 61940 36688
rect 61996 36728 62036 36737
rect 62188 36728 62228 36737
rect 62036 36688 62188 36728
rect 61996 36679 62036 36688
rect 62188 36679 62228 36688
rect 62379 36728 62421 36737
rect 62379 36688 62380 36728
rect 62420 36688 62421 36728
rect 62379 36679 62421 36688
rect 62476 36728 62516 36737
rect 62380 36594 62420 36679
rect 62284 36140 62324 36149
rect 62476 36140 62516 36688
rect 62324 36100 62516 36140
rect 62284 36091 62324 36100
rect 62572 36056 62612 37939
rect 62380 36016 62612 36056
rect 61899 35972 61941 35981
rect 61899 35932 61900 35972
rect 61940 35932 61941 35972
rect 61899 35923 61941 35932
rect 61708 35092 61844 35132
rect 61611 35048 61653 35057
rect 61611 35008 61612 35048
rect 61652 35008 61653 35048
rect 61611 34999 61653 35008
rect 61515 34376 61557 34385
rect 61515 34336 61516 34376
rect 61556 34336 61557 34376
rect 61515 34327 61557 34336
rect 61612 34376 61652 34999
rect 61708 34721 61748 35092
rect 61900 35057 61940 35923
rect 61996 35888 62036 35897
rect 61899 35048 61941 35057
rect 61899 35008 61900 35048
rect 61940 35008 61941 35048
rect 61899 34999 61941 35008
rect 61996 34973 62036 35848
rect 62092 35888 62132 35897
rect 62284 35888 62324 35897
rect 61803 34964 61845 34973
rect 61803 34924 61804 34964
rect 61844 34924 61845 34964
rect 61803 34915 61845 34924
rect 61995 34964 62037 34973
rect 61995 34924 61996 34964
rect 62036 34924 62037 34964
rect 61995 34915 62037 34924
rect 61707 34712 61749 34721
rect 61707 34672 61708 34712
rect 61748 34672 61749 34712
rect 61707 34663 61749 34672
rect 61516 34242 61556 34327
rect 61612 33965 61652 34336
rect 61708 34376 61748 34663
rect 61611 33956 61653 33965
rect 61611 33916 61612 33956
rect 61652 33916 61653 33956
rect 61611 33907 61653 33916
rect 60459 33704 60501 33713
rect 60459 33664 60460 33704
rect 60500 33664 60501 33704
rect 60459 33655 60501 33664
rect 61612 33140 61652 33907
rect 61708 33797 61748 34336
rect 61804 34376 61844 34915
rect 62092 34796 62132 35848
rect 61804 34327 61844 34336
rect 61900 34756 62132 34796
rect 62188 35848 62284 35888
rect 61707 33788 61749 33797
rect 61707 33748 61708 33788
rect 61748 33748 61749 33788
rect 61707 33739 61749 33748
rect 61900 33713 61940 34756
rect 61996 34553 62036 34638
rect 62188 34628 62228 35848
rect 62284 35839 62324 35848
rect 62283 34964 62325 34973
rect 62283 34924 62284 34964
rect 62324 34924 62325 34964
rect 62283 34915 62325 34924
rect 62284 34830 62324 34915
rect 62092 34588 62228 34628
rect 61995 34544 62037 34553
rect 61995 34504 61996 34544
rect 62036 34504 62037 34544
rect 61995 34495 62037 34504
rect 61995 34376 62037 34385
rect 61995 34336 61996 34376
rect 62036 34336 62037 34376
rect 61995 34327 62037 34336
rect 61996 34242 62036 34327
rect 62092 34124 62132 34588
rect 62187 34376 62229 34385
rect 62187 34336 62188 34376
rect 62228 34336 62229 34376
rect 62187 34327 62229 34336
rect 62284 34376 62324 34385
rect 62188 34242 62228 34327
rect 62187 34124 62229 34133
rect 62092 34084 62188 34124
rect 62228 34084 62229 34124
rect 62187 34075 62229 34084
rect 61995 34040 62037 34049
rect 61995 34000 61996 34040
rect 62036 34000 62037 34040
rect 61995 33991 62037 34000
rect 61899 33704 61941 33713
rect 61899 33664 61900 33704
rect 61940 33664 61941 33704
rect 61899 33655 61941 33664
rect 61996 33536 62036 33991
rect 62188 33704 62228 34075
rect 62284 33872 62324 34336
rect 62380 34049 62420 36016
rect 62476 34964 62516 34973
rect 62516 34924 62612 34964
rect 62476 34915 62516 34924
rect 62379 34040 62421 34049
rect 62379 34000 62380 34040
rect 62420 34000 62421 34040
rect 62379 33991 62421 34000
rect 62284 33823 62324 33832
rect 62188 33655 62228 33664
rect 62379 33704 62421 33713
rect 62379 33664 62380 33704
rect 62420 33664 62421 33704
rect 62379 33655 62421 33664
rect 62476 33704 62516 33713
rect 62572 33704 62612 34924
rect 62668 34376 62708 38116
rect 63436 37400 63476 38284
rect 63532 38240 63572 38249
rect 63532 37988 63572 38200
rect 63628 38240 63668 38249
rect 67467 38240 67509 38249
rect 63668 38200 64340 38240
rect 63628 38191 63668 38200
rect 64204 38072 64244 38081
rect 63532 37948 64052 37988
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 63724 37400 63764 37409
rect 63436 37360 63724 37400
rect 63724 37351 63764 37360
rect 63532 37232 63572 37241
rect 63340 37192 63532 37232
rect 63340 36821 63380 37192
rect 63532 37183 63572 37192
rect 64012 37148 64052 37948
rect 64108 37400 64148 37409
rect 64204 37400 64244 38032
rect 64148 37360 64244 37400
rect 64108 37351 64148 37360
rect 63916 37108 64052 37148
rect 63916 36821 63956 37108
rect 63339 36812 63381 36821
rect 63339 36772 63340 36812
rect 63380 36772 63381 36812
rect 63339 36763 63381 36772
rect 63915 36812 63957 36821
rect 63915 36772 63916 36812
rect 63956 36772 63957 36812
rect 63915 36763 63957 36772
rect 64300 36812 64340 38200
rect 67467 38200 67468 38240
rect 67508 38200 67509 38240
rect 67467 38191 67509 38200
rect 67660 38240 67700 38249
rect 67083 38156 67125 38165
rect 67083 38116 67084 38156
rect 67124 38116 67125 38156
rect 67083 38107 67125 38116
rect 66508 38072 66548 38081
rect 66548 38032 66740 38072
rect 66508 38023 66548 38032
rect 66315 37988 66357 37997
rect 66315 37948 66316 37988
rect 66356 37948 66357 37988
rect 66315 37939 66357 37948
rect 64971 37400 65013 37409
rect 64971 37360 64972 37400
rect 65012 37360 65013 37400
rect 64971 37351 65013 37360
rect 65643 37400 65685 37409
rect 65643 37360 65644 37400
rect 65684 37360 65685 37400
rect 65643 37351 65685 37360
rect 66316 37400 66356 37939
rect 66316 37351 66356 37360
rect 66700 37400 66740 38032
rect 67084 38022 67124 38107
rect 67468 38106 67508 38191
rect 67660 37997 67700 38200
rect 67756 38240 67796 38249
rect 67947 38240 67989 38249
rect 67796 38200 67892 38240
rect 67756 38191 67796 38200
rect 66700 37351 66740 37360
rect 67276 37988 67316 37997
rect 64972 37266 65012 37351
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 64300 36763 64340 36772
rect 62956 36728 62996 36739
rect 62956 36653 62996 36688
rect 63244 36728 63284 36737
rect 62955 36644 62997 36653
rect 62955 36604 62956 36644
rect 62996 36604 62997 36644
rect 62955 36595 62997 36604
rect 63147 36644 63189 36653
rect 63147 36604 63148 36644
rect 63188 36604 63189 36644
rect 63147 36595 63189 36604
rect 62764 35216 62804 35225
rect 62764 34973 62804 35176
rect 62859 35216 62901 35225
rect 62859 35176 62860 35216
rect 62900 35176 62901 35216
rect 62859 35167 62901 35176
rect 63148 35216 63188 36595
rect 63244 36485 63284 36688
rect 63340 36678 63380 36763
rect 63820 36728 63860 36737
rect 63628 36560 63668 36569
rect 63820 36560 63860 36688
rect 63916 36678 63956 36763
rect 64011 36728 64053 36737
rect 64011 36688 64012 36728
rect 64052 36688 64053 36728
rect 64011 36679 64053 36688
rect 64204 36728 64244 36737
rect 64012 36594 64052 36679
rect 63668 36520 63860 36560
rect 63628 36511 63668 36520
rect 63243 36476 63285 36485
rect 63243 36436 63244 36476
rect 63284 36436 63285 36476
rect 63243 36427 63285 36436
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 62860 35082 62900 35167
rect 62763 34964 62805 34973
rect 62763 34924 62764 34964
rect 62804 34924 62805 34964
rect 62763 34915 62805 34924
rect 63148 34637 63188 35176
rect 63628 35048 63668 35057
rect 63436 35008 63628 35048
rect 63147 34628 63189 34637
rect 63147 34588 63148 34628
rect 63188 34588 63189 34628
rect 63147 34579 63189 34588
rect 62860 34385 62900 34470
rect 62956 34420 63284 34460
rect 62668 33881 62708 34336
rect 62859 34376 62901 34385
rect 62859 34336 62860 34376
rect 62900 34336 62901 34376
rect 62859 34327 62901 34336
rect 62956 34376 62996 34420
rect 62956 34327 62996 34336
rect 62763 34292 62805 34301
rect 62763 34252 62764 34292
rect 62804 34252 62805 34292
rect 62763 34243 62805 34252
rect 62764 34158 62804 34243
rect 62860 34040 62900 34327
rect 63147 34292 63189 34301
rect 63147 34252 63148 34292
rect 63188 34252 63189 34292
rect 63147 34243 63189 34252
rect 63148 34158 63188 34243
rect 62764 34000 62900 34040
rect 62667 33872 62709 33881
rect 62667 33832 62668 33872
rect 62708 33832 62709 33872
rect 62667 33823 62709 33832
rect 62764 33788 62804 34000
rect 63244 33872 63284 34420
rect 63436 34376 63476 35008
rect 63628 34999 63668 35008
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 64011 34628 64053 34637
rect 64011 34588 64012 34628
rect 64052 34588 64053 34628
rect 64011 34579 64053 34588
rect 63532 34376 63572 34385
rect 63436 34336 63532 34376
rect 63532 34327 63572 34336
rect 62764 33739 62804 33748
rect 63148 33832 63284 33872
rect 63148 33788 63188 33832
rect 63148 33739 63188 33748
rect 62668 33704 62708 33713
rect 62572 33664 62668 33704
rect 62380 33570 62420 33655
rect 61900 33496 62036 33536
rect 60939 33116 60981 33125
rect 60939 33076 60940 33116
rect 60980 33076 60981 33116
rect 61612 33100 61844 33140
rect 60939 33067 60981 33076
rect 60940 32982 60980 33067
rect 61132 33032 61172 33041
rect 60940 32696 60980 32705
rect 60940 32453 60980 32656
rect 60939 32444 60981 32453
rect 60939 32404 60940 32444
rect 60980 32404 60981 32444
rect 60939 32395 60981 32404
rect 60268 31555 60308 31564
rect 60364 32192 60404 32201
rect 60075 31520 60117 31529
rect 60075 31480 60076 31520
rect 60116 31480 60117 31520
rect 60075 31471 60117 31480
rect 60076 31436 60116 31471
rect 60076 31385 60116 31396
rect 60364 31277 60404 32152
rect 60748 32192 60788 32201
rect 61132 32192 61172 32992
rect 61323 32780 61365 32789
rect 61323 32740 61324 32780
rect 61364 32740 61365 32780
rect 61323 32731 61365 32740
rect 60788 32152 61172 32192
rect 60748 32143 60788 32152
rect 60747 31940 60789 31949
rect 60747 31900 60748 31940
rect 60788 31900 60789 31940
rect 60747 31891 60789 31900
rect 60651 31436 60693 31445
rect 60651 31396 60652 31436
rect 60692 31396 60693 31436
rect 60651 31387 60693 31396
rect 60363 31268 60405 31277
rect 60363 31228 60364 31268
rect 60404 31228 60405 31268
rect 60363 31219 60405 31228
rect 60268 31184 60308 31193
rect 60268 31109 60308 31144
rect 60555 31184 60597 31193
rect 60555 31144 60556 31184
rect 60596 31144 60597 31184
rect 60555 31135 60597 31144
rect 60267 31100 60309 31109
rect 60267 31060 60268 31100
rect 60308 31060 60309 31100
rect 60267 31051 60309 31060
rect 59595 30808 59596 30848
rect 59636 30808 59637 30848
rect 59595 30799 59637 30808
rect 59884 30808 60020 30848
rect 60075 30848 60117 30857
rect 60075 30808 60076 30848
rect 60116 30808 60117 30848
rect 59595 30596 59637 30605
rect 59500 30556 59596 30596
rect 59636 30556 59637 30596
rect 59595 30547 59637 30556
rect 59404 29924 59444 29933
rect 59404 29513 59444 29884
rect 59212 29464 59348 29504
rect 59403 29504 59445 29513
rect 59403 29464 59404 29504
rect 59444 29464 59445 29504
rect 59115 29252 59157 29261
rect 59115 29212 59116 29252
rect 59156 29212 59157 29252
rect 59115 29203 59157 29212
rect 59116 29084 59156 29203
rect 59212 29168 59252 29464
rect 59403 29455 59445 29464
rect 59308 29336 59348 29345
rect 59596 29336 59636 30547
rect 59691 29924 59733 29933
rect 59691 29884 59692 29924
rect 59732 29884 59733 29924
rect 59691 29875 59733 29884
rect 59692 29840 59732 29875
rect 59692 29789 59732 29800
rect 59884 29345 59924 30808
rect 60075 30799 60117 30808
rect 59979 30680 60021 30689
rect 59979 30640 59980 30680
rect 60020 30640 60021 30680
rect 59979 30631 60021 30640
rect 59980 30546 60020 30631
rect 59979 30092 60021 30101
rect 59979 30052 59980 30092
rect 60020 30052 60021 30092
rect 59979 30043 60021 30052
rect 59980 29840 60020 30043
rect 59980 29791 60020 29800
rect 60076 29840 60116 30799
rect 60268 30605 60308 31051
rect 60364 30680 60404 30689
rect 60267 30596 60309 30605
rect 60267 30556 60268 30596
rect 60308 30556 60309 30596
rect 60267 30547 60309 30556
rect 60364 30512 60404 30640
rect 60556 30680 60596 31135
rect 60556 30631 60596 30640
rect 60556 30512 60596 30521
rect 60364 30472 60556 30512
rect 60556 30463 60596 30472
rect 60267 30428 60309 30437
rect 60267 30388 60268 30428
rect 60308 30388 60309 30428
rect 60267 30379 60309 30388
rect 59883 29336 59925 29345
rect 59348 29296 59732 29336
rect 59308 29287 59348 29296
rect 59500 29168 59540 29177
rect 59212 29128 59500 29168
rect 59116 29035 59156 29044
rect 59020 28708 59156 28748
rect 59019 28580 59061 28589
rect 59019 28540 59020 28580
rect 59060 28540 59061 28580
rect 59019 28531 59061 28540
rect 59020 28446 59060 28531
rect 59020 28160 59060 28169
rect 59020 26900 59060 28120
rect 59116 26909 59156 28708
rect 59404 28589 59444 29128
rect 59500 29119 59540 29128
rect 59692 29168 59732 29296
rect 59883 29296 59884 29336
rect 59924 29296 59925 29336
rect 59883 29287 59925 29296
rect 59692 29119 59732 29128
rect 59788 29168 59828 29177
rect 60076 29168 60116 29800
rect 60171 29504 60213 29513
rect 60171 29464 60172 29504
rect 60212 29464 60213 29504
rect 60171 29455 60213 29464
rect 59828 29128 60116 29168
rect 59788 29119 59828 29128
rect 59500 28916 59540 28925
rect 59403 28580 59445 28589
rect 59403 28540 59404 28580
rect 59444 28540 59445 28580
rect 59403 28531 59445 28540
rect 59212 28328 59252 28337
rect 59212 27833 59252 28288
rect 59404 28328 59444 28337
rect 59307 28160 59349 28169
rect 59307 28120 59308 28160
rect 59348 28120 59349 28160
rect 59404 28160 59444 28288
rect 59500 28328 59540 28876
rect 60172 28580 60212 29455
rect 60268 29168 60308 30379
rect 60363 30008 60405 30017
rect 60363 29968 60364 30008
rect 60404 29968 60405 30008
rect 60363 29959 60405 29968
rect 60364 29874 60404 29959
rect 60556 29756 60596 29765
rect 60460 29336 60500 29345
rect 60556 29336 60596 29716
rect 60500 29296 60596 29336
rect 60460 29287 60500 29296
rect 60268 29119 60308 29128
rect 60363 29168 60405 29177
rect 60363 29128 60364 29168
rect 60404 29128 60405 29168
rect 60363 29119 60405 29128
rect 60556 29168 60596 29179
rect 60364 29034 60404 29119
rect 60556 29093 60596 29128
rect 60555 29084 60597 29093
rect 60555 29044 60556 29084
rect 60596 29044 60597 29084
rect 60555 29035 60597 29044
rect 60172 28540 60596 28580
rect 59788 28496 59828 28505
rect 59500 28279 59540 28288
rect 59596 28456 59788 28496
rect 59828 28456 60308 28496
rect 59596 28160 59636 28456
rect 59788 28447 59828 28456
rect 59404 28120 59636 28160
rect 59692 28328 59732 28337
rect 59307 28111 59349 28120
rect 59308 28026 59348 28111
rect 59692 27992 59732 28288
rect 59883 28328 59925 28337
rect 59883 28288 59884 28328
rect 59924 28288 59925 28328
rect 59883 28279 59925 28288
rect 60076 28328 60116 28337
rect 59404 27952 59732 27992
rect 59211 27824 59253 27833
rect 59211 27784 59212 27824
rect 59252 27784 59253 27824
rect 59211 27775 59253 27784
rect 59307 27656 59349 27665
rect 59307 27616 59308 27656
rect 59348 27616 59349 27656
rect 59307 27607 59349 27616
rect 59020 26851 59060 26860
rect 59115 26900 59157 26909
rect 59115 26860 59116 26900
rect 59156 26860 59157 26900
rect 59115 26851 59157 26860
rect 59308 26816 59348 27607
rect 59404 27068 59444 27952
rect 59884 27833 59924 28279
rect 59691 27824 59733 27833
rect 59691 27784 59692 27824
rect 59732 27784 59733 27824
rect 59691 27775 59733 27784
rect 59883 27824 59925 27833
rect 59883 27784 59884 27824
rect 59924 27784 59925 27824
rect 59883 27775 59925 27784
rect 59692 27690 59732 27775
rect 59788 27656 59828 27667
rect 59788 27581 59828 27616
rect 59884 27656 59924 27665
rect 59787 27572 59829 27581
rect 59787 27532 59788 27572
rect 59828 27532 59829 27572
rect 59787 27523 59829 27532
rect 59499 27404 59541 27413
rect 59499 27364 59500 27404
rect 59540 27364 59541 27404
rect 59499 27355 59541 27364
rect 59404 27019 59444 27028
rect 59308 26776 59444 26816
rect 59115 26648 59157 26657
rect 59115 26608 59116 26648
rect 59156 26608 59157 26648
rect 59115 26599 59157 26608
rect 58923 26480 58965 26489
rect 58923 26440 58924 26480
rect 58964 26440 58965 26480
rect 58923 26431 58965 26440
rect 58828 26095 58868 26104
rect 58828 25976 58868 25985
rect 58636 25936 58828 25976
rect 58828 25927 58868 25936
rect 58924 25817 58964 26431
rect 59019 26312 59061 26321
rect 59019 26272 59020 26312
rect 59060 26272 59061 26312
rect 59019 26263 59061 26272
rect 59020 26144 59060 26263
rect 59020 26095 59060 26104
rect 59116 26144 59156 26599
rect 59307 26396 59349 26405
rect 59307 26356 59308 26396
rect 59348 26356 59349 26396
rect 59307 26347 59349 26356
rect 59116 26095 59156 26104
rect 58923 25808 58965 25817
rect 58923 25768 58924 25808
rect 58964 25768 58965 25808
rect 58923 25759 58965 25768
rect 58731 25640 58773 25649
rect 58731 25600 58732 25640
rect 58772 25600 58773 25640
rect 58731 25591 58773 25600
rect 58635 25304 58677 25313
rect 58444 25264 58636 25304
rect 58676 25264 58677 25304
rect 58635 25255 58677 25264
rect 58443 25136 58485 25145
rect 58443 25096 58444 25136
rect 58484 25096 58485 25136
rect 58443 25087 58485 25096
rect 58348 24800 58388 24809
rect 58252 24760 58348 24800
rect 58348 24751 58388 24760
rect 58156 24583 58196 24592
rect 58252 24632 58292 24641
rect 58444 24632 58484 25087
rect 58636 24641 58676 25255
rect 58292 24592 58484 24632
rect 58635 24632 58677 24641
rect 58635 24592 58636 24632
rect 58676 24592 58677 24632
rect 58252 24583 58292 24592
rect 58635 24583 58677 24592
rect 58732 24128 58772 25591
rect 58828 24548 58868 24557
rect 58924 24548 58964 25759
rect 59211 25220 59253 25229
rect 59211 25180 59212 25220
rect 59252 25180 59253 25220
rect 59211 25171 59253 25180
rect 59020 24800 59060 24809
rect 59020 24641 59060 24760
rect 59019 24632 59061 24641
rect 59019 24592 59020 24632
rect 59060 24592 59061 24632
rect 59019 24583 59061 24592
rect 58868 24508 58964 24548
rect 58828 24499 58868 24508
rect 59212 24464 59252 25171
rect 59308 24968 59348 26347
rect 59404 26144 59444 26776
rect 59500 26657 59540 27355
rect 59787 27236 59829 27245
rect 59787 27196 59788 27236
rect 59828 27196 59829 27236
rect 59787 27187 59829 27196
rect 59788 26816 59828 27187
rect 59884 27077 59924 27616
rect 59980 27656 60020 27665
rect 59980 27413 60020 27616
rect 59979 27404 60021 27413
rect 59979 27364 59980 27404
rect 60020 27364 60021 27404
rect 59979 27355 60021 27364
rect 59883 27068 59925 27077
rect 59883 27028 59884 27068
rect 59924 27028 59925 27068
rect 59883 27019 59925 27028
rect 60076 26984 60116 28288
rect 60268 28328 60308 28456
rect 60268 28279 60308 28288
rect 60363 28328 60405 28337
rect 60363 28288 60364 28328
rect 60404 28288 60405 28328
rect 60363 28279 60405 28288
rect 60556 28328 60596 28540
rect 60652 28505 60692 31387
rect 60748 31016 60788 31891
rect 60843 31604 60885 31613
rect 60843 31564 60844 31604
rect 60884 31564 60885 31604
rect 60843 31555 60885 31564
rect 60844 31470 60884 31555
rect 60844 31184 60884 31193
rect 61035 31184 61077 31193
rect 60884 31144 60980 31184
rect 60844 31135 60884 31144
rect 60748 30976 60884 31016
rect 60748 30680 60788 30689
rect 60748 30176 60788 30640
rect 60844 30680 60884 30976
rect 60844 30631 60884 30640
rect 60940 30512 60980 31144
rect 61035 31144 61036 31184
rect 61076 31144 61077 31184
rect 61035 31135 61077 31144
rect 61036 30689 61076 31135
rect 61035 30680 61077 30689
rect 61035 30640 61036 30680
rect 61076 30640 61077 30680
rect 61035 30631 61077 30640
rect 61228 30680 61268 30689
rect 60940 30472 61076 30512
rect 60939 30260 60981 30269
rect 60939 30220 60940 30260
rect 60980 30220 60981 30260
rect 60939 30211 60981 30220
rect 60748 30136 60884 30176
rect 60747 30008 60789 30017
rect 60747 29968 60748 30008
rect 60788 29968 60789 30008
rect 60747 29959 60789 29968
rect 60748 29168 60788 29959
rect 60844 29252 60884 30136
rect 60940 29840 60980 30211
rect 60940 29791 60980 29800
rect 60844 29177 60884 29212
rect 60748 29119 60788 29128
rect 60843 29168 60885 29177
rect 60843 29128 60844 29168
rect 60884 29128 60885 29168
rect 60843 29119 60885 29128
rect 60940 29168 60980 29177
rect 61036 29168 61076 30472
rect 61131 30428 61173 30437
rect 61131 30388 61132 30428
rect 61172 30388 61173 30428
rect 61131 30379 61173 30388
rect 61132 30294 61172 30379
rect 61228 30101 61268 30640
rect 61227 30092 61269 30101
rect 61227 30052 61228 30092
rect 61268 30052 61269 30092
rect 61227 30043 61269 30052
rect 61324 29420 61364 32731
rect 61804 32696 61844 33100
rect 61900 32873 61940 33496
rect 61995 33368 62037 33377
rect 61995 33328 61996 33368
rect 62036 33328 62037 33368
rect 61995 33319 62037 33328
rect 61996 33140 62036 33319
rect 62476 33140 62516 33664
rect 62668 33655 62708 33664
rect 62860 33704 62900 33713
rect 61996 33100 62228 33140
rect 62476 33100 62708 33140
rect 61899 32864 61941 32873
rect 61899 32824 61900 32864
rect 61940 32824 61941 32864
rect 61899 32815 61941 32824
rect 61804 32656 61940 32696
rect 61611 32192 61653 32201
rect 61611 32152 61612 32192
rect 61652 32152 61653 32192
rect 61611 32143 61653 32152
rect 61803 32192 61845 32201
rect 61803 32152 61804 32192
rect 61844 32152 61845 32192
rect 61803 32143 61845 32152
rect 61612 32058 61652 32143
rect 61420 30512 61460 30521
rect 61420 30269 61460 30472
rect 61419 30260 61461 30269
rect 61419 30220 61420 30260
rect 61460 30220 61461 30260
rect 61419 30211 61461 30220
rect 61804 29840 61844 32143
rect 61900 31361 61940 32656
rect 61995 32612 62037 32621
rect 61995 32572 61996 32612
rect 62036 32572 62037 32612
rect 61995 32563 62037 32572
rect 61996 31529 62036 32563
rect 61995 31520 62037 31529
rect 61995 31480 61996 31520
rect 62036 31480 62037 31520
rect 61995 31471 62037 31480
rect 61899 31352 61941 31361
rect 61899 31312 61900 31352
rect 61940 31312 61941 31352
rect 61899 31303 61941 31312
rect 61804 29791 61844 29800
rect 60980 29128 61076 29168
rect 61132 29380 61364 29420
rect 61132 29336 61172 29380
rect 60940 29119 60980 29128
rect 60844 29088 60884 29119
rect 61132 29093 61172 29296
rect 61131 29084 61173 29093
rect 61131 29044 61132 29084
rect 61172 29044 61173 29084
rect 61131 29035 61173 29044
rect 61324 29084 61364 29093
rect 61035 28832 61077 28841
rect 61035 28792 61036 28832
rect 61076 28792 61077 28832
rect 61035 28783 61077 28792
rect 60651 28496 60693 28505
rect 60651 28456 60652 28496
rect 60692 28456 60693 28496
rect 60651 28447 60693 28456
rect 60940 28412 60980 28421
rect 60364 28194 60404 28279
rect 60172 28160 60212 28169
rect 60172 27740 60212 28120
rect 60460 27740 60500 27749
rect 60172 27700 60460 27740
rect 60460 27691 60500 27700
rect 60267 27572 60309 27581
rect 60267 27532 60268 27572
rect 60308 27532 60309 27572
rect 60267 27523 60309 27532
rect 60076 26944 60212 26984
rect 59979 26900 60021 26909
rect 59979 26860 59980 26900
rect 60020 26860 60021 26900
rect 59979 26851 60021 26860
rect 59788 26767 59828 26776
rect 59692 26732 59732 26743
rect 59692 26657 59732 26692
rect 59499 26648 59541 26657
rect 59499 26608 59500 26648
rect 59540 26608 59541 26648
rect 59499 26599 59541 26608
rect 59691 26648 59733 26657
rect 59691 26608 59692 26648
rect 59732 26608 59733 26648
rect 59691 26599 59733 26608
rect 59691 26480 59733 26489
rect 59691 26440 59692 26480
rect 59732 26440 59733 26480
rect 59691 26431 59733 26440
rect 59404 25985 59444 26104
rect 59499 26144 59541 26153
rect 59499 26104 59500 26144
rect 59540 26104 59541 26144
rect 59499 26095 59541 26104
rect 59596 26144 59636 26153
rect 59500 26010 59540 26095
rect 59403 25976 59445 25985
rect 59403 25936 59404 25976
rect 59444 25936 59445 25976
rect 59403 25927 59445 25936
rect 59499 25220 59541 25229
rect 59596 25220 59636 26104
rect 59692 25229 59732 26431
rect 59788 26144 59828 26153
rect 59788 25304 59828 26104
rect 59883 26144 59925 26153
rect 59883 26104 59884 26144
rect 59924 26104 59925 26144
rect 59883 26095 59925 26104
rect 59884 26010 59924 26095
rect 59788 25264 59924 25304
rect 59499 25180 59500 25220
rect 59540 25180 59636 25220
rect 59691 25220 59733 25229
rect 59691 25180 59692 25220
rect 59732 25180 59733 25220
rect 59499 25171 59541 25180
rect 59691 25171 59733 25180
rect 59308 24928 59444 24968
rect 59307 24800 59349 24809
rect 59307 24760 59308 24800
rect 59348 24760 59349 24800
rect 59307 24751 59349 24760
rect 59212 24415 59252 24424
rect 58732 24088 58868 24128
rect 58059 23792 58101 23801
rect 58059 23752 58060 23792
rect 58100 23752 58101 23792
rect 58059 23743 58101 23752
rect 58347 23792 58389 23801
rect 58347 23752 58348 23792
rect 58388 23752 58389 23792
rect 58347 23743 58389 23752
rect 58444 23792 58484 23803
rect 58060 23658 58100 23743
rect 58156 23624 58196 23633
rect 57963 23540 58005 23549
rect 57963 23500 57964 23540
rect 58004 23500 58005 23540
rect 57963 23491 58005 23500
rect 58059 23456 58101 23465
rect 58059 23416 58060 23456
rect 58100 23416 58101 23456
rect 58059 23407 58101 23416
rect 58060 23060 58100 23407
rect 57772 23020 57985 23060
rect 57655 22596 57695 23020
rect 57945 22596 57985 23020
rect 58055 23020 58100 23060
rect 58055 22596 58095 23020
rect 58156 22784 58196 23584
rect 58348 23060 58388 23743
rect 58444 23717 58484 23752
rect 58828 23792 58868 24088
rect 59308 23792 59348 24751
rect 59404 24380 59444 24928
rect 59595 24800 59637 24809
rect 59595 24760 59596 24800
rect 59636 24760 59637 24800
rect 59595 24751 59637 24760
rect 59499 24716 59541 24725
rect 59499 24676 59500 24716
rect 59540 24676 59541 24716
rect 59499 24667 59541 24676
rect 59500 24582 59540 24667
rect 59596 24632 59636 24751
rect 59692 24641 59732 25171
rect 59788 25136 59828 25145
rect 59788 24725 59828 25096
rect 59884 24977 59924 25264
rect 59883 24968 59925 24977
rect 59883 24928 59884 24968
rect 59924 24928 59925 24968
rect 59883 24919 59925 24928
rect 59787 24716 59829 24725
rect 59787 24676 59788 24716
rect 59828 24676 59829 24716
rect 59787 24667 59829 24676
rect 59596 24583 59636 24592
rect 59691 24632 59733 24641
rect 59691 24592 59692 24632
rect 59732 24592 59733 24632
rect 59691 24583 59733 24592
rect 59883 24632 59925 24641
rect 59883 24592 59884 24632
rect 59924 24592 59925 24632
rect 59883 24583 59925 24592
rect 59884 24498 59924 24583
rect 59980 24389 60020 26851
rect 60076 26816 60116 26825
rect 60076 26489 60116 26776
rect 60075 26480 60117 26489
rect 60075 26440 60076 26480
rect 60116 26440 60117 26480
rect 60075 26431 60117 26440
rect 60075 26144 60117 26153
rect 60172 26144 60212 26944
rect 60268 26732 60308 27523
rect 60459 27488 60501 27497
rect 60459 27448 60460 27488
rect 60500 27448 60501 27488
rect 60459 27439 60501 27448
rect 60363 27152 60405 27161
rect 60363 27112 60364 27152
rect 60404 27112 60405 27152
rect 60363 27103 60405 27112
rect 60364 26900 60404 27103
rect 60364 26851 60404 26860
rect 60268 26692 60404 26732
rect 60267 26312 60309 26321
rect 60267 26272 60268 26312
rect 60308 26272 60309 26312
rect 60267 26263 60309 26272
rect 60075 26104 60076 26144
rect 60116 26104 60212 26144
rect 60075 26095 60117 26104
rect 60076 26010 60116 26095
rect 60268 26060 60308 26263
rect 60268 26011 60308 26020
rect 60076 25892 60116 25901
rect 60116 25852 60308 25892
rect 60076 25843 60116 25852
rect 60268 25304 60308 25852
rect 60268 25255 60308 25264
rect 60364 25145 60404 26692
rect 60460 26321 60500 27439
rect 60556 27068 60596 28288
rect 60651 28328 60693 28337
rect 60651 28288 60652 28328
rect 60692 28288 60693 28328
rect 60651 28279 60693 28288
rect 60748 28328 60788 28337
rect 60652 28194 60692 28279
rect 60748 27245 60788 28288
rect 60940 27917 60980 28372
rect 60939 27908 60981 27917
rect 60939 27868 60940 27908
rect 60980 27868 60981 27908
rect 60939 27859 60981 27868
rect 60843 27656 60885 27665
rect 60843 27616 60844 27656
rect 60884 27616 60885 27656
rect 60843 27607 60885 27616
rect 60844 27522 60884 27607
rect 60939 27320 60981 27329
rect 60939 27280 60940 27320
rect 60980 27280 60981 27320
rect 60939 27271 60981 27280
rect 60747 27236 60789 27245
rect 60747 27196 60748 27236
rect 60788 27196 60789 27236
rect 60747 27187 60789 27196
rect 60748 27068 60788 27077
rect 60556 27028 60748 27068
rect 60748 27019 60788 27028
rect 60843 26900 60885 26909
rect 60843 26860 60844 26900
rect 60884 26860 60885 26900
rect 60843 26851 60885 26860
rect 60940 26900 60980 27271
rect 60940 26851 60980 26860
rect 60555 26732 60597 26741
rect 60555 26692 60556 26732
rect 60596 26692 60597 26732
rect 60555 26683 60597 26692
rect 60556 26648 60596 26683
rect 60459 26312 60501 26321
rect 60459 26272 60460 26312
rect 60500 26272 60501 26312
rect 60459 26263 60501 26272
rect 60459 26144 60501 26153
rect 60459 26104 60460 26144
rect 60500 26104 60501 26144
rect 60459 26095 60501 26104
rect 60460 25976 60500 26095
rect 60363 25136 60405 25145
rect 60363 25096 60364 25136
rect 60404 25096 60405 25136
rect 60363 25087 60405 25096
rect 60460 25061 60500 25936
rect 60459 25052 60501 25061
rect 60459 25012 60460 25052
rect 60500 25012 60501 25052
rect 60459 25003 60501 25012
rect 60267 24968 60309 24977
rect 60267 24928 60268 24968
rect 60308 24928 60309 24968
rect 60267 24919 60309 24928
rect 60171 24716 60213 24725
rect 60171 24676 60172 24716
rect 60212 24676 60213 24716
rect 60171 24667 60213 24676
rect 60268 24716 60308 24919
rect 60363 24800 60405 24809
rect 60363 24760 60364 24800
rect 60404 24760 60405 24800
rect 60363 24751 60405 24760
rect 60268 24667 60308 24676
rect 60172 24632 60212 24667
rect 60172 24581 60212 24592
rect 60364 24632 60404 24751
rect 60364 24583 60404 24592
rect 60459 24632 60501 24641
rect 60459 24592 60460 24632
rect 60500 24592 60501 24632
rect 60459 24583 60501 24592
rect 59979 24380 60021 24389
rect 59404 24340 59732 24380
rect 59692 23792 59732 24340
rect 59979 24340 59980 24380
rect 60020 24340 60021 24380
rect 59979 24331 60021 24340
rect 60363 24380 60405 24389
rect 60363 24340 60364 24380
rect 60404 24340 60405 24380
rect 60460 24380 60500 24583
rect 60556 24548 60596 26608
rect 60748 26648 60788 26657
rect 60651 26228 60693 26237
rect 60651 26188 60652 26228
rect 60692 26188 60693 26228
rect 60651 26179 60693 26188
rect 60652 26060 60692 26179
rect 60652 26011 60692 26020
rect 60748 25901 60788 26608
rect 60844 25976 60884 26851
rect 61036 26228 61076 28783
rect 61132 28160 61172 28169
rect 61172 28120 61268 28160
rect 61132 28111 61172 28120
rect 61131 27656 61173 27665
rect 61131 27616 61132 27656
rect 61172 27616 61173 27656
rect 61131 27607 61173 27616
rect 61132 26984 61172 27607
rect 61228 27329 61268 28120
rect 61324 27497 61364 29044
rect 61707 28328 61749 28337
rect 61707 28288 61708 28328
rect 61748 28288 61749 28328
rect 61707 28279 61749 28288
rect 61708 27656 61748 28279
rect 61900 28244 61940 28253
rect 61900 27833 61940 28204
rect 61899 27824 61941 27833
rect 61899 27784 61900 27824
rect 61940 27784 61941 27824
rect 61899 27775 61941 27784
rect 61708 27607 61748 27616
rect 61323 27488 61365 27497
rect 61323 27448 61324 27488
rect 61364 27448 61365 27488
rect 61323 27439 61365 27448
rect 61227 27320 61269 27329
rect 61227 27280 61228 27320
rect 61268 27280 61269 27320
rect 61227 27271 61269 27280
rect 61996 27077 62036 31471
rect 61995 27068 62037 27077
rect 61995 27028 61996 27068
rect 62036 27028 62037 27068
rect 61995 27019 62037 27028
rect 61132 26935 61172 26944
rect 62092 26984 62132 26993
rect 61323 26564 61365 26573
rect 61323 26524 61324 26564
rect 61364 26524 61365 26564
rect 61323 26515 61365 26524
rect 61227 26312 61269 26321
rect 61227 26272 61228 26312
rect 61268 26272 61269 26312
rect 61227 26263 61269 26272
rect 60747 25892 60789 25901
rect 60747 25852 60748 25892
rect 60788 25852 60789 25892
rect 60747 25843 60789 25852
rect 60652 25304 60692 25313
rect 60652 25145 60692 25264
rect 60651 25136 60693 25145
rect 60651 25096 60652 25136
rect 60692 25096 60693 25136
rect 60651 25087 60693 25096
rect 60748 24725 60788 25843
rect 60844 25817 60884 25936
rect 60940 26188 61076 26228
rect 60843 25808 60885 25817
rect 60843 25768 60844 25808
rect 60884 25768 60885 25808
rect 60843 25759 60885 25768
rect 60940 25388 60980 26188
rect 61228 26069 61268 26263
rect 61035 26060 61077 26069
rect 61035 26020 61036 26060
rect 61076 26020 61077 26060
rect 61035 26011 61077 26020
rect 61227 26060 61269 26069
rect 61227 26020 61228 26060
rect 61268 26020 61269 26060
rect 61227 26011 61269 26020
rect 61036 25926 61076 26011
rect 61131 25976 61173 25985
rect 61131 25936 61132 25976
rect 61172 25936 61173 25976
rect 61131 25927 61173 25936
rect 60940 25348 61076 25388
rect 60939 25136 60981 25145
rect 60939 25096 60940 25136
rect 60980 25096 60981 25136
rect 60939 25087 60981 25096
rect 60747 24716 60789 24725
rect 60747 24676 60748 24716
rect 60788 24676 60789 24716
rect 60747 24667 60789 24676
rect 60748 24548 60788 24557
rect 60556 24508 60748 24548
rect 60748 24499 60788 24508
rect 60940 24464 60980 25087
rect 60940 24415 60980 24424
rect 60556 24380 60596 24389
rect 60460 24340 60556 24380
rect 60363 24331 60405 24340
rect 60556 24331 60596 24340
rect 60076 23792 60116 23801
rect 58868 23752 59060 23792
rect 58828 23743 58868 23752
rect 58443 23708 58485 23717
rect 58443 23668 58444 23708
rect 58484 23668 58485 23708
rect 59020 23708 59060 23752
rect 59348 23752 59636 23792
rect 59308 23743 59348 23752
rect 59020 23668 59252 23708
rect 58443 23659 58485 23668
rect 58540 23624 58580 23633
rect 58540 23060 58580 23584
rect 58924 23624 58964 23633
rect 58964 23584 59156 23624
rect 58924 23575 58964 23584
rect 58348 23020 58495 23060
rect 58540 23020 58785 23060
rect 58156 22744 58385 22784
rect 58345 22596 58385 22744
rect 58455 22596 58495 23020
rect 58745 22596 58785 23020
rect 58854 22868 58896 22877
rect 58854 22828 58855 22868
rect 58895 22828 58896 22868
rect 58854 22819 58896 22828
rect 58855 22596 58895 22819
rect 59116 22784 59156 23584
rect 59212 23060 59252 23668
rect 59404 23624 59444 23633
rect 59404 23060 59444 23584
rect 59596 23060 59636 23752
rect 59732 23752 60020 23792
rect 59692 23743 59732 23752
rect 59788 23624 59828 23633
rect 59788 23060 59828 23584
rect 59980 23060 60020 23752
rect 60364 23792 60404 24331
rect 60460 23792 60500 23801
rect 60844 23792 60884 23801
rect 61036 23792 61076 25348
rect 61132 24641 61172 25927
rect 61131 24632 61173 24641
rect 61131 24592 61132 24632
rect 61172 24592 61173 24632
rect 61131 24583 61173 24592
rect 61324 23792 61364 26515
rect 61611 26228 61653 26237
rect 61611 26188 61612 26228
rect 61652 26188 61653 26228
rect 61611 26179 61653 26188
rect 61612 26094 61652 26179
rect 61996 26144 62036 26153
rect 62092 26144 62132 26944
rect 62036 26104 62132 26144
rect 61996 26095 62036 26104
rect 61515 25304 61557 25313
rect 61515 25264 61516 25304
rect 61556 25264 61557 25304
rect 61515 25255 61557 25264
rect 61516 25170 61556 25255
rect 61707 24968 61749 24977
rect 61707 24928 61708 24968
rect 61748 24928 61749 24968
rect 61707 24919 61749 24928
rect 61708 23792 61748 24919
rect 62188 24137 62228 33100
rect 62476 32873 62516 32958
rect 62475 32864 62517 32873
rect 62475 32824 62476 32864
rect 62516 32824 62517 32864
rect 62475 32815 62517 32824
rect 62572 32864 62612 32873
rect 62380 32696 62420 32705
rect 62420 32656 62516 32696
rect 62380 32647 62420 32656
rect 62283 31856 62325 31865
rect 62283 31816 62284 31856
rect 62324 31816 62325 31856
rect 62283 31807 62325 31816
rect 62284 30932 62324 31807
rect 62476 31352 62516 32656
rect 62572 32621 62612 32824
rect 62668 32864 62708 33100
rect 62860 33032 62900 33664
rect 63052 33704 63092 33713
rect 63052 33545 63092 33664
rect 63243 33704 63285 33713
rect 63243 33664 63244 33704
rect 63284 33664 63285 33704
rect 63243 33655 63285 33664
rect 63147 33620 63189 33629
rect 63147 33580 63148 33620
rect 63188 33580 63189 33620
rect 63147 33571 63189 33580
rect 63051 33536 63093 33545
rect 63051 33496 63052 33536
rect 63092 33496 63093 33536
rect 63051 33487 63093 33496
rect 63148 33284 63188 33571
rect 63244 33570 63284 33655
rect 63724 33536 63764 33545
rect 63436 33496 63724 33536
rect 63148 33244 63284 33284
rect 62860 32992 63092 33032
rect 62571 32612 62613 32621
rect 62571 32572 62572 32612
rect 62612 32572 62613 32612
rect 62571 32563 62613 32572
rect 62668 32360 62708 32824
rect 62860 32864 62900 32873
rect 62764 32360 62804 32369
rect 62668 32320 62764 32360
rect 62571 32276 62613 32285
rect 62571 32236 62572 32276
rect 62612 32236 62708 32276
rect 62571 32227 62613 32236
rect 62476 31303 62516 31312
rect 62668 31352 62708 32236
rect 62764 32117 62804 32320
rect 62763 32108 62805 32117
rect 62763 32068 62764 32108
rect 62804 32068 62805 32108
rect 62763 32059 62805 32068
rect 62860 32024 62900 32824
rect 63052 32864 63092 32992
rect 63244 32957 63284 33244
rect 63436 33140 63476 33496
rect 63724 33487 63764 33496
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 64012 33140 64052 34579
rect 63436 33100 63668 33140
rect 63243 32948 63285 32957
rect 63243 32908 63244 32948
rect 63284 32908 63285 32948
rect 63243 32899 63285 32908
rect 62956 32780 62996 32789
rect 62956 32705 62996 32740
rect 62955 32696 62997 32705
rect 62955 32656 62956 32696
rect 62996 32656 62997 32696
rect 62955 32647 62997 32656
rect 62956 32285 62996 32647
rect 62955 32276 62997 32285
rect 62955 32236 62956 32276
rect 62996 32236 62997 32276
rect 62955 32227 62997 32236
rect 62956 32024 62996 32033
rect 62860 31984 62956 32024
rect 62956 31975 62996 31984
rect 63052 31697 63092 32824
rect 63147 32864 63189 32873
rect 63147 32824 63148 32864
rect 63188 32824 63189 32864
rect 63147 32815 63189 32824
rect 63628 32864 63668 33100
rect 63628 32815 63668 32824
rect 63820 33100 64052 33140
rect 64204 33140 64244 36688
rect 64396 36728 64436 36739
rect 64396 36653 64436 36688
rect 65355 36728 65397 36737
rect 65355 36688 65356 36728
rect 65396 36688 65397 36728
rect 65355 36679 65397 36688
rect 64395 36644 64437 36653
rect 64395 36604 64396 36644
rect 64436 36604 64437 36644
rect 64395 36595 64437 36604
rect 64491 36056 64533 36065
rect 64491 36016 64492 36056
rect 64532 36016 64533 36056
rect 64491 36007 64533 36016
rect 64395 35888 64437 35897
rect 64395 35848 64396 35888
rect 64436 35848 64437 35888
rect 64395 35839 64437 35848
rect 64396 35754 64436 35839
rect 64396 34376 64436 34385
rect 64492 34376 64532 36007
rect 64780 35888 64820 35897
rect 64780 35720 64820 35848
rect 64684 35680 64820 35720
rect 64684 35384 64724 35680
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 64684 35344 64916 35384
rect 64876 35048 64916 35344
rect 64876 34999 64916 35008
rect 64436 34336 64532 34376
rect 64396 34327 64436 34336
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 64204 33100 64724 33140
rect 63148 31865 63188 32815
rect 63244 32780 63284 32789
rect 63244 32369 63284 32740
rect 63339 32612 63381 32621
rect 63339 32572 63340 32612
rect 63380 32572 63381 32612
rect 63339 32563 63381 32572
rect 63243 32360 63285 32369
rect 63243 32320 63244 32360
rect 63284 32320 63285 32360
rect 63243 32311 63285 32320
rect 63340 32219 63380 32563
rect 63435 32276 63477 32285
rect 63435 32236 63436 32276
rect 63476 32236 63477 32276
rect 63435 32227 63477 32236
rect 63244 32192 63284 32203
rect 63340 32170 63380 32179
rect 63244 32117 63284 32152
rect 63243 32108 63285 32117
rect 63243 32068 63244 32108
rect 63284 32068 63285 32108
rect 63243 32059 63285 32068
rect 63436 31940 63476 32227
rect 63244 31900 63476 31940
rect 63628 32192 63668 32201
rect 63628 31940 63668 32152
rect 63820 31940 63860 33100
rect 64492 32864 64532 32873
rect 63915 32780 63957 32789
rect 63915 32740 63916 32780
rect 63956 32740 63957 32780
rect 63915 32731 63957 32740
rect 63916 32192 63956 32731
rect 64107 32696 64149 32705
rect 64107 32656 64108 32696
rect 64148 32656 64149 32696
rect 64107 32647 64149 32656
rect 64011 32360 64053 32369
rect 64011 32320 64012 32360
rect 64052 32320 64053 32360
rect 64011 32311 64053 32320
rect 64012 32226 64052 32311
rect 63916 32143 63956 32152
rect 64108 32192 64148 32647
rect 64299 32276 64341 32285
rect 64299 32236 64300 32276
rect 64340 32236 64436 32276
rect 64299 32227 64341 32236
rect 64108 32143 64148 32152
rect 64204 32192 64244 32201
rect 64204 32024 64244 32152
rect 64396 32192 64436 32236
rect 64492 32201 64532 32824
rect 64587 32612 64629 32621
rect 64587 32572 64588 32612
rect 64628 32572 64629 32612
rect 64587 32563 64629 32572
rect 64396 32143 64436 32152
rect 64491 32192 64533 32201
rect 64491 32152 64492 32192
rect 64532 32152 64533 32192
rect 64491 32143 64533 32152
rect 64588 32192 64628 32563
rect 64588 32143 64628 32152
rect 64492 32024 64532 32033
rect 64204 31984 64492 32024
rect 64492 31975 64532 31984
rect 63628 31900 64052 31940
rect 63147 31856 63189 31865
rect 63147 31816 63148 31856
rect 63188 31816 63189 31856
rect 63147 31807 63189 31816
rect 63051 31688 63093 31697
rect 63051 31648 63052 31688
rect 63092 31648 63093 31688
rect 63051 31639 63093 31648
rect 63052 31520 63092 31529
rect 62668 31303 62708 31312
rect 62764 31480 63052 31520
rect 62764 31352 62804 31480
rect 63052 31471 63092 31480
rect 63147 31352 63189 31361
rect 62764 31303 62804 31312
rect 63051 31314 63092 31337
rect 63051 31277 63052 31314
rect 62571 31268 62613 31277
rect 62571 31228 62572 31268
rect 62612 31228 62613 31268
rect 62571 31219 62613 31228
rect 63050 31274 63052 31277
rect 63147 31312 63148 31352
rect 63188 31312 63189 31352
rect 63147 31303 63189 31312
rect 63244 31352 63284 31900
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 63532 31520 63572 31529
rect 63050 31268 63092 31274
rect 63050 31228 63051 31268
rect 63091 31228 63092 31268
rect 62572 31134 62612 31219
rect 63050 31198 63092 31228
rect 62284 30892 62612 30932
rect 62475 30764 62517 30773
rect 62475 30724 62476 30764
rect 62516 30724 62517 30764
rect 62475 30715 62517 30724
rect 62380 29000 62420 29009
rect 62284 28328 62324 28337
rect 62380 28328 62420 28960
rect 62324 28288 62420 28328
rect 62284 28279 62324 28288
rect 62283 27068 62325 27077
rect 62283 27028 62284 27068
rect 62324 27028 62325 27068
rect 62283 27019 62325 27028
rect 62284 26909 62324 27019
rect 62283 26900 62325 26909
rect 62283 26860 62284 26900
rect 62324 26860 62325 26900
rect 62283 26851 62325 26860
rect 62283 24464 62325 24473
rect 62283 24424 62284 24464
rect 62324 24424 62325 24464
rect 62283 24415 62325 24424
rect 62187 24128 62229 24137
rect 62187 24088 62188 24128
rect 62228 24088 62229 24128
rect 62187 24079 62229 24088
rect 62284 24053 62324 24415
rect 62476 24389 62516 30715
rect 62572 24473 62612 30892
rect 63052 30680 63092 30689
rect 62859 30428 62901 30437
rect 62859 30388 62860 30428
rect 62900 30388 62901 30428
rect 62859 30379 62901 30388
rect 62860 29840 62900 30379
rect 63052 30269 63092 30640
rect 63051 30260 63093 30269
rect 63051 30220 63052 30260
rect 63092 30220 63093 30260
rect 63051 30211 63093 30220
rect 62955 30092 62997 30101
rect 62955 30052 62956 30092
rect 62996 30052 62997 30092
rect 62955 30043 62997 30052
rect 62956 29958 62996 30043
rect 63148 29924 63188 31303
rect 63244 31193 63284 31312
rect 63340 31337 63380 31346
rect 63243 31184 63285 31193
rect 63243 31144 63244 31184
rect 63284 31144 63285 31184
rect 63243 31135 63285 31144
rect 63340 30932 63380 31297
rect 63244 30892 63380 30932
rect 63244 30176 63284 30892
rect 63436 30680 63476 30689
rect 63532 30680 63572 31480
rect 63476 30640 63572 30680
rect 63436 30631 63476 30640
rect 63435 30260 63477 30269
rect 63435 30220 63436 30260
rect 63476 30220 63477 30260
rect 63435 30211 63477 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 63339 30176 63381 30185
rect 63244 30136 63340 30176
rect 63380 30136 63381 30176
rect 63244 30008 63284 30136
rect 63339 30127 63381 30136
rect 63340 30108 63380 30127
rect 63436 30092 63476 30211
rect 63628 30092 63668 30101
rect 63436 30052 63628 30092
rect 63628 30043 63668 30052
rect 63244 29968 63476 30008
rect 63148 29884 63284 29924
rect 63244 29840 63284 29884
rect 62860 29800 63092 29840
rect 62956 29672 62996 29681
rect 62956 29009 62996 29632
rect 62955 29000 62997 29009
rect 62955 28960 62956 29000
rect 62996 28960 62997 29000
rect 62955 28951 62997 28960
rect 63052 28916 63092 29800
rect 63436 29840 63476 29968
rect 64012 29933 64052 31900
rect 64107 31856 64149 31865
rect 64107 31816 64108 31856
rect 64148 31816 64149 31856
rect 64107 31807 64149 31816
rect 64011 29924 64053 29933
rect 64011 29884 64012 29924
rect 64052 29884 64053 29924
rect 64011 29875 64053 29884
rect 63244 29791 63284 29800
rect 63340 29819 63380 29828
rect 63436 29791 63476 29800
rect 63627 29840 63669 29849
rect 63627 29800 63628 29840
rect 63668 29800 63669 29840
rect 63627 29791 63669 29800
rect 63819 29840 63861 29849
rect 63819 29800 63820 29840
rect 63860 29800 63861 29840
rect 63819 29791 63861 29800
rect 63916 29840 63956 29849
rect 63147 29756 63189 29765
rect 63147 29716 63148 29756
rect 63188 29716 63189 29756
rect 63147 29707 63189 29716
rect 63148 29622 63188 29707
rect 63340 29681 63380 29779
rect 63628 29706 63668 29791
rect 63820 29706 63860 29791
rect 63339 29672 63381 29681
rect 63339 29632 63340 29672
rect 63380 29632 63381 29672
rect 63339 29623 63381 29632
rect 63436 29336 63476 29345
rect 63916 29336 63956 29800
rect 64108 29336 64148 31807
rect 64684 30689 64724 33100
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 65259 32192 65301 32201
rect 65259 32152 65260 32192
rect 65300 32152 65301 32192
rect 65259 32143 65301 32152
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 64300 30680 64340 30689
rect 64683 30680 64725 30689
rect 64340 30640 64436 30680
rect 64300 30631 64340 30640
rect 63476 29296 63956 29336
rect 64012 29296 64148 29336
rect 63436 29287 63476 29296
rect 63531 29168 63573 29177
rect 63340 29157 63380 29166
rect 63531 29128 63532 29168
rect 63572 29128 63573 29168
rect 63531 29119 63573 29128
rect 63628 29168 63668 29177
rect 63820 29168 63860 29177
rect 63668 29128 63820 29168
rect 63628 29119 63668 29128
rect 63340 28916 63380 29117
rect 63435 29084 63477 29093
rect 63435 29044 63436 29084
rect 63476 29044 63477 29084
rect 63435 29035 63477 29044
rect 63052 28876 63380 28916
rect 63147 28328 63189 28337
rect 63147 28288 63148 28328
rect 63188 28288 63189 28328
rect 63147 28279 63189 28288
rect 63148 28194 63188 28279
rect 62860 27404 62900 27413
rect 62860 27245 62900 27364
rect 62859 27236 62901 27245
rect 62859 27196 62860 27236
rect 62900 27196 62901 27236
rect 62859 27187 62901 27196
rect 62860 26573 62900 27187
rect 63244 26825 63284 28876
rect 63436 27581 63476 29035
rect 63532 29034 63572 29119
rect 63820 28916 63860 29128
rect 63915 29168 63957 29177
rect 63915 29128 63916 29168
rect 63956 29128 63957 29168
rect 63915 29119 63957 29128
rect 64012 29168 64052 29296
rect 63916 29034 63956 29119
rect 64012 29093 64052 29128
rect 64108 29168 64148 29177
rect 64011 29084 64053 29093
rect 64011 29044 64012 29084
rect 64052 29044 64053 29084
rect 64011 29035 64053 29044
rect 64012 29004 64052 29035
rect 63820 28876 64052 28916
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 63723 28496 63765 28505
rect 63723 28456 63724 28496
rect 63764 28456 63765 28496
rect 63723 28447 63765 28456
rect 63531 27992 63573 28001
rect 63531 27952 63532 27992
rect 63572 27952 63573 27992
rect 63531 27943 63573 27952
rect 63435 27572 63477 27581
rect 63435 27532 63436 27572
rect 63476 27532 63477 27572
rect 63435 27523 63477 27532
rect 63532 27404 63572 27943
rect 63724 27413 63764 28447
rect 64012 28253 64052 28876
rect 64011 28244 64053 28253
rect 64011 28204 64012 28244
rect 64052 28204 64053 28244
rect 64011 28195 64053 28204
rect 64011 27824 64053 27833
rect 64011 27784 64012 27824
rect 64052 27784 64053 27824
rect 64011 27775 64053 27784
rect 64012 27690 64052 27775
rect 63820 27656 63860 27665
rect 63436 27364 63572 27404
rect 63723 27404 63765 27413
rect 63723 27364 63724 27404
rect 63764 27364 63765 27404
rect 63820 27404 63860 27616
rect 63915 27656 63957 27665
rect 63915 27616 63916 27656
rect 63956 27616 63957 27656
rect 63915 27607 63957 27616
rect 64108 27656 64148 29128
rect 64203 29168 64245 29177
rect 64203 29128 64204 29168
rect 64244 29128 64245 29168
rect 64203 29119 64245 29128
rect 64108 27607 64148 27616
rect 63916 27522 63956 27607
rect 63820 27364 64052 27404
rect 63243 26816 63285 26825
rect 63243 26776 63244 26816
rect 63284 26776 63285 26816
rect 63243 26767 63285 26776
rect 62859 26564 62901 26573
rect 62859 26524 62860 26564
rect 62900 26524 62901 26564
rect 62859 26515 62901 26524
rect 62860 26144 62900 26153
rect 62860 25313 62900 26104
rect 63436 25481 63476 27364
rect 63723 27355 63765 27364
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 63820 27068 63860 27077
rect 64012 27068 64052 27364
rect 64204 27152 64244 29119
rect 64396 28337 64436 30640
rect 64683 30640 64684 30680
rect 64724 30640 64725 30680
rect 64683 30631 64725 30640
rect 64587 29756 64629 29765
rect 64587 29716 64588 29756
rect 64628 29716 64629 29756
rect 64587 29707 64629 29716
rect 64588 28337 64628 29707
rect 64684 28505 64724 30631
rect 65260 30260 65300 32143
rect 65356 31445 65396 36679
rect 65644 36065 65684 37351
rect 66124 37232 66164 37241
rect 66124 36653 66164 37192
rect 67276 36905 67316 37948
rect 67467 37988 67509 37997
rect 67467 37948 67468 37988
rect 67508 37948 67509 37988
rect 67467 37939 67509 37948
rect 67659 37988 67701 37997
rect 67659 37948 67660 37988
rect 67700 37948 67701 37988
rect 67659 37939 67701 37948
rect 67468 37854 67508 37939
rect 67563 37400 67605 37409
rect 67563 37360 67564 37400
rect 67604 37360 67605 37400
rect 67563 37351 67605 37360
rect 67564 37266 67604 37351
rect 67275 36896 67317 36905
rect 67275 36856 67276 36896
rect 67316 36856 67317 36896
rect 67275 36847 67317 36856
rect 67755 36896 67797 36905
rect 67755 36856 67756 36896
rect 67796 36856 67797 36896
rect 67755 36847 67797 36856
rect 66508 36728 66548 36737
rect 66700 36728 66740 36737
rect 66548 36688 66644 36728
rect 66508 36679 66548 36688
rect 66123 36644 66165 36653
rect 66123 36604 66124 36644
rect 66164 36604 66165 36644
rect 66123 36595 66165 36604
rect 66508 36476 66548 36485
rect 65643 36056 65685 36065
rect 65643 36016 65644 36056
rect 65684 36016 65685 36056
rect 65643 36007 65685 36016
rect 65644 35888 65684 36007
rect 66508 35897 66548 36436
rect 66604 36149 66644 36688
rect 66603 36140 66645 36149
rect 66603 36100 66604 36140
rect 66644 36100 66645 36140
rect 66603 36091 66645 36100
rect 65644 35839 65684 35848
rect 66507 35888 66549 35897
rect 66507 35848 66508 35888
rect 66548 35848 66549 35888
rect 66507 35839 66549 35848
rect 65643 35720 65685 35729
rect 65643 35680 65644 35720
rect 65684 35680 65685 35720
rect 65643 35671 65685 35680
rect 65644 35057 65684 35671
rect 66700 35561 66740 36688
rect 66796 36728 66836 36737
rect 66796 36560 66836 36688
rect 67180 36728 67220 36737
rect 67372 36728 67412 36737
rect 67220 36688 67316 36728
rect 67180 36679 67220 36688
rect 67180 36560 67220 36569
rect 66796 36520 67180 36560
rect 67180 36511 67220 36520
rect 67276 36308 67316 36688
rect 67372 36392 67412 36688
rect 67467 36728 67509 36737
rect 67467 36688 67468 36728
rect 67508 36688 67509 36728
rect 67467 36679 67509 36688
rect 67468 36594 67508 36679
rect 67756 36644 67796 36847
rect 67756 36595 67796 36604
rect 67372 36352 67508 36392
rect 67276 36268 67412 36308
rect 67275 36140 67317 36149
rect 67275 36100 67276 36140
rect 67316 36100 67317 36140
rect 67275 36091 67317 36100
rect 67180 35897 67220 35982
rect 66988 35888 67028 35897
rect 66796 35720 66836 35729
rect 66988 35720 67028 35848
rect 66836 35680 67028 35720
rect 67084 35888 67124 35897
rect 67084 35720 67124 35848
rect 67179 35888 67221 35897
rect 67179 35848 67180 35888
rect 67220 35848 67221 35888
rect 67179 35839 67221 35848
rect 67276 35888 67316 36091
rect 67372 35897 67412 36268
rect 67276 35839 67316 35848
rect 67371 35888 67413 35897
rect 67371 35848 67372 35888
rect 67412 35848 67413 35888
rect 67371 35839 67413 35848
rect 67084 35680 67220 35720
rect 66027 35552 66069 35561
rect 66027 35512 66028 35552
rect 66068 35512 66069 35552
rect 66027 35503 66069 35512
rect 66699 35552 66741 35561
rect 66699 35512 66700 35552
rect 66740 35512 66741 35552
rect 66699 35503 66741 35512
rect 66028 35300 66068 35503
rect 66796 35384 66836 35680
rect 67083 35552 67125 35561
rect 67083 35512 67084 35552
rect 67124 35512 67125 35552
rect 67083 35503 67125 35512
rect 66028 35251 66068 35260
rect 66604 35344 66836 35384
rect 65932 35216 65972 35225
rect 65643 35048 65685 35057
rect 65643 35008 65644 35048
rect 65684 35008 65685 35048
rect 65643 34999 65685 35008
rect 65548 34208 65588 34217
rect 65452 34168 65548 34208
rect 65452 33797 65492 34168
rect 65548 34159 65588 34168
rect 65451 33788 65493 33797
rect 65451 33748 65452 33788
rect 65492 33748 65493 33788
rect 65451 33739 65493 33748
rect 65452 31949 65492 33739
rect 65547 33704 65589 33713
rect 65547 33664 65548 33704
rect 65588 33664 65589 33704
rect 65547 33655 65589 33664
rect 65451 31940 65493 31949
rect 65451 31900 65452 31940
rect 65492 31900 65493 31940
rect 65451 31891 65493 31900
rect 65548 31772 65588 33655
rect 65644 32873 65684 34999
rect 65835 34880 65877 34889
rect 65835 34840 65836 34880
rect 65876 34840 65877 34880
rect 65835 34831 65877 34840
rect 65836 34721 65876 34831
rect 65835 34712 65877 34721
rect 65835 34672 65836 34712
rect 65876 34672 65877 34712
rect 65835 34663 65877 34672
rect 65739 34208 65781 34217
rect 65739 34168 65740 34208
rect 65780 34168 65781 34208
rect 65739 34159 65781 34168
rect 65643 32864 65685 32873
rect 65643 32824 65644 32864
rect 65684 32824 65685 32864
rect 65643 32815 65685 32824
rect 65644 32696 65684 32707
rect 65644 32621 65684 32656
rect 65643 32612 65685 32621
rect 65643 32572 65644 32612
rect 65684 32572 65685 32612
rect 65643 32563 65685 32572
rect 65740 32192 65780 34159
rect 65836 33536 65876 34663
rect 65932 33881 65972 35176
rect 66124 35216 66164 35225
rect 66124 35048 66164 35176
rect 66604 35216 66644 35344
rect 66316 35048 66356 35057
rect 66124 35008 66316 35048
rect 66316 34999 66356 35008
rect 66316 34385 66356 34470
rect 66124 34376 66164 34385
rect 66124 34133 66164 34336
rect 66315 34376 66357 34385
rect 66315 34336 66316 34376
rect 66356 34336 66357 34376
rect 66315 34327 66357 34336
rect 66412 34376 66452 34385
rect 66604 34376 66644 35176
rect 66700 35216 66740 35225
rect 66988 35216 67028 35225
rect 66700 34973 66740 35176
rect 66796 35176 66988 35216
rect 66699 34964 66741 34973
rect 66699 34924 66700 34964
rect 66740 34924 66741 34964
rect 66699 34915 66741 34924
rect 66452 34336 66644 34376
rect 66412 34327 66452 34336
rect 66220 34208 66260 34217
rect 66316 34208 66356 34327
rect 66796 34217 66836 35176
rect 66988 35167 67028 35176
rect 66891 34712 66933 34721
rect 66891 34672 66892 34712
rect 66932 34672 66933 34712
rect 66891 34663 66933 34672
rect 66892 34628 66932 34663
rect 66892 34577 66932 34588
rect 66892 34376 66932 34385
rect 66795 34208 66837 34217
rect 66316 34168 66548 34208
rect 66123 34124 66165 34133
rect 66123 34084 66124 34124
rect 66164 34084 66165 34124
rect 66123 34075 66165 34084
rect 66220 33956 66260 34168
rect 66220 33916 66452 33956
rect 65931 33872 65973 33881
rect 65931 33832 65932 33872
rect 65972 33832 65973 33872
rect 65931 33823 65973 33832
rect 66220 33788 66260 33797
rect 66124 33704 66164 33713
rect 66124 33536 66164 33664
rect 65836 33496 65972 33536
rect 65835 33368 65877 33377
rect 65835 33328 65836 33368
rect 65876 33328 65877 33368
rect 65835 33319 65877 33328
rect 65836 32864 65876 33319
rect 65932 33140 65972 33496
rect 66028 33496 66164 33536
rect 66028 33377 66068 33496
rect 66027 33368 66069 33377
rect 66027 33328 66028 33368
rect 66068 33328 66069 33368
rect 66027 33319 66069 33328
rect 65932 33100 66068 33140
rect 65836 32815 65876 32824
rect 65931 32864 65973 32873
rect 65931 32824 65932 32864
rect 65972 32824 65973 32864
rect 65931 32815 65973 32824
rect 66028 32864 66068 33100
rect 66028 32815 66068 32824
rect 66124 32864 66164 32873
rect 66220 32864 66260 33748
rect 66316 33704 66356 33713
rect 66316 33140 66356 33664
rect 66412 33704 66452 33916
rect 66412 33655 66452 33664
rect 66508 33545 66548 34168
rect 66795 34168 66796 34208
rect 66836 34168 66837 34208
rect 66795 34159 66837 34168
rect 66603 33704 66645 33713
rect 66603 33664 66604 33704
rect 66644 33664 66645 33704
rect 66603 33655 66645 33664
rect 66796 33704 66836 33713
rect 66604 33570 66644 33655
rect 66507 33536 66549 33545
rect 66507 33496 66508 33536
rect 66548 33496 66549 33536
rect 66507 33487 66549 33496
rect 66700 33452 66740 33461
rect 66700 33140 66740 33412
rect 66316 33100 66740 33140
rect 66316 32864 66356 32873
rect 66220 32824 66316 32864
rect 65932 32730 65972 32815
rect 66124 32696 66164 32824
rect 66316 32815 66356 32824
rect 66219 32696 66261 32705
rect 66124 32656 66220 32696
rect 66260 32656 66261 32696
rect 66219 32647 66261 32656
rect 66220 32276 66260 32647
rect 66220 32227 66260 32236
rect 65835 32192 65877 32201
rect 65740 32152 65836 32192
rect 65876 32152 65877 32192
rect 65835 32143 65877 32152
rect 66124 32192 66164 32201
rect 65836 32058 65876 32143
rect 66124 31772 66164 32152
rect 66315 32192 66357 32201
rect 66315 32152 66316 32192
rect 66356 32152 66357 32192
rect 66315 32143 66357 32152
rect 65548 31732 65684 31772
rect 66124 31732 66260 31772
rect 65644 31613 65684 31732
rect 65643 31604 65685 31613
rect 65643 31564 65644 31604
rect 65684 31564 65685 31604
rect 65643 31555 65685 31564
rect 65355 31436 65397 31445
rect 65355 31396 65356 31436
rect 65396 31396 65397 31436
rect 65355 31387 65397 31396
rect 65164 30220 65300 30260
rect 65164 29840 65204 30220
rect 65164 29765 65204 29800
rect 65163 29756 65205 29765
rect 65163 29716 65164 29756
rect 65204 29716 65205 29756
rect 65163 29707 65205 29716
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 64972 29168 65012 29179
rect 64972 29093 65012 29128
rect 65164 29168 65204 29177
rect 65204 29128 65300 29168
rect 65164 29119 65204 29128
rect 64971 29084 65013 29093
rect 64971 29044 64972 29084
rect 65012 29044 65013 29084
rect 64971 29035 65013 29044
rect 65068 28916 65108 28925
rect 65108 28876 65204 28916
rect 65068 28867 65108 28876
rect 64683 28496 64725 28505
rect 64683 28456 64684 28496
rect 64724 28456 64725 28496
rect 64683 28447 64725 28456
rect 64395 28328 64437 28337
rect 64395 28288 64396 28328
rect 64436 28288 64437 28328
rect 64395 28279 64437 28288
rect 64587 28328 64629 28337
rect 64587 28288 64588 28328
rect 64628 28288 64629 28328
rect 64587 28279 64629 28288
rect 64876 28328 64916 28337
rect 64299 28244 64341 28253
rect 64299 28204 64300 28244
rect 64340 28204 64341 28244
rect 64299 28195 64341 28204
rect 64300 28160 64340 28195
rect 64300 28109 64340 28120
rect 64396 27413 64436 28279
rect 64588 28194 64628 28279
rect 64876 28169 64916 28288
rect 64971 28244 65013 28253
rect 64971 28204 64972 28244
rect 65012 28204 65013 28244
rect 64971 28195 65013 28204
rect 64875 28160 64917 28169
rect 64875 28120 64876 28160
rect 64916 28120 64917 28160
rect 64875 28111 64917 28120
rect 64972 28110 65012 28195
rect 65164 28160 65204 28876
rect 65260 28580 65300 29128
rect 65356 29093 65396 31387
rect 65644 30701 65684 31555
rect 65739 31436 65781 31445
rect 65739 31396 65740 31436
rect 65780 31396 65781 31436
rect 65739 31387 65781 31396
rect 65644 30652 65684 30661
rect 65740 30596 65780 31387
rect 66220 31361 66260 31732
rect 66316 31604 66356 32143
rect 66316 31555 66356 31564
rect 66315 31436 66357 31445
rect 66315 31396 66316 31436
rect 66356 31396 66357 31436
rect 66315 31387 66357 31396
rect 66219 31352 66261 31361
rect 66219 31312 66220 31352
rect 66260 31312 66261 31352
rect 66219 31303 66261 31312
rect 66316 31352 66356 31387
rect 66412 31352 66452 33100
rect 66796 33032 66836 33664
rect 66508 32992 66836 33032
rect 66508 32402 66548 32992
rect 66699 32864 66741 32873
rect 66699 32824 66700 32864
rect 66740 32824 66741 32864
rect 66699 32815 66741 32824
rect 66700 32730 66740 32815
rect 66508 32353 66548 32362
rect 66699 32192 66741 32201
rect 66699 32152 66700 32192
rect 66740 32152 66741 32192
rect 66699 32143 66741 32152
rect 66700 32058 66740 32143
rect 66892 31697 66932 34336
rect 67084 34376 67124 35503
rect 67180 34889 67220 35680
rect 67276 35216 67316 35225
rect 67179 34880 67221 34889
rect 67179 34840 67180 34880
rect 67220 34840 67221 34880
rect 67179 34831 67221 34840
rect 67276 34721 67316 35176
rect 67468 34721 67508 36352
rect 67755 36056 67797 36065
rect 67755 36016 67756 36056
rect 67796 36016 67797 36056
rect 67755 36007 67797 36016
rect 67660 35216 67700 35225
rect 67563 34964 67605 34973
rect 67563 34924 67564 34964
rect 67604 34924 67605 34964
rect 67563 34915 67605 34924
rect 67275 34712 67317 34721
rect 67275 34672 67276 34712
rect 67316 34672 67317 34712
rect 67275 34663 67317 34672
rect 67467 34712 67509 34721
rect 67467 34672 67468 34712
rect 67508 34672 67509 34712
rect 67467 34663 67509 34672
rect 67468 34544 67508 34553
rect 67084 34327 67124 34336
rect 67180 34504 67468 34544
rect 67180 34376 67220 34504
rect 67468 34495 67508 34504
rect 67180 34327 67220 34336
rect 67371 34376 67413 34385
rect 67371 34336 67372 34376
rect 67412 34336 67413 34376
rect 67371 34327 67413 34336
rect 67564 34376 67604 34915
rect 67660 34889 67700 35176
rect 67659 34880 67701 34889
rect 67659 34840 67660 34880
rect 67700 34840 67701 34880
rect 67659 34831 67701 34840
rect 67756 34712 67796 36007
rect 67852 35813 67892 38200
rect 67947 38200 67948 38240
rect 67988 38200 67989 38240
rect 67947 38191 67989 38200
rect 68044 38240 68084 38249
rect 67948 38106 67988 38191
rect 67948 36896 67988 36905
rect 68044 36896 68084 38200
rect 67988 36856 68084 36896
rect 68140 38240 68180 38249
rect 67948 36847 67988 36856
rect 68043 36644 68085 36653
rect 68043 36604 68044 36644
rect 68084 36604 68085 36644
rect 68043 36595 68085 36604
rect 67948 36476 67988 36485
rect 67948 35981 67988 36436
rect 67947 35972 67989 35981
rect 67947 35932 67948 35972
rect 67988 35932 67989 35972
rect 67947 35923 67989 35932
rect 67851 35804 67893 35813
rect 67851 35764 67852 35804
rect 67892 35764 67893 35804
rect 67851 35755 67893 35764
rect 67851 34880 67893 34889
rect 67851 34840 67852 34880
rect 67892 34840 67893 34880
rect 67851 34831 67893 34840
rect 67564 34327 67604 34336
rect 67660 34672 67796 34712
rect 66988 33536 67028 33545
rect 66988 32873 67028 33496
rect 66987 32864 67029 32873
rect 66987 32824 66988 32864
rect 67028 32824 67029 32864
rect 66987 32815 67029 32824
rect 67084 32192 67124 32201
rect 67124 32152 67220 32192
rect 67084 32143 67124 32152
rect 66891 31688 66933 31697
rect 66891 31648 66892 31688
rect 66932 31648 66933 31688
rect 66891 31639 66933 31648
rect 66892 31520 66932 31529
rect 66604 31480 66892 31520
rect 66508 31352 66548 31361
rect 66412 31312 66508 31352
rect 66316 31301 66356 31312
rect 66508 31303 66548 31312
rect 66604 31352 66644 31480
rect 66892 31471 66932 31480
rect 67180 31520 67220 32152
rect 67180 31471 67220 31480
rect 66988 31361 67028 31446
rect 66604 31303 66644 31312
rect 66796 31352 66836 31361
rect 66796 31184 66836 31312
rect 66987 31352 67029 31361
rect 66987 31312 66988 31352
rect 67028 31312 67029 31352
rect 66987 31303 67029 31312
rect 67372 31184 67412 34327
rect 67660 33140 67700 34672
rect 67756 34544 67796 34553
rect 67852 34544 67892 34831
rect 67796 34504 67892 34544
rect 67756 34495 67796 34504
rect 67564 33100 67700 33140
rect 68044 33140 68084 36595
rect 68140 35393 68180 38200
rect 68236 38240 68276 38249
rect 68236 37241 68276 38200
rect 69291 38240 69333 38249
rect 69291 38200 69292 38240
rect 69332 38200 69333 38240
rect 69291 38191 69333 38200
rect 70635 38240 70677 38249
rect 70635 38200 70636 38240
rect 70676 38200 70677 38240
rect 70635 38191 70677 38200
rect 71020 38240 71060 38251
rect 68907 38156 68949 38165
rect 68907 38116 68908 38156
rect 68948 38116 68949 38156
rect 68907 38107 68949 38116
rect 68427 37400 68469 37409
rect 68427 37360 68428 37400
rect 68468 37360 68469 37400
rect 68427 37351 68469 37360
rect 68235 37232 68277 37241
rect 68235 37192 68236 37232
rect 68276 37192 68277 37232
rect 68235 37183 68277 37192
rect 68236 36728 68276 36737
rect 68236 35477 68276 36688
rect 68428 36065 68468 37351
rect 68619 37232 68661 37241
rect 68716 37232 68756 37241
rect 68619 37192 68620 37232
rect 68660 37192 68716 37232
rect 68619 37183 68661 37192
rect 68716 37183 68756 37192
rect 68523 36812 68565 36821
rect 68523 36772 68524 36812
rect 68564 36772 68565 36812
rect 68523 36763 68565 36772
rect 68524 36728 68564 36763
rect 68620 36737 68660 37183
rect 68524 36677 68564 36688
rect 68619 36728 68661 36737
rect 68619 36688 68620 36728
rect 68660 36688 68661 36728
rect 68619 36679 68661 36688
rect 68811 36728 68853 36737
rect 68811 36688 68812 36728
rect 68852 36688 68853 36728
rect 68811 36679 68853 36688
rect 68620 36594 68660 36679
rect 68427 36056 68469 36065
rect 68427 36016 68428 36056
rect 68468 36016 68469 36056
rect 68427 36007 68469 36016
rect 68235 35468 68277 35477
rect 68235 35428 68236 35468
rect 68276 35428 68277 35468
rect 68235 35419 68277 35428
rect 68139 35384 68181 35393
rect 68139 35344 68140 35384
rect 68180 35344 68181 35384
rect 68139 35335 68181 35344
rect 68428 35216 68468 36007
rect 68524 35216 68564 35225
rect 68428 35176 68524 35216
rect 68524 35167 68564 35176
rect 68812 34889 68852 36679
rect 68908 36560 68948 38107
rect 69100 37988 69140 37997
rect 69100 37409 69140 37948
rect 69099 37400 69141 37409
rect 69099 37360 69100 37400
rect 69140 37360 69141 37400
rect 69099 37351 69141 37360
rect 69196 37316 69236 37325
rect 69196 37232 69236 37276
rect 69100 37192 69236 37232
rect 69100 36980 69140 37192
rect 69292 37148 69332 38191
rect 70636 38106 70676 38191
rect 71020 38165 71060 38200
rect 71212 38240 71252 38249
rect 74283 38240 74325 38249
rect 71252 38200 71732 38240
rect 71212 38191 71252 38200
rect 71019 38156 71061 38165
rect 71019 38116 71020 38156
rect 71060 38116 71061 38156
rect 71019 38107 71061 38116
rect 71404 38072 71444 38081
rect 69387 37988 69429 37997
rect 69387 37948 69388 37988
rect 69428 37948 69429 37988
rect 69387 37939 69429 37948
rect 70060 37988 70100 37997
rect 68908 36511 68948 36520
rect 69004 36940 69140 36980
rect 69196 37108 69332 37148
rect 69004 36476 69044 36940
rect 69100 36737 69140 36822
rect 69099 36728 69141 36737
rect 69099 36688 69100 36728
rect 69140 36688 69141 36728
rect 69099 36679 69141 36688
rect 69100 36476 69140 36485
rect 69004 36436 69100 36476
rect 69100 36427 69140 36436
rect 69099 35888 69141 35897
rect 69099 35848 69100 35888
rect 69140 35848 69141 35888
rect 69099 35839 69141 35848
rect 68811 34880 68853 34889
rect 68811 34840 68812 34880
rect 68852 34840 68853 34880
rect 68811 34831 68853 34840
rect 68811 34628 68853 34637
rect 68811 34588 68812 34628
rect 68852 34588 68853 34628
rect 68811 34579 68853 34588
rect 68812 34494 68852 34579
rect 68044 33100 68564 33140
rect 69100 33125 69140 35839
rect 69196 33965 69236 37108
rect 69388 37064 69428 37939
rect 69580 37400 69620 37409
rect 69580 37241 69620 37360
rect 69579 37232 69621 37241
rect 69579 37192 69580 37232
rect 69620 37192 69621 37232
rect 69579 37183 69621 37192
rect 69292 37024 69428 37064
rect 69292 36728 69332 37024
rect 69579 36812 69621 36821
rect 69579 36772 69580 36812
rect 69620 36772 69621 36812
rect 69579 36763 69621 36772
rect 69292 36679 69332 36688
rect 69388 36728 69428 36737
rect 69388 36560 69428 36688
rect 69580 36728 69620 36763
rect 69580 36677 69620 36688
rect 69772 36728 69812 36737
rect 69676 36560 69716 36569
rect 69388 36520 69676 36560
rect 69676 36511 69716 36520
rect 69483 36056 69525 36065
rect 69772 36056 69812 36688
rect 69483 36016 69484 36056
rect 69524 36016 69525 36056
rect 69483 36007 69525 36016
rect 69580 36016 69812 36056
rect 69484 35922 69524 36007
rect 69580 35645 69620 36016
rect 69675 35888 69717 35897
rect 69675 35848 69676 35888
rect 69716 35848 69717 35888
rect 69675 35839 69717 35848
rect 69868 35888 69908 35897
rect 69676 35754 69716 35839
rect 69771 35804 69813 35813
rect 69771 35764 69772 35804
rect 69812 35764 69813 35804
rect 69771 35755 69813 35764
rect 69772 35670 69812 35755
rect 69868 35729 69908 35848
rect 69963 35888 70005 35897
rect 69963 35848 69964 35888
rect 70004 35848 70005 35888
rect 69963 35839 70005 35848
rect 69964 35754 70004 35839
rect 69867 35720 69909 35729
rect 69867 35680 69868 35720
rect 69908 35680 69909 35720
rect 69867 35671 69909 35680
rect 69291 35636 69333 35645
rect 69291 35596 69292 35636
rect 69332 35596 69333 35636
rect 69291 35587 69333 35596
rect 69579 35636 69621 35645
rect 69579 35596 69580 35636
rect 69620 35596 69621 35636
rect 69579 35587 69621 35596
rect 69195 33956 69237 33965
rect 69195 33916 69196 33956
rect 69236 33916 69237 33956
rect 69195 33907 69237 33916
rect 67564 32864 67604 33100
rect 67564 32815 67604 32824
rect 67947 32192 67989 32201
rect 67947 32152 67948 32192
rect 67988 32152 67989 32192
rect 67947 32143 67989 32152
rect 67948 32058 67988 32143
rect 66796 31144 67412 31184
rect 68235 30764 68277 30773
rect 68235 30724 68236 30764
rect 68276 30724 68277 30764
rect 68235 30715 68277 30724
rect 65644 30556 65780 30596
rect 65836 30680 65876 30689
rect 65452 30428 65492 30437
rect 65452 30185 65492 30388
rect 65451 30176 65493 30185
rect 65451 30136 65452 30176
rect 65492 30136 65588 30176
rect 65451 30127 65493 30136
rect 65452 29840 65492 29849
rect 65452 29681 65492 29800
rect 65548 29840 65588 30136
rect 65548 29791 65588 29800
rect 65451 29672 65493 29681
rect 65451 29632 65452 29672
rect 65492 29632 65493 29672
rect 65451 29623 65493 29632
rect 65644 29168 65684 30556
rect 65740 30428 65780 30437
rect 65740 29849 65780 30388
rect 65836 30092 65876 30640
rect 66027 30680 66069 30689
rect 66027 30640 66028 30680
rect 66068 30640 66069 30680
rect 66027 30631 66069 30640
rect 66220 30680 66260 30689
rect 66028 30546 66068 30631
rect 66124 30428 66164 30437
rect 65836 30043 65876 30052
rect 65932 30388 66124 30428
rect 65739 29840 65781 29849
rect 65739 29800 65740 29840
rect 65780 29800 65876 29840
rect 65739 29791 65781 29800
rect 65740 29706 65780 29791
rect 65355 29084 65397 29093
rect 65355 29044 65356 29084
rect 65396 29044 65397 29084
rect 65355 29035 65397 29044
rect 65547 29084 65589 29093
rect 65547 29044 65548 29084
rect 65588 29044 65589 29084
rect 65547 29035 65589 29044
rect 65260 28531 65300 28540
rect 65164 28120 65396 28160
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 65163 27824 65205 27833
rect 65163 27784 65164 27824
rect 65204 27784 65205 27824
rect 65163 27775 65205 27784
rect 65164 27656 65204 27775
rect 65259 27740 65301 27749
rect 65259 27700 65260 27740
rect 65300 27700 65301 27740
rect 65259 27691 65301 27700
rect 65164 27607 65204 27616
rect 65260 27606 65300 27691
rect 65356 27665 65396 28120
rect 65355 27656 65397 27665
rect 65355 27616 65356 27656
rect 65396 27616 65397 27656
rect 65355 27607 65397 27616
rect 65452 27656 65492 27667
rect 64491 27572 64533 27581
rect 64491 27532 64492 27572
rect 64532 27532 64533 27572
rect 64491 27523 64533 27532
rect 64395 27404 64437 27413
rect 64395 27364 64396 27404
rect 64436 27364 64437 27404
rect 64395 27355 64437 27364
rect 64492 27236 64532 27523
rect 65356 27522 65396 27607
rect 65452 27581 65492 27616
rect 65451 27572 65493 27581
rect 65451 27532 65452 27572
rect 65492 27532 65493 27572
rect 65451 27523 65493 27532
rect 65259 27404 65301 27413
rect 65259 27364 65260 27404
rect 65300 27364 65301 27404
rect 65259 27355 65301 27364
rect 64396 27196 64532 27236
rect 64299 27152 64341 27161
rect 64204 27112 64300 27152
rect 64340 27112 64341 27152
rect 64299 27103 64341 27112
rect 63860 27028 64052 27068
rect 63820 27019 63860 27028
rect 63819 26816 63861 26825
rect 64012 26816 64052 26825
rect 63819 26776 63820 26816
rect 63860 26776 63861 26816
rect 63819 26767 63861 26776
rect 63916 26776 64012 26816
rect 63820 26153 63860 26767
rect 63819 26144 63861 26153
rect 63819 26104 63820 26144
rect 63860 26104 63861 26144
rect 63819 26095 63861 26104
rect 63916 25901 63956 26776
rect 64012 26767 64052 26776
rect 64108 26816 64148 26825
rect 63915 25892 63957 25901
rect 63915 25852 63916 25892
rect 63956 25852 63957 25892
rect 63915 25843 63957 25852
rect 64012 25892 64052 25901
rect 64108 25892 64148 26776
rect 64204 26144 64244 26153
rect 64204 25892 64244 26104
rect 64300 26144 64340 27103
rect 64300 26095 64340 26104
rect 64396 26144 64436 27196
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 64779 26228 64821 26237
rect 64779 26188 64780 26228
rect 64820 26188 64821 26228
rect 64779 26179 64821 26188
rect 64396 26095 64436 26104
rect 64492 26144 64532 26153
rect 64492 26060 64532 26104
rect 64684 26133 64724 26142
rect 64780 26094 64820 26179
rect 64876 26144 64916 26153
rect 64684 26060 64724 26093
rect 64492 26020 64724 26060
rect 64052 25852 64244 25892
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 64012 25565 64052 25852
rect 63531 25556 63573 25565
rect 63531 25516 63532 25556
rect 63572 25516 63573 25556
rect 63531 25507 63573 25516
rect 64011 25556 64053 25565
rect 64011 25516 64012 25556
rect 64052 25516 64053 25556
rect 64011 25507 64053 25516
rect 63435 25472 63477 25481
rect 63435 25432 63436 25472
rect 63476 25432 63477 25472
rect 63435 25423 63477 25432
rect 62859 25304 62901 25313
rect 62859 25264 62860 25304
rect 62900 25264 62901 25304
rect 62859 25255 62901 25264
rect 63148 25304 63188 25315
rect 63148 25229 63188 25264
rect 63436 25304 63476 25313
rect 63147 25220 63189 25229
rect 63147 25180 63148 25220
rect 63188 25180 63189 25220
rect 63147 25171 63189 25180
rect 62668 25136 62708 25145
rect 62668 24809 62708 25096
rect 63436 25061 63476 25264
rect 63532 25304 63572 25507
rect 63723 25472 63765 25481
rect 63723 25432 63724 25472
rect 63764 25432 63765 25472
rect 63723 25423 63765 25432
rect 63820 25472 63860 25481
rect 63627 25388 63669 25397
rect 63627 25348 63628 25388
rect 63668 25348 63669 25388
rect 63627 25339 63669 25348
rect 63532 25255 63572 25264
rect 63435 25052 63477 25061
rect 63435 25012 63436 25052
rect 63476 25012 63477 25052
rect 63435 25003 63477 25012
rect 62667 24800 62709 24809
rect 62667 24760 62668 24800
rect 62708 24760 62709 24800
rect 62667 24751 62709 24760
rect 62571 24464 62613 24473
rect 62571 24424 62572 24464
rect 62612 24424 62613 24464
rect 62571 24415 62613 24424
rect 63051 24464 63093 24473
rect 63051 24424 63052 24464
rect 63092 24424 63093 24464
rect 63051 24415 63093 24424
rect 62475 24380 62517 24389
rect 62475 24340 62476 24380
rect 62516 24340 62517 24380
rect 62475 24331 62517 24340
rect 62955 24296 62997 24305
rect 62955 24256 62956 24296
rect 62996 24256 62997 24296
rect 62955 24247 62997 24256
rect 62859 24212 62901 24221
rect 62859 24172 62860 24212
rect 62900 24172 62901 24212
rect 62859 24163 62901 24172
rect 62091 24044 62133 24053
rect 62091 24004 62092 24044
rect 62132 24004 62133 24044
rect 62091 23995 62133 24004
rect 62283 24044 62325 24053
rect 62283 24004 62284 24044
rect 62324 24004 62325 24044
rect 62283 23995 62325 24004
rect 62092 23792 62132 23995
rect 62475 23876 62517 23885
rect 62475 23836 62476 23876
rect 62516 23836 62517 23876
rect 62475 23827 62517 23836
rect 62763 23876 62805 23885
rect 62763 23836 62764 23876
rect 62804 23836 62805 23876
rect 62763 23827 62805 23836
rect 62476 23792 62516 23827
rect 60364 23752 60460 23792
rect 60500 23752 60692 23792
rect 60076 23549 60116 23752
rect 60460 23743 60500 23752
rect 60172 23624 60212 23633
rect 60075 23540 60117 23549
rect 60075 23500 60076 23540
rect 60116 23500 60117 23540
rect 60075 23491 60117 23500
rect 60172 23060 60212 23584
rect 60556 23624 60596 23633
rect 59212 23020 59295 23060
rect 59404 23020 59540 23060
rect 59596 23020 59695 23060
rect 59788 23020 59924 23060
rect 59980 23020 60095 23060
rect 60172 23020 60385 23060
rect 59116 22744 59185 22784
rect 59145 22596 59185 22744
rect 59255 22596 59295 23020
rect 59500 22784 59540 23020
rect 59500 22744 59585 22784
rect 59545 22596 59585 22744
rect 59655 22596 59695 23020
rect 59884 22784 59924 23020
rect 59884 22744 59985 22784
rect 59945 22596 59985 22744
rect 60055 22596 60095 23020
rect 60345 22596 60385 23020
rect 60454 22784 60496 22793
rect 60556 22784 60596 23584
rect 60652 23060 60692 23752
rect 60884 23752 61268 23792
rect 60844 23743 60884 23752
rect 60940 23624 60980 23633
rect 60940 23060 60980 23584
rect 61228 23060 61268 23752
rect 61364 23752 61652 23792
rect 61324 23743 61364 23752
rect 61420 23624 61460 23633
rect 61420 23060 61460 23584
rect 61612 23060 61652 23752
rect 61748 23752 62036 23792
rect 61708 23743 61748 23752
rect 61804 23624 61844 23633
rect 61804 23060 61844 23584
rect 61996 23060 62036 23752
rect 62132 23752 62420 23792
rect 62092 23743 62132 23752
rect 62188 23624 62228 23633
rect 62188 23060 62228 23584
rect 62380 23060 62420 23752
rect 62476 23741 62516 23752
rect 62572 23624 62612 23633
rect 62572 23060 62612 23584
rect 62764 23060 62804 23827
rect 62860 23792 62900 24163
rect 62956 23885 62996 24247
rect 63052 23969 63092 24415
rect 63051 23960 63093 23969
rect 63051 23920 63052 23960
rect 63092 23920 63093 23960
rect 63051 23911 63093 23920
rect 62955 23876 62997 23885
rect 62955 23836 62956 23876
rect 62996 23836 62997 23876
rect 62955 23827 62997 23836
rect 62860 23465 62900 23752
rect 63244 23792 63284 23801
rect 63244 23633 63284 23752
rect 63628 23792 63668 25339
rect 63724 24464 63764 25423
rect 63820 24641 63860 25432
rect 64396 25304 64436 25313
rect 64436 25264 64724 25304
rect 64396 25255 64436 25264
rect 64012 25220 64052 25229
rect 63915 25136 63957 25145
rect 63915 25096 63916 25136
rect 63956 25096 63957 25136
rect 63915 25087 63957 25096
rect 63819 24632 63861 24641
rect 63819 24592 63820 24632
rect 63860 24592 63861 24632
rect 63819 24583 63861 24592
rect 63916 24632 63956 25087
rect 64012 24800 64052 25180
rect 64587 25052 64629 25061
rect 64587 25012 64588 25052
rect 64628 25012 64629 25052
rect 64587 25003 64629 25012
rect 64012 24751 64052 24760
rect 64204 24760 64532 24800
rect 64107 24716 64149 24725
rect 64107 24676 64108 24716
rect 64148 24676 64149 24716
rect 64107 24667 64149 24676
rect 63916 24583 63956 24592
rect 64108 24632 64148 24667
rect 64108 24581 64148 24592
rect 64204 24632 64244 24760
rect 64492 24716 64532 24760
rect 64492 24667 64532 24676
rect 64204 24583 64244 24592
rect 64396 24632 64436 24643
rect 64396 24557 64436 24592
rect 64588 24632 64628 25003
rect 64588 24583 64628 24592
rect 64395 24548 64437 24557
rect 64395 24508 64396 24548
rect 64436 24508 64437 24548
rect 64395 24499 64437 24508
rect 64684 24473 64724 25264
rect 64876 25136 64916 26104
rect 64972 26144 65012 26153
rect 64972 25985 65012 26104
rect 64971 25976 65013 25985
rect 64971 25936 64972 25976
rect 65012 25936 65013 25976
rect 64971 25927 65013 25936
rect 65260 25304 65300 27355
rect 65548 26321 65588 29035
rect 65644 27833 65684 29128
rect 65740 29252 65780 29261
rect 65740 29000 65780 29212
rect 65836 29168 65876 29800
rect 65836 29119 65876 29128
rect 65932 29168 65972 30388
rect 66124 30379 66164 30388
rect 66220 30260 66260 30640
rect 68236 30630 68276 30715
rect 66508 30512 66548 30521
rect 66220 30220 66261 30260
rect 66221 30176 66261 30220
rect 66220 30136 66261 30176
rect 65932 29119 65972 29128
rect 66028 29756 66068 29765
rect 66028 29000 66068 29716
rect 66220 29681 66260 30136
rect 66412 29840 66452 29849
rect 66508 29840 66548 30472
rect 66603 30344 66645 30353
rect 66603 30304 66604 30344
rect 66644 30304 66645 30344
rect 66603 30295 66645 30304
rect 66452 29800 66548 29840
rect 66412 29791 66452 29800
rect 66219 29672 66261 29681
rect 66219 29632 66220 29672
rect 66260 29632 66261 29672
rect 66219 29623 66261 29632
rect 65740 28960 66068 29000
rect 66124 28328 66164 28337
rect 65740 28244 65780 28253
rect 65643 27824 65685 27833
rect 65643 27784 65644 27824
rect 65684 27784 65685 27824
rect 65643 27775 65685 27784
rect 65740 27749 65780 28204
rect 65835 28160 65877 28169
rect 65835 28120 65836 28160
rect 65876 28120 65877 28160
rect 65835 28111 65877 28120
rect 65739 27740 65781 27749
rect 65739 27700 65740 27740
rect 65780 27700 65781 27740
rect 65739 27691 65781 27700
rect 65644 27656 65684 27665
rect 65355 26312 65397 26321
rect 65355 26272 65356 26312
rect 65396 26272 65397 26312
rect 65355 26263 65397 26272
rect 65547 26312 65589 26321
rect 65547 26272 65548 26312
rect 65588 26272 65589 26312
rect 65547 26263 65589 26272
rect 65260 25255 65300 25264
rect 64876 25096 65300 25136
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 65260 24725 65300 25096
rect 64875 24716 64917 24725
rect 64875 24676 64876 24716
rect 64916 24676 64917 24716
rect 64875 24667 64917 24676
rect 65259 24716 65301 24725
rect 65259 24676 65260 24716
rect 65300 24676 65301 24716
rect 65259 24667 65301 24676
rect 64779 24632 64821 24641
rect 64779 24592 64780 24632
rect 64820 24592 64821 24632
rect 64779 24583 64821 24592
rect 64780 24498 64820 24583
rect 64876 24582 64916 24667
rect 65356 24641 65396 26263
rect 65452 26153 65492 26238
rect 65451 26144 65493 26153
rect 65451 26104 65452 26144
rect 65492 26104 65493 26144
rect 65451 26095 65493 26104
rect 65644 26144 65684 27616
rect 65836 27656 65876 28111
rect 65931 27824 65973 27833
rect 65931 27784 65932 27824
rect 65972 27784 65973 27824
rect 65931 27775 65973 27784
rect 65836 27607 65876 27616
rect 65739 27572 65781 27581
rect 65739 27532 65740 27572
rect 65780 27532 65781 27572
rect 65739 27523 65781 27532
rect 65740 27438 65780 27523
rect 65740 26648 65780 26657
rect 65740 26153 65780 26608
rect 65451 25976 65493 25985
rect 65451 25936 65452 25976
rect 65492 25936 65493 25976
rect 65451 25927 65493 25936
rect 65452 25842 65492 25927
rect 65644 25901 65684 26104
rect 65739 26144 65781 26153
rect 65739 26104 65740 26144
rect 65780 26104 65781 26144
rect 65739 26095 65781 26104
rect 65740 26010 65780 26095
rect 65643 25892 65685 25901
rect 65643 25852 65644 25892
rect 65684 25852 65685 25892
rect 65643 25843 65685 25852
rect 64971 24632 65013 24641
rect 64971 24592 64972 24632
rect 65012 24592 65013 24632
rect 64971 24583 65013 24592
rect 65355 24632 65397 24641
rect 65355 24592 65356 24632
rect 65396 24592 65397 24632
rect 65355 24583 65397 24592
rect 64972 24498 65012 24583
rect 65644 24557 65684 25843
rect 65932 25145 65972 27775
rect 66124 27488 66164 28288
rect 66220 27488 66260 27497
rect 66124 27448 66220 27488
rect 66220 27439 66260 27448
rect 66411 26816 66453 26825
rect 66411 26776 66412 26816
rect 66452 26776 66453 26816
rect 66411 26767 66453 26776
rect 66412 25976 66452 26767
rect 66412 25927 66452 25936
rect 65931 25136 65973 25145
rect 65931 25096 65932 25136
rect 65972 25096 65973 25136
rect 65931 25087 65973 25096
rect 66412 25136 66452 25145
rect 65932 24641 65972 25087
rect 66412 25061 66452 25096
rect 66411 25052 66453 25061
rect 66411 25012 66412 25052
rect 66452 25012 66453 25052
rect 66411 25003 66453 25012
rect 66412 24725 66452 25003
rect 66411 24716 66453 24725
rect 66411 24676 66412 24716
rect 66452 24676 66453 24716
rect 66411 24667 66453 24676
rect 65931 24632 65973 24641
rect 65931 24592 65932 24632
rect 65972 24592 65973 24632
rect 65931 24583 65973 24592
rect 65643 24548 65685 24557
rect 65643 24508 65644 24548
rect 65684 24508 65685 24548
rect 65643 24499 65685 24508
rect 64683 24464 64725 24473
rect 63724 24424 64148 24464
rect 64108 23792 64148 24424
rect 64683 24424 64684 24464
rect 64724 24424 64725 24464
rect 64683 24415 64725 24424
rect 65163 24464 65205 24473
rect 65163 24424 65164 24464
rect 65204 24424 65205 24464
rect 65163 24415 65205 24424
rect 65164 24330 65204 24415
rect 66123 24380 66165 24389
rect 66123 24340 66124 24380
rect 66164 24340 66165 24380
rect 66123 24331 66165 24340
rect 65739 24128 65781 24137
rect 65739 24088 65740 24128
rect 65780 24088 65781 24128
rect 65739 24079 65781 24088
rect 65259 24044 65301 24053
rect 65259 24004 65260 24044
rect 65300 24004 65301 24044
rect 65259 23995 65301 24004
rect 65643 24044 65685 24053
rect 65643 24004 65644 24044
rect 65684 24004 65685 24044
rect 65643 23995 65685 24004
rect 64875 23960 64917 23969
rect 64875 23920 64876 23960
rect 64916 23920 64917 23960
rect 64875 23911 64917 23920
rect 65163 23960 65205 23969
rect 65163 23920 65164 23960
rect 65204 23920 65205 23960
rect 65163 23911 65205 23920
rect 64491 23876 64533 23885
rect 64491 23836 64492 23876
rect 64532 23836 64533 23876
rect 64491 23827 64533 23836
rect 64779 23876 64821 23885
rect 64779 23836 64780 23876
rect 64820 23836 64821 23876
rect 64779 23827 64821 23836
rect 64492 23792 64532 23827
rect 63668 23752 64052 23792
rect 63628 23743 63668 23752
rect 62956 23624 62996 23633
rect 62859 23456 62901 23465
rect 62859 23416 62860 23456
rect 62900 23416 62901 23456
rect 62859 23407 62901 23416
rect 62956 23060 62996 23584
rect 63243 23624 63285 23633
rect 63243 23584 63244 23624
rect 63284 23584 63285 23624
rect 63243 23575 63285 23584
rect 63340 23624 63380 23633
rect 63627 23624 63669 23633
rect 63380 23584 63476 23624
rect 63340 23575 63380 23584
rect 63243 23456 63285 23465
rect 63243 23416 63244 23456
rect 63284 23416 63285 23456
rect 63243 23407 63285 23416
rect 63244 23060 63284 23407
rect 63436 23060 63476 23584
rect 63627 23584 63628 23624
rect 63668 23584 63669 23624
rect 63627 23575 63669 23584
rect 63724 23624 63764 23633
rect 63764 23584 63956 23624
rect 63724 23575 63764 23584
rect 63628 23060 63668 23575
rect 60652 23020 60895 23060
rect 60940 23020 61185 23060
rect 61228 23020 61295 23060
rect 61420 23020 61556 23060
rect 61612 23020 61695 23060
rect 61804 23020 61940 23060
rect 61996 23020 62095 23060
rect 62188 23020 62324 23060
rect 62380 23020 62495 23060
rect 62572 23020 62708 23060
rect 62764 23020 62895 23060
rect 62956 23020 63185 23060
rect 63244 23020 63295 23060
rect 63436 23020 63585 23060
rect 63628 23020 63695 23060
rect 60454 22744 60455 22784
rect 60495 22744 60500 22784
rect 60556 22744 60785 22784
rect 60454 22735 60500 22744
rect 60460 22280 60500 22735
rect 60745 22596 60785 22744
rect 60855 22596 60895 23020
rect 61145 22596 61185 23020
rect 61255 22596 61295 23020
rect 61516 22784 61556 23020
rect 61516 22744 61585 22784
rect 61545 22596 61585 22744
rect 61655 22596 61695 23020
rect 61900 22784 61940 23020
rect 61900 22744 61985 22784
rect 61945 22596 61985 22744
rect 62055 22596 62095 23020
rect 62284 22784 62324 23020
rect 62284 22744 62385 22784
rect 62345 22596 62385 22744
rect 62455 22596 62495 23020
rect 62668 22784 62708 23020
rect 62668 22744 62785 22784
rect 62745 22596 62785 22744
rect 62855 22596 62895 23020
rect 63145 22596 63185 23020
rect 63255 22596 63295 23020
rect 63545 22596 63585 23020
rect 63655 22596 63695 23020
rect 63916 22784 63956 23584
rect 64012 23060 64052 23752
rect 64148 23752 64436 23792
rect 64108 23743 64148 23752
rect 64204 23624 64244 23633
rect 64204 23060 64244 23584
rect 64396 23060 64436 23752
rect 64492 23741 64532 23752
rect 64588 23624 64628 23633
rect 64588 23060 64628 23584
rect 64780 23060 64820 23827
rect 64876 23792 64916 23911
rect 64876 23743 64916 23752
rect 64972 23624 65012 23633
rect 64972 23060 65012 23584
rect 65164 23060 65204 23911
rect 65260 23792 65300 23995
rect 65260 23743 65300 23752
rect 65356 23624 65396 23633
rect 65356 23060 65396 23584
rect 65644 23060 65684 23995
rect 65740 23792 65780 24079
rect 66124 23792 66164 24331
rect 66508 23792 66548 23801
rect 66604 23792 66644 30295
rect 67276 29840 67316 29849
rect 66795 28664 66837 28673
rect 66795 28624 66796 28664
rect 66836 28624 66837 28664
rect 66795 28615 66837 28624
rect 66796 23792 66836 28615
rect 67276 28337 67316 29800
rect 68427 29672 68469 29681
rect 68427 29632 68428 29672
rect 68468 29632 68469 29672
rect 68427 29623 68469 29632
rect 67755 29252 67797 29261
rect 67755 29212 67756 29252
rect 67796 29212 67797 29252
rect 67755 29203 67797 29212
rect 67756 29118 67796 29203
rect 68140 29168 68180 29177
rect 68140 28496 68180 29128
rect 68428 29093 68468 29623
rect 68427 29084 68469 29093
rect 68427 29044 68428 29084
rect 68468 29044 68469 29084
rect 68427 29035 68469 29044
rect 68427 28580 68469 28589
rect 68427 28540 68428 28580
rect 68468 28540 68469 28580
rect 68427 28531 68469 28540
rect 68332 28496 68372 28505
rect 68140 28456 68332 28496
rect 68332 28447 68372 28456
rect 66987 28328 67029 28337
rect 66892 28288 66988 28328
rect 67028 28288 67029 28328
rect 66892 27413 66932 28288
rect 66987 28279 67029 28288
rect 67275 28328 67317 28337
rect 67275 28288 67276 28328
rect 67316 28288 67317 28328
rect 67275 28279 67317 28288
rect 66988 28194 67028 28279
rect 68139 28160 68181 28169
rect 68139 28120 68140 28160
rect 68180 28120 68181 28160
rect 68139 28111 68181 28120
rect 68140 28026 68180 28111
rect 68331 27824 68373 27833
rect 68331 27784 68332 27824
rect 68372 27784 68373 27824
rect 68331 27775 68373 27784
rect 67564 27572 67604 27581
rect 66891 27404 66933 27413
rect 67372 27404 67412 27413
rect 66891 27364 66892 27404
rect 66932 27364 66933 27404
rect 66891 27355 66933 27364
rect 67276 27364 67372 27404
rect 66892 26816 66932 27355
rect 66892 26767 66932 26776
rect 67276 26237 67316 27364
rect 67372 27355 67412 27364
rect 67564 26993 67604 27532
rect 67659 27320 67701 27329
rect 67659 27280 67660 27320
rect 67700 27280 67701 27320
rect 67659 27271 67701 27280
rect 67563 26984 67605 26993
rect 67563 26944 67564 26984
rect 67604 26944 67605 26984
rect 67563 26935 67605 26944
rect 67660 26657 67700 27271
rect 67755 26816 67797 26825
rect 67755 26776 67756 26816
rect 67796 26776 67797 26816
rect 67755 26767 67797 26776
rect 68332 26816 68372 27775
rect 68428 27749 68468 28531
rect 68427 27740 68469 27749
rect 68427 27700 68428 27740
rect 68468 27700 68469 27740
rect 68427 27691 68469 27700
rect 68428 27572 68468 27691
rect 68428 27523 68468 27532
rect 68524 26984 68564 33100
rect 69099 33116 69141 33125
rect 69099 33076 69100 33116
rect 69140 33076 69236 33116
rect 69099 33067 69141 33076
rect 69196 32875 69236 33076
rect 68908 32864 68948 32873
rect 68908 32705 68948 32824
rect 69003 32864 69045 32873
rect 69003 32824 69004 32864
rect 69044 32824 69045 32864
rect 69196 32826 69236 32835
rect 69003 32815 69045 32824
rect 69004 32730 69044 32815
rect 69292 32780 69332 35587
rect 69580 35132 69620 35587
rect 69963 35384 70005 35393
rect 69963 35344 69964 35384
rect 70004 35344 70005 35384
rect 69963 35335 70005 35344
rect 69580 35092 69812 35132
rect 69675 34964 69717 34973
rect 69675 34924 69676 34964
rect 69716 34924 69717 34964
rect 69675 34915 69717 34924
rect 69676 34830 69716 34915
rect 69772 34889 69812 35092
rect 69771 34880 69813 34889
rect 69771 34840 69772 34880
rect 69812 34840 69813 34880
rect 69771 34831 69813 34840
rect 69579 34796 69621 34805
rect 69579 34756 69580 34796
rect 69620 34756 69621 34796
rect 69579 34747 69621 34756
rect 69196 32740 69332 32780
rect 69388 32780 69428 32789
rect 68715 32696 68757 32705
rect 68715 32656 68716 32696
rect 68756 32656 68757 32696
rect 68715 32647 68757 32656
rect 68907 32696 68949 32705
rect 68907 32656 68908 32696
rect 68948 32656 68949 32696
rect 68907 32647 68949 32656
rect 69099 32696 69141 32705
rect 69099 32656 69100 32696
rect 69140 32656 69141 32696
rect 69099 32647 69141 32656
rect 68716 32562 68756 32647
rect 69100 32562 69140 32647
rect 68811 32444 68853 32453
rect 68811 32404 68812 32444
rect 68852 32404 68853 32444
rect 68811 32395 68853 32404
rect 68716 31520 68756 31529
rect 68620 31480 68716 31520
rect 68620 30680 68660 31480
rect 68716 31471 68756 31480
rect 68620 30631 68660 30640
rect 68619 27824 68661 27833
rect 68619 27784 68620 27824
rect 68660 27784 68661 27824
rect 68619 27775 68661 27784
rect 68620 27690 68660 27775
rect 68524 26944 68756 26984
rect 68332 26767 68372 26776
rect 68524 26816 68564 26825
rect 67756 26682 67796 26767
rect 68140 26732 68180 26741
rect 67852 26692 68140 26732
rect 67659 26648 67701 26657
rect 67659 26608 67660 26648
rect 67700 26608 67701 26648
rect 67659 26599 67701 26608
rect 67371 26396 67413 26405
rect 67371 26356 67372 26396
rect 67412 26356 67413 26396
rect 67371 26347 67413 26356
rect 67275 26228 67317 26237
rect 67275 26188 67276 26228
rect 67316 26188 67317 26228
rect 67275 26179 67317 26188
rect 67179 26144 67221 26153
rect 67179 26104 67180 26144
rect 67220 26104 67221 26144
rect 67179 26095 67221 26104
rect 67276 26144 67316 26179
rect 67180 25976 67220 26095
rect 67276 26093 67316 26104
rect 67372 26144 67412 26347
rect 67756 26312 67796 26321
rect 67852 26312 67892 26692
rect 68140 26683 68180 26692
rect 68428 26648 68468 26657
rect 68236 26608 68428 26648
rect 68236 26396 68276 26608
rect 68428 26599 68468 26608
rect 68427 26480 68469 26489
rect 68427 26440 68428 26480
rect 68468 26440 68469 26480
rect 68427 26431 68469 26440
rect 67796 26272 67892 26312
rect 67948 26356 68276 26396
rect 67756 26263 67796 26272
rect 67372 26095 67412 26104
rect 67468 26144 67508 26153
rect 67660 26144 67700 26153
rect 67508 26104 67660 26144
rect 67468 26095 67508 26104
rect 67660 26095 67700 26104
rect 67852 26144 67892 26153
rect 67180 25936 67508 25976
rect 67084 25304 67124 25315
rect 67084 25229 67124 25264
rect 67372 25304 67412 25313
rect 67083 25220 67125 25229
rect 67083 25180 67084 25220
rect 67124 25180 67125 25220
rect 67083 25171 67125 25180
rect 67372 25145 67412 25264
rect 67468 25304 67508 25936
rect 67852 25892 67892 26104
rect 67948 26144 67988 26356
rect 68235 26228 68277 26237
rect 67948 26095 67988 26104
rect 68140 26188 68236 26228
rect 68276 26188 68277 26228
rect 68140 26144 68180 26188
rect 68235 26179 68277 26188
rect 68140 26095 68180 26104
rect 68332 26144 68372 26153
rect 68236 25892 68276 25901
rect 67852 25852 68236 25892
rect 67852 25724 67892 25852
rect 68236 25843 68276 25852
rect 67468 25255 67508 25264
rect 67660 25684 67892 25724
rect 67371 25136 67413 25145
rect 67371 25096 67372 25136
rect 67412 25096 67413 25136
rect 67371 25087 67413 25096
rect 67660 25061 67700 25684
rect 67756 25556 67796 25565
rect 68332 25556 68372 26104
rect 67796 25516 68372 25556
rect 67756 25507 67796 25516
rect 68332 25313 68372 25398
rect 68331 25304 68373 25313
rect 68331 25264 68332 25304
rect 68372 25264 68373 25304
rect 68331 25255 68373 25264
rect 67948 25220 67988 25229
rect 67756 25180 67948 25220
rect 67659 25052 67701 25061
rect 67659 25012 67660 25052
rect 67700 25012 67701 25052
rect 67659 25003 67701 25012
rect 67563 24800 67605 24809
rect 67563 24760 67564 24800
rect 67604 24760 67605 24800
rect 67563 24751 67605 24760
rect 67756 24800 67796 25180
rect 67948 25171 67988 25180
rect 67851 25052 67893 25061
rect 67851 25012 67852 25052
rect 67892 25012 67893 25052
rect 67851 25003 67893 25012
rect 68331 25052 68373 25061
rect 68331 25012 68332 25052
rect 68372 25012 68373 25052
rect 68331 25003 68373 25012
rect 67756 24751 67796 24760
rect 67564 23960 67604 24751
rect 67659 24632 67701 24641
rect 67659 24592 67660 24632
rect 67700 24592 67701 24632
rect 67659 24583 67701 24592
rect 67852 24632 67892 25003
rect 67852 24583 67892 24592
rect 67948 24760 68276 24800
rect 67948 24632 67988 24760
rect 68236 24716 68276 24760
rect 68236 24667 68276 24676
rect 67948 24583 67988 24592
rect 68139 24632 68181 24641
rect 68139 24592 68140 24632
rect 68180 24592 68181 24632
rect 68139 24583 68181 24592
rect 68332 24632 68372 25003
rect 68332 24583 68372 24592
rect 67660 24498 67700 24583
rect 68140 24498 68180 24583
rect 67564 23920 67700 23960
rect 66892 23792 66932 23801
rect 67275 23792 67317 23801
rect 65780 23752 66068 23792
rect 65740 23743 65780 23752
rect 65836 23624 65876 23633
rect 65836 23060 65876 23584
rect 66028 23060 66068 23752
rect 66164 23752 66452 23792
rect 66124 23743 66164 23752
rect 66220 23624 66260 23633
rect 66220 23060 66260 23584
rect 66412 23060 66452 23752
rect 66548 23752 66740 23792
rect 66796 23752 66892 23792
rect 66932 23752 67220 23792
rect 66508 23743 66548 23752
rect 66604 23624 66644 23633
rect 66604 23060 66644 23584
rect 66700 23204 66740 23752
rect 66892 23743 66932 23752
rect 66988 23624 67028 23633
rect 66700 23164 66836 23204
rect 66796 23060 66836 23164
rect 66988 23060 67028 23584
rect 67180 23060 67220 23752
rect 67275 23752 67276 23792
rect 67316 23752 67317 23792
rect 67275 23743 67317 23752
rect 67563 23792 67605 23801
rect 67563 23752 67564 23792
rect 67604 23752 67605 23792
rect 67563 23743 67605 23752
rect 67660 23792 67700 23920
rect 67276 23658 67316 23743
rect 67372 23624 67412 23633
rect 67372 23060 67412 23584
rect 67564 23060 67604 23743
rect 67660 23717 67700 23752
rect 68140 23792 68180 23801
rect 68428 23792 68468 26431
rect 68524 25976 68564 26776
rect 68619 26816 68661 26825
rect 68619 26776 68620 26816
rect 68660 26776 68661 26816
rect 68619 26767 68661 26776
rect 68620 26682 68660 26767
rect 68619 26564 68661 26573
rect 68619 26524 68620 26564
rect 68660 26524 68661 26564
rect 68619 26515 68661 26524
rect 68620 26237 68660 26515
rect 68619 26228 68661 26237
rect 68619 26188 68620 26228
rect 68660 26188 68661 26228
rect 68619 26179 68661 26188
rect 68619 25976 68661 25985
rect 68524 25936 68620 25976
rect 68660 25936 68661 25976
rect 68619 25927 68661 25936
rect 68620 25842 68660 25927
rect 68523 25304 68565 25313
rect 68523 25264 68524 25304
rect 68564 25264 68565 25304
rect 68523 25255 68565 25264
rect 68524 24464 68564 25255
rect 68524 24415 68564 24424
rect 68523 23960 68565 23969
rect 68523 23920 68524 23960
rect 68564 23920 68565 23960
rect 68523 23911 68565 23920
rect 68180 23752 68468 23792
rect 68140 23743 68180 23752
rect 67659 23708 67701 23717
rect 67659 23668 67660 23708
rect 67700 23668 67701 23708
rect 67659 23659 67701 23668
rect 68043 23708 68085 23717
rect 68043 23668 68044 23708
rect 68084 23668 68085 23708
rect 68043 23659 68085 23668
rect 67660 23628 67700 23659
rect 67756 23624 67796 23633
rect 67756 23060 67796 23584
rect 68044 23060 68084 23659
rect 68236 23624 68276 23633
rect 68236 23060 68276 23584
rect 68428 23060 68468 23752
rect 68524 23792 68564 23911
rect 68716 23801 68756 26944
rect 68812 26489 68852 32395
rect 69003 32192 69045 32201
rect 69003 32152 69004 32192
rect 69044 32152 69045 32192
rect 69003 32143 69045 32152
rect 69004 29168 69044 32143
rect 69100 31940 69140 31949
rect 69100 31361 69140 31900
rect 69099 31352 69141 31361
rect 69099 31312 69100 31352
rect 69140 31312 69141 31352
rect 69099 31303 69141 31312
rect 69100 31193 69140 31303
rect 69099 31184 69141 31193
rect 69099 31144 69100 31184
rect 69140 31144 69141 31184
rect 69099 31135 69141 31144
rect 69004 29119 69044 29128
rect 69100 29924 69140 29933
rect 68907 29000 68949 29009
rect 68907 28960 68908 29000
rect 68948 28960 68949 29000
rect 68907 28951 68949 28960
rect 68811 26480 68853 26489
rect 68811 26440 68812 26480
rect 68852 26440 68853 26480
rect 68811 26431 68853 26440
rect 68811 26228 68853 26237
rect 68811 26188 68812 26228
rect 68852 26188 68853 26228
rect 68811 26179 68853 26188
rect 68812 26060 68852 26179
rect 68812 26011 68852 26020
rect 68908 23969 68948 28951
rect 69100 28580 69140 29884
rect 69004 28540 69140 28580
rect 69004 27833 69044 28540
rect 69196 28496 69236 32740
rect 69291 32108 69333 32117
rect 69291 32068 69292 32108
rect 69332 32068 69333 32108
rect 69291 32059 69333 32068
rect 69292 30092 69332 32059
rect 69388 32033 69428 32740
rect 69483 32192 69525 32201
rect 69483 32152 69484 32192
rect 69524 32152 69525 32192
rect 69483 32143 69525 32152
rect 69387 32024 69429 32033
rect 69387 31984 69388 32024
rect 69428 31984 69429 32024
rect 69387 31975 69429 31984
rect 69484 30680 69524 32143
rect 69484 30631 69524 30640
rect 69292 29849 69332 30052
rect 69580 30008 69620 34747
rect 69964 34376 70004 35335
rect 69964 34327 70004 34336
rect 69963 33704 70005 33713
rect 69963 33664 69964 33704
rect 70004 33664 70005 33704
rect 69963 33655 70005 33664
rect 69868 33536 69908 33545
rect 69868 33140 69908 33496
rect 69772 33100 69908 33140
rect 69772 32864 69812 33100
rect 69772 32815 69812 32824
rect 69771 32696 69813 32705
rect 69964 32696 70004 33655
rect 69771 32656 69772 32696
rect 69812 32656 69813 32696
rect 69771 32647 69813 32656
rect 69868 32656 70004 32696
rect 69772 32192 69812 32647
rect 69772 32143 69812 32152
rect 69868 32192 69908 32656
rect 70060 32360 70100 37948
rect 71115 37988 71157 37997
rect 71115 37948 71116 37988
rect 71156 37948 71157 37988
rect 71115 37939 71157 37948
rect 71116 37854 71156 37939
rect 70443 37400 70485 37409
rect 70443 37360 70444 37400
rect 70484 37360 70485 37400
rect 70443 37351 70485 37360
rect 70444 36737 70484 37351
rect 71404 37241 71444 38032
rect 71403 37232 71445 37241
rect 71403 37192 71404 37232
rect 71444 37192 71445 37232
rect 71403 37183 71445 37192
rect 71596 37232 71636 37241
rect 70731 36896 70773 36905
rect 70731 36856 70732 36896
rect 70772 36856 70773 36896
rect 70731 36847 70773 36856
rect 70443 36728 70485 36737
rect 70443 36688 70444 36728
rect 70484 36688 70485 36728
rect 70443 36679 70485 36688
rect 70251 35972 70293 35981
rect 70251 35932 70252 35972
rect 70292 35932 70293 35972
rect 70251 35923 70293 35932
rect 70252 35141 70292 35923
rect 70347 35888 70389 35897
rect 70347 35848 70348 35888
rect 70388 35848 70389 35888
rect 70347 35839 70389 35848
rect 70348 35309 70388 35839
rect 70444 35393 70484 36679
rect 70443 35384 70485 35393
rect 70443 35344 70444 35384
rect 70484 35344 70485 35384
rect 70443 35335 70485 35344
rect 70347 35300 70389 35309
rect 70347 35260 70348 35300
rect 70388 35260 70389 35300
rect 70347 35251 70389 35260
rect 70348 35216 70388 35251
rect 70251 35132 70293 35141
rect 70251 35092 70252 35132
rect 70292 35092 70293 35132
rect 70251 35083 70293 35092
rect 70252 33140 70292 35083
rect 70348 34637 70388 35176
rect 70443 35216 70485 35225
rect 70443 35176 70444 35216
rect 70484 35176 70485 35216
rect 70443 35167 70485 35176
rect 70540 35216 70580 35227
rect 70347 34628 70389 34637
rect 70347 34588 70348 34628
rect 70388 34588 70389 34628
rect 70347 34579 70389 34588
rect 70252 33100 70388 33140
rect 69868 32143 69908 32152
rect 69964 32320 70100 32360
rect 69964 32024 70004 32320
rect 70060 32192 70100 32201
rect 70252 32192 70292 32201
rect 70100 32152 70252 32192
rect 70060 32143 70100 32152
rect 70252 32143 70292 32152
rect 70348 32192 70388 33100
rect 69868 31984 70004 32024
rect 70059 32024 70101 32033
rect 70059 31984 70060 32024
rect 70100 31984 70101 32024
rect 69675 30092 69717 30101
rect 69675 30052 69676 30092
rect 69716 30052 69717 30092
rect 69675 30043 69717 30052
rect 69388 29968 69620 30008
rect 69291 29840 69333 29849
rect 69291 29800 69292 29840
rect 69332 29800 69333 29840
rect 69291 29791 69333 29800
rect 69100 28456 69236 28496
rect 69003 27824 69045 27833
rect 69003 27784 69004 27824
rect 69044 27784 69045 27824
rect 69003 27775 69045 27784
rect 69100 27581 69140 28456
rect 69195 28328 69237 28337
rect 69195 28288 69196 28328
rect 69236 28288 69237 28328
rect 69195 28279 69237 28288
rect 69099 27572 69141 27581
rect 69099 27532 69100 27572
rect 69140 27532 69141 27572
rect 69099 27523 69141 27532
rect 69099 27404 69141 27413
rect 69099 27364 69100 27404
rect 69140 27364 69141 27404
rect 69099 27355 69141 27364
rect 69100 26816 69140 27355
rect 69100 26767 69140 26776
rect 69003 26480 69045 26489
rect 69003 26440 69004 26480
rect 69044 26440 69045 26480
rect 69003 26431 69045 26440
rect 68907 23960 68949 23969
rect 68812 23920 68908 23960
rect 68948 23920 68949 23960
rect 68524 23743 68564 23752
rect 68715 23792 68757 23801
rect 68715 23752 68716 23792
rect 68756 23752 68757 23792
rect 68715 23743 68757 23752
rect 68620 23624 68660 23633
rect 68620 23060 68660 23584
rect 68812 23060 68852 23920
rect 68907 23911 68949 23920
rect 68908 23792 68948 23801
rect 69004 23792 69044 26431
rect 69099 26312 69141 26321
rect 69099 26272 69100 26312
rect 69140 26272 69141 26312
rect 69099 26263 69141 26272
rect 69100 25136 69140 26263
rect 69196 25901 69236 28279
rect 69388 27656 69428 29968
rect 69483 29840 69525 29849
rect 69483 29800 69484 29840
rect 69524 29800 69525 29840
rect 69483 29791 69525 29800
rect 69676 29840 69716 30043
rect 69676 29791 69716 29800
rect 69771 29840 69813 29849
rect 69771 29800 69772 29840
rect 69812 29800 69813 29840
rect 69771 29791 69813 29800
rect 69484 29706 69524 29791
rect 69579 29756 69621 29765
rect 69579 29716 69580 29756
rect 69620 29716 69621 29756
rect 69579 29707 69621 29716
rect 69580 29622 69620 29707
rect 69772 29706 69812 29791
rect 69771 29168 69813 29177
rect 69771 29128 69772 29168
rect 69812 29128 69813 29168
rect 69771 29119 69813 29128
rect 69772 28160 69812 29119
rect 69868 28337 69908 31984
rect 70059 31975 70101 31984
rect 70060 31890 70100 31975
rect 70251 31940 70293 31949
rect 70251 31900 70252 31940
rect 70292 31900 70293 31940
rect 70251 31891 70293 31900
rect 70252 30008 70292 31891
rect 70348 30428 70388 32152
rect 70444 32192 70484 35167
rect 70540 35141 70580 35176
rect 70635 35216 70677 35225
rect 70635 35176 70636 35216
rect 70676 35176 70677 35216
rect 70635 35167 70677 35176
rect 70539 35132 70581 35141
rect 70539 35092 70540 35132
rect 70580 35092 70581 35132
rect 70539 35083 70581 35092
rect 70636 35082 70676 35167
rect 70635 34880 70677 34889
rect 70635 34840 70636 34880
rect 70676 34840 70677 34880
rect 70635 34831 70677 34840
rect 70636 33965 70676 34831
rect 70732 34469 70772 36847
rect 71596 36821 71636 37192
rect 71595 36812 71637 36821
rect 71595 36772 71596 36812
rect 71636 36772 71637 36812
rect 71595 36763 71637 36772
rect 71596 36569 71636 36763
rect 71595 36560 71637 36569
rect 71595 36520 71596 36560
rect 71636 36520 71637 36560
rect 71595 36511 71637 36520
rect 70923 36476 70965 36485
rect 70923 36436 70924 36476
rect 70964 36436 70965 36476
rect 70923 36427 70965 36436
rect 70924 36342 70964 36427
rect 70827 36056 70869 36065
rect 70827 36016 70828 36056
rect 70868 36016 70869 36056
rect 70827 36007 70869 36016
rect 70731 34460 70773 34469
rect 70731 34420 70732 34460
rect 70772 34420 70773 34460
rect 70731 34411 70773 34420
rect 70828 34376 70868 36007
rect 71500 35888 71540 35897
rect 71403 35804 71445 35813
rect 71403 35764 71404 35804
rect 71444 35764 71445 35804
rect 71403 35755 71445 35764
rect 70923 35468 70965 35477
rect 70923 35428 70924 35468
rect 70964 35428 70965 35468
rect 70923 35419 70965 35428
rect 70828 34327 70868 34336
rect 70924 35216 70964 35419
rect 71307 35300 71349 35309
rect 71307 35260 71308 35300
rect 71348 35260 71349 35300
rect 71307 35251 71349 35260
rect 71212 35216 71252 35225
rect 70924 34208 70964 35176
rect 70732 34168 70964 34208
rect 71116 35176 71212 35216
rect 70635 33956 70677 33965
rect 70635 33916 70636 33956
rect 70676 33916 70677 33956
rect 70635 33907 70677 33916
rect 70636 32864 70676 32873
rect 70539 32276 70581 32285
rect 70539 32236 70540 32276
rect 70580 32236 70581 32276
rect 70539 32227 70581 32236
rect 70444 30680 70484 32152
rect 70540 32192 70580 32227
rect 70636 32201 70676 32824
rect 70732 32369 70772 34168
rect 71019 33956 71061 33965
rect 71019 33916 71020 33956
rect 71060 33916 71061 33956
rect 71019 33907 71061 33916
rect 71020 33140 71060 33907
rect 71116 33545 71156 35176
rect 71212 35167 71252 35176
rect 71308 35166 71348 35251
rect 71211 34544 71253 34553
rect 71211 34504 71212 34544
rect 71252 34504 71253 34544
rect 71211 34495 71253 34504
rect 71212 34376 71252 34495
rect 71307 34460 71349 34469
rect 71307 34420 71308 34460
rect 71348 34420 71349 34460
rect 71307 34411 71349 34420
rect 71212 34327 71252 34336
rect 71115 33536 71157 33545
rect 71115 33496 71116 33536
rect 71156 33496 71157 33536
rect 71115 33487 71157 33496
rect 71308 33140 71348 34411
rect 71404 33704 71444 35755
rect 71500 35048 71540 35848
rect 71692 35888 71732 38200
rect 74283 38200 74284 38240
rect 74324 38200 74325 38240
rect 74283 38191 74325 38200
rect 75244 38240 75284 38249
rect 76972 38240 77012 38249
rect 75284 38200 75380 38240
rect 75244 38191 75284 38200
rect 74284 38106 74324 38191
rect 71980 38072 72020 38081
rect 72020 38032 72404 38072
rect 71980 38023 72020 38032
rect 72075 36728 72117 36737
rect 72075 36688 72076 36728
rect 72116 36688 72117 36728
rect 72364 36728 72404 38032
rect 73323 37568 73365 37577
rect 74284 37568 74324 37577
rect 73323 37528 73324 37568
rect 73364 37528 73365 37568
rect 73323 37519 73365 37528
rect 74188 37528 74284 37568
rect 73131 37484 73173 37493
rect 73131 37444 73132 37484
rect 73172 37444 73173 37484
rect 73131 37435 73173 37444
rect 72844 37400 72884 37409
rect 72844 36896 72884 37360
rect 72940 37400 72980 37409
rect 72940 37157 72980 37360
rect 73036 37400 73076 37409
rect 72939 37148 72981 37157
rect 72939 37108 72940 37148
rect 72980 37108 72981 37148
rect 72939 37099 72981 37108
rect 73036 37073 73076 37360
rect 73132 37400 73172 37435
rect 73132 37349 73172 37360
rect 73227 37400 73269 37409
rect 73227 37360 73228 37400
rect 73268 37360 73269 37400
rect 73227 37351 73269 37360
rect 73324 37400 73364 37519
rect 73707 37484 73749 37493
rect 73707 37444 73708 37484
rect 73748 37444 73844 37484
rect 73707 37435 73749 37444
rect 73324 37351 73364 37360
rect 73515 37400 73557 37409
rect 73515 37360 73516 37400
rect 73556 37360 73557 37400
rect 73515 37351 73557 37360
rect 73612 37400 73652 37409
rect 73035 37064 73077 37073
rect 73035 37024 73036 37064
rect 73076 37024 73077 37064
rect 73035 37015 73077 37024
rect 72844 36856 73076 36896
rect 72940 36728 72980 36737
rect 72364 36688 72940 36728
rect 72075 36679 72117 36688
rect 72940 36679 72980 36688
rect 72076 36594 72116 36679
rect 72939 36560 72981 36569
rect 72939 36520 72940 36560
rect 72980 36520 72981 36560
rect 72939 36511 72981 36520
rect 72171 36476 72213 36485
rect 72171 36436 72172 36476
rect 72212 36436 72213 36476
rect 72171 36427 72213 36436
rect 72172 36065 72212 36427
rect 72171 36056 72213 36065
rect 72171 36016 72172 36056
rect 72212 36016 72213 36056
rect 72171 36007 72213 36016
rect 72076 35897 72116 35982
rect 71596 35804 71636 35813
rect 71596 35384 71636 35764
rect 71692 35561 71732 35848
rect 71883 35888 71925 35897
rect 71883 35848 71884 35888
rect 71924 35848 71925 35888
rect 71883 35839 71925 35848
rect 72075 35888 72117 35897
rect 72075 35848 72076 35888
rect 72116 35848 72117 35888
rect 72075 35839 72117 35848
rect 72172 35888 72212 36007
rect 72172 35839 72212 35848
rect 72844 35888 72884 35897
rect 71884 35754 71924 35839
rect 71980 35720 72020 35729
rect 72020 35680 72116 35720
rect 71980 35671 72020 35680
rect 71691 35552 71733 35561
rect 71691 35512 71692 35552
rect 71732 35512 71733 35552
rect 71691 35503 71733 35512
rect 71596 35344 72020 35384
rect 71787 35216 71829 35225
rect 71787 35176 71788 35216
rect 71828 35176 71829 35216
rect 71787 35167 71829 35176
rect 71788 35082 71828 35167
rect 71596 35048 71636 35057
rect 71500 35008 71596 35048
rect 71596 34999 71636 35008
rect 71788 34964 71828 34973
rect 71692 34924 71788 34964
rect 71499 34796 71541 34805
rect 71499 34756 71500 34796
rect 71540 34756 71541 34796
rect 71499 34747 71541 34756
rect 71500 34049 71540 34747
rect 71692 34553 71732 34924
rect 71788 34915 71828 34924
rect 71884 34712 71924 35344
rect 71980 35216 72020 35344
rect 71980 35167 72020 35176
rect 72076 35216 72116 35680
rect 72651 35552 72693 35561
rect 72651 35512 72652 35552
rect 72692 35512 72693 35552
rect 72651 35503 72693 35512
rect 72076 35167 72116 35176
rect 71788 34672 71924 34712
rect 72556 35048 72596 35057
rect 71691 34544 71733 34553
rect 71691 34504 71692 34544
rect 71732 34504 71733 34544
rect 71691 34495 71733 34504
rect 71596 34376 71636 34385
rect 71499 34040 71541 34049
rect 71499 34000 71500 34040
rect 71540 34000 71541 34040
rect 71499 33991 71541 34000
rect 71596 33872 71636 34336
rect 71692 34376 71732 34385
rect 71788 34376 71828 34672
rect 71884 34544 71924 34553
rect 71924 34504 72116 34544
rect 71884 34495 71924 34504
rect 71732 34336 71828 34376
rect 71884 34376 71924 34385
rect 71692 34327 71732 34336
rect 71884 34292 71924 34336
rect 71979 34376 72021 34385
rect 71979 34336 71980 34376
rect 72020 34336 72021 34376
rect 71979 34327 72021 34336
rect 72076 34376 72116 34504
rect 72076 34327 72116 34336
rect 72460 34376 72500 34385
rect 72556 34376 72596 35008
rect 72500 34336 72596 34376
rect 72460 34327 72500 34336
rect 71788 34252 71924 34292
rect 71788 34049 71828 34252
rect 71980 34208 72020 34327
rect 71884 34168 72020 34208
rect 71787 34040 71829 34049
rect 71787 34000 71788 34040
rect 71828 34000 71829 34040
rect 71787 33991 71829 34000
rect 71596 33832 71732 33872
rect 71692 33788 71732 33832
rect 71692 33739 71732 33748
rect 71596 33704 71636 33713
rect 71404 33664 71596 33704
rect 71020 33100 71252 33140
rect 71308 33100 71444 33140
rect 70923 32864 70965 32873
rect 70923 32824 70924 32864
rect 70964 32824 70965 32864
rect 70923 32815 70965 32824
rect 70731 32360 70773 32369
rect 70731 32320 70732 32360
rect 70772 32320 70773 32360
rect 70731 32311 70773 32320
rect 70540 32141 70580 32152
rect 70635 32192 70677 32201
rect 70635 32152 70636 32192
rect 70676 32152 70677 32192
rect 70635 32143 70677 32152
rect 70732 32192 70772 32203
rect 70732 32117 70772 32152
rect 70924 32192 70964 32815
rect 71115 32612 71157 32621
rect 71020 32572 71116 32612
rect 71156 32572 71157 32612
rect 71020 32285 71060 32572
rect 71115 32563 71157 32572
rect 71019 32276 71061 32285
rect 71019 32236 71020 32276
rect 71060 32236 71061 32276
rect 71019 32227 71061 32236
rect 70924 32143 70964 32152
rect 71020 32192 71060 32227
rect 71020 32142 71060 32152
rect 70731 32108 70773 32117
rect 70731 32068 70732 32108
rect 70772 32068 70773 32108
rect 71212 32108 71252 33100
rect 71212 32068 71348 32108
rect 70731 32059 70773 32068
rect 70732 31940 70772 31949
rect 71211 31940 71253 31949
rect 70772 31900 70868 31940
rect 70732 31891 70772 31900
rect 70731 31520 70773 31529
rect 70731 31480 70732 31520
rect 70772 31480 70773 31520
rect 70731 31471 70773 31480
rect 70540 31352 70580 31361
rect 70540 30857 70580 31312
rect 70732 31352 70772 31471
rect 70732 31303 70772 31312
rect 70828 31352 70868 31900
rect 71211 31900 71212 31940
rect 71252 31900 71253 31940
rect 71211 31891 71253 31900
rect 71115 31520 71157 31529
rect 71115 31480 71116 31520
rect 71156 31480 71157 31520
rect 71115 31471 71157 31480
rect 71116 31386 71156 31471
rect 70828 31303 70868 31312
rect 71020 31352 71060 31361
rect 70636 31184 70676 31193
rect 70539 30848 70581 30857
rect 70539 30808 70540 30848
rect 70580 30808 70581 30848
rect 70539 30799 70581 30808
rect 70636 30773 70676 31144
rect 71020 31109 71060 31312
rect 71212 31352 71252 31891
rect 70731 31100 70773 31109
rect 70731 31060 70732 31100
rect 70772 31060 70773 31100
rect 70731 31051 70773 31060
rect 71019 31100 71061 31109
rect 71019 31060 71020 31100
rect 71060 31060 71061 31100
rect 71019 31051 71061 31060
rect 70635 30764 70677 30773
rect 70635 30724 70636 30764
rect 70676 30724 70677 30764
rect 70635 30715 70677 30724
rect 70539 30680 70581 30689
rect 70444 30640 70540 30680
rect 70580 30640 70581 30680
rect 70539 30631 70581 30640
rect 70443 30428 70485 30437
rect 70348 30388 70444 30428
rect 70484 30388 70485 30428
rect 70443 30379 70485 30388
rect 70252 29968 70388 30008
rect 69964 29840 70004 29851
rect 69964 29765 70004 29800
rect 70060 29840 70100 29849
rect 69963 29756 70005 29765
rect 69963 29716 69964 29756
rect 70004 29716 70005 29756
rect 69963 29707 70005 29716
rect 69963 29504 70005 29513
rect 69963 29464 69964 29504
rect 70004 29464 70005 29504
rect 69963 29455 70005 29464
rect 69964 28580 70004 29455
rect 70060 28841 70100 29800
rect 70252 29840 70292 29849
rect 70156 29672 70196 29681
rect 70156 29261 70196 29632
rect 70252 29336 70292 29800
rect 70348 29513 70388 29968
rect 70347 29504 70389 29513
rect 70347 29464 70348 29504
rect 70388 29464 70389 29504
rect 70347 29455 70389 29464
rect 70348 29336 70388 29345
rect 70252 29296 70348 29336
rect 70348 29287 70388 29296
rect 70155 29252 70197 29261
rect 70155 29212 70156 29252
rect 70196 29212 70197 29252
rect 70155 29203 70197 29212
rect 70444 29168 70484 30379
rect 70540 29177 70580 30631
rect 70636 30428 70676 30437
rect 70636 29849 70676 30388
rect 70732 30092 70772 31051
rect 70827 30848 70869 30857
rect 70827 30808 70828 30848
rect 70868 30808 70869 30848
rect 70827 30799 70869 30808
rect 70828 30714 70868 30799
rect 71020 30689 71060 30774
rect 70924 30680 70964 30689
rect 70924 30437 70964 30640
rect 71019 30680 71061 30689
rect 71019 30640 71020 30680
rect 71060 30640 71061 30680
rect 71019 30631 71061 30640
rect 71116 30680 71156 30689
rect 71019 30512 71061 30521
rect 71019 30472 71020 30512
rect 71060 30472 71061 30512
rect 71019 30463 71061 30472
rect 70923 30428 70965 30437
rect 70923 30388 70924 30428
rect 70964 30388 70965 30428
rect 70923 30379 70965 30388
rect 71020 30260 71060 30463
rect 70732 30043 70772 30052
rect 70924 30220 71060 30260
rect 70635 29840 70677 29849
rect 70635 29800 70636 29840
rect 70676 29800 70677 29840
rect 70635 29791 70677 29800
rect 70827 29504 70869 29513
rect 70827 29464 70828 29504
rect 70868 29464 70869 29504
rect 70827 29455 70869 29464
rect 70828 29336 70868 29455
rect 70828 29287 70868 29296
rect 70444 29119 70484 29128
rect 70539 29168 70581 29177
rect 70539 29128 70540 29168
rect 70580 29128 70581 29168
rect 70539 29119 70581 29128
rect 70636 29168 70676 29179
rect 70155 29084 70197 29093
rect 70155 29044 70156 29084
rect 70196 29044 70197 29084
rect 70155 29035 70197 29044
rect 70156 28950 70196 29035
rect 70540 29034 70580 29119
rect 70636 29093 70676 29128
rect 70635 29084 70677 29093
rect 70924 29084 70964 30220
rect 71116 30176 71156 30640
rect 71020 30136 71156 30176
rect 71020 29849 71060 30136
rect 71115 30008 71157 30017
rect 71115 29968 71116 30008
rect 71156 29968 71157 30008
rect 71115 29959 71157 29968
rect 71019 29840 71061 29849
rect 71019 29800 71020 29840
rect 71060 29800 71061 29840
rect 71019 29791 71061 29800
rect 71116 29840 71156 29959
rect 71116 29791 71156 29800
rect 71020 29706 71060 29791
rect 71212 29336 71252 31312
rect 71308 30857 71348 32068
rect 71404 31781 71444 33100
rect 71500 32873 71540 33664
rect 71596 33655 71636 33664
rect 71788 33704 71828 33713
rect 71788 33545 71828 33664
rect 71787 33536 71829 33545
rect 71787 33496 71788 33536
rect 71828 33496 71829 33536
rect 71787 33487 71829 33496
rect 71499 32864 71541 32873
rect 71499 32824 71500 32864
rect 71540 32824 71541 32864
rect 71499 32815 71541 32824
rect 71787 32696 71829 32705
rect 71787 32656 71788 32696
rect 71828 32656 71829 32696
rect 71787 32647 71829 32656
rect 71788 32562 71828 32647
rect 71499 32360 71541 32369
rect 71499 32320 71500 32360
rect 71540 32320 71541 32360
rect 71499 32311 71541 32320
rect 71691 32360 71733 32369
rect 71691 32320 71692 32360
rect 71732 32320 71733 32360
rect 71691 32311 71733 32320
rect 71403 31772 71445 31781
rect 71403 31732 71404 31772
rect 71444 31732 71445 31772
rect 71403 31723 71445 31732
rect 71403 31604 71445 31613
rect 71403 31564 71404 31604
rect 71444 31564 71445 31604
rect 71403 31555 71445 31564
rect 71404 31470 71444 31555
rect 71403 31352 71445 31361
rect 71403 31312 71404 31352
rect 71444 31312 71445 31352
rect 71403 31303 71445 31312
rect 71404 31218 71444 31303
rect 71500 31016 71540 32311
rect 71692 32192 71732 32311
rect 71692 32143 71732 32152
rect 71691 31772 71733 31781
rect 71691 31732 71692 31772
rect 71732 31732 71733 31772
rect 71691 31723 71733 31732
rect 71595 31520 71637 31529
rect 71595 31480 71596 31520
rect 71636 31480 71637 31520
rect 71595 31471 71637 31480
rect 71596 31352 71636 31471
rect 71692 31436 71732 31723
rect 71884 31697 71924 34168
rect 71979 34040 72021 34049
rect 71979 34000 71980 34040
rect 72020 34000 72021 34040
rect 71979 33991 72021 34000
rect 71980 33704 72020 33991
rect 71980 33629 72020 33664
rect 72171 33704 72213 33713
rect 72171 33664 72172 33704
rect 72212 33664 72213 33704
rect 72171 33655 72213 33664
rect 72268 33704 72308 33713
rect 71979 33620 72021 33629
rect 71979 33580 71980 33620
rect 72020 33580 72021 33620
rect 71979 33571 72021 33580
rect 72172 33570 72212 33655
rect 71980 33452 72020 33461
rect 71980 33140 72020 33412
rect 71980 33100 72212 33140
rect 72172 32864 72212 33100
rect 72172 32815 72212 32824
rect 71979 32696 72021 32705
rect 71979 32656 71980 32696
rect 72020 32656 72021 32696
rect 71979 32647 72021 32656
rect 71980 32444 72020 32647
rect 71980 32404 72116 32444
rect 71979 32276 72021 32285
rect 71979 32236 71980 32276
rect 72020 32236 72021 32276
rect 71979 32227 72021 32236
rect 72076 32276 72116 32404
rect 72076 32227 72116 32236
rect 71980 32192 72020 32227
rect 71980 32141 72020 32152
rect 71979 32024 72021 32033
rect 71979 31984 71980 32024
rect 72020 31984 72021 32024
rect 71979 31975 72021 31984
rect 71883 31688 71925 31697
rect 71883 31648 71884 31688
rect 71924 31648 71925 31688
rect 71883 31639 71925 31648
rect 71884 31436 71924 31445
rect 71692 31396 71884 31436
rect 71884 31387 71924 31396
rect 71596 31303 71636 31312
rect 71692 31337 71732 31346
rect 71692 31268 71732 31297
rect 71692 31228 71828 31268
rect 71691 31100 71733 31109
rect 71691 31060 71692 31100
rect 71732 31060 71733 31100
rect 71691 31051 71733 31060
rect 71404 30976 71540 31016
rect 71595 31016 71637 31025
rect 71595 30976 71596 31016
rect 71636 30976 71637 31016
rect 71307 30848 71349 30857
rect 71307 30808 71308 30848
rect 71348 30808 71349 30848
rect 71307 30799 71349 30808
rect 71307 30596 71349 30605
rect 71307 30556 71308 30596
rect 71348 30556 71349 30596
rect 71307 30547 71349 30556
rect 71308 30462 71348 30547
rect 71404 29840 71444 30976
rect 71595 30967 71637 30976
rect 71499 30848 71541 30857
rect 71499 30808 71500 30848
rect 71540 30808 71541 30848
rect 71499 30799 71541 30808
rect 71500 30714 71540 30799
rect 71500 30428 71540 30437
rect 71500 29933 71540 30388
rect 71499 29924 71541 29933
rect 71499 29884 71500 29924
rect 71540 29884 71541 29924
rect 71499 29875 71541 29884
rect 71404 29513 71444 29800
rect 71403 29504 71445 29513
rect 71403 29464 71404 29504
rect 71444 29464 71445 29504
rect 71596 29504 71636 30967
rect 71692 30764 71732 31051
rect 71692 30715 71732 30724
rect 71788 30269 71828 31228
rect 71787 30260 71829 30269
rect 71787 30220 71788 30260
rect 71828 30220 71829 30260
rect 71787 30211 71829 30220
rect 71691 30092 71733 30101
rect 71980 30092 72020 31975
rect 72268 31856 72308 33664
rect 72460 33704 72500 33713
rect 72460 33140 72500 33664
rect 72555 33704 72597 33713
rect 72555 33664 72556 33704
rect 72596 33664 72597 33704
rect 72555 33655 72597 33664
rect 72652 33704 72692 35503
rect 72844 34385 72884 35848
rect 72843 34376 72885 34385
rect 72843 34336 72844 34376
rect 72884 34336 72885 34376
rect 72843 34327 72885 34336
rect 72556 33570 72596 33655
rect 72364 33100 72500 33140
rect 72364 32024 72404 33100
rect 72652 33041 72692 33664
rect 72844 33536 72884 33545
rect 72651 33032 72693 33041
rect 72651 32992 72652 33032
rect 72692 32992 72693 33032
rect 72651 32983 72693 32992
rect 72459 32864 72501 32873
rect 72459 32824 72460 32864
rect 72500 32824 72501 32864
rect 72459 32815 72501 32824
rect 72556 32864 72596 32873
rect 72844 32864 72884 33496
rect 72940 33140 72980 36511
rect 73036 36065 73076 36856
rect 73228 36644 73268 37351
rect 73516 37266 73556 37351
rect 73323 37232 73365 37241
rect 73323 37192 73324 37232
rect 73364 37192 73365 37232
rect 73323 37183 73365 37192
rect 73420 37232 73460 37241
rect 73324 36812 73364 37183
rect 73420 36896 73460 37192
rect 73420 36856 73556 36896
rect 73324 36763 73364 36772
rect 73516 36812 73556 36856
rect 73516 36763 73556 36772
rect 73228 36604 73556 36644
rect 73516 36224 73556 36604
rect 73324 36184 73556 36224
rect 73035 36056 73077 36065
rect 73035 36016 73036 36056
rect 73076 36016 73077 36056
rect 73035 36007 73077 36016
rect 73227 36056 73269 36065
rect 73227 36016 73228 36056
rect 73268 36016 73269 36056
rect 73227 36007 73269 36016
rect 73131 35888 73173 35897
rect 73131 35848 73132 35888
rect 73172 35848 73173 35888
rect 73131 35839 73173 35848
rect 73228 35888 73268 36007
rect 73228 35839 73268 35848
rect 73132 35754 73172 35839
rect 73227 35552 73269 35561
rect 73227 35512 73228 35552
rect 73268 35512 73269 35552
rect 73324 35552 73364 36184
rect 73612 36140 73652 37360
rect 73804 37400 73844 37444
rect 73804 37351 73844 37360
rect 73995 37400 74037 37409
rect 73995 37360 73996 37400
rect 74036 37360 74037 37400
rect 73995 37351 74037 37360
rect 74092 37400 74132 37409
rect 74188 37400 74228 37528
rect 74284 37519 74324 37528
rect 74132 37360 74228 37400
rect 74284 37400 74324 37409
rect 74092 37351 74132 37360
rect 73996 37266 74036 37351
rect 73899 37232 73941 37241
rect 73899 37192 73900 37232
rect 73940 37192 73941 37232
rect 73899 37183 73941 37192
rect 73900 37098 73940 37183
rect 73900 36728 73940 36737
rect 73940 36688 74132 36728
rect 73900 36679 73940 36688
rect 73804 36140 73844 36149
rect 73612 36100 73804 36140
rect 73804 36091 73844 36100
rect 73516 36056 73556 36065
rect 73324 35512 73460 35552
rect 73227 35503 73269 35512
rect 73228 35300 73268 35503
rect 73420 35300 73460 35512
rect 73228 35260 73364 35300
rect 72940 33100 73172 33140
rect 73035 33032 73077 33041
rect 73035 32992 73036 33032
rect 73076 32992 73077 33032
rect 73035 32983 73077 32992
rect 72596 32824 72884 32864
rect 72556 32815 72596 32824
rect 72460 32192 72500 32815
rect 72747 32276 72789 32285
rect 72747 32236 72748 32276
rect 72788 32236 72789 32276
rect 72747 32227 72789 32236
rect 72556 32192 72596 32201
rect 72460 32152 72556 32192
rect 72460 32033 72500 32152
rect 72556 32143 72596 32152
rect 72748 32192 72788 32227
rect 72748 32141 72788 32152
rect 72939 32192 72981 32201
rect 72939 32152 72940 32192
rect 72980 32152 72981 32192
rect 72939 32143 72981 32152
rect 72364 31975 72404 31984
rect 72459 32024 72501 32033
rect 72459 31984 72460 32024
rect 72500 31984 72501 32024
rect 72459 31975 72501 31984
rect 72652 31940 72692 31949
rect 72652 31856 72692 31900
rect 72268 31816 72692 31856
rect 72075 31604 72117 31613
rect 72075 31564 72076 31604
rect 72116 31564 72117 31604
rect 72075 31555 72117 31564
rect 72076 31470 72116 31555
rect 72268 31520 72308 31529
rect 72076 30680 72116 30689
rect 72268 30680 72308 31480
rect 72116 30640 72308 30680
rect 72940 30680 72980 32143
rect 73036 31949 73076 32983
rect 73035 31940 73077 31949
rect 73035 31900 73036 31940
rect 73076 31900 73077 31940
rect 73035 31891 73077 31900
rect 72076 30631 72116 30640
rect 72940 30631 72980 30640
rect 72171 30260 72213 30269
rect 72171 30220 72172 30260
rect 72212 30220 72213 30260
rect 72171 30211 72213 30220
rect 72172 30092 72212 30211
rect 71691 30052 71692 30092
rect 71732 30052 72116 30092
rect 71691 30043 71733 30052
rect 71692 29958 71732 30043
rect 71883 29924 71925 29933
rect 71883 29884 71884 29924
rect 71924 29884 71925 29924
rect 71883 29875 71925 29884
rect 71884 29790 71924 29875
rect 72076 29840 72116 30052
rect 72172 30043 72212 30052
rect 72267 30008 72309 30017
rect 72267 29968 72268 30008
rect 72308 29968 72309 30008
rect 72267 29959 72309 29968
rect 72076 29791 72116 29800
rect 72268 29840 72308 29959
rect 72268 29791 72308 29800
rect 71596 29464 71924 29504
rect 71403 29455 71445 29464
rect 71692 29336 71732 29345
rect 71212 29296 71692 29336
rect 71692 29287 71732 29296
rect 71308 29168 71348 29177
rect 71116 29128 71308 29168
rect 71019 29084 71061 29093
rect 70635 29044 70636 29084
rect 70676 29044 70772 29084
rect 70924 29044 71020 29084
rect 71060 29044 71061 29084
rect 70635 29035 70677 29044
rect 70347 28916 70389 28925
rect 70347 28876 70348 28916
rect 70388 28876 70389 28916
rect 70347 28867 70389 28876
rect 70059 28832 70101 28841
rect 70059 28792 70060 28832
rect 70100 28792 70101 28832
rect 70059 28783 70101 28792
rect 69964 28540 70196 28580
rect 70060 28412 70100 28421
rect 69867 28328 69909 28337
rect 69867 28288 69868 28328
rect 69908 28288 69909 28328
rect 69867 28279 69909 28288
rect 69868 28160 69908 28169
rect 69772 28120 69868 28160
rect 69868 28111 69908 28120
rect 70060 28001 70100 28372
rect 70059 27992 70101 28001
rect 70059 27952 70060 27992
rect 70100 27952 70101 27992
rect 70059 27943 70101 27952
rect 70059 27824 70101 27833
rect 70059 27784 70060 27824
rect 70100 27784 70101 27824
rect 70059 27775 70101 27784
rect 69772 27665 69812 27750
rect 69292 27616 69428 27656
rect 69580 27656 69620 27665
rect 69771 27656 69813 27665
rect 69620 27616 69716 27656
rect 69292 26984 69332 27616
rect 69580 27607 69620 27616
rect 69388 27488 69428 27497
rect 69428 27448 69524 27488
rect 69388 27439 69428 27448
rect 69292 26944 69428 26984
rect 69291 26816 69333 26825
rect 69291 26776 69292 26816
rect 69332 26776 69333 26816
rect 69291 26767 69333 26776
rect 69292 26237 69332 26767
rect 69388 26321 69428 26944
rect 69484 26816 69524 27448
rect 69579 27404 69621 27413
rect 69579 27364 69580 27404
rect 69620 27364 69621 27404
rect 69579 27355 69621 27364
rect 69580 27270 69620 27355
rect 69484 26767 69524 26776
rect 69483 26396 69525 26405
rect 69483 26356 69484 26396
rect 69524 26356 69525 26396
rect 69483 26347 69525 26356
rect 69387 26312 69429 26321
rect 69387 26272 69388 26312
rect 69428 26272 69429 26312
rect 69387 26263 69429 26272
rect 69291 26228 69333 26237
rect 69291 26188 69292 26228
rect 69332 26188 69333 26228
rect 69291 26179 69333 26188
rect 69292 26144 69332 26179
rect 69292 26094 69332 26104
rect 69387 26144 69429 26153
rect 69387 26104 69388 26144
rect 69428 26104 69429 26144
rect 69387 26095 69429 26104
rect 69484 26144 69524 26347
rect 69580 26312 69620 26321
rect 69676 26312 69716 27616
rect 69771 27616 69772 27656
rect 69812 27616 69813 27656
rect 69771 27607 69813 27616
rect 69868 27656 69908 27665
rect 69771 27488 69813 27497
rect 69771 27448 69772 27488
rect 69812 27448 69813 27488
rect 69868 27488 69908 27616
rect 70060 27656 70100 27775
rect 70060 27607 70100 27616
rect 70060 27488 70100 27497
rect 69868 27448 70060 27488
rect 69771 27439 69813 27448
rect 70060 27439 70100 27448
rect 69620 26272 69716 26312
rect 69580 26263 69620 26272
rect 69484 26095 69524 26104
rect 69388 26010 69428 26095
rect 69195 25892 69237 25901
rect 69195 25852 69196 25892
rect 69236 25852 69237 25892
rect 69195 25843 69237 25852
rect 69196 25304 69236 25843
rect 69196 25255 69236 25264
rect 69100 25096 69332 25136
rect 69292 23792 69332 25096
rect 69676 23792 69716 23801
rect 69772 23792 69812 27439
rect 70156 23969 70196 28540
rect 70251 28496 70293 28505
rect 70251 28456 70252 28496
rect 70292 28456 70293 28496
rect 70251 28447 70293 28456
rect 70252 27656 70292 28447
rect 70348 28328 70388 28867
rect 70635 28580 70677 28589
rect 70635 28540 70636 28580
rect 70676 28540 70677 28580
rect 70635 28531 70677 28540
rect 70348 28279 70388 28288
rect 70636 28328 70676 28531
rect 70636 28279 70676 28288
rect 70732 28328 70772 29044
rect 71019 29035 71061 29044
rect 71020 28950 71060 29035
rect 70827 28916 70869 28925
rect 70827 28876 70828 28916
rect 70868 28876 70869 28916
rect 70827 28867 70869 28876
rect 70828 28782 70868 28867
rect 71116 28505 71156 29128
rect 71308 29119 71348 29128
rect 71500 29168 71540 29177
rect 71404 28916 71444 28925
rect 71308 28876 71404 28916
rect 71211 28832 71253 28841
rect 71211 28792 71212 28832
rect 71252 28792 71253 28832
rect 71211 28783 71253 28792
rect 71020 28496 71060 28505
rect 70732 28160 70772 28288
rect 70252 27497 70292 27616
rect 70348 28120 70772 28160
rect 70828 28456 71020 28496
rect 70348 27656 70388 28120
rect 70539 27992 70581 28001
rect 70539 27952 70540 27992
rect 70580 27952 70581 27992
rect 70539 27943 70581 27952
rect 70731 27992 70773 28001
rect 70731 27952 70732 27992
rect 70772 27952 70773 27992
rect 70731 27943 70773 27952
rect 70348 27607 70388 27616
rect 70251 27488 70293 27497
rect 70251 27448 70252 27488
rect 70292 27448 70293 27488
rect 70251 27439 70293 27448
rect 70348 26816 70388 26825
rect 70348 25901 70388 26776
rect 70540 26153 70580 27943
rect 70635 27824 70677 27833
rect 70635 27784 70636 27824
rect 70676 27784 70677 27824
rect 70635 27775 70677 27784
rect 70636 27656 70676 27775
rect 70732 27740 70772 27943
rect 70732 27691 70772 27700
rect 70636 27607 70676 27616
rect 70828 27656 70868 28456
rect 71020 28447 71060 28456
rect 71115 28496 71157 28505
rect 71115 28456 71116 28496
rect 71156 28456 71157 28496
rect 71115 28447 71157 28456
rect 71019 28328 71061 28337
rect 71019 28288 71020 28328
rect 71060 28288 71061 28328
rect 71019 28279 71061 28288
rect 70828 27607 70868 27616
rect 71020 27656 71060 28279
rect 71212 28001 71252 28783
rect 71211 27992 71253 28001
rect 71211 27952 71212 27992
rect 71252 27952 71253 27992
rect 71211 27943 71253 27952
rect 70635 27488 70677 27497
rect 70635 27448 70636 27488
rect 70676 27448 70677 27488
rect 70635 27439 70677 27448
rect 70539 26144 70581 26153
rect 70539 26104 70540 26144
rect 70580 26104 70581 26144
rect 70539 26095 70581 26104
rect 70636 26069 70676 27439
rect 71020 27404 71060 27616
rect 71116 27740 71156 27749
rect 71116 27488 71156 27700
rect 71212 27656 71252 27943
rect 71212 27607 71252 27616
rect 71308 27656 71348 28876
rect 71404 28867 71444 28876
rect 71500 28589 71540 29128
rect 71595 29084 71637 29093
rect 71595 29044 71596 29084
rect 71636 29044 71637 29084
rect 71595 29035 71637 29044
rect 71884 29084 71924 29464
rect 71924 29044 72020 29084
rect 71884 29035 71924 29044
rect 71499 28580 71541 28589
rect 71499 28540 71500 28580
rect 71540 28540 71541 28580
rect 71499 28531 71541 28540
rect 71308 27607 71348 27616
rect 71404 28244 71444 28253
rect 71404 27488 71444 28204
rect 71499 28160 71541 28169
rect 71499 28120 71500 28160
rect 71540 28120 71541 28160
rect 71499 28111 71541 28120
rect 71116 27448 71444 27488
rect 71500 27404 71540 28111
rect 70828 27364 71060 27404
rect 71404 27364 71540 27404
rect 70443 26060 70485 26069
rect 70443 26020 70444 26060
rect 70484 26020 70485 26060
rect 70443 26011 70485 26020
rect 70635 26060 70677 26069
rect 70635 26020 70636 26060
rect 70676 26020 70677 26060
rect 70635 26011 70677 26020
rect 70444 25926 70484 26011
rect 70539 25976 70581 25985
rect 70539 25936 70540 25976
rect 70580 25936 70581 25976
rect 70539 25927 70581 25936
rect 70347 25892 70389 25901
rect 70347 25852 70348 25892
rect 70388 25852 70389 25892
rect 70347 25843 70389 25852
rect 70348 25136 70388 25147
rect 70348 25061 70388 25096
rect 70347 25052 70389 25061
rect 70347 25012 70348 25052
rect 70388 25012 70389 25052
rect 70347 25003 70389 25012
rect 70540 24977 70580 25927
rect 70636 25892 70676 25901
rect 70828 25892 70868 27364
rect 71115 27320 71157 27329
rect 71115 27280 71116 27320
rect 71156 27280 71157 27320
rect 71115 27271 71157 27280
rect 70923 27152 70965 27161
rect 70923 27112 70924 27152
rect 70964 27112 70965 27152
rect 70923 27103 70965 27112
rect 70924 26144 70964 27103
rect 71019 26312 71061 26321
rect 71019 26272 71020 26312
rect 71060 26272 71061 26312
rect 71019 26263 71061 26272
rect 70924 26095 70964 26104
rect 71020 25976 71060 26263
rect 70676 25852 70868 25892
rect 70924 25936 71060 25976
rect 70636 25843 70676 25852
rect 70732 25565 70772 25852
rect 70731 25556 70773 25565
rect 70731 25516 70732 25556
rect 70772 25516 70773 25556
rect 70731 25507 70773 25516
rect 70636 25220 70676 25229
rect 70539 24968 70581 24977
rect 70539 24928 70540 24968
rect 70580 24928 70581 24968
rect 70539 24919 70581 24928
rect 70636 24464 70676 25180
rect 70732 24632 70772 25507
rect 70732 24583 70772 24592
rect 70924 24632 70964 25936
rect 71020 25304 71060 25313
rect 71020 24809 71060 25264
rect 71019 24800 71061 24809
rect 71019 24760 71020 24800
rect 71060 24760 71061 24800
rect 71019 24751 71061 24760
rect 70924 24583 70964 24592
rect 71019 24632 71061 24641
rect 71019 24592 71020 24632
rect 71060 24592 71061 24632
rect 71019 24583 71061 24592
rect 71020 24498 71060 24583
rect 70732 24464 70772 24473
rect 70636 24424 70732 24464
rect 70732 24415 70772 24424
rect 70155 23960 70197 23969
rect 70155 23920 70156 23960
rect 70196 23920 70197 23960
rect 70155 23911 70197 23920
rect 70539 23960 70581 23969
rect 70539 23920 70540 23960
rect 70580 23920 70581 23960
rect 70539 23911 70581 23920
rect 70827 23960 70869 23969
rect 70827 23920 70828 23960
rect 70868 23920 70869 23960
rect 70827 23911 70869 23920
rect 70155 23792 70197 23801
rect 68948 23752 69236 23792
rect 68908 23743 68948 23752
rect 69004 23624 69044 23633
rect 69004 23060 69044 23584
rect 69196 23060 69236 23752
rect 69332 23752 69620 23792
rect 69292 23743 69332 23752
rect 69388 23624 69428 23633
rect 69388 23060 69428 23584
rect 69580 23060 69620 23752
rect 69716 23752 70004 23792
rect 69676 23743 69716 23752
rect 69772 23624 69812 23633
rect 69772 23060 69812 23584
rect 69964 23060 70004 23752
rect 70155 23752 70156 23792
rect 70196 23752 70197 23792
rect 70155 23743 70197 23752
rect 70443 23792 70485 23801
rect 70443 23752 70444 23792
rect 70484 23752 70485 23792
rect 70443 23743 70485 23752
rect 70540 23792 70580 23911
rect 70540 23743 70580 23752
rect 70156 23658 70196 23743
rect 70252 23624 70292 23633
rect 70252 23060 70292 23584
rect 70444 23060 70484 23743
rect 70636 23624 70676 23633
rect 70636 23060 70676 23584
rect 70828 23060 70868 23911
rect 70924 23792 70964 23801
rect 71116 23792 71156 27271
rect 71307 26228 71349 26237
rect 71307 26188 71308 26228
rect 71348 26188 71349 26228
rect 71307 26179 71349 26188
rect 71212 26144 71252 26153
rect 71212 25481 71252 26104
rect 71308 26094 71348 26179
rect 71404 25808 71444 27364
rect 71596 27161 71636 29035
rect 71692 28916 71732 28925
rect 71692 27833 71732 28876
rect 71788 28328 71828 28337
rect 71828 28288 71924 28328
rect 71788 28279 71828 28288
rect 71691 27824 71733 27833
rect 71691 27784 71692 27824
rect 71732 27784 71733 27824
rect 71691 27775 71733 27784
rect 71787 27656 71829 27665
rect 71787 27616 71788 27656
rect 71828 27616 71829 27656
rect 71787 27607 71829 27616
rect 71595 27152 71637 27161
rect 71595 27112 71596 27152
rect 71636 27112 71637 27152
rect 71595 27103 71637 27112
rect 71691 27068 71733 27077
rect 71691 27028 71692 27068
rect 71732 27028 71733 27068
rect 71691 27019 71733 27028
rect 71692 26900 71732 27019
rect 71692 26851 71732 26860
rect 71500 26648 71540 26657
rect 71500 26237 71540 26608
rect 71788 26321 71828 27607
rect 71884 27488 71924 28288
rect 71884 27439 71924 27448
rect 71883 27152 71925 27161
rect 71883 27112 71884 27152
rect 71924 27112 71925 27152
rect 71883 27103 71925 27112
rect 71884 27068 71924 27103
rect 71884 27017 71924 27028
rect 71980 27068 72020 29044
rect 72652 28328 72692 28337
rect 72076 27068 72116 27077
rect 71980 27028 72076 27068
rect 71883 26648 71925 26657
rect 71883 26608 71884 26648
rect 71924 26608 71925 26648
rect 71883 26599 71925 26608
rect 71884 26514 71924 26599
rect 71980 26489 72020 27028
rect 72076 27019 72116 27028
rect 72268 26900 72308 26909
rect 72268 26741 72308 26860
rect 72267 26732 72309 26741
rect 72267 26692 72268 26732
rect 72308 26692 72309 26732
rect 72267 26683 72309 26692
rect 71979 26480 72021 26489
rect 71979 26440 71980 26480
rect 72020 26440 72021 26480
rect 71979 26431 72021 26440
rect 71787 26312 71829 26321
rect 71787 26272 71788 26312
rect 71828 26272 71924 26312
rect 71787 26263 71829 26272
rect 71499 26228 71541 26237
rect 71499 26188 71500 26228
rect 71540 26188 71541 26228
rect 71499 26179 71541 26188
rect 71884 26228 71924 26272
rect 71884 26179 71924 26188
rect 71788 26144 71828 26153
rect 71596 25976 71636 25985
rect 71788 25976 71828 26104
rect 71980 26144 72020 26431
rect 71980 26095 72020 26104
rect 71636 25936 71828 25976
rect 71596 25927 71636 25936
rect 72652 25901 72692 28288
rect 73035 26900 73077 26909
rect 73035 26860 73036 26900
rect 73076 26860 73077 26900
rect 73035 26851 73077 26860
rect 73036 26816 73076 26851
rect 73036 26765 73076 26776
rect 71979 25892 72021 25901
rect 71979 25852 71980 25892
rect 72020 25852 72021 25892
rect 71979 25843 72021 25852
rect 72651 25892 72693 25901
rect 72651 25852 72652 25892
rect 72692 25852 72693 25892
rect 72651 25843 72693 25852
rect 71404 25768 71732 25808
rect 71211 25472 71253 25481
rect 71211 25432 71212 25472
rect 71252 25432 71253 25472
rect 71211 25423 71253 25432
rect 71403 25136 71445 25145
rect 71403 25096 71404 25136
rect 71444 25096 71445 25136
rect 71403 25087 71445 25096
rect 71211 24968 71253 24977
rect 71211 24928 71212 24968
rect 71252 24928 71253 24968
rect 71211 24919 71253 24928
rect 71212 24632 71252 24919
rect 71212 24583 71252 24592
rect 71307 24632 71349 24641
rect 71307 24592 71308 24632
rect 71348 24592 71349 24632
rect 71307 24583 71349 24592
rect 71404 24632 71444 25087
rect 71595 24800 71637 24809
rect 71595 24760 71596 24800
rect 71636 24760 71637 24800
rect 71595 24751 71637 24760
rect 71404 24583 71444 24592
rect 71308 24498 71348 24583
rect 71596 24464 71636 24751
rect 71596 24415 71636 24424
rect 71308 23792 71348 23801
rect 71692 23792 71732 25768
rect 71884 25304 71924 25313
rect 71980 25304 72020 25843
rect 71924 25264 72020 25304
rect 71884 25255 71924 25264
rect 72843 25136 72885 25145
rect 72843 25096 72844 25136
rect 72884 25096 72885 25136
rect 72843 25087 72885 25096
rect 73035 25136 73077 25145
rect 73035 25096 73036 25136
rect 73076 25096 73077 25136
rect 73035 25087 73077 25096
rect 72459 25052 72501 25061
rect 72459 25012 72460 25052
rect 72500 25012 72501 25052
rect 72459 25003 72501 25012
rect 72075 24716 72117 24725
rect 72075 24676 72076 24716
rect 72116 24676 72117 24716
rect 72075 24667 72117 24676
rect 72076 23792 72116 24667
rect 72460 23792 72500 25003
rect 72844 23792 72884 25087
rect 73036 25002 73076 25087
rect 73132 23969 73172 33100
rect 73228 31025 73268 35260
rect 73324 35216 73364 35260
rect 73420 35251 73460 35260
rect 73324 35167 73364 35176
rect 73516 35216 73556 36016
rect 74092 36056 74132 36688
rect 74092 36007 74132 36016
rect 74284 35981 74324 37360
rect 74476 37400 74516 37409
rect 74476 35981 74516 37360
rect 74572 37400 74612 37411
rect 74572 37325 74612 37360
rect 74956 37400 74996 37411
rect 74956 37325 74996 37360
rect 75052 37400 75092 37409
rect 74571 37316 74613 37325
rect 74571 37276 74572 37316
rect 74612 37276 74613 37316
rect 74571 37267 74613 37276
rect 74955 37316 74997 37325
rect 74955 37276 74956 37316
rect 74996 37276 74997 37316
rect 74955 37267 74997 37276
rect 75052 37157 75092 37360
rect 75148 37400 75188 37409
rect 75051 37148 75093 37157
rect 75051 37108 75052 37148
rect 75092 37108 75093 37148
rect 75051 37099 75093 37108
rect 74763 36728 74805 36737
rect 74763 36688 74764 36728
rect 74804 36688 74805 36728
rect 74763 36679 74805 36688
rect 74764 36594 74804 36679
rect 75052 36065 75092 37099
rect 75148 37073 75188 37360
rect 75243 37232 75285 37241
rect 75243 37192 75244 37232
rect 75284 37192 75285 37232
rect 75243 37183 75285 37192
rect 75244 37098 75284 37183
rect 75147 37064 75189 37073
rect 75147 37024 75148 37064
rect 75188 37024 75189 37064
rect 75147 37015 75189 37024
rect 75051 36056 75093 36065
rect 75051 36016 75052 36056
rect 75092 36016 75093 36056
rect 75051 36007 75093 36016
rect 74283 35972 74325 35981
rect 74283 35932 74284 35972
rect 74324 35932 74325 35972
rect 74283 35923 74325 35932
rect 74475 35972 74517 35981
rect 74475 35932 74476 35972
rect 74516 35932 74517 35972
rect 74475 35923 74517 35932
rect 73708 35888 73748 35897
rect 73708 35729 73748 35848
rect 73899 35888 73941 35897
rect 73899 35848 73900 35888
rect 73940 35848 73941 35888
rect 73899 35839 73941 35848
rect 73900 35754 73940 35839
rect 73707 35720 73749 35729
rect 73707 35680 73708 35720
rect 73748 35680 73749 35720
rect 73707 35671 73749 35680
rect 73516 35167 73556 35176
rect 74187 35216 74229 35225
rect 74187 35176 74188 35216
rect 74228 35176 74229 35216
rect 74187 35167 74229 35176
rect 74188 35082 74228 35167
rect 73324 34376 73364 34385
rect 73364 34336 73556 34376
rect 73324 34327 73364 34336
rect 73516 33140 73556 34336
rect 73516 33100 73652 33140
rect 73612 32873 73652 33100
rect 73419 32864 73461 32873
rect 73419 32824 73420 32864
rect 73460 32824 73461 32864
rect 73419 32815 73461 32824
rect 73611 32864 73653 32873
rect 73611 32824 73612 32864
rect 73652 32824 73653 32864
rect 73611 32815 73653 32824
rect 73420 32730 73460 32815
rect 73612 32201 73652 32815
rect 73899 32276 73941 32285
rect 73899 32236 73900 32276
rect 73940 32236 73941 32276
rect 73899 32227 73941 32236
rect 73611 32192 73653 32201
rect 73611 32152 73612 32192
rect 73652 32152 73653 32192
rect 73611 32143 73653 32152
rect 73612 31268 73652 31277
rect 73227 31016 73269 31025
rect 73227 30976 73228 31016
rect 73268 30976 73269 31016
rect 73227 30967 73269 30976
rect 73612 30857 73652 31228
rect 73611 30848 73653 30857
rect 73611 30808 73612 30848
rect 73652 30808 73653 30848
rect 73611 30799 73653 30808
rect 73900 30176 73940 32227
rect 74092 32024 74132 32033
rect 73996 31984 74092 32024
rect 73996 31352 74036 31984
rect 74092 31975 74132 31984
rect 73996 31303 74036 31312
rect 74092 30428 74132 30437
rect 73900 30136 74036 30176
rect 73707 30008 73749 30017
rect 73707 29968 73708 30008
rect 73748 29968 73749 30008
rect 73707 29959 73749 29968
rect 73900 30008 73940 30017
rect 73420 29126 73460 29135
rect 73420 28757 73460 29086
rect 73419 28748 73461 28757
rect 73419 28708 73420 28748
rect 73460 28708 73461 28748
rect 73419 28699 73461 28708
rect 73516 27488 73556 27497
rect 73516 27152 73556 27448
rect 73420 27112 73556 27152
rect 73420 26852 73460 27112
rect 73420 26803 73460 26812
rect 73227 25976 73269 25985
rect 73227 25936 73228 25976
rect 73268 25936 73269 25976
rect 73227 25927 73269 25936
rect 73420 25934 73460 25943
rect 73228 25304 73268 25927
rect 73420 25640 73460 25894
rect 73420 25600 73556 25640
rect 73516 25304 73556 25600
rect 73612 25304 73652 25313
rect 73516 25264 73612 25304
rect 73228 25255 73268 25264
rect 73612 25255 73652 25264
rect 73131 23960 73173 23969
rect 73131 23920 73132 23960
rect 73172 23920 73173 23960
rect 73131 23911 73173 23920
rect 73323 23960 73365 23969
rect 73323 23920 73324 23960
rect 73364 23920 73365 23960
rect 73323 23911 73365 23920
rect 73611 23960 73653 23969
rect 73611 23920 73612 23960
rect 73652 23920 73653 23960
rect 73611 23911 73653 23920
rect 73324 23792 73364 23911
rect 71116 23752 71308 23792
rect 71348 23752 71636 23792
rect 70924 23633 70964 23752
rect 71308 23743 71348 23752
rect 70923 23624 70965 23633
rect 70923 23584 70924 23624
rect 70964 23584 70965 23624
rect 70923 23575 70965 23584
rect 71020 23624 71060 23633
rect 71020 23060 71060 23584
rect 71211 23624 71253 23633
rect 71211 23584 71212 23624
rect 71252 23584 71253 23624
rect 71211 23575 71253 23584
rect 71404 23624 71444 23633
rect 71212 23060 71252 23575
rect 71404 23060 71444 23584
rect 71596 23060 71636 23752
rect 71732 23752 72020 23792
rect 71692 23743 71732 23752
rect 71788 23624 71828 23633
rect 71788 23060 71828 23584
rect 71980 23060 72020 23752
rect 72116 23752 72404 23792
rect 72076 23743 72116 23752
rect 72172 23624 72212 23633
rect 72172 23060 72212 23584
rect 72364 23060 72404 23752
rect 72500 23752 72692 23792
rect 72460 23743 72500 23752
rect 72556 23624 72596 23633
rect 64012 23020 64095 23060
rect 64204 23020 64340 23060
rect 64396 23020 64495 23060
rect 64588 23020 64724 23060
rect 64780 23020 64895 23060
rect 64972 23020 65108 23060
rect 65164 23020 65295 23060
rect 65356 23020 65585 23060
rect 65644 23020 65695 23060
rect 65836 23020 65985 23060
rect 66028 23020 66095 23060
rect 66220 23020 66356 23060
rect 66412 23020 66495 23060
rect 66604 23020 66740 23060
rect 66796 23020 66895 23060
rect 66988 23020 67124 23060
rect 67180 23020 67295 23060
rect 67372 23020 67508 23060
rect 67564 23020 67700 23060
rect 67756 23020 67985 23060
rect 68044 23020 68095 23060
rect 68236 23020 68385 23060
rect 68428 23020 68495 23060
rect 68620 23020 68756 23060
rect 68812 23020 68895 23060
rect 69004 23020 69140 23060
rect 69196 23020 69295 23060
rect 69388 23020 69524 23060
rect 69580 23020 69695 23060
rect 69772 23020 69908 23060
rect 69964 23020 70095 23060
rect 70252 23020 70385 23060
rect 70444 23020 70495 23060
rect 70636 23020 70785 23060
rect 70828 23020 70895 23060
rect 71020 23020 71156 23060
rect 71212 23020 71295 23060
rect 71404 23020 71540 23060
rect 71596 23020 71695 23060
rect 71788 23020 71924 23060
rect 71980 23020 72095 23060
rect 72172 23020 72308 23060
rect 72364 23020 72495 23060
rect 63916 22744 63985 22784
rect 63945 22596 63985 22744
rect 64055 22596 64095 23020
rect 64300 22784 64340 23020
rect 64300 22744 64385 22784
rect 64345 22596 64385 22744
rect 64455 22596 64495 23020
rect 64684 22784 64724 23020
rect 64684 22744 64785 22784
rect 64745 22596 64785 22744
rect 64855 22596 64895 23020
rect 65068 22784 65108 23020
rect 65068 22744 65185 22784
rect 65145 22596 65185 22744
rect 65255 22596 65295 23020
rect 65545 22596 65585 23020
rect 65655 22596 65695 23020
rect 65945 22596 65985 23020
rect 66055 22596 66095 23020
rect 66316 22784 66356 23020
rect 66316 22744 66385 22784
rect 66345 22596 66385 22744
rect 66455 22596 66495 23020
rect 66700 22784 66740 23020
rect 66700 22744 66785 22784
rect 66745 22596 66785 22744
rect 66855 22596 66895 23020
rect 67084 22784 67124 23020
rect 67084 22744 67185 22784
rect 67145 22596 67185 22744
rect 67255 22596 67295 23020
rect 67468 22784 67508 23020
rect 67660 22784 67700 23020
rect 67468 22744 67585 22784
rect 67545 22596 67585 22744
rect 67655 22744 67700 22784
rect 67655 22596 67695 22744
rect 67945 22596 67985 23020
rect 68055 22596 68095 23020
rect 68345 22596 68385 23020
rect 68455 22596 68495 23020
rect 68716 22784 68756 23020
rect 68716 22744 68785 22784
rect 68745 22596 68785 22744
rect 68855 22596 68895 23020
rect 69100 22784 69140 23020
rect 69100 22744 69185 22784
rect 69145 22596 69185 22744
rect 69255 22596 69295 23020
rect 69484 22784 69524 23020
rect 69484 22744 69585 22784
rect 69545 22596 69585 22744
rect 69655 22596 69695 23020
rect 69868 22784 69908 23020
rect 69868 22744 69985 22784
rect 69945 22596 69985 22744
rect 70055 22596 70095 23020
rect 70345 22596 70385 23020
rect 70455 22596 70495 23020
rect 70745 22596 70785 23020
rect 70855 22596 70895 23020
rect 71116 22784 71156 23020
rect 71116 22744 71185 22784
rect 71145 22596 71185 22744
rect 71255 22596 71295 23020
rect 71500 22784 71540 23020
rect 71500 22744 71585 22784
rect 71545 22596 71585 22744
rect 71655 22596 71695 23020
rect 71884 22784 71924 23020
rect 71884 22744 71985 22784
rect 71945 22596 71985 22744
rect 72055 22596 72095 23020
rect 72268 22784 72308 23020
rect 72268 22744 72385 22784
rect 72345 22596 72385 22744
rect 72455 22596 72495 23020
rect 72556 22784 72596 23584
rect 72652 23060 72692 23752
rect 72884 23752 73268 23792
rect 72844 23743 72884 23752
rect 72940 23624 72980 23633
rect 72940 23060 72980 23584
rect 73228 23060 73268 23752
rect 73324 23743 73364 23752
rect 73420 23624 73460 23633
rect 73460 23584 73556 23624
rect 73420 23556 73460 23584
rect 72652 23020 72895 23060
rect 72940 23020 73185 23060
rect 73228 23020 73295 23060
rect 72556 22744 72785 22784
rect 72745 22596 72785 22744
rect 72855 22596 72895 23020
rect 73145 22596 73185 23020
rect 73255 22596 73295 23020
rect 73516 22784 73556 23584
rect 73612 23060 73652 23911
rect 73708 23792 73748 29959
rect 73804 29168 73844 29177
rect 73900 29168 73940 29968
rect 73844 29128 73940 29168
rect 73804 29119 73844 29128
rect 73803 28580 73845 28589
rect 73803 28540 73804 28580
rect 73844 28540 73845 28580
rect 73803 28531 73845 28540
rect 73804 28446 73844 28531
rect 73804 28160 73844 28169
rect 73804 23969 73844 28120
rect 73803 23960 73845 23969
rect 73803 23920 73804 23960
rect 73844 23920 73845 23960
rect 73803 23911 73845 23920
rect 73996 23876 74036 30136
rect 74092 30017 74132 30388
rect 74091 30008 74133 30017
rect 74091 29968 74092 30008
rect 74132 29968 74133 30008
rect 74091 29959 74133 29968
rect 74284 28001 74324 35923
rect 74572 35216 74612 35225
rect 75340 35216 75380 38200
rect 75916 38072 75956 38081
rect 75820 38032 75916 38072
rect 75820 37400 75860 38032
rect 75916 38023 75956 38032
rect 75820 37351 75860 37360
rect 76587 37400 76629 37409
rect 76587 37360 76588 37400
rect 76628 37360 76629 37400
rect 76587 37351 76629 37360
rect 76684 37400 76724 37409
rect 75436 37316 75476 37325
rect 75476 37276 75668 37316
rect 75436 37267 75476 37276
rect 75531 37064 75573 37073
rect 75531 37024 75532 37064
rect 75572 37024 75573 37064
rect 75531 37015 75573 37024
rect 75436 35216 75476 35225
rect 74612 35176 74708 35216
rect 75340 35176 75436 35216
rect 74572 35167 74612 35176
rect 74379 34964 74421 34973
rect 74379 34924 74380 34964
rect 74420 34924 74421 34964
rect 74379 34915 74421 34924
rect 74283 27992 74325 28001
rect 74283 27952 74284 27992
rect 74324 27952 74325 27992
rect 74283 27943 74325 27952
rect 74380 26984 74420 34915
rect 74668 34544 74708 35176
rect 74668 34495 74708 34504
rect 75339 34376 75381 34385
rect 75339 34336 75340 34376
rect 75380 34336 75381 34376
rect 75339 34327 75381 34336
rect 74476 34208 74516 34217
rect 74476 33545 74516 34168
rect 74475 33536 74517 33545
rect 74475 33496 74476 33536
rect 74516 33496 74517 33536
rect 74475 33487 74517 33496
rect 75148 33536 75188 33545
rect 74763 33452 74805 33461
rect 74763 33412 74764 33452
rect 74804 33412 74805 33452
rect 74763 33403 74805 33412
rect 74764 32864 74804 33403
rect 74764 32815 74804 32824
rect 74859 32864 74901 32873
rect 74859 32824 74860 32864
rect 74900 32824 74901 32864
rect 74859 32815 74901 32824
rect 75148 32864 75188 33496
rect 75148 32815 75188 32824
rect 74572 32696 74612 32705
rect 74572 32285 74612 32656
rect 74571 32276 74613 32285
rect 74571 32236 74572 32276
rect 74612 32236 74613 32276
rect 74571 32227 74613 32236
rect 74860 31352 74900 32815
rect 75147 32696 75189 32705
rect 75147 32656 75148 32696
rect 75188 32656 75189 32696
rect 75147 32647 75189 32656
rect 74668 31312 74860 31352
rect 74571 31184 74613 31193
rect 74571 31144 74572 31184
rect 74612 31144 74613 31184
rect 74571 31135 74613 31144
rect 74092 26944 74420 26984
rect 74092 24053 74132 26944
rect 74284 26816 74324 26825
rect 74324 26776 74420 26816
rect 74284 26767 74324 26776
rect 74188 26144 74228 26153
rect 74188 24800 74228 26104
rect 74284 26144 74324 26153
rect 74284 25565 74324 26104
rect 74380 25901 74420 26776
rect 74476 26153 74516 26238
rect 74475 26144 74517 26153
rect 74475 26104 74476 26144
rect 74516 26104 74517 26144
rect 74475 26095 74517 26104
rect 74475 25976 74517 25985
rect 74475 25936 74476 25976
rect 74516 25936 74517 25976
rect 74475 25927 74517 25936
rect 74379 25892 74421 25901
rect 74379 25852 74380 25892
rect 74420 25852 74421 25892
rect 74379 25843 74421 25852
rect 74283 25556 74325 25565
rect 74283 25516 74284 25556
rect 74324 25516 74325 25556
rect 74283 25507 74325 25516
rect 74380 25304 74420 25843
rect 74476 25842 74516 25927
rect 74475 25304 74517 25313
rect 74380 25264 74476 25304
rect 74516 25264 74517 25304
rect 74475 25255 74517 25264
rect 74476 25170 74516 25255
rect 74572 25052 74612 31135
rect 74668 29168 74708 31312
rect 74860 31303 74900 31312
rect 74859 31016 74901 31025
rect 74859 30976 74860 31016
rect 74900 30976 74901 31016
rect 74859 30967 74901 30976
rect 74860 30848 74900 30967
rect 75148 30890 75188 32647
rect 75340 31100 75380 34327
rect 75436 32873 75476 35176
rect 75532 34385 75572 37015
rect 75628 36644 75668 37276
rect 76107 37232 76149 37241
rect 76107 37192 76108 37232
rect 76148 37192 76149 37232
rect 76107 37183 76149 37192
rect 76108 36728 76148 37183
rect 76299 36812 76341 36821
rect 76299 36772 76300 36812
rect 76340 36772 76341 36812
rect 76299 36763 76341 36772
rect 76108 36679 76148 36688
rect 76300 36728 76340 36763
rect 76300 36677 76340 36688
rect 76396 36728 76436 36737
rect 75628 36604 76052 36644
rect 76012 36560 76052 36604
rect 76108 36560 76148 36569
rect 76012 36520 76108 36560
rect 76108 36511 76148 36520
rect 75916 36476 75956 36485
rect 75723 36056 75765 36065
rect 75723 36016 75724 36056
rect 75764 36016 75765 36056
rect 75723 36007 75765 36016
rect 75531 34376 75573 34385
rect 75628 34376 75668 34385
rect 75531 34336 75532 34376
rect 75572 34336 75628 34376
rect 75531 34327 75573 34336
rect 75628 34327 75668 34336
rect 75724 34376 75764 36007
rect 75916 35897 75956 36436
rect 76396 36056 76436 36688
rect 76588 36728 76628 37351
rect 76684 36737 76724 37360
rect 76875 37316 76917 37325
rect 76875 37276 76876 37316
rect 76916 37276 76917 37316
rect 76875 37267 76917 37276
rect 76779 36812 76821 36821
rect 76779 36772 76780 36812
rect 76820 36772 76821 36812
rect 76779 36763 76821 36772
rect 76588 36679 76628 36688
rect 76683 36728 76725 36737
rect 76683 36688 76684 36728
rect 76724 36688 76725 36728
rect 76683 36679 76725 36688
rect 76780 36728 76820 36763
rect 76780 36677 76820 36688
rect 76876 36728 76916 37267
rect 76876 36679 76916 36688
rect 76587 36560 76629 36569
rect 76587 36520 76588 36560
rect 76628 36520 76629 36560
rect 76587 36511 76629 36520
rect 76588 36426 76628 36511
rect 76779 36392 76821 36401
rect 76779 36352 76780 36392
rect 76820 36352 76821 36392
rect 76779 36343 76821 36352
rect 76300 36016 76436 36056
rect 75915 35888 75957 35897
rect 75915 35848 75916 35888
rect 75956 35848 75957 35888
rect 75915 35839 75957 35848
rect 76203 35888 76245 35897
rect 76203 35848 76204 35888
rect 76244 35848 76245 35888
rect 76203 35839 76245 35848
rect 75820 34385 75860 34470
rect 75531 34208 75573 34217
rect 75531 34168 75532 34208
rect 75572 34168 75573 34208
rect 75531 34159 75573 34168
rect 75532 34074 75572 34159
rect 75724 34124 75764 34336
rect 75819 34376 75861 34385
rect 75819 34336 75820 34376
rect 75860 34336 75861 34376
rect 75819 34327 75861 34336
rect 75628 34084 75764 34124
rect 75628 33140 75668 34084
rect 75819 33788 75861 33797
rect 75819 33748 75820 33788
rect 75860 33748 75861 33788
rect 75819 33739 75861 33748
rect 75532 33100 75668 33140
rect 75724 33704 75764 33713
rect 75435 32864 75477 32873
rect 75435 32824 75436 32864
rect 75476 32824 75477 32864
rect 75435 32815 75477 32824
rect 75532 31277 75572 33100
rect 75724 32360 75764 33664
rect 75820 33704 75860 33739
rect 75820 33653 75860 33664
rect 75916 32705 75956 35839
rect 76204 35754 76244 35839
rect 76300 35804 76340 36016
rect 76395 35888 76437 35897
rect 76395 35848 76396 35888
rect 76436 35848 76437 35888
rect 76395 35839 76437 35848
rect 76492 35888 76532 35897
rect 76300 35755 76340 35764
rect 76011 35216 76053 35225
rect 76011 35176 76012 35216
rect 76052 35176 76053 35216
rect 76011 35167 76053 35176
rect 76012 34544 76052 35167
rect 76396 34637 76436 35839
rect 76492 35384 76532 35848
rect 76588 35384 76628 35393
rect 76492 35344 76588 35384
rect 76588 35335 76628 35344
rect 76588 34964 76628 34973
rect 76628 34924 76724 34964
rect 76588 34915 76628 34924
rect 76587 34712 76629 34721
rect 76587 34672 76588 34712
rect 76628 34672 76629 34712
rect 76587 34663 76629 34672
rect 76395 34628 76437 34637
rect 76395 34588 76396 34628
rect 76436 34588 76437 34628
rect 76395 34579 76437 34588
rect 76012 34495 76052 34504
rect 76203 34544 76245 34553
rect 76203 34504 76204 34544
rect 76244 34504 76245 34544
rect 76203 34495 76245 34504
rect 76012 34376 76052 34385
rect 76012 34217 76052 34336
rect 76204 34376 76244 34495
rect 76588 34469 76628 34663
rect 76587 34460 76629 34469
rect 76587 34420 76588 34460
rect 76628 34420 76629 34460
rect 76587 34411 76629 34420
rect 76204 34327 76244 34336
rect 76300 34376 76340 34385
rect 76011 34208 76053 34217
rect 76011 34168 76012 34208
rect 76052 34168 76053 34208
rect 76011 34159 76053 34168
rect 76300 33881 76340 34336
rect 76588 34376 76628 34411
rect 76684 34385 76724 34924
rect 76588 34326 76628 34336
rect 76683 34376 76725 34385
rect 76683 34336 76684 34376
rect 76724 34336 76725 34376
rect 76683 34327 76725 34336
rect 76299 33872 76341 33881
rect 76299 33832 76300 33872
rect 76340 33832 76341 33872
rect 76299 33823 76341 33832
rect 76684 33713 76724 33798
rect 76012 33704 76052 33713
rect 76204 33704 76244 33713
rect 76052 33664 76204 33704
rect 76012 33655 76052 33664
rect 76204 33655 76244 33664
rect 76300 33704 76340 33713
rect 76203 33536 76245 33545
rect 76203 33496 76204 33536
rect 76244 33496 76245 33536
rect 76203 33487 76245 33496
rect 76011 33452 76053 33461
rect 76011 33412 76012 33452
rect 76052 33412 76053 33452
rect 76011 33403 76053 33412
rect 76012 33318 76052 33403
rect 76011 32864 76053 32873
rect 76011 32824 76012 32864
rect 76052 32824 76053 32864
rect 76011 32815 76053 32824
rect 76012 32730 76052 32815
rect 75915 32696 75957 32705
rect 75915 32656 75916 32696
rect 75956 32656 75957 32696
rect 75915 32647 75957 32656
rect 75916 32360 75956 32369
rect 75724 32320 75916 32360
rect 75916 32311 75956 32320
rect 75819 32192 75861 32201
rect 75819 32152 75820 32192
rect 75860 32152 75861 32192
rect 75819 32143 75861 32152
rect 76012 32192 76052 32201
rect 75531 31268 75573 31277
rect 75531 31228 75532 31268
rect 75572 31228 75573 31268
rect 75531 31219 75573 31228
rect 75340 31060 75764 31100
rect 75339 30932 75381 30941
rect 75339 30892 75340 30932
rect 75380 30892 75381 30932
rect 75148 30850 75284 30890
rect 75339 30883 75381 30892
rect 75531 30932 75573 30941
rect 75531 30892 75532 30932
rect 75572 30892 75573 30932
rect 75531 30883 75573 30892
rect 74860 30799 74900 30808
rect 74763 30680 74805 30689
rect 74955 30680 74997 30689
rect 74763 30640 74764 30680
rect 74804 30640 74900 30680
rect 74763 30631 74805 30640
rect 74860 30521 74900 30640
rect 74955 30640 74956 30680
rect 74996 30640 74997 30680
rect 74955 30631 74997 30640
rect 75052 30680 75092 30689
rect 74859 30512 74901 30521
rect 74859 30472 74860 30512
rect 74900 30472 74901 30512
rect 74859 30463 74901 30472
rect 74956 30437 74996 30631
rect 75052 30521 75092 30640
rect 75147 30680 75189 30689
rect 75147 30640 75148 30680
rect 75188 30640 75189 30680
rect 75147 30631 75189 30640
rect 75148 30546 75188 30631
rect 75051 30512 75093 30521
rect 75051 30472 75052 30512
rect 75092 30472 75093 30512
rect 75051 30463 75093 30472
rect 74955 30428 74997 30437
rect 74955 30388 74956 30428
rect 74996 30388 74997 30428
rect 74955 30379 74997 30388
rect 74956 30269 74996 30379
rect 74955 30260 74997 30269
rect 74955 30220 74956 30260
rect 74996 30220 74997 30260
rect 74955 30211 74997 30220
rect 75244 30092 75284 30850
rect 75340 30680 75380 30883
rect 75435 30848 75477 30857
rect 75435 30808 75436 30848
rect 75476 30808 75477 30848
rect 75435 30799 75477 30808
rect 75436 30714 75476 30799
rect 75340 30631 75380 30640
rect 75532 30680 75572 30883
rect 75532 30631 75572 30640
rect 75628 30680 75668 30689
rect 75435 30512 75477 30521
rect 75435 30472 75436 30512
rect 75476 30472 75477 30512
rect 75435 30463 75477 30472
rect 75339 30260 75381 30269
rect 75339 30220 75340 30260
rect 75380 30220 75381 30260
rect 75339 30211 75381 30220
rect 74956 30052 75284 30092
rect 74859 29756 74901 29765
rect 74859 29716 74860 29756
rect 74900 29716 74901 29756
rect 74859 29707 74901 29716
rect 74860 29672 74900 29707
rect 74860 29621 74900 29632
rect 74668 29119 74708 29128
rect 74860 27656 74900 27665
rect 74764 27616 74860 27656
rect 74667 27068 74709 27077
rect 74667 27028 74668 27068
rect 74708 27028 74709 27068
rect 74667 27019 74709 27028
rect 74668 26648 74708 27019
rect 74764 26825 74804 27616
rect 74860 27607 74900 27616
rect 74860 27404 74900 27413
rect 74860 26909 74900 27364
rect 74859 26900 74901 26909
rect 74859 26860 74860 26900
rect 74900 26860 74901 26900
rect 74859 26851 74901 26860
rect 74763 26816 74805 26825
rect 74763 26776 74764 26816
rect 74804 26776 74805 26816
rect 74763 26767 74805 26776
rect 74859 26732 74901 26741
rect 74859 26692 74860 26732
rect 74900 26692 74901 26732
rect 74859 26683 74901 26692
rect 74668 26608 74804 26648
rect 74764 26405 74804 26608
rect 74763 26396 74805 26405
rect 74763 26356 74764 26396
rect 74804 26356 74805 26396
rect 74763 26347 74805 26356
rect 74667 26144 74709 26153
rect 74667 26104 74668 26144
rect 74708 26104 74709 26144
rect 74667 26095 74709 26104
rect 74764 26144 74804 26347
rect 74860 26237 74900 26683
rect 74956 26312 74996 30052
rect 75051 29924 75093 29933
rect 75051 29884 75052 29924
rect 75092 29884 75093 29924
rect 75051 29875 75093 29884
rect 75052 29790 75092 29875
rect 75340 29840 75380 30211
rect 75340 29791 75380 29800
rect 75436 29840 75476 30463
rect 75531 30260 75573 30269
rect 75531 30220 75532 30260
rect 75572 30220 75573 30260
rect 75531 30211 75573 30220
rect 75532 30008 75572 30211
rect 75628 30092 75668 30640
rect 75724 30269 75764 31060
rect 75723 30260 75765 30269
rect 75723 30220 75724 30260
rect 75764 30220 75765 30260
rect 75723 30211 75765 30220
rect 75724 30092 75764 30101
rect 75628 30052 75724 30092
rect 75724 30043 75764 30052
rect 75532 29968 75668 30008
rect 75436 29791 75476 29800
rect 75531 29840 75573 29849
rect 75531 29800 75532 29840
rect 75572 29800 75573 29840
rect 75531 29791 75573 29800
rect 75532 29706 75572 29791
rect 75244 29672 75284 29681
rect 75244 28328 75284 29632
rect 75339 28748 75381 28757
rect 75339 28708 75340 28748
rect 75380 28708 75381 28748
rect 75339 28699 75381 28708
rect 75244 28279 75284 28288
rect 75340 28244 75380 28699
rect 75435 28328 75477 28337
rect 75435 28288 75436 28328
rect 75476 28288 75477 28328
rect 75435 28279 75477 28288
rect 75532 28328 75572 28337
rect 75340 28195 75380 28204
rect 75436 28194 75476 28279
rect 75435 27992 75477 28001
rect 75435 27952 75436 27992
rect 75476 27952 75477 27992
rect 75435 27943 75477 27952
rect 75051 27656 75093 27665
rect 75051 27616 75052 27656
rect 75092 27616 75093 27656
rect 75051 27607 75093 27616
rect 75148 27656 75188 27665
rect 75436 27656 75476 27943
rect 75532 27824 75572 28288
rect 75628 27824 75668 29968
rect 75820 29924 75860 32143
rect 76012 31781 76052 32152
rect 76108 32192 76148 32201
rect 76011 31772 76053 31781
rect 76011 31732 76012 31772
rect 76052 31732 76053 31772
rect 76011 31723 76053 31732
rect 76012 31604 76052 31613
rect 76108 31604 76148 32152
rect 76052 31564 76148 31604
rect 76012 31555 76052 31564
rect 75915 31520 75957 31529
rect 75915 31480 75916 31520
rect 75956 31480 75957 31520
rect 75915 31471 75957 31480
rect 75916 30437 75956 31471
rect 76012 31184 76052 31193
rect 76012 30689 76052 31144
rect 76204 30848 76244 33487
rect 76108 30808 76244 30848
rect 76011 30680 76053 30689
rect 76011 30640 76012 30680
rect 76052 30640 76053 30680
rect 76011 30631 76053 30640
rect 75915 30428 75957 30437
rect 75915 30388 75916 30428
rect 75956 30388 75957 30428
rect 75915 30379 75957 30388
rect 75724 29884 75860 29924
rect 75724 29840 75764 29884
rect 75724 29791 75764 29800
rect 75916 29840 75956 29851
rect 75916 29765 75956 29800
rect 76011 29840 76053 29849
rect 76011 29800 76012 29840
rect 76052 29800 76053 29840
rect 76011 29791 76053 29800
rect 75915 29756 75957 29765
rect 75915 29716 75916 29756
rect 75956 29716 75957 29756
rect 75915 29707 75957 29716
rect 76012 29513 76052 29791
rect 76011 29504 76053 29513
rect 75820 29464 76012 29504
rect 76052 29464 76053 29504
rect 75820 29336 75860 29464
rect 76011 29455 76053 29464
rect 76108 29336 76148 30808
rect 76300 30773 76340 33664
rect 76396 33704 76436 33713
rect 76299 30764 76341 30773
rect 76299 30724 76300 30764
rect 76340 30724 76341 30764
rect 76299 30715 76341 30724
rect 76204 30680 76244 30689
rect 76204 30437 76244 30640
rect 76396 30521 76436 33664
rect 76492 33704 76532 33713
rect 76492 33461 76532 33664
rect 76587 33704 76629 33713
rect 76587 33664 76588 33704
rect 76628 33664 76629 33704
rect 76587 33655 76629 33664
rect 76683 33704 76725 33713
rect 76683 33664 76684 33704
rect 76724 33664 76725 33704
rect 76683 33655 76725 33664
rect 76491 33452 76533 33461
rect 76491 33412 76492 33452
rect 76532 33412 76533 33452
rect 76491 33403 76533 33412
rect 76588 32201 76628 33655
rect 76684 33452 76724 33463
rect 76684 33377 76724 33412
rect 76683 33368 76725 33377
rect 76683 33328 76684 33368
rect 76724 33328 76725 33368
rect 76683 33319 76725 33328
rect 76587 32192 76629 32201
rect 76587 32152 76588 32192
rect 76628 32152 76629 32192
rect 76587 32143 76629 32152
rect 76683 32024 76725 32033
rect 76683 31984 76684 32024
rect 76724 31984 76725 32024
rect 76683 31975 76725 31984
rect 76491 31100 76533 31109
rect 76491 31060 76492 31100
rect 76532 31060 76533 31100
rect 76491 31051 76533 31060
rect 76492 30680 76532 31051
rect 76492 30631 76532 30640
rect 76587 30680 76629 30689
rect 76587 30640 76588 30680
rect 76628 30640 76629 30680
rect 76587 30631 76629 30640
rect 76588 30546 76628 30631
rect 76395 30512 76437 30521
rect 76395 30472 76396 30512
rect 76436 30472 76437 30512
rect 76395 30463 76437 30472
rect 76203 30428 76245 30437
rect 76684 30428 76724 31975
rect 76203 30388 76204 30428
rect 76244 30388 76245 30428
rect 76203 30379 76245 30388
rect 76492 30388 76724 30428
rect 76204 29345 76244 30379
rect 76299 30344 76341 30353
rect 76299 30304 76300 30344
rect 76340 30304 76341 30344
rect 76299 30295 76341 30304
rect 75820 29287 75860 29296
rect 76012 29296 76148 29336
rect 76203 29336 76245 29345
rect 76203 29296 76204 29336
rect 76244 29296 76245 29336
rect 75628 27784 75860 27824
rect 75532 27775 75572 27784
rect 75052 27522 75092 27607
rect 75051 27404 75093 27413
rect 75051 27364 75052 27404
rect 75092 27364 75093 27404
rect 75051 27355 75093 27364
rect 75052 26396 75092 27355
rect 75148 26648 75188 27616
rect 75244 27616 75436 27656
rect 75244 27413 75284 27616
rect 75436 27607 75476 27616
rect 75628 27656 75668 27665
rect 75628 27488 75668 27616
rect 75340 27448 75668 27488
rect 75724 27656 75764 27665
rect 75243 27404 75285 27413
rect 75243 27364 75244 27404
rect 75284 27364 75285 27404
rect 75243 27355 75285 27364
rect 75148 26608 75292 26648
rect 75252 26396 75292 26608
rect 75052 26356 75185 26396
rect 75145 26312 75185 26356
rect 75244 26356 75292 26396
rect 75244 26312 75284 26356
rect 74956 26272 75092 26312
rect 75145 26272 75188 26312
rect 74859 26228 74901 26237
rect 74859 26188 74860 26228
rect 74900 26188 74901 26228
rect 74859 26179 74901 26188
rect 74764 26095 74804 26104
rect 74860 26144 74900 26179
rect 74668 26010 74708 26095
rect 74860 26094 74900 26104
rect 74955 26144 74997 26153
rect 74955 26104 74956 26144
rect 74996 26104 74997 26144
rect 74955 26095 74997 26104
rect 74956 26010 74996 26095
rect 74763 25976 74805 25985
rect 74763 25936 74764 25976
rect 74804 25936 74805 25976
rect 74763 25927 74805 25936
rect 74572 25012 74708 25052
rect 74475 24968 74517 24977
rect 74475 24928 74476 24968
rect 74516 24928 74517 24968
rect 74475 24919 74517 24928
rect 74380 24800 74420 24809
rect 74188 24760 74380 24800
rect 74380 24751 74420 24760
rect 74283 24632 74325 24641
rect 74283 24592 74284 24632
rect 74324 24592 74325 24632
rect 74283 24583 74325 24592
rect 74476 24632 74516 24919
rect 74571 24884 74613 24893
rect 74571 24844 74572 24884
rect 74612 24844 74613 24884
rect 74571 24835 74613 24844
rect 74284 24498 74324 24583
rect 74476 24557 74516 24592
rect 74572 24632 74612 24835
rect 74572 24583 74612 24592
rect 74475 24548 74517 24557
rect 74475 24508 74476 24548
rect 74516 24508 74517 24548
rect 74475 24499 74517 24508
rect 74476 24468 74516 24499
rect 74091 24044 74133 24053
rect 74091 24004 74092 24044
rect 74132 24004 74133 24044
rect 74091 23995 74133 24004
rect 73996 23836 74132 23876
rect 74092 23792 74132 23836
rect 74476 23792 74516 23801
rect 74668 23792 74708 25012
rect 74764 24641 74804 25927
rect 74763 24632 74805 24641
rect 74763 24592 74764 24632
rect 74804 24592 74805 24632
rect 74763 24583 74805 24592
rect 74859 24044 74901 24053
rect 74859 24004 74860 24044
rect 74900 24004 74901 24044
rect 74859 23995 74901 24004
rect 73748 23752 74036 23792
rect 73708 23743 73748 23752
rect 73804 23624 73844 23633
rect 73804 23060 73844 23584
rect 73996 23060 74036 23752
rect 74132 23752 74420 23792
rect 74092 23743 74132 23752
rect 74188 23624 74228 23633
rect 74188 23060 74228 23584
rect 74380 23060 74420 23752
rect 74516 23752 74708 23792
rect 74476 23743 74516 23752
rect 74572 23624 74612 23633
rect 74572 23060 74612 23584
rect 74668 23204 74708 23752
rect 74860 23792 74900 23995
rect 75052 23801 75092 26272
rect 75148 26144 75188 26272
rect 75244 26263 75284 26272
rect 75148 25985 75188 26104
rect 75340 26144 75380 27448
rect 75627 26984 75669 26993
rect 75724 26984 75764 27616
rect 75820 27077 75860 27784
rect 75819 27068 75861 27077
rect 75819 27028 75820 27068
rect 75860 27028 75861 27068
rect 75819 27019 75861 27028
rect 75627 26944 75628 26984
rect 75668 26944 75764 26984
rect 75627 26935 75669 26944
rect 75435 26900 75477 26909
rect 75820 26900 75860 27019
rect 75435 26860 75436 26900
rect 75476 26860 75477 26900
rect 75435 26851 75477 26860
rect 75724 26860 75860 26900
rect 75436 26766 75476 26851
rect 75627 26816 75669 26825
rect 75627 26776 75628 26816
rect 75668 26776 75669 26816
rect 75627 26767 75669 26776
rect 75724 26816 75764 26860
rect 75915 26816 75957 26825
rect 75724 26767 75764 26776
rect 75820 26795 75860 26804
rect 75628 26682 75668 26767
rect 75915 26776 75916 26816
rect 75956 26776 75957 26816
rect 75915 26767 75957 26776
rect 75820 26741 75860 26755
rect 75819 26732 75861 26741
rect 75819 26692 75820 26732
rect 75860 26692 75861 26732
rect 75819 26683 75861 26692
rect 75820 26660 75860 26683
rect 75916 26682 75956 26767
rect 75723 26648 75765 26657
rect 75723 26608 75724 26648
rect 75764 26608 75765 26648
rect 75723 26599 75765 26608
rect 75147 25976 75189 25985
rect 75147 25936 75148 25976
rect 75188 25936 75189 25976
rect 75147 25927 75189 25936
rect 75340 24557 75380 26104
rect 75435 26144 75477 26153
rect 75435 26104 75436 26144
rect 75476 26104 75668 26144
rect 75435 26095 75477 26104
rect 75436 26010 75476 26095
rect 75628 25556 75668 26104
rect 75628 25507 75668 25516
rect 75724 25388 75764 26599
rect 75819 26480 75861 26489
rect 75819 26440 75820 26480
rect 75860 26440 75861 26480
rect 75819 26431 75861 26440
rect 75820 26153 75860 26431
rect 75819 26144 75861 26153
rect 75819 26104 75820 26144
rect 75860 26104 75861 26144
rect 75819 26095 75861 26104
rect 75436 25348 75764 25388
rect 75436 24632 75476 25348
rect 75820 25304 75860 26095
rect 75916 25565 75956 25650
rect 75915 25556 75957 25565
rect 75915 25516 75916 25556
rect 75956 25516 75957 25556
rect 75915 25507 75957 25516
rect 76012 25472 76052 29296
rect 76203 29287 76245 29296
rect 76108 29168 76148 29177
rect 76204 29168 76244 29287
rect 76148 29128 76244 29168
rect 76108 29119 76148 29128
rect 76204 26816 76244 26825
rect 76204 26657 76244 26776
rect 76300 26741 76340 30295
rect 76492 29840 76532 30388
rect 76492 29791 76532 29800
rect 76684 29840 76724 29849
rect 76588 29756 76628 29765
rect 76491 29504 76533 29513
rect 76491 29464 76492 29504
rect 76532 29464 76533 29504
rect 76491 29455 76533 29464
rect 76492 29252 76532 29455
rect 76492 29203 76532 29212
rect 76396 29168 76436 29177
rect 76396 28421 76436 29128
rect 76395 28412 76437 28421
rect 76395 28372 76396 28412
rect 76436 28372 76437 28412
rect 76395 28363 76437 28372
rect 76588 28337 76628 29716
rect 76684 29000 76724 29800
rect 76780 29168 76820 36343
rect 76972 35468 77012 38200
rect 77260 38240 77300 38249
rect 77260 37157 77300 38200
rect 77356 38240 77396 38249
rect 77356 37241 77396 38200
rect 77644 37988 77684 37997
rect 77451 37400 77493 37409
rect 77451 37360 77452 37400
rect 77492 37360 77493 37400
rect 77451 37351 77493 37360
rect 77355 37232 77397 37241
rect 77355 37192 77356 37232
rect 77396 37192 77397 37232
rect 77355 37183 77397 37192
rect 77259 37148 77301 37157
rect 77259 37108 77260 37148
rect 77300 37108 77301 37148
rect 77259 37099 77301 37108
rect 77068 36728 77108 36737
rect 77068 36569 77108 36688
rect 77067 36560 77109 36569
rect 77067 36520 77068 36560
rect 77108 36520 77109 36560
rect 77067 36511 77109 36520
rect 77260 36401 77300 37099
rect 77452 36728 77492 37351
rect 77547 36812 77589 36821
rect 77547 36772 77548 36812
rect 77588 36772 77589 36812
rect 77547 36763 77589 36772
rect 77452 36679 77492 36688
rect 77259 36392 77301 36401
rect 77259 36352 77260 36392
rect 77300 36352 77301 36392
rect 77259 36343 77301 36352
rect 77548 36140 77588 36763
rect 77548 36091 77588 36100
rect 77067 35888 77109 35897
rect 77067 35848 77068 35888
rect 77108 35848 77109 35888
rect 77067 35839 77109 35848
rect 77260 35888 77300 35897
rect 77068 35561 77108 35839
rect 77164 35804 77204 35813
rect 77067 35552 77109 35561
rect 77067 35512 77068 35552
rect 77108 35512 77109 35552
rect 77067 35503 77109 35512
rect 76876 35428 77012 35468
rect 76876 34721 76916 35428
rect 77164 35384 77204 35764
rect 76972 35344 77204 35384
rect 76875 34712 76917 34721
rect 76875 34672 76876 34712
rect 76916 34672 76917 34712
rect 76875 34663 76917 34672
rect 76972 34553 77012 35344
rect 77068 35216 77108 35225
rect 77108 35176 77204 35216
rect 77068 35167 77108 35176
rect 77067 34628 77109 34637
rect 77067 34588 77068 34628
rect 77108 34588 77109 34628
rect 77067 34579 77109 34588
rect 76971 34544 77013 34553
rect 76971 34504 76972 34544
rect 77012 34504 77013 34544
rect 76971 34495 77013 34504
rect 76876 34376 76916 34387
rect 76876 34301 76916 34336
rect 76971 34376 77013 34385
rect 76971 34336 76972 34376
rect 77012 34336 77013 34376
rect 76971 34327 77013 34336
rect 76875 34292 76917 34301
rect 76875 34252 76876 34292
rect 76916 34252 76917 34292
rect 76875 34243 76917 34252
rect 76972 34242 77012 34327
rect 77068 33956 77108 34579
rect 77164 34460 77204 35176
rect 77260 34628 77300 35848
rect 77451 35888 77493 35897
rect 77451 35848 77452 35888
rect 77492 35848 77493 35888
rect 77451 35839 77493 35848
rect 77644 35888 77684 37948
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 78412 37568 78452 37577
rect 78412 37409 78452 37528
rect 78028 37400 78068 37409
rect 77932 37360 78028 37400
rect 77835 37232 77877 37241
rect 77835 37192 77836 37232
rect 77876 37192 77877 37232
rect 77835 37183 77877 37192
rect 77836 37098 77876 37183
rect 77836 36056 77876 36065
rect 77644 35839 77684 35848
rect 77740 36016 77836 36056
rect 77452 35754 77492 35839
rect 77452 35216 77492 35225
rect 77740 35216 77780 36016
rect 77836 36007 77876 36016
rect 77932 35729 77972 37360
rect 78028 37351 78068 37360
rect 78220 37400 78260 37409
rect 78123 37316 78165 37325
rect 78123 37276 78124 37316
rect 78164 37276 78165 37316
rect 78123 37267 78165 37276
rect 78124 37182 78164 37267
rect 78220 37157 78260 37360
rect 78411 37400 78453 37409
rect 78411 37360 78412 37400
rect 78452 37360 78453 37400
rect 78411 37351 78453 37360
rect 78219 37148 78261 37157
rect 78219 37108 78220 37148
rect 78260 37108 78261 37148
rect 78219 37099 78261 37108
rect 79467 37148 79509 37157
rect 79467 37108 79468 37148
rect 79508 37108 79509 37148
rect 79467 37099 79509 37108
rect 79468 36896 79508 37099
rect 79468 36847 79508 36856
rect 78315 36728 78357 36737
rect 78315 36688 78316 36728
rect 78356 36688 78357 36728
rect 78315 36679 78357 36688
rect 78316 36594 78356 36679
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 77931 35720 77973 35729
rect 77931 35680 77932 35720
rect 77972 35680 77973 35720
rect 77931 35671 77973 35680
rect 77492 35176 77780 35216
rect 77452 35167 77492 35176
rect 77260 34579 77300 34588
rect 77452 34544 77492 34553
rect 77356 34504 77452 34544
rect 77356 34460 77396 34504
rect 77452 34495 77492 34504
rect 77643 34544 77685 34553
rect 77643 34504 77644 34544
rect 77684 34504 77685 34544
rect 77643 34495 77685 34504
rect 77164 34420 77396 34460
rect 77452 34376 77492 34385
rect 76886 33916 77108 33956
rect 77356 34336 77452 34376
rect 76886 33872 76926 33916
rect 76876 33832 76926 33872
rect 76876 33704 76916 33832
rect 76876 31697 76916 33664
rect 76972 33704 77012 33713
rect 76972 33461 77012 33664
rect 77259 33704 77301 33713
rect 77356 33704 77396 34336
rect 77452 34327 77492 34336
rect 77644 34376 77684 34495
rect 77644 34327 77684 34336
rect 77740 34376 77780 34385
rect 77740 34208 77780 34336
rect 77932 34376 77972 35671
rect 78316 35216 78356 35225
rect 77932 34327 77972 34336
rect 78123 34376 78165 34385
rect 78123 34336 78124 34376
rect 78164 34336 78165 34376
rect 78123 34327 78165 34336
rect 78028 34292 78068 34301
rect 78028 34208 78068 34252
rect 77740 34168 78068 34208
rect 77259 33664 77260 33704
rect 77300 33664 77396 33704
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77259 33655 77301 33664
rect 77451 33655 77493 33664
rect 77548 33704 77588 33713
rect 77588 33664 77972 33704
rect 77548 33655 77588 33664
rect 77260 33570 77300 33655
rect 77452 33570 77492 33655
rect 77355 33536 77397 33545
rect 77355 33496 77356 33536
rect 77396 33496 77397 33536
rect 77355 33487 77397 33496
rect 77836 33536 77876 33545
rect 76971 33452 77013 33461
rect 76971 33412 76972 33452
rect 77012 33412 77013 33452
rect 76971 33403 77013 33412
rect 77163 33452 77205 33461
rect 77163 33412 77164 33452
rect 77204 33412 77205 33452
rect 77163 33403 77205 33412
rect 77260 33452 77300 33461
rect 77164 33116 77204 33403
rect 77164 33041 77204 33076
rect 77163 33032 77205 33041
rect 77163 32992 77164 33032
rect 77204 32992 77205 33032
rect 77163 32983 77205 32992
rect 77164 32952 77204 32983
rect 76971 32360 77013 32369
rect 77260 32360 77300 33412
rect 76971 32320 76972 32360
rect 77012 32320 77013 32360
rect 76971 32311 77013 32320
rect 77068 32320 77300 32360
rect 76875 31688 76917 31697
rect 76875 31648 76876 31688
rect 76916 31648 76917 31688
rect 76875 31639 76917 31648
rect 76972 31529 77012 32311
rect 77068 32276 77108 32320
rect 77068 32227 77108 32236
rect 77163 32024 77205 32033
rect 77163 31984 77164 32024
rect 77204 31984 77205 32024
rect 77163 31975 77205 31984
rect 76971 31520 77013 31529
rect 76971 31480 76972 31520
rect 77012 31480 77013 31520
rect 76971 31471 77013 31480
rect 76972 31352 77012 31361
rect 76876 31312 76972 31352
rect 76876 30890 76916 31312
rect 76972 31303 77012 31312
rect 77164 31352 77204 31975
rect 77356 31520 77396 33487
rect 77836 33140 77876 33496
rect 77548 33100 77876 33140
rect 77452 32864 77492 32873
rect 77452 32369 77492 32824
rect 77451 32360 77493 32369
rect 77451 32320 77452 32360
rect 77492 32320 77493 32360
rect 77451 32311 77493 32320
rect 77452 32192 77492 32201
rect 77548 32192 77588 33100
rect 77739 33032 77781 33041
rect 77739 32992 77740 33032
rect 77780 32992 77876 33032
rect 77739 32983 77781 32992
rect 77740 32864 77780 32873
rect 77740 32705 77780 32824
rect 77836 32864 77876 32992
rect 77836 32815 77876 32824
rect 77739 32696 77781 32705
rect 77739 32656 77740 32696
rect 77780 32656 77781 32696
rect 77739 32647 77781 32656
rect 77492 32152 77588 32192
rect 77452 32143 77492 32152
rect 77932 31604 77972 33664
rect 78124 33545 78164 34327
rect 78123 33536 78165 33545
rect 78123 33496 78124 33536
rect 78164 33496 78165 33536
rect 78123 33487 78165 33496
rect 78316 33140 78356 35176
rect 79468 34964 79508 34973
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 79468 34385 79508 34924
rect 79467 34376 79509 34385
rect 79467 34336 79468 34376
rect 79508 34336 79509 34376
rect 79467 34327 79509 34336
rect 78411 33704 78453 33713
rect 78411 33664 78412 33704
rect 78452 33664 78453 33704
rect 78411 33655 78453 33664
rect 78220 33100 78356 33140
rect 78412 33116 78452 33655
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 78123 33032 78165 33041
rect 78123 32992 78124 33032
rect 78164 32992 78165 33032
rect 78123 32983 78165 32992
rect 78124 32898 78164 32983
rect 78220 32873 78260 33100
rect 78412 33067 78452 33076
rect 78507 33032 78549 33041
rect 78507 32992 78508 33032
rect 78548 32992 78549 33032
rect 78507 32983 78549 32992
rect 78219 32864 78261 32873
rect 78219 32824 78220 32864
rect 78260 32824 78261 32864
rect 78219 32815 78261 32824
rect 78316 32864 78356 32873
rect 78508 32864 78548 32983
rect 78356 32824 78452 32864
rect 78316 32815 78356 32824
rect 78027 32696 78069 32705
rect 78027 32656 78028 32696
rect 78068 32656 78069 32696
rect 78027 32647 78069 32656
rect 78028 31949 78068 32647
rect 78220 32192 78260 32815
rect 78316 32192 78356 32201
rect 78220 32152 78316 32192
rect 78027 31940 78069 31949
rect 78027 31900 78028 31940
rect 78068 31900 78069 31940
rect 78027 31891 78069 31900
rect 77932 31555 77972 31564
rect 77356 31480 77780 31520
rect 77164 31303 77204 31312
rect 77451 31352 77493 31361
rect 77451 31312 77452 31352
rect 77492 31312 77493 31352
rect 77451 31303 77493 31312
rect 77644 31352 77684 31361
rect 77068 31268 77108 31277
rect 77068 30941 77108 31228
rect 77452 31025 77492 31303
rect 77548 31268 77588 31277
rect 77451 31016 77493 31025
rect 77451 30976 77452 31016
rect 77492 30976 77493 31016
rect 77451 30967 77493 30976
rect 77067 30932 77109 30941
rect 77067 30892 77068 30932
rect 77108 30892 77300 30932
rect 77067 30883 77109 30892
rect 76876 30841 76916 30850
rect 77068 30680 77108 30689
rect 76971 30260 77013 30269
rect 76971 30220 76972 30260
rect 77012 30220 77013 30260
rect 76971 30211 77013 30220
rect 76972 29840 77012 30211
rect 77068 30092 77108 30640
rect 77163 30680 77205 30689
rect 77163 30640 77164 30680
rect 77204 30640 77205 30680
rect 77163 30631 77205 30640
rect 77068 30043 77108 30052
rect 77068 29840 77108 29849
rect 76972 29800 77068 29840
rect 76780 29128 76916 29168
rect 76780 29000 76820 29009
rect 76684 28960 76780 29000
rect 76780 28951 76820 28960
rect 76683 28664 76725 28673
rect 76683 28624 76684 28664
rect 76724 28624 76725 28664
rect 76683 28615 76725 28624
rect 76684 28580 76724 28615
rect 76684 28529 76724 28540
rect 76876 28496 76916 29128
rect 76780 28456 76916 28496
rect 76972 28496 77012 29800
rect 77068 29791 77108 29800
rect 77164 29765 77204 30631
rect 77260 29840 77300 30892
rect 77548 30848 77588 31228
rect 77644 31109 77684 31312
rect 77643 31100 77685 31109
rect 77643 31060 77644 31100
rect 77684 31060 77685 31100
rect 77643 31051 77685 31060
rect 77644 30857 77684 31051
rect 77260 29791 77300 29800
rect 77356 30808 77588 30848
rect 77643 30848 77685 30857
rect 77643 30808 77644 30848
rect 77684 30808 77685 30848
rect 77356 29840 77396 30808
rect 77643 30799 77685 30808
rect 77452 30680 77492 30689
rect 77492 30640 77684 30680
rect 77452 30631 77492 30640
rect 77547 30512 77589 30521
rect 77547 30472 77548 30512
rect 77588 30472 77589 30512
rect 77547 30463 77589 30472
rect 77548 29840 77588 30463
rect 77644 30008 77684 30640
rect 77644 29959 77684 29968
rect 77548 29800 77684 29840
rect 77356 29791 77396 29800
rect 77163 29756 77205 29765
rect 77163 29716 77164 29756
rect 77204 29716 77205 29756
rect 77163 29707 77205 29716
rect 77068 29168 77108 29177
rect 77068 28673 77108 29128
rect 77067 28664 77109 28673
rect 77067 28624 77068 28664
rect 77108 28624 77109 28664
rect 77067 28615 77109 28624
rect 76972 28456 77108 28496
rect 76587 28328 76629 28337
rect 76587 28288 76588 28328
rect 76628 28288 76629 28328
rect 76587 28279 76629 28288
rect 76684 28328 76724 28337
rect 76684 28085 76724 28288
rect 76683 28076 76725 28085
rect 76683 28036 76684 28076
rect 76724 28036 76725 28076
rect 76683 28027 76725 28036
rect 76780 27824 76820 28456
rect 76875 28328 76917 28337
rect 76875 28288 76876 28328
rect 76916 28288 76917 28328
rect 76875 28279 76917 28288
rect 76972 28328 77012 28339
rect 76876 28194 76916 28279
rect 76972 28253 77012 28288
rect 76971 28244 77013 28253
rect 76971 28204 76972 28244
rect 77012 28204 77013 28244
rect 76971 28195 77013 28204
rect 77068 28085 77108 28456
rect 77164 28328 77204 29707
rect 77452 29168 77492 29177
rect 77452 28496 77492 29128
rect 77548 28496 77588 28505
rect 77452 28456 77548 28496
rect 77548 28447 77588 28456
rect 77164 28279 77204 28288
rect 77355 28328 77397 28337
rect 77355 28288 77356 28328
rect 77396 28288 77397 28328
rect 77355 28279 77397 28288
rect 77259 28244 77301 28253
rect 77259 28204 77260 28244
rect 77300 28204 77301 28244
rect 77259 28195 77301 28204
rect 77163 28160 77205 28169
rect 77163 28120 77164 28160
rect 77204 28120 77205 28160
rect 77163 28111 77205 28120
rect 77067 28076 77109 28085
rect 77067 28036 77068 28076
rect 77108 28036 77109 28076
rect 77067 28027 77109 28036
rect 76684 27784 76820 27824
rect 76492 26816 76532 26825
rect 76299 26732 76341 26741
rect 76299 26692 76300 26732
rect 76340 26692 76341 26732
rect 76299 26683 76341 26692
rect 76492 26657 76532 26776
rect 76587 26816 76629 26825
rect 76587 26776 76588 26816
rect 76628 26776 76629 26816
rect 76587 26767 76629 26776
rect 76588 26682 76628 26767
rect 76203 26648 76245 26657
rect 76203 26608 76204 26648
rect 76244 26608 76245 26648
rect 76203 26599 76245 26608
rect 76491 26648 76533 26657
rect 76491 26608 76492 26648
rect 76532 26608 76533 26648
rect 76491 26599 76533 26608
rect 76299 25556 76341 25565
rect 76299 25516 76300 25556
rect 76340 25516 76341 25556
rect 76684 25556 76724 27784
rect 76780 27656 76820 27665
rect 76780 26153 76820 27616
rect 76875 27656 76917 27665
rect 76875 27616 76876 27656
rect 76916 27616 76917 27656
rect 76875 27607 76917 27616
rect 76972 27656 77012 27665
rect 76876 27522 76916 27607
rect 76876 27068 76916 27077
rect 76972 27068 77012 27616
rect 77067 27656 77109 27665
rect 77067 27616 77068 27656
rect 77108 27616 77109 27656
rect 77067 27607 77109 27616
rect 77164 27656 77204 28111
rect 77260 28110 77300 28195
rect 77356 28194 77396 28279
rect 77164 27607 77204 27616
rect 77356 27656 77396 27665
rect 76916 27028 77012 27068
rect 76876 27019 76916 27028
rect 77068 26900 77108 27607
rect 77260 27404 77300 27413
rect 77068 26860 77204 26900
rect 77068 26732 77108 26741
rect 76972 26692 77068 26732
rect 76972 26312 77012 26692
rect 77068 26683 77108 26692
rect 77164 26312 77204 26860
rect 76972 26263 77012 26272
rect 77068 26272 77204 26312
rect 76779 26144 76821 26153
rect 76779 26104 76780 26144
rect 76820 26104 76821 26144
rect 76779 26095 76821 26104
rect 76876 26144 76916 26153
rect 76876 25976 76916 26104
rect 77068 26144 77108 26272
rect 77068 26095 77108 26104
rect 77164 26144 77204 26153
rect 77260 26144 77300 27364
rect 77356 26657 77396 27616
rect 77548 27488 77588 27497
rect 77452 27448 77548 27488
rect 77452 26816 77492 27448
rect 77548 27439 77588 27448
rect 77452 26767 77492 26776
rect 77355 26648 77397 26657
rect 77355 26608 77356 26648
rect 77396 26608 77397 26648
rect 77355 26599 77397 26608
rect 77204 26104 77300 26144
rect 77355 26144 77397 26153
rect 77355 26104 77356 26144
rect 77396 26104 77397 26144
rect 77164 26095 77204 26104
rect 77355 26095 77397 26104
rect 76876 25936 76926 25976
rect 76886 25892 76926 25936
rect 76876 25852 76926 25892
rect 76684 25516 76820 25556
rect 76299 25507 76341 25516
rect 76012 25432 76148 25472
rect 76005 25319 76045 25328
rect 75820 25255 75860 25264
rect 75916 25279 76005 25319
rect 75628 25136 75668 25145
rect 75668 25096 75860 25136
rect 75628 25087 75668 25096
rect 75820 24716 75860 25096
rect 75820 24667 75860 24676
rect 75436 24583 75476 24592
rect 75723 24632 75765 24641
rect 75723 24592 75724 24632
rect 75764 24592 75765 24632
rect 75723 24583 75765 24592
rect 75339 24548 75381 24557
rect 75339 24508 75340 24548
rect 75380 24508 75381 24548
rect 75339 24499 75381 24508
rect 75724 24498 75764 24583
rect 75916 24473 75956 25279
rect 76005 25270 76045 25279
rect 76108 25220 76148 25432
rect 76012 25180 76148 25220
rect 76204 25304 76244 25313
rect 75915 24464 75957 24473
rect 75915 24424 75916 24464
rect 75956 24424 75957 24464
rect 75915 24415 75957 24424
rect 75243 23876 75285 23885
rect 75243 23836 75244 23876
rect 75284 23836 75285 23876
rect 75243 23827 75285 23836
rect 75531 23876 75573 23885
rect 75531 23836 75532 23876
rect 75572 23836 75573 23876
rect 75531 23827 75573 23836
rect 74860 23633 74900 23752
rect 75051 23792 75093 23801
rect 75051 23752 75052 23792
rect 75092 23752 75093 23792
rect 75051 23743 75093 23752
rect 75244 23792 75284 23827
rect 75244 23741 75284 23752
rect 74859 23624 74901 23633
rect 74859 23584 74860 23624
rect 74900 23584 74901 23624
rect 74859 23575 74901 23584
rect 74956 23624 74996 23633
rect 74668 23164 74900 23204
rect 73612 23020 73695 23060
rect 73804 23020 73940 23060
rect 73996 23020 74095 23060
rect 74188 23020 74324 23060
rect 74380 23020 74495 23060
rect 74572 23020 74785 23060
rect 73516 22744 73585 22784
rect 73545 22596 73585 22744
rect 73655 22596 73695 23020
rect 73900 22784 73940 23020
rect 73900 22744 73985 22784
rect 73945 22596 73985 22744
rect 74055 22596 74095 23020
rect 74284 22784 74324 23020
rect 74284 22744 74385 22784
rect 74345 22596 74385 22744
rect 74455 22596 74495 23020
rect 74745 22596 74785 23020
rect 74860 22868 74900 23164
rect 74956 23060 74996 23584
rect 75243 23624 75285 23633
rect 75243 23584 75244 23624
rect 75284 23584 75285 23624
rect 75243 23575 75285 23584
rect 75340 23624 75380 23633
rect 75244 23060 75284 23575
rect 75340 23060 75380 23584
rect 75532 23204 75572 23827
rect 75628 23792 75668 23801
rect 76012 23792 76052 25180
rect 76204 24800 76244 25264
rect 76300 25304 76340 25507
rect 76492 25472 76532 25481
rect 76532 25432 76724 25472
rect 76492 25423 76532 25432
rect 76300 25255 76340 25264
rect 76492 25304 76532 25315
rect 76492 25229 76532 25264
rect 76684 25304 76724 25432
rect 76684 25255 76724 25264
rect 76491 25220 76533 25229
rect 76491 25180 76492 25220
rect 76532 25180 76533 25220
rect 76491 25171 76533 25180
rect 76204 24760 76532 24800
rect 76492 24716 76532 24760
rect 76492 24667 76532 24676
rect 76396 24632 76436 24643
rect 76396 24557 76436 24592
rect 76587 24632 76629 24641
rect 76587 24592 76588 24632
rect 76628 24592 76629 24632
rect 76587 24583 76629 24592
rect 76395 24548 76437 24557
rect 76395 24508 76396 24548
rect 76436 24508 76437 24548
rect 76395 24499 76437 24508
rect 76588 24498 76628 24583
rect 76107 24464 76149 24473
rect 76107 24424 76108 24464
rect 76148 24424 76149 24464
rect 76107 24415 76149 24424
rect 76108 24330 76148 24415
rect 75668 23752 76052 23792
rect 75628 23743 75668 23752
rect 75724 23624 75764 23633
rect 75764 23584 75956 23624
rect 75724 23575 75764 23584
rect 75532 23164 75668 23204
rect 75628 23060 75668 23164
rect 74956 23020 75185 23060
rect 75244 23020 75295 23060
rect 75340 23020 75585 23060
rect 75628 23020 75695 23060
rect 74855 22828 74900 22868
rect 74855 22596 74895 22828
rect 75145 22596 75185 23020
rect 75255 22596 75295 23020
rect 75545 22596 75585 23020
rect 75655 22596 75695 23020
rect 75916 22784 75956 23584
rect 76012 23060 76052 23752
rect 76107 23792 76149 23801
rect 76107 23752 76108 23792
rect 76148 23752 76149 23792
rect 76107 23743 76149 23752
rect 76491 23792 76533 23801
rect 76491 23752 76492 23792
rect 76532 23752 76533 23792
rect 76780 23792 76820 25516
rect 76876 25229 76916 25852
rect 77068 25304 77108 25313
rect 76875 25220 76917 25229
rect 76875 25180 76876 25220
rect 76916 25180 76917 25220
rect 76875 25171 76917 25180
rect 77068 24464 77108 25264
rect 77164 24464 77204 24473
rect 77068 24424 77164 24464
rect 77164 24415 77204 24424
rect 76972 23792 77012 23801
rect 76780 23752 76972 23792
rect 76491 23743 76533 23752
rect 76108 23658 76148 23743
rect 76204 23624 76244 23633
rect 76204 23060 76244 23584
rect 76492 23060 76532 23743
rect 76876 23624 76916 23633
rect 76780 23584 76876 23624
rect 76780 23060 76820 23584
rect 76876 23575 76916 23584
rect 76972 23060 77012 23752
rect 77260 23792 77300 23801
rect 77356 23792 77396 26095
rect 77300 23752 77396 23792
rect 77548 23792 77588 23801
rect 77644 23792 77684 29800
rect 77740 26153 77780 31480
rect 77835 31352 77877 31361
rect 77835 31312 77836 31352
rect 77876 31312 77877 31352
rect 77835 31303 77877 31312
rect 78028 31352 78068 31891
rect 77836 31218 77876 31303
rect 77835 30848 77877 30857
rect 77835 30808 77836 30848
rect 77876 30808 77877 30848
rect 77835 30799 77877 30808
rect 77739 26144 77781 26153
rect 77739 26104 77740 26144
rect 77780 26104 77781 26144
rect 77739 26095 77781 26104
rect 77836 25976 77876 30799
rect 78028 30521 78068 31312
rect 78316 30680 78356 32152
rect 78412 32033 78452 32824
rect 78508 32815 78548 32824
rect 78411 32024 78453 32033
rect 78411 31984 78412 32024
rect 78452 31984 78453 32024
rect 78411 31975 78453 31984
rect 79467 31940 79509 31949
rect 79467 31900 79468 31940
rect 79508 31900 79509 31940
rect 79467 31891 79509 31900
rect 79468 31806 79508 31891
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 79467 30848 79509 30857
rect 79467 30808 79468 30848
rect 79508 30808 79509 30848
rect 79467 30799 79509 30808
rect 79468 30714 79508 30799
rect 78027 30512 78069 30521
rect 78027 30472 78028 30512
rect 78068 30472 78069 30512
rect 78027 30463 78069 30472
rect 78316 29168 78356 30640
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 78316 29119 78356 29128
rect 79468 28916 79508 28925
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 79468 28337 79508 28876
rect 78123 28328 78165 28337
rect 78123 28288 78124 28328
rect 78164 28288 78165 28328
rect 78123 28279 78165 28288
rect 79467 28328 79509 28337
rect 79467 28288 79468 28328
rect 79508 28288 79509 28328
rect 79467 28279 79509 28288
rect 77588 23752 77684 23792
rect 77164 23624 77204 23633
rect 77164 23060 77204 23584
rect 77260 23060 77300 23752
rect 77548 23743 77588 23752
rect 76012 23020 76095 23060
rect 76204 23020 76385 23060
rect 75916 22744 75985 22784
rect 75945 22596 75985 22744
rect 76055 22596 76095 23020
rect 76345 22596 76385 23020
rect 76455 23020 76532 23060
rect 76745 23020 76820 23060
rect 76876 23020 77012 23060
rect 77145 23020 77204 23060
rect 77255 23020 77300 23060
rect 77452 23624 77492 23633
rect 77452 23060 77492 23584
rect 77644 23060 77684 23752
rect 77740 25936 77876 25976
rect 77740 23792 77780 25936
rect 77931 25304 77973 25313
rect 77931 25264 77932 25304
rect 77972 25264 77973 25304
rect 77931 25255 77973 25264
rect 77932 25170 77972 25255
rect 78124 23792 78164 28279
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 78316 26816 78356 26825
rect 78316 25313 78356 26776
rect 78507 26648 78549 26657
rect 78507 26608 78508 26648
rect 78548 26608 78549 26648
rect 78507 26599 78549 26608
rect 79467 26648 79509 26657
rect 79467 26608 79468 26648
rect 79508 26608 79509 26648
rect 79467 26599 79509 26608
rect 78315 25304 78357 25313
rect 78315 25264 78316 25304
rect 78356 25264 78357 25304
rect 78315 25255 78357 25264
rect 78508 23792 78548 26599
rect 79468 26514 79508 26599
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79084 25136 79124 25145
rect 78988 25096 79084 25136
rect 78988 24641 79028 25096
rect 79084 25087 79124 25096
rect 78987 24632 79029 24641
rect 78987 24592 78988 24632
rect 79028 24592 79029 24632
rect 78987 24583 79029 24592
rect 77780 23752 78068 23792
rect 77740 23743 77780 23752
rect 77836 23624 77876 23633
rect 77836 23060 77876 23584
rect 78028 23060 78068 23752
rect 78164 23752 78452 23792
rect 78124 23743 78164 23752
rect 78220 23624 78260 23633
rect 78220 23060 78260 23584
rect 77452 23020 77585 23060
rect 77644 23020 77695 23060
rect 77836 23020 77985 23060
rect 78028 23020 78095 23060
rect 78220 23020 78356 23060
rect 76455 22596 76495 23020
rect 76745 22596 76785 23020
rect 76876 22784 76916 23020
rect 76855 22744 76916 22784
rect 76855 22596 76895 22744
rect 77145 22596 77185 23020
rect 77255 22596 77295 23020
rect 77545 22596 77585 23020
rect 77655 22596 77695 23020
rect 77945 22596 77985 23020
rect 78055 22596 78095 23020
rect 78316 22784 78356 23020
rect 78412 22868 78452 23752
rect 78508 23060 78548 23752
rect 78796 23792 78836 23801
rect 78988 23792 79028 24583
rect 78836 23752 79028 23792
rect 79083 23792 79125 23801
rect 79083 23752 79084 23792
rect 79124 23752 79125 23792
rect 78604 23624 78644 23633
rect 78644 23584 78740 23624
rect 78604 23575 78644 23584
rect 78700 23060 78740 23584
rect 78796 23465 78836 23752
rect 79083 23743 79125 23752
rect 79372 23792 79412 23801
rect 79084 23658 79124 23743
rect 78892 23624 78932 23633
rect 78795 23456 78837 23465
rect 78795 23416 78796 23456
rect 78836 23416 78837 23456
rect 78795 23407 78837 23416
rect 78892 23060 78932 23584
rect 79180 23624 79220 23633
rect 79372 23624 79412 23752
rect 79220 23584 79412 23624
rect 79180 23575 79220 23584
rect 79275 23456 79317 23465
rect 79275 23416 79276 23456
rect 79316 23416 79317 23456
rect 79275 23407 79317 23416
rect 79276 23060 79316 23407
rect 78508 23020 78644 23060
rect 78700 23020 78785 23060
rect 78892 23020 79185 23060
rect 78412 22828 78495 22868
rect 78316 22744 78385 22784
rect 78345 22596 78385 22744
rect 78455 22596 78495 22828
rect 78604 22793 78644 23020
rect 78603 22784 78645 22793
rect 78603 22744 78604 22784
rect 78644 22744 78645 22784
rect 78603 22735 78645 22744
rect 78745 22596 78785 23020
rect 78854 22784 78896 22793
rect 78854 22744 78855 22784
rect 78895 22744 78896 22784
rect 78854 22735 78896 22744
rect 78855 22596 78895 22735
rect 79145 22596 79185 23020
rect 79255 23020 79316 23060
rect 79372 23060 79412 23584
rect 79468 23624 79508 23633
rect 79508 23584 79700 23624
rect 79468 23575 79508 23584
rect 79660 23060 79700 23584
rect 79372 23020 79585 23060
rect 79255 22596 79295 23020
rect 79545 22596 79585 23020
rect 79655 23020 79700 23060
rect 79655 22596 79695 23020
rect 60457 22269 60500 22280
rect 60455 22240 60500 22269
rect 60455 22229 60497 22240
rect 60455 22176 60495 22229
rect 53067 17660 53109 17669
rect 53067 17620 53068 17660
rect 53108 17620 53109 17660
rect 53067 17611 53109 17620
rect 53545 17333 53585 17472
rect 53544 17324 53586 17333
rect 53544 17284 53545 17324
rect 53585 17284 53586 17324
rect 53544 17275 53586 17284
rect 53655 17249 53695 17472
rect 53945 17249 53985 17472
rect 53654 17240 53696 17249
rect 53654 17200 53655 17240
rect 53695 17200 53696 17240
rect 53654 17191 53696 17200
rect 53944 17240 53986 17249
rect 53944 17200 53945 17240
rect 53985 17200 53986 17240
rect 53944 17191 53986 17200
rect 52875 17156 52917 17165
rect 52875 17116 52876 17156
rect 52916 17116 52917 17156
rect 52875 17107 52917 17116
rect 54055 17072 54095 17472
rect 54345 17165 54385 17472
rect 54455 17165 54495 17472
rect 54344 17156 54386 17165
rect 54344 17116 54345 17156
rect 54385 17116 54386 17156
rect 54344 17107 54386 17116
rect 54454 17156 54496 17165
rect 54745 17156 54785 17472
rect 54454 17116 54455 17156
rect 54495 17116 54496 17156
rect 54454 17107 54496 17116
rect 54700 17116 54785 17156
rect 52588 17021 52628 17032
rect 54028 17032 54095 17072
rect 52491 16988 52533 16997
rect 52491 16948 52492 16988
rect 52532 16948 52533 16988
rect 52491 16939 52533 16948
rect 54028 16829 54068 17032
rect 52395 16820 52437 16829
rect 52395 16780 52396 16820
rect 52436 16780 52437 16820
rect 52395 16771 52437 16780
rect 54027 16820 54069 16829
rect 54027 16780 54028 16820
rect 54068 16780 54069 16820
rect 54027 16771 54069 16780
rect 52396 16686 52436 16771
rect 53067 16736 53109 16745
rect 53067 16696 53068 16736
rect 53108 16696 53109 16736
rect 53067 16687 53109 16696
rect 52491 16652 52533 16661
rect 52491 16612 52492 16652
rect 52532 16612 52533 16652
rect 52491 16603 52533 16612
rect 52108 16400 52148 16409
rect 52148 16360 52340 16400
rect 52108 16351 52148 16360
rect 52012 16207 52148 16247
rect 52011 15392 52053 15401
rect 52011 15352 52012 15392
rect 52052 15352 52053 15392
rect 52011 15343 52053 15352
rect 52012 14720 52052 15343
rect 52012 14671 52052 14680
rect 51916 14512 52052 14552
rect 52012 13712 52052 14512
rect 52108 13889 52148 16207
rect 52300 14048 52340 16360
rect 52395 16232 52437 16241
rect 52395 16192 52396 16232
rect 52436 16192 52437 16232
rect 52395 16183 52437 16192
rect 52492 16232 52532 16603
rect 52779 16568 52821 16577
rect 52779 16528 52780 16568
rect 52820 16528 52821 16568
rect 52779 16519 52821 16528
rect 52780 16325 52820 16519
rect 52779 16316 52821 16325
rect 52779 16276 52780 16316
rect 52820 16276 52821 16316
rect 52779 16267 52821 16276
rect 52492 16183 52532 16192
rect 52780 16232 52820 16267
rect 53068 16241 53108 16687
rect 53739 16652 53781 16661
rect 53739 16612 53740 16652
rect 53780 16612 53781 16652
rect 53739 16603 53781 16612
rect 53740 16409 53780 16603
rect 53644 16400 53684 16409
rect 53356 16360 53644 16400
rect 52396 14981 52436 16183
rect 52780 16181 52820 16192
rect 53067 16232 53109 16241
rect 53067 16183 53068 16232
rect 53108 16183 53109 16232
rect 53356 16232 53396 16360
rect 53644 16351 53684 16360
rect 53739 16400 53781 16409
rect 53739 16360 53740 16400
rect 53780 16360 53781 16400
rect 53739 16351 53781 16360
rect 53932 16400 53972 16409
rect 54316 16400 54356 16409
rect 53260 16190 53300 16199
rect 53068 16169 53108 16178
rect 53356 16183 53396 16192
rect 53548 16232 53588 16241
rect 53164 16064 53204 16073
rect 53068 15644 53108 15653
rect 53164 15644 53204 16024
rect 53108 15604 53204 15644
rect 53068 15595 53108 15604
rect 52683 15560 52725 15569
rect 53260 15560 53300 16150
rect 53548 16064 53588 16192
rect 53740 16232 53780 16351
rect 53740 16183 53780 16192
rect 52683 15520 52684 15560
rect 52724 15520 52725 15560
rect 52683 15511 52725 15520
rect 53164 15520 53300 15560
rect 53356 16024 53588 16064
rect 52684 15426 52724 15511
rect 53164 15392 53204 15520
rect 53068 15352 53204 15392
rect 52395 14972 52437 14981
rect 52395 14932 52396 14972
rect 52436 14932 52437 14972
rect 52395 14923 52437 14932
rect 52683 14300 52725 14309
rect 52683 14260 52684 14300
rect 52724 14260 52725 14300
rect 52683 14251 52725 14260
rect 52587 14216 52629 14225
rect 52587 14176 52588 14216
rect 52628 14176 52629 14216
rect 52587 14167 52629 14176
rect 52588 14132 52628 14167
rect 52588 14081 52628 14092
rect 52684 14057 52724 14251
rect 53068 14225 53108 15352
rect 53163 14972 53205 14981
rect 53163 14932 53164 14972
rect 53204 14932 53205 14972
rect 53163 14923 53205 14932
rect 53164 14838 53204 14923
rect 53164 14552 53204 14561
rect 53164 14468 53204 14512
rect 53164 14428 53290 14468
rect 53067 14216 53109 14225
rect 53067 14176 53068 14216
rect 53108 14176 53109 14216
rect 53067 14167 53109 14176
rect 53250 14063 53290 14428
rect 52492 14048 52532 14057
rect 52300 14008 52492 14048
rect 52492 13999 52532 14008
rect 52683 14048 52725 14057
rect 52683 14008 52684 14048
rect 52724 14008 52725 14048
rect 53250 14014 53290 14023
rect 53356 14048 53396 16024
rect 53932 15980 53972 16360
rect 54220 16360 54316 16400
rect 54027 16232 54069 16241
rect 54027 16192 54028 16232
rect 54068 16192 54069 16232
rect 54027 16183 54069 16192
rect 53452 15940 53972 15980
rect 53452 15560 53492 15940
rect 53643 15728 53685 15737
rect 53643 15688 53644 15728
rect 53684 15688 53685 15728
rect 53643 15679 53685 15688
rect 53452 15511 53492 15520
rect 53452 14720 53492 14729
rect 53644 14720 53684 15679
rect 54028 14813 54068 16183
rect 54027 14804 54069 14813
rect 54027 14764 54028 14804
rect 54068 14764 54069 14804
rect 54027 14755 54069 14764
rect 53492 14680 53684 14720
rect 53452 14671 53492 14680
rect 53643 14552 53685 14561
rect 53643 14512 53644 14552
rect 53684 14512 53685 14552
rect 53643 14503 53685 14512
rect 53451 14132 53493 14141
rect 53451 14092 53452 14132
rect 53492 14092 53493 14132
rect 53451 14083 53493 14092
rect 52683 13999 52725 14008
rect 52684 13914 52724 13999
rect 53356 13973 53396 14008
rect 53355 13964 53397 13973
rect 53355 13924 53356 13964
rect 53396 13924 53397 13964
rect 53355 13915 53397 13924
rect 53452 13964 53492 14083
rect 53548 14048 53588 14057
rect 53548 13964 53588 14008
rect 53452 13924 53588 13964
rect 52107 13880 52149 13889
rect 52107 13840 52108 13880
rect 52148 13840 52149 13880
rect 52107 13831 52149 13840
rect 52012 13672 52244 13712
rect 51915 13628 51957 13637
rect 51915 13588 51916 13628
rect 51956 13588 51957 13628
rect 51915 13579 51957 13588
rect 51916 13208 51956 13579
rect 52107 13292 52149 13301
rect 52107 13252 52108 13292
rect 52148 13252 52149 13292
rect 52107 13243 52149 13252
rect 51916 12965 51956 13168
rect 52108 13208 52148 13243
rect 52108 13157 52148 13168
rect 52012 13124 52052 13133
rect 52012 12980 52052 13084
rect 51915 12956 51957 12965
rect 51915 12916 51916 12956
rect 51956 12916 51957 12956
rect 52012 12940 52148 12980
rect 51915 12907 51957 12916
rect 51668 12412 51860 12452
rect 52012 12536 52052 12545
rect 51628 12403 51668 12412
rect 51820 12284 51860 12293
rect 50859 11864 50901 11873
rect 50956 11864 50996 12244
rect 50859 11824 50860 11864
rect 50900 11824 50996 11864
rect 51148 12244 51284 12284
rect 51628 12244 51820 12284
rect 50859 11815 50901 11824
rect 50860 11696 50900 11815
rect 50860 11647 50900 11656
rect 51148 11696 51188 12244
rect 51532 11864 51572 11873
rect 51532 11705 51572 11824
rect 51628 11780 51668 12244
rect 51820 12235 51860 12244
rect 51724 11948 51764 11957
rect 52012 11948 52052 12496
rect 51764 11908 52052 11948
rect 51724 11899 51764 11908
rect 51723 11780 51765 11789
rect 51628 11740 51724 11780
rect 51764 11740 51765 11780
rect 51723 11731 51765 11740
rect 51148 11647 51188 11656
rect 51531 11696 51573 11705
rect 51531 11656 51532 11696
rect 51572 11656 51573 11696
rect 51531 11647 51573 11656
rect 51724 11696 51764 11731
rect 51724 11645 51764 11656
rect 51916 11696 51956 11707
rect 51916 11621 51956 11656
rect 52012 11696 52052 11705
rect 52108 11696 52148 12940
rect 52204 12116 52244 13672
rect 52492 13376 52532 13385
rect 53356 13376 53396 13915
rect 52492 12980 52532 13336
rect 53269 13336 53396 13376
rect 53269 13301 53309 13336
rect 53259 13292 53309 13301
rect 53259 13252 53260 13292
rect 53300 13252 53309 13292
rect 53259 13243 53301 13252
rect 53260 13137 53300 13243
rect 53355 13208 53397 13217
rect 53355 13168 53356 13208
rect 53396 13168 53397 13208
rect 53355 13159 53397 13168
rect 52396 12940 52532 12980
rect 52396 12536 52436 12940
rect 53356 12620 53396 13159
rect 53452 13133 53492 13924
rect 53548 13796 53588 13805
rect 53548 13217 53588 13756
rect 53644 13385 53684 14503
rect 53740 14048 53780 14057
rect 53740 13880 53780 14008
rect 54124 14048 54164 14057
rect 54220 14048 54260 16360
rect 54316 16351 54356 16360
rect 54700 16241 54740 17116
rect 54855 17072 54895 17472
rect 55145 17249 55185 17472
rect 54987 17240 55029 17249
rect 54987 17200 54988 17240
rect 55028 17200 55029 17240
rect 54987 17191 55029 17200
rect 55144 17240 55186 17249
rect 55144 17200 55145 17240
rect 55185 17200 55186 17240
rect 55144 17191 55186 17200
rect 54796 17032 54895 17072
rect 54796 16484 54836 17032
rect 54796 16435 54836 16444
rect 54699 16232 54741 16241
rect 54699 16192 54700 16232
rect 54740 16192 54741 16232
rect 54699 16183 54741 16192
rect 54988 16232 55028 17191
rect 55255 17072 55295 17472
rect 55545 17249 55585 17472
rect 55544 17240 55586 17249
rect 55544 17200 55545 17240
rect 55585 17200 55586 17240
rect 55544 17191 55586 17200
rect 55655 17072 55695 17472
rect 55945 17249 55985 17472
rect 55944 17240 55986 17249
rect 55944 17200 55945 17240
rect 55985 17200 55986 17240
rect 55944 17191 55986 17200
rect 56055 17072 56095 17472
rect 56345 17156 56385 17472
rect 55084 17032 55295 17072
rect 55372 17032 55695 17072
rect 55756 17032 56095 17072
rect 56332 17116 56385 17156
rect 55084 16484 55124 17032
rect 55084 16435 55124 16444
rect 55372 16484 55412 17032
rect 55372 16435 55412 16444
rect 55563 16484 55605 16493
rect 55563 16444 55564 16484
rect 55604 16444 55605 16484
rect 55563 16435 55605 16444
rect 55756 16484 55796 17032
rect 55756 16435 55796 16444
rect 55467 16400 55509 16409
rect 55467 16360 55468 16400
rect 55508 16360 55509 16400
rect 55467 16351 55509 16360
rect 55083 16316 55125 16325
rect 55083 16276 55084 16316
rect 55124 16276 55125 16316
rect 55083 16267 55125 16276
rect 54988 16183 55028 16192
rect 54700 16098 54740 16183
rect 54315 15560 54357 15569
rect 54315 15520 54316 15560
rect 54356 15520 54357 15560
rect 54315 15511 54357 15520
rect 54987 15560 55029 15569
rect 54987 15520 54988 15560
rect 55028 15520 55029 15560
rect 54987 15511 55029 15520
rect 54316 15426 54356 15511
rect 54699 14720 54741 14729
rect 54892 14720 54932 14729
rect 54699 14680 54700 14720
rect 54740 14680 54892 14720
rect 54699 14671 54741 14680
rect 54892 14671 54932 14680
rect 54164 14008 54260 14048
rect 54124 13999 54164 14008
rect 53740 13840 54644 13880
rect 54507 13712 54549 13721
rect 54507 13672 54508 13712
rect 54548 13672 54549 13712
rect 54507 13663 54549 13672
rect 54315 13628 54357 13637
rect 54315 13588 54316 13628
rect 54356 13588 54357 13628
rect 54315 13579 54357 13588
rect 54316 13385 54356 13579
rect 53643 13376 53685 13385
rect 53643 13336 53644 13376
rect 53684 13336 53685 13376
rect 53643 13327 53685 13336
rect 54315 13376 54357 13385
rect 54315 13336 54316 13376
rect 54356 13336 54357 13376
rect 54315 13327 54357 13336
rect 53547 13208 53589 13217
rect 53547 13168 53548 13208
rect 53588 13168 53589 13208
rect 53547 13159 53589 13168
rect 53451 13124 53493 13133
rect 53451 13084 53452 13124
rect 53492 13084 53493 13124
rect 53451 13075 53493 13084
rect 54316 12704 54356 13327
rect 54411 13208 54453 13217
rect 54411 13168 54412 13208
rect 54452 13168 54453 13208
rect 54411 13159 54453 13168
rect 54508 13208 54548 13663
rect 54508 13159 54548 13168
rect 54412 13074 54452 13159
rect 54604 13124 54644 13840
rect 54700 13460 54740 14671
rect 54988 14477 55028 15511
rect 54987 14468 55029 14477
rect 54987 14428 54988 14468
rect 55028 14428 55029 14468
rect 54987 14419 55029 14428
rect 54988 14048 55028 14419
rect 54988 13999 55028 14008
rect 55084 13964 55124 16267
rect 55275 16232 55317 16241
rect 55275 16192 55276 16232
rect 55316 16192 55317 16232
rect 55275 16183 55317 16192
rect 55276 16098 55316 16183
rect 55179 16064 55221 16073
rect 55179 16024 55180 16064
rect 55220 16024 55221 16064
rect 55179 16015 55221 16024
rect 55180 14048 55220 16015
rect 55468 15728 55508 16351
rect 55564 15905 55604 16435
rect 55659 16232 55701 16241
rect 56044 16232 56084 16241
rect 56332 16232 56372 17116
rect 56455 17072 56495 17472
rect 56745 17156 56785 17472
rect 55659 16192 55660 16232
rect 55700 16192 55701 16232
rect 55659 16183 55701 16192
rect 55852 16192 56044 16232
rect 56084 16192 56372 16232
rect 56428 17032 56495 17072
rect 56620 17116 56785 17156
rect 55660 16098 55700 16183
rect 55755 16064 55797 16073
rect 55755 16024 55756 16064
rect 55796 16024 55797 16064
rect 55755 16015 55797 16024
rect 55563 15896 55605 15905
rect 55563 15856 55564 15896
rect 55604 15856 55605 15896
rect 55563 15847 55605 15856
rect 55468 15679 55508 15688
rect 55180 14008 55316 14048
rect 55084 13924 55220 13964
rect 54700 13420 54836 13460
rect 54700 13217 54740 13302
rect 54699 13208 54741 13217
rect 54699 13168 54700 13208
rect 54740 13168 54741 13208
rect 54699 13159 54741 13168
rect 54604 13075 54644 13084
rect 54796 13040 54836 13420
rect 55180 13301 55220 13924
rect 55179 13292 55221 13301
rect 55179 13252 55180 13292
rect 55220 13252 55221 13292
rect 55179 13243 55221 13252
rect 55083 13208 55125 13217
rect 55083 13168 55084 13208
rect 55124 13168 55125 13208
rect 55083 13159 55125 13168
rect 55180 13208 55220 13243
rect 55084 13074 55124 13159
rect 55180 13158 55220 13168
rect 55276 13208 55316 14008
rect 55756 13469 55796 16015
rect 55852 13805 55892 16192
rect 56044 16183 56084 16192
rect 56140 16064 56180 16073
rect 56428 16064 56468 17032
rect 56620 16988 56660 17116
rect 56855 17072 56895 17472
rect 57145 17156 57185 17472
rect 56524 16948 56660 16988
rect 56812 17032 56895 17072
rect 57100 17116 57185 17156
rect 56524 16232 56564 16948
rect 56812 16736 56852 17032
rect 56620 16696 56852 16736
rect 56620 16484 56660 16696
rect 56620 16435 56660 16444
rect 56908 16232 56948 16241
rect 57100 16232 57140 17116
rect 57255 17072 57295 17472
rect 57545 17324 57585 17472
rect 56524 16157 56564 16192
rect 56812 16192 56908 16232
rect 56948 16192 57140 16232
rect 57196 17032 57295 17072
rect 57388 17284 57585 17324
rect 57655 17324 57695 17472
rect 57655 17284 57716 17324
rect 56523 16148 56565 16157
rect 56523 16108 56524 16148
rect 56564 16108 56565 16148
rect 56523 16099 56565 16108
rect 56524 16097 56564 16099
rect 56180 16024 56468 16064
rect 56140 16015 56180 16024
rect 56043 15896 56085 15905
rect 56043 15856 56044 15896
rect 56084 15856 56085 15896
rect 56043 15847 56085 15856
rect 56044 14720 56084 15847
rect 56716 14888 56756 14897
rect 56620 14848 56716 14888
rect 56044 14671 56084 14680
rect 56331 14720 56373 14729
rect 56331 14680 56332 14720
rect 56372 14680 56373 14720
rect 56331 14671 56373 14680
rect 56332 14586 56372 14671
rect 56428 14636 56468 14645
rect 55947 14468 55989 14477
rect 55947 14428 55948 14468
rect 55988 14428 55989 14468
rect 55947 14419 55989 14428
rect 55851 13796 55893 13805
rect 55851 13756 55852 13796
rect 55892 13756 55893 13796
rect 55851 13747 55893 13756
rect 55755 13460 55797 13469
rect 55755 13420 55756 13460
rect 55796 13420 55797 13460
rect 55755 13411 55797 13420
rect 55276 13049 55316 13168
rect 55371 13208 55413 13217
rect 55371 13168 55372 13208
rect 55412 13168 55413 13208
rect 55371 13159 55413 13168
rect 55372 13074 55412 13159
rect 54700 13000 54836 13040
rect 55275 13040 55317 13049
rect 55275 13000 55276 13040
rect 55316 13000 55317 13040
rect 54700 12980 54740 13000
rect 55275 12991 55317 13000
rect 54604 12940 54740 12980
rect 55948 12980 55988 14419
rect 56428 14300 56468 14596
rect 56140 14260 56468 14300
rect 56140 14216 56180 14260
rect 56140 14167 56180 14176
rect 56427 14132 56469 14141
rect 56427 14092 56428 14132
rect 56468 14092 56469 14132
rect 56427 14083 56469 14092
rect 56428 14048 56468 14083
rect 56235 13964 56277 13973
rect 56235 13924 56236 13964
rect 56276 13924 56277 13964
rect 56235 13915 56277 13924
rect 56140 13796 56180 13805
rect 56044 13756 56140 13796
rect 56044 13217 56084 13756
rect 56140 13747 56180 13756
rect 56043 13208 56085 13217
rect 56043 13168 56044 13208
rect 56084 13168 56085 13208
rect 56043 13159 56085 13168
rect 56140 13208 56180 13217
rect 56236 13208 56276 13915
rect 56428 13637 56468 14008
rect 56620 14048 56660 14848
rect 56716 14839 56756 14848
rect 56620 13999 56660 14008
rect 56523 13796 56565 13805
rect 56523 13756 56524 13796
rect 56564 13756 56565 13796
rect 56523 13747 56565 13756
rect 56524 13662 56564 13747
rect 56427 13628 56469 13637
rect 56427 13588 56428 13628
rect 56468 13588 56469 13628
rect 56427 13579 56469 13588
rect 56812 13553 56852 16192
rect 56908 16183 56948 16192
rect 57004 16064 57044 16073
rect 57196 16064 57236 17032
rect 57388 16988 57428 17284
rect 57044 16024 57236 16064
rect 57292 16948 57428 16988
rect 57292 16232 57332 16948
rect 57676 16736 57716 17284
rect 57945 17165 57985 17472
rect 57944 17156 57986 17165
rect 57944 17116 57945 17156
rect 57985 17116 58004 17156
rect 57944 17107 58004 17116
rect 57388 16696 57716 16736
rect 57388 16484 57428 16696
rect 57388 16435 57428 16444
rect 57580 16400 57620 16409
rect 57004 16015 57044 16024
rect 57292 15989 57332 16192
rect 57484 16360 57580 16400
rect 57291 15980 57333 15989
rect 57291 15940 57292 15980
rect 57332 15940 57333 15980
rect 57291 15931 57333 15940
rect 57100 15560 57140 15569
rect 56908 15520 57100 15560
rect 56908 14972 56948 15520
rect 57100 15511 57140 15520
rect 57484 15560 57524 16360
rect 57580 16351 57620 16360
rect 57964 16232 58004 17107
rect 58055 17072 58095 17472
rect 58345 17249 58385 17472
rect 58344 17240 58386 17249
rect 58344 17200 58345 17240
rect 58385 17200 58386 17240
rect 58344 17191 58386 17200
rect 58455 17072 58495 17472
rect 58745 17156 58785 17472
rect 58055 17032 58100 17072
rect 58060 16484 58100 17032
rect 58060 16435 58100 16444
rect 58348 17032 58495 17072
rect 58540 17116 58785 17156
rect 58348 16484 58388 17032
rect 58348 16435 58388 16444
rect 58540 16241 58580 17116
rect 58855 17072 58895 17472
rect 59145 17156 59185 17472
rect 58636 17032 58895 17072
rect 59116 17116 59185 17156
rect 58636 16484 58676 17032
rect 59116 16988 59156 17116
rect 59255 17072 59295 17472
rect 59545 17156 59585 17472
rect 58636 16435 58676 16444
rect 58924 16948 59156 16988
rect 59212 17032 59295 17072
rect 59500 17116 59585 17156
rect 57964 16183 58004 16192
rect 58251 16232 58293 16241
rect 58251 16192 58252 16232
rect 58292 16192 58293 16232
rect 58251 16183 58293 16192
rect 58539 16232 58581 16241
rect 58539 16192 58540 16232
rect 58580 16192 58581 16232
rect 58539 16183 58581 16192
rect 58924 16232 58964 16948
rect 59212 16736 59252 17032
rect 59020 16696 59252 16736
rect 59020 16484 59060 16696
rect 59020 16435 59060 16444
rect 59308 16232 59348 16241
rect 59500 16232 59540 17116
rect 59655 17072 59695 17472
rect 59945 17156 59985 17472
rect 58252 16098 58292 16183
rect 58540 16098 58580 16183
rect 57867 15896 57909 15905
rect 57867 15856 57868 15896
rect 57908 15856 57909 15896
rect 57867 15847 57909 15856
rect 57484 15511 57524 15520
rect 56908 14923 56948 14932
rect 57484 14888 57524 14897
rect 57196 14848 57484 14888
rect 56908 14813 56948 14844
rect 56907 14804 56949 14813
rect 56907 14764 56908 14804
rect 56948 14764 56949 14804
rect 56907 14755 56949 14764
rect 56908 14720 56948 14755
rect 56908 13721 56948 14680
rect 57100 14720 57140 14729
rect 57100 13805 57140 14680
rect 57196 14720 57236 14848
rect 57484 14839 57524 14848
rect 57196 14671 57236 14680
rect 57388 14720 57428 14729
rect 57388 13973 57428 14680
rect 57579 14720 57621 14729
rect 57579 14680 57580 14720
rect 57620 14680 57621 14720
rect 57579 14671 57621 14680
rect 57580 14586 57620 14671
rect 57675 14468 57717 14477
rect 57675 14428 57676 14468
rect 57716 14428 57717 14468
rect 57675 14419 57717 14428
rect 57387 13964 57429 13973
rect 57387 13924 57388 13964
rect 57428 13924 57429 13964
rect 57387 13915 57429 13924
rect 57099 13796 57141 13805
rect 57099 13756 57100 13796
rect 57140 13756 57141 13796
rect 57099 13747 57141 13756
rect 56907 13712 56949 13721
rect 56907 13672 56908 13712
rect 56948 13672 56949 13712
rect 56907 13663 56949 13672
rect 56811 13544 56853 13553
rect 56811 13504 56812 13544
rect 56852 13504 56853 13544
rect 56811 13495 56853 13504
rect 56332 13376 56372 13385
rect 56372 13336 56756 13376
rect 56332 13327 56372 13336
rect 56716 13292 56756 13336
rect 56716 13252 56852 13292
rect 56180 13168 56276 13208
rect 56332 13208 56372 13219
rect 56140 13159 56180 13168
rect 56044 13074 56084 13159
rect 56332 13133 56372 13168
rect 56427 13208 56469 13217
rect 56427 13168 56428 13208
rect 56468 13168 56469 13208
rect 56427 13159 56469 13168
rect 56524 13208 56564 13217
rect 56331 13124 56373 13133
rect 56331 13084 56332 13124
rect 56372 13084 56373 13124
rect 56331 13075 56373 13084
rect 55948 12940 56084 12980
rect 54412 12704 54452 12713
rect 54316 12664 54412 12704
rect 54412 12655 54452 12664
rect 52396 12487 52436 12496
rect 53293 12580 53396 12620
rect 53293 12536 53333 12580
rect 53293 12293 53333 12496
rect 53292 12284 53334 12293
rect 53292 12244 53293 12284
rect 53333 12244 53334 12284
rect 53292 12235 53334 12244
rect 52204 12076 52436 12116
rect 52396 11705 52436 12076
rect 52587 11864 52629 11873
rect 52587 11824 52588 11864
rect 52628 11824 52629 11864
rect 52587 11815 52629 11824
rect 52052 11656 52148 11696
rect 52203 11696 52245 11705
rect 52203 11656 52204 11696
rect 52244 11656 52245 11696
rect 52012 11647 52052 11656
rect 52203 11647 52245 11656
rect 52395 11696 52437 11705
rect 52395 11656 52396 11696
rect 52436 11656 52437 11696
rect 52395 11647 52437 11656
rect 50763 11612 50805 11621
rect 50763 11572 50764 11612
rect 50804 11572 50805 11612
rect 50763 11563 50805 11572
rect 51243 11612 51285 11621
rect 51243 11572 51244 11612
rect 51284 11572 51285 11612
rect 51243 11563 51285 11572
rect 51435 11612 51477 11621
rect 51435 11572 51436 11612
rect 51476 11572 51477 11612
rect 51435 11563 51477 11572
rect 51915 11612 51957 11621
rect 51915 11572 51916 11612
rect 51956 11572 51957 11612
rect 51915 11563 51957 11572
rect 50572 11024 50612 11033
rect 50572 10856 50612 10984
rect 50667 11024 50709 11033
rect 50667 10984 50668 11024
rect 50708 10984 50709 11024
rect 50667 10975 50709 10984
rect 50764 11024 50804 11563
rect 51244 11478 51284 11563
rect 50955 11192 50997 11201
rect 50955 11152 50956 11192
rect 50996 11152 50997 11192
rect 50955 11143 50997 11152
rect 50860 11033 50900 11118
rect 50764 10975 50804 10984
rect 50859 11024 50901 11033
rect 50859 10984 50860 11024
rect 50900 10984 50901 11024
rect 50859 10975 50901 10984
rect 50956 11024 50996 11143
rect 50956 10975 50996 10984
rect 51052 11024 51092 11033
rect 51244 11024 51284 11033
rect 51092 10984 51244 11024
rect 51052 10975 51092 10984
rect 51244 10975 51284 10984
rect 51436 11024 51476 11563
rect 52204 11562 52244 11647
rect 52299 11612 52341 11621
rect 52299 11572 52300 11612
rect 52340 11572 52341 11612
rect 52299 11563 52341 11572
rect 52300 11478 52340 11563
rect 52396 11562 52436 11647
rect 52107 11192 52149 11201
rect 52107 11152 52108 11192
rect 52148 11152 52149 11192
rect 52107 11143 52149 11152
rect 51436 10975 51476 10984
rect 51532 11024 51572 11033
rect 51244 10856 51284 10865
rect 50572 10816 51244 10856
rect 51244 10807 51284 10816
rect 51052 10184 51092 10193
rect 50283 9512 50325 9521
rect 50283 9472 50284 9512
rect 50324 9472 50325 9512
rect 50283 9463 50325 9472
rect 50380 9344 50420 9353
rect 50188 9304 50380 9344
rect 50380 9295 50420 9304
rect 50956 8840 50996 8849
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 50476 8000 50516 8009
rect 49612 7748 49652 7757
rect 49612 7169 49652 7708
rect 50476 7505 50516 7960
rect 50860 8000 50900 8009
rect 50956 8000 50996 8800
rect 50900 7960 50996 8000
rect 50860 7951 50900 7960
rect 50475 7496 50517 7505
rect 50475 7456 50476 7496
rect 50516 7456 50517 7496
rect 50475 7447 50517 7456
rect 51052 7169 51092 10144
rect 51532 9680 51572 10984
rect 51915 10940 51957 10949
rect 51915 10900 51916 10940
rect 51956 10900 51957 10940
rect 51915 10891 51957 10900
rect 51916 10806 51956 10891
rect 51724 10772 51764 10781
rect 51532 9631 51572 9640
rect 51628 10732 51724 10772
rect 51435 9512 51477 9521
rect 51435 9472 51436 9512
rect 51476 9472 51477 9512
rect 51435 9463 51477 9472
rect 51628 9512 51668 10732
rect 51724 10723 51764 10732
rect 52011 9680 52053 9689
rect 52011 9640 52012 9680
rect 52052 9640 52053 9680
rect 52011 9631 52053 9640
rect 51436 9378 51476 9463
rect 51628 9437 51668 9472
rect 51723 9512 51765 9521
rect 51723 9472 51724 9512
rect 51764 9472 51765 9512
rect 51723 9463 51765 9472
rect 51627 9428 51669 9437
rect 51627 9388 51628 9428
rect 51668 9388 51669 9428
rect 51627 9379 51669 9388
rect 51628 9348 51668 9379
rect 51724 9378 51764 9463
rect 51147 8168 51189 8177
rect 51147 8128 51148 8168
rect 51188 8128 51189 8168
rect 51147 8119 51189 8128
rect 51148 7412 51188 8119
rect 51148 7363 51188 7372
rect 51724 8000 51764 8009
rect 51724 7169 51764 7960
rect 51916 7328 51956 7337
rect 51820 7288 51916 7328
rect 49611 7160 49653 7169
rect 49611 7120 49612 7160
rect 49652 7120 49653 7160
rect 49611 7111 49653 7120
rect 49995 7160 50037 7169
rect 49995 7120 49996 7160
rect 50036 7120 50037 7160
rect 49995 7111 50037 7120
rect 50187 7160 50229 7169
rect 50187 7120 50188 7160
rect 50228 7120 50229 7160
rect 50187 7111 50229 7120
rect 50859 7160 50901 7169
rect 50859 7120 50860 7160
rect 50900 7120 50901 7160
rect 50859 7111 50901 7120
rect 51051 7160 51093 7169
rect 51051 7120 51052 7160
rect 51092 7120 51093 7160
rect 51051 7111 51093 7120
rect 51723 7160 51765 7169
rect 51723 7120 51724 7160
rect 51764 7120 51765 7160
rect 51723 7111 51765 7120
rect 49996 7026 50036 7111
rect 49036 6952 49172 6992
rect 49516 6952 49652 6992
rect 48844 6488 48884 6497
rect 48884 6448 49076 6488
rect 48844 6439 48884 6448
rect 48939 6320 48981 6329
rect 48939 6280 48940 6320
rect 48980 6280 48981 6320
rect 48939 6271 48981 6280
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 48844 5816 48884 5825
rect 48459 5648 48501 5657
rect 48459 5608 48460 5648
rect 48500 5608 48501 5648
rect 48459 5599 48501 5608
rect 48460 5514 48500 5599
rect 48556 5564 48596 5573
rect 48268 5356 48500 5396
rect 48267 4976 48309 4985
rect 48267 4936 48268 4976
rect 48308 4936 48309 4976
rect 48267 4927 48309 4936
rect 48460 4976 48500 5356
rect 48556 5069 48596 5524
rect 48844 5396 48884 5776
rect 48652 5356 48884 5396
rect 48555 5060 48597 5069
rect 48555 5020 48556 5060
rect 48596 5020 48597 5060
rect 48555 5011 48597 5020
rect 48460 4927 48500 4936
rect 48652 4976 48692 5356
rect 48652 4927 48692 4936
rect 48843 4976 48885 4985
rect 48843 4936 48844 4976
rect 48884 4936 48885 4976
rect 48843 4927 48885 4936
rect 48940 4976 48980 6271
rect 49036 5900 49076 6448
rect 49036 5851 49076 5860
rect 49036 5648 49076 5657
rect 49132 5648 49172 6952
rect 49228 6488 49268 6497
rect 49268 6448 49556 6488
rect 49228 6439 49268 6448
rect 49516 5816 49556 6448
rect 49516 5767 49556 5776
rect 49076 5608 49172 5648
rect 49228 5648 49268 5657
rect 49036 5599 49076 5608
rect 49131 5480 49173 5489
rect 49131 5440 49132 5480
rect 49172 5440 49173 5480
rect 49131 5431 49173 5440
rect 48940 4927 48980 4936
rect 49132 4976 49172 5431
rect 49132 4927 49172 4936
rect 48268 4724 48308 4927
rect 48556 4817 48596 4902
rect 48844 4842 48884 4927
rect 49228 4901 49268 5608
rect 49324 5648 49364 5657
rect 49612 5648 49652 6952
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 50092 6488 50132 6497
rect 50188 6488 50228 7111
rect 50132 6448 50228 6488
rect 50092 6439 50132 6448
rect 49900 5648 49940 5657
rect 49612 5608 49900 5648
rect 49324 5480 49364 5608
rect 49900 5599 49940 5608
rect 50091 5648 50133 5657
rect 50091 5608 50092 5648
rect 50132 5608 50133 5648
rect 50091 5599 50133 5608
rect 49996 5564 50036 5573
rect 49996 5480 50036 5524
rect 50092 5514 50132 5599
rect 49324 5440 50036 5480
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 49227 4892 49269 4901
rect 49227 4852 49228 4892
rect 49268 4852 49269 4892
rect 49227 4843 49269 4852
rect 48555 4808 48597 4817
rect 50188 4808 50228 4817
rect 48555 4768 48556 4808
rect 48596 4768 48597 4808
rect 48555 4759 48597 4768
rect 49996 4768 50188 4808
rect 47596 4087 47636 4096
rect 47692 4136 47732 4145
rect 48268 4136 48308 4684
rect 49132 4724 49172 4733
rect 49172 4684 49556 4724
rect 49132 4675 49172 4684
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 47732 4096 48308 4136
rect 47692 4087 47732 4096
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49516 3464 49556 4684
rect 49996 4136 50036 4768
rect 50188 4759 50228 4768
rect 50763 4220 50805 4229
rect 50763 4180 50764 4220
rect 50804 4180 50805 4220
rect 50763 4171 50805 4180
rect 49996 4087 50036 4096
rect 49612 4052 49652 4061
rect 49612 3968 49652 4012
rect 49612 3928 50324 3968
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 50187 3800 50229 3809
rect 50187 3760 50188 3800
rect 50228 3760 50229 3800
rect 50187 3751 50229 3760
rect 50092 3464 50132 3473
rect 49516 3424 50092 3464
rect 50092 3415 50132 3424
rect 50188 3464 50228 3751
rect 50284 3632 50324 3928
rect 50284 3583 50324 3592
rect 50188 3415 50228 3424
rect 50380 3464 50420 3473
rect 50668 3464 50708 3473
rect 50420 3424 50668 3464
rect 50380 3415 50420 3424
rect 50668 3415 50708 3424
rect 50764 3464 50804 4171
rect 50860 4136 50900 7111
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51820 6488 51860 7288
rect 51916 7279 51956 7288
rect 51820 6439 51860 6448
rect 51436 6354 51476 6439
rect 51244 6236 51284 6247
rect 51244 6161 51284 6196
rect 51243 6152 51285 6161
rect 51243 6112 51244 6152
rect 51284 6112 51285 6152
rect 51243 6103 51285 6112
rect 51244 5657 51284 6103
rect 51243 5648 51285 5657
rect 51243 5608 51244 5648
rect 51284 5608 51285 5648
rect 51243 5599 51285 5608
rect 52012 5573 52052 9631
rect 52108 9605 52148 11143
rect 52299 11024 52341 11033
rect 52492 11024 52532 11033
rect 52299 10984 52300 11024
rect 52340 10984 52341 11024
rect 52299 10975 52341 10984
rect 52396 10984 52492 11024
rect 52203 10100 52245 10109
rect 52203 10060 52204 10100
rect 52244 10060 52245 10100
rect 52203 10051 52245 10060
rect 52204 10016 52244 10051
rect 52107 9596 52149 9605
rect 52107 9556 52108 9596
rect 52148 9556 52149 9596
rect 52107 9547 52149 9556
rect 52204 9521 52244 9976
rect 52203 9512 52245 9521
rect 52203 9472 52204 9512
rect 52244 9472 52245 9512
rect 52203 9463 52245 9472
rect 52300 9512 52340 10975
rect 52396 9680 52436 10984
rect 52492 10975 52532 10984
rect 52492 10772 52532 10781
rect 52492 10193 52532 10732
rect 52491 10184 52533 10193
rect 52491 10144 52492 10184
rect 52532 10144 52533 10184
rect 52491 10135 52533 10144
rect 52588 10184 52628 11815
rect 53739 11780 53781 11789
rect 53739 11740 53740 11780
rect 53780 11740 53781 11780
rect 53739 11731 53781 11740
rect 53643 11696 53685 11705
rect 53643 11656 53644 11696
rect 53684 11656 53685 11696
rect 53643 11647 53685 11656
rect 52683 11024 52725 11033
rect 52683 10984 52684 11024
rect 52724 10984 52725 11024
rect 52683 10975 52725 10984
rect 52780 11024 52820 11033
rect 53068 11024 53108 11033
rect 52820 10984 52916 11024
rect 52780 10975 52820 10984
rect 52684 10890 52724 10975
rect 52780 10184 52820 10193
rect 52588 10144 52780 10184
rect 52492 9680 52532 9689
rect 52396 9640 52492 9680
rect 52492 9631 52532 9640
rect 52204 9378 52244 9463
rect 52300 8093 52340 9472
rect 52395 9512 52437 9521
rect 52395 9472 52396 9512
rect 52436 9472 52437 9512
rect 52395 9463 52437 9472
rect 52396 9378 52436 9463
rect 52588 9092 52628 10144
rect 52780 10135 52820 10144
rect 52683 9680 52725 9689
rect 52683 9640 52684 9680
rect 52724 9640 52725 9680
rect 52683 9631 52725 9640
rect 52780 9680 52820 9689
rect 52876 9680 52916 10984
rect 53068 10865 53108 10984
rect 53163 11024 53205 11033
rect 53163 10984 53164 11024
rect 53204 10984 53205 11024
rect 53451 11024 53493 11033
rect 53163 10975 53205 10984
rect 53260 11001 53300 11010
rect 53164 10890 53204 10975
rect 53451 10984 53452 11024
rect 53492 10984 53493 11024
rect 53451 10975 53493 10984
rect 53548 11024 53588 11033
rect 53067 10856 53109 10865
rect 53067 10816 53068 10856
rect 53108 10816 53109 10856
rect 53067 10807 53109 10816
rect 53068 10184 53108 10807
rect 53260 10604 53300 10961
rect 53452 10890 53492 10975
rect 53548 10949 53588 10984
rect 53547 10940 53589 10949
rect 53547 10900 53548 10940
rect 53588 10900 53589 10940
rect 53547 10891 53589 10900
rect 53260 10564 53396 10604
rect 53068 10135 53108 10144
rect 53163 10100 53205 10109
rect 53163 10060 53164 10100
rect 53204 10060 53205 10100
rect 53163 10051 53205 10060
rect 53164 9966 53204 10051
rect 52820 9640 52916 9680
rect 52780 9631 52820 9640
rect 52684 9512 52724 9631
rect 52684 9463 52724 9472
rect 52876 9512 52916 9523
rect 53356 9521 53396 10564
rect 53548 10436 53588 10891
rect 53644 10604 53684 11647
rect 53740 11192 53780 11731
rect 53740 11152 54068 11192
rect 53740 11024 53780 11152
rect 53740 10975 53780 10984
rect 53932 11024 53972 11033
rect 53740 10856 53780 10865
rect 53932 10856 53972 10984
rect 53780 10816 53972 10856
rect 53740 10807 53780 10816
rect 53644 10564 53876 10604
rect 53740 10436 53780 10445
rect 53548 10396 53740 10436
rect 53740 10387 53780 10396
rect 53452 10352 53492 10361
rect 53492 10312 53684 10352
rect 53452 10303 53492 10312
rect 53644 10184 53684 10312
rect 53836 10184 53876 10564
rect 53644 10135 53684 10144
rect 53740 10144 53836 10184
rect 53451 9764 53493 9773
rect 53451 9724 53452 9764
rect 53492 9724 53493 9764
rect 53451 9715 53493 9724
rect 52876 9437 52916 9472
rect 52972 9512 53012 9521
rect 52875 9428 52917 9437
rect 52875 9388 52876 9428
rect 52916 9388 52917 9428
rect 52875 9379 52917 9388
rect 52683 9092 52725 9101
rect 52588 9052 52684 9092
rect 52724 9052 52725 9092
rect 52683 9043 52725 9052
rect 52299 8084 52341 8093
rect 52299 8044 52300 8084
rect 52340 8044 52341 8084
rect 52299 8035 52341 8044
rect 52587 8084 52629 8093
rect 52587 8044 52588 8084
rect 52628 8044 52629 8084
rect 52587 8035 52629 8044
rect 52395 6740 52437 6749
rect 52395 6700 52396 6740
rect 52436 6700 52437 6740
rect 52395 6691 52437 6700
rect 52300 5648 52340 5657
rect 52011 5564 52053 5573
rect 52011 5524 52012 5564
rect 52052 5524 52053 5564
rect 52011 5515 52053 5524
rect 52204 5144 52244 5153
rect 52300 5144 52340 5608
rect 52396 5648 52436 6691
rect 52491 6488 52533 6497
rect 52491 6448 52492 6488
rect 52532 6448 52533 6488
rect 52491 6439 52533 6448
rect 52396 5599 52436 5608
rect 52492 5564 52532 6439
rect 52588 5909 52628 8035
rect 52684 6992 52724 9043
rect 52972 8597 53012 9472
rect 53067 9512 53109 9521
rect 53067 9472 53068 9512
rect 53108 9472 53109 9512
rect 53067 9463 53109 9472
rect 53355 9512 53397 9521
rect 53355 9472 53356 9512
rect 53396 9472 53397 9512
rect 53355 9463 53397 9472
rect 52971 8588 53013 8597
rect 52971 8548 52972 8588
rect 53012 8548 53013 8588
rect 52971 8539 53013 8548
rect 52876 8168 52916 8177
rect 52972 8168 53012 8539
rect 52916 8128 53012 8168
rect 53068 8168 53108 9463
rect 53163 9092 53205 9101
rect 53163 9052 53164 9092
rect 53204 9052 53205 9092
rect 53163 9043 53205 9052
rect 53164 8672 53204 9043
rect 53164 8623 53204 8632
rect 53452 8672 53492 9715
rect 53452 8623 53492 8632
rect 53644 9512 53684 9521
rect 53740 9512 53780 10144
rect 53836 10135 53876 10144
rect 53684 9472 53780 9512
rect 53836 9512 53876 9521
rect 53355 8588 53397 8597
rect 53355 8548 53356 8588
rect 53396 8548 53397 8588
rect 53355 8539 53397 8548
rect 53547 8588 53589 8597
rect 53547 8548 53548 8588
rect 53588 8548 53589 8588
rect 53547 8539 53589 8548
rect 53068 8128 53204 8168
rect 52876 8119 52916 8128
rect 53068 8000 53108 8009
rect 52780 7960 53068 8000
rect 52780 7160 52820 7960
rect 53068 7951 53108 7960
rect 53164 8000 53204 8128
rect 53259 8084 53301 8093
rect 53259 8044 53260 8084
rect 53300 8044 53301 8084
rect 53259 8035 53301 8044
rect 52971 7832 53013 7841
rect 52971 7792 52972 7832
rect 53012 7792 53013 7832
rect 52971 7783 53013 7792
rect 52875 7496 52917 7505
rect 52875 7456 52876 7496
rect 52916 7456 52917 7496
rect 52875 7447 52917 7456
rect 52780 7111 52820 7120
rect 52876 7076 52916 7447
rect 52972 7160 53012 7783
rect 52972 7111 53012 7120
rect 53068 7160 53108 7169
rect 53068 7085 53108 7120
rect 52876 7027 52916 7036
rect 53066 7076 53108 7085
rect 53066 7036 53067 7076
rect 53107 7036 53108 7076
rect 53066 7027 53108 7036
rect 52684 6952 52820 6992
rect 52683 6488 52725 6497
rect 52683 6448 52684 6488
rect 52724 6448 52725 6488
rect 52683 6439 52725 6448
rect 52684 6354 52724 6439
rect 52587 5900 52629 5909
rect 52587 5860 52588 5900
rect 52628 5860 52629 5900
rect 52587 5851 52629 5860
rect 52780 5825 52820 6952
rect 53164 6908 53204 7960
rect 53260 8021 53300 8035
rect 53260 7949 53300 7981
rect 53356 8000 53396 8539
rect 53548 8454 53588 8539
rect 53356 7951 53396 7960
rect 53644 7337 53684 9472
rect 53740 9260 53780 9269
rect 53740 8093 53780 9220
rect 53836 8924 53876 9472
rect 54028 9017 54068 11152
rect 54316 11024 54356 11033
rect 54316 10352 54356 10984
rect 54412 10352 54452 10361
rect 54316 10312 54412 10352
rect 54412 10303 54452 10312
rect 54123 9764 54165 9773
rect 54123 9724 54124 9764
rect 54164 9724 54165 9764
rect 54123 9715 54165 9724
rect 54124 9512 54164 9715
rect 54124 9463 54164 9472
rect 54315 9512 54357 9521
rect 54315 9472 54316 9512
rect 54356 9472 54452 9512
rect 54315 9463 54357 9472
rect 54316 9378 54356 9463
rect 54220 9260 54260 9269
rect 54027 9008 54069 9017
rect 54027 8968 54028 9008
rect 54068 8968 54069 9008
rect 54027 8959 54069 8968
rect 53836 8875 53876 8884
rect 54028 8252 54068 8959
rect 53932 8212 54068 8252
rect 53739 8084 53781 8093
rect 53739 8044 53740 8084
rect 53780 8044 53781 8084
rect 53739 8035 53781 8044
rect 53740 7841 53780 8035
rect 53932 8000 53972 8212
rect 53739 7832 53781 7841
rect 53739 7792 53740 7832
rect 53780 7792 53781 7832
rect 53739 7783 53781 7792
rect 53643 7328 53685 7337
rect 53643 7288 53644 7328
rect 53684 7288 53685 7328
rect 53932 7328 53972 7960
rect 54028 8084 54068 8093
rect 54028 7832 54068 8044
rect 54123 8084 54165 8093
rect 54123 8044 54124 8084
rect 54164 8044 54165 8084
rect 54123 8035 54165 8044
rect 54124 8000 54164 8035
rect 54124 7949 54164 7960
rect 54220 8000 54260 9220
rect 54220 7951 54260 7960
rect 54316 8588 54356 8597
rect 54316 7832 54356 8548
rect 54028 7792 54356 7832
rect 54412 7337 54452 9472
rect 54604 7925 54644 12940
rect 54795 12620 54837 12629
rect 54795 12580 54796 12620
rect 54836 12580 54837 12620
rect 54795 12571 54837 12580
rect 54796 12486 54836 12571
rect 55180 12536 55220 12545
rect 56044 12536 56084 12940
rect 55220 12496 55316 12536
rect 55180 12487 55220 12496
rect 55179 12284 55221 12293
rect 55179 12244 55180 12284
rect 55220 12244 55221 12284
rect 55179 12235 55221 12244
rect 55180 11024 55220 12235
rect 55276 11864 55316 12496
rect 56044 12487 56084 12496
rect 55276 11815 55316 11824
rect 56332 11864 56372 11873
rect 56332 11444 56372 11824
rect 56428 11528 56468 13159
rect 56524 11696 56564 13168
rect 56619 13208 56661 13217
rect 56812 13208 56852 13252
rect 56619 13168 56620 13208
rect 56660 13194 56756 13208
rect 56660 13168 56716 13194
rect 56619 13159 56661 13168
rect 56812 13159 56852 13168
rect 56716 13145 56756 13154
rect 56620 13040 56660 13049
rect 56620 12629 56660 13000
rect 56715 12956 56757 12965
rect 56715 12916 56716 12956
rect 56756 12916 56757 12956
rect 56715 12907 56757 12916
rect 56619 12620 56661 12629
rect 56619 12580 56620 12620
rect 56660 12580 56661 12620
rect 56619 12571 56661 12580
rect 56524 11647 56564 11656
rect 56620 11696 56660 11705
rect 56620 11528 56660 11656
rect 56716 11696 56756 12907
rect 57388 12881 57428 13915
rect 57483 13124 57525 13133
rect 57483 13084 57484 13124
rect 57524 13084 57525 13124
rect 57483 13075 57525 13084
rect 57484 12980 57524 13075
rect 57676 13049 57716 14419
rect 57771 14300 57813 14309
rect 57771 14260 57772 14300
rect 57812 14260 57813 14300
rect 57771 14251 57813 14260
rect 57772 14069 57812 14251
rect 57772 14020 57812 14029
rect 57868 13964 57908 15847
rect 58348 15560 58388 15569
rect 58348 14477 58388 15520
rect 58636 14888 58676 14897
rect 58540 14848 58636 14888
rect 58347 14468 58389 14477
rect 58347 14428 58348 14468
rect 58388 14428 58389 14468
rect 58347 14419 58389 14428
rect 57963 14300 58005 14309
rect 57963 14260 57964 14300
rect 58004 14260 58005 14300
rect 57963 14251 58005 14260
rect 57772 13924 57908 13964
rect 57964 14048 58004 14251
rect 57772 13208 57812 13924
rect 57868 13796 57908 13805
rect 57868 13469 57908 13756
rect 57867 13460 57909 13469
rect 57867 13420 57868 13460
rect 57908 13420 57909 13460
rect 57867 13411 57909 13420
rect 57867 13292 57909 13301
rect 57867 13252 57868 13292
rect 57908 13252 57909 13292
rect 57867 13243 57909 13252
rect 57772 13159 57812 13168
rect 57675 13040 57717 13049
rect 57675 13000 57676 13040
rect 57716 13000 57717 13040
rect 57675 12991 57717 13000
rect 57868 12980 57908 13243
rect 57964 13208 58004 14008
rect 58156 14048 58196 14057
rect 58156 13880 58196 14008
rect 58540 14048 58580 14848
rect 58636 14839 58676 14848
rect 58924 14561 58964 16192
rect 59212 16192 59308 16232
rect 59348 16192 59540 16232
rect 59596 17032 59695 17072
rect 59884 17116 59985 17156
rect 58923 14552 58965 14561
rect 58923 14512 58924 14552
rect 58964 14512 58965 14552
rect 58923 14503 58965 14512
rect 58540 13999 58580 14008
rect 58156 13840 58964 13880
rect 58827 13712 58869 13721
rect 58827 13672 58828 13712
rect 58868 13672 58869 13712
rect 58827 13663 58869 13672
rect 58251 13628 58293 13637
rect 58251 13588 58252 13628
rect 58292 13588 58293 13628
rect 58251 13579 58293 13588
rect 58060 13208 58100 13217
rect 57964 13168 58060 13208
rect 58060 13159 58100 13168
rect 58156 13124 58196 13133
rect 58059 13040 58101 13049
rect 58059 13000 58060 13040
rect 58100 13000 58101 13040
rect 58059 12991 58101 13000
rect 57484 12940 57620 12980
rect 57868 12940 58004 12980
rect 57387 12872 57429 12881
rect 57387 12832 57388 12872
rect 57428 12832 57429 12872
rect 57387 12823 57429 12832
rect 57195 12704 57237 12713
rect 57195 12664 57196 12704
rect 57236 12664 57237 12704
rect 57195 12655 57237 12664
rect 57196 12570 57236 12655
rect 57483 11948 57525 11957
rect 57483 11908 57484 11948
rect 57524 11908 57525 11948
rect 57483 11899 57525 11908
rect 56811 11864 56853 11873
rect 56811 11824 56812 11864
rect 56852 11824 56853 11864
rect 56811 11815 56853 11824
rect 57292 11864 57332 11873
rect 56716 11647 56756 11656
rect 56812 11696 56852 11815
rect 57292 11705 57332 11824
rect 57484 11780 57524 11899
rect 57484 11731 57524 11740
rect 56812 11647 56852 11656
rect 57291 11696 57333 11705
rect 57291 11656 57292 11696
rect 57332 11656 57333 11696
rect 57580 11696 57620 12940
rect 57867 12872 57909 12881
rect 57867 12832 57868 12872
rect 57908 12832 57909 12872
rect 57867 12823 57909 12832
rect 57675 12704 57717 12713
rect 57675 12664 57676 12704
rect 57716 12664 57717 12704
rect 57675 12655 57717 12664
rect 57676 11873 57716 12655
rect 57771 12452 57813 12461
rect 57771 12412 57772 12452
rect 57812 12412 57813 12452
rect 57771 12403 57813 12412
rect 57772 12318 57812 12403
rect 57675 11864 57717 11873
rect 57675 11824 57676 11864
rect 57716 11824 57717 11864
rect 57675 11815 57717 11824
rect 57676 11696 57716 11705
rect 57580 11656 57676 11696
rect 57291 11647 57333 11656
rect 57676 11647 57716 11656
rect 57868 11696 57908 12823
rect 57964 12704 58004 12940
rect 57964 12655 58004 12664
rect 57964 12284 58004 12295
rect 57964 12209 58004 12244
rect 57963 12200 58005 12209
rect 57963 12160 57964 12200
rect 58004 12160 58005 12200
rect 57963 12151 58005 12160
rect 57963 11864 58005 11873
rect 57963 11824 57964 11864
rect 58004 11824 58005 11864
rect 57963 11815 58005 11824
rect 57868 11647 57908 11656
rect 57964 11696 58004 11815
rect 57964 11647 58004 11656
rect 56428 11488 56660 11528
rect 56332 11404 56660 11444
rect 56331 11276 56373 11285
rect 56331 11236 56332 11276
rect 56372 11236 56373 11276
rect 56331 11227 56373 11236
rect 55180 10975 55220 10984
rect 56332 11192 56372 11227
rect 56332 10865 56372 11152
rect 56524 11024 56564 11033
rect 56620 11024 56660 11404
rect 56908 11024 56948 11033
rect 56620 10984 56908 11024
rect 56331 10856 56373 10865
rect 56331 10816 56332 10856
rect 56372 10816 56373 10856
rect 56331 10807 56373 10816
rect 56524 10445 56564 10984
rect 56908 10975 56948 10984
rect 56523 10436 56565 10445
rect 56523 10396 56524 10436
rect 56564 10396 56565 10436
rect 56523 10387 56565 10396
rect 56715 9764 56757 9773
rect 56715 9724 56716 9764
rect 56756 9724 56757 9764
rect 56715 9715 56757 9724
rect 54796 9344 54836 9353
rect 54700 8672 54740 8681
rect 54796 8672 54836 9304
rect 56428 9344 56468 9353
rect 54740 8632 54836 8672
rect 55564 8672 55604 8681
rect 54700 8623 54740 8632
rect 54603 7916 54645 7925
rect 54603 7876 54604 7916
rect 54644 7876 54645 7916
rect 54603 7867 54645 7876
rect 54219 7328 54261 7337
rect 53932 7288 54164 7328
rect 53452 7253 53492 7284
rect 53643 7279 53685 7288
rect 53451 7244 53493 7253
rect 53451 7204 53452 7244
rect 53492 7204 53493 7244
rect 53451 7195 53493 7204
rect 53452 7160 53492 7195
rect 52876 6868 53204 6908
rect 53260 7118 53300 7127
rect 52779 5816 52821 5825
rect 52779 5776 52780 5816
rect 52820 5776 52821 5816
rect 52779 5767 52821 5776
rect 52588 5648 52628 5657
rect 52780 5648 52820 5657
rect 52628 5608 52780 5648
rect 52588 5599 52628 5608
rect 52780 5599 52820 5608
rect 52876 5648 52916 6868
rect 53260 6740 53300 7078
rect 53355 7076 53397 7085
rect 53355 7036 53356 7076
rect 53396 7036 53397 7076
rect 53355 7027 53397 7036
rect 53356 6942 53396 7027
rect 53260 6700 53396 6740
rect 52971 5900 53013 5909
rect 53356 5900 53396 6700
rect 52971 5860 52972 5900
rect 53012 5860 53013 5900
rect 52971 5851 53013 5860
rect 53164 5860 53396 5900
rect 52492 5515 52532 5524
rect 52395 5480 52437 5489
rect 52395 5440 52396 5480
rect 52436 5440 52437 5480
rect 52395 5431 52437 5440
rect 52244 5104 52340 5144
rect 52204 5095 52244 5104
rect 51532 4976 51572 4985
rect 51532 4397 51572 4936
rect 51628 4976 51668 4985
rect 51531 4388 51573 4397
rect 51531 4348 51532 4388
rect 51572 4348 51573 4388
rect 51531 4339 51573 4348
rect 51628 4313 51668 4936
rect 51819 4976 51861 4985
rect 51819 4936 51820 4976
rect 51860 4936 51861 4976
rect 51819 4927 51861 4936
rect 52012 4976 52052 4985
rect 51820 4842 51860 4927
rect 51819 4724 51861 4733
rect 51819 4684 51820 4724
rect 51860 4684 51861 4724
rect 51819 4675 51861 4684
rect 51820 4590 51860 4675
rect 51723 4472 51765 4481
rect 51723 4432 51724 4472
rect 51764 4432 51765 4472
rect 51723 4423 51765 4432
rect 51627 4304 51669 4313
rect 51627 4264 51628 4304
rect 51668 4264 51669 4304
rect 51627 4255 51669 4264
rect 50860 4087 50900 4096
rect 50859 3968 50901 3977
rect 50859 3928 50860 3968
rect 50900 3928 50901 3968
rect 50859 3919 50901 3928
rect 50764 3415 50804 3424
rect 50860 3464 50900 3919
rect 51628 3809 51668 4255
rect 51627 3800 51669 3809
rect 51627 3760 51628 3800
rect 51668 3760 51669 3800
rect 51627 3751 51669 3760
rect 50860 3415 50900 3424
rect 50955 3464 50997 3473
rect 50955 3424 50956 3464
rect 50996 3424 50997 3464
rect 50955 3415 50997 3424
rect 51724 3464 51764 4423
rect 52012 4388 52052 4936
rect 52012 4339 52052 4348
rect 52108 4976 52148 4985
rect 52108 4145 52148 4936
rect 52300 4976 52340 4985
rect 52396 4976 52436 5431
rect 52340 4936 52436 4976
rect 52492 4976 52532 4985
rect 52107 4136 52149 4145
rect 52107 4096 52108 4136
rect 52148 4096 52149 4136
rect 52107 4087 52149 4096
rect 52012 3968 52052 3977
rect 52052 3928 52148 3968
rect 52012 3919 52052 3928
rect 52108 3557 52148 3928
rect 52107 3548 52149 3557
rect 52107 3508 52108 3548
rect 52148 3508 52149 3548
rect 52107 3499 52149 3508
rect 51724 3415 51764 3424
rect 52011 3464 52053 3473
rect 52011 3424 52012 3464
rect 52052 3424 52053 3464
rect 52011 3415 52053 3424
rect 50956 3330 50996 3415
rect 52012 3330 52052 3415
rect 52108 3414 52148 3499
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 52300 2717 52340 4936
rect 52395 4724 52437 4733
rect 52395 4684 52396 4724
rect 52436 4684 52437 4724
rect 52395 4675 52437 4684
rect 52396 4136 52436 4675
rect 52396 4087 52436 4096
rect 52396 3296 52436 3305
rect 52492 3296 52532 4936
rect 52683 4976 52725 4985
rect 52876 4976 52916 5608
rect 52683 4936 52684 4976
rect 52724 4936 52725 4976
rect 52683 4927 52725 4936
rect 52780 4936 52916 4976
rect 52972 5648 53012 5851
rect 52684 4842 52724 4927
rect 52588 4724 52628 4733
rect 52588 4313 52628 4684
rect 52683 4388 52725 4397
rect 52683 4348 52684 4388
rect 52724 4348 52725 4388
rect 52683 4339 52725 4348
rect 52587 4304 52629 4313
rect 52587 4264 52588 4304
rect 52628 4264 52629 4304
rect 52587 4255 52629 4264
rect 52587 4136 52629 4145
rect 52587 4096 52588 4136
rect 52628 4096 52629 4136
rect 52587 4087 52629 4096
rect 52588 3464 52628 4087
rect 52684 3548 52724 4339
rect 52780 4313 52820 4936
rect 52876 4808 52916 4817
rect 52779 4304 52821 4313
rect 52779 4264 52780 4304
rect 52820 4264 52821 4304
rect 52779 4255 52821 4264
rect 52780 4136 52820 4145
rect 52876 4136 52916 4768
rect 52820 4096 52916 4136
rect 52780 4087 52820 4096
rect 52972 3977 53012 5608
rect 53067 5648 53109 5657
rect 53067 5608 53068 5648
rect 53108 5608 53109 5648
rect 53067 5599 53109 5608
rect 53068 5514 53108 5599
rect 53164 5573 53204 5860
rect 53452 5816 53492 7120
rect 53356 5776 53492 5816
rect 53548 7160 53588 7169
rect 53163 5564 53205 5573
rect 53163 5524 53164 5564
rect 53204 5524 53205 5564
rect 53163 5515 53205 5524
rect 53259 4136 53301 4145
rect 53356 4136 53396 5776
rect 53548 5657 53588 7120
rect 53547 5648 53589 5657
rect 53547 5608 53548 5648
rect 53588 5608 53589 5648
rect 53547 5599 53589 5608
rect 53644 4901 53684 7279
rect 54124 6488 54164 7288
rect 54219 7288 54220 7328
rect 54260 7288 54261 7328
rect 54219 7279 54261 7288
rect 54411 7328 54453 7337
rect 54411 7288 54412 7328
rect 54452 7288 54453 7328
rect 54411 7279 54453 7288
rect 55276 7328 55316 7337
rect 54220 7160 54260 7279
rect 54891 7244 54933 7253
rect 54891 7204 54892 7244
rect 54932 7204 54933 7244
rect 54891 7195 54933 7204
rect 54220 7111 54260 7120
rect 54412 7160 54452 7169
rect 54452 7120 54548 7160
rect 54412 7111 54452 7120
rect 54316 7076 54356 7085
rect 54316 6749 54356 7036
rect 54315 6740 54357 6749
rect 54315 6700 54316 6740
rect 54356 6700 54357 6740
rect 54315 6691 54357 6700
rect 54219 6572 54261 6581
rect 54219 6532 54220 6572
rect 54260 6532 54261 6572
rect 54219 6523 54261 6532
rect 54028 6448 54124 6488
rect 53836 6236 53876 6245
rect 53740 6196 53836 6236
rect 53740 5657 53780 6196
rect 53836 6187 53876 6196
rect 53836 5741 53876 5772
rect 53835 5732 53877 5741
rect 53835 5692 53836 5732
rect 53876 5692 53877 5732
rect 53835 5683 53877 5692
rect 53739 5648 53781 5657
rect 53739 5608 53740 5648
rect 53780 5608 53781 5648
rect 53739 5599 53781 5608
rect 53836 5648 53876 5683
rect 53643 4892 53685 4901
rect 53643 4852 53644 4892
rect 53684 4852 53685 4892
rect 53643 4843 53685 4852
rect 53836 4481 53876 5608
rect 54028 4985 54068 6448
rect 54124 6439 54164 6448
rect 54220 6438 54260 6523
rect 54316 6488 54356 6691
rect 54316 6439 54356 6448
rect 54412 6488 54452 6497
rect 54412 5825 54452 6448
rect 54508 5900 54548 7120
rect 54892 7110 54932 7195
rect 55084 6992 55124 7001
rect 54892 6952 55084 6992
rect 54603 6572 54645 6581
rect 54603 6532 54604 6572
rect 54644 6532 54645 6572
rect 54603 6523 54645 6532
rect 54604 6438 54644 6523
rect 54508 5851 54548 5860
rect 54411 5816 54453 5825
rect 54411 5776 54412 5816
rect 54452 5776 54453 5816
rect 54411 5767 54453 5776
rect 54795 5816 54837 5825
rect 54795 5776 54796 5816
rect 54836 5776 54837 5816
rect 54795 5767 54837 5776
rect 54123 5732 54165 5741
rect 54123 5692 54124 5732
rect 54164 5692 54165 5732
rect 54123 5683 54165 5692
rect 54699 5732 54741 5741
rect 54699 5692 54700 5732
rect 54740 5692 54741 5732
rect 54699 5683 54741 5692
rect 54796 5732 54836 5767
rect 54124 5648 54164 5683
rect 54124 5597 54164 5608
rect 54219 5648 54261 5657
rect 54219 5608 54220 5648
rect 54260 5608 54261 5648
rect 54219 5599 54261 5608
rect 54700 5648 54740 5683
rect 54796 5681 54836 5692
rect 54892 5657 54932 6952
rect 55084 6943 55124 6952
rect 55276 6824 55316 7288
rect 55564 7169 55604 8632
rect 55947 8588 55989 8597
rect 55947 8548 55948 8588
rect 55988 8548 55989 8588
rect 55947 8539 55989 8548
rect 55948 8084 55988 8539
rect 55948 8035 55988 8044
rect 56332 8000 56372 8009
rect 56428 8000 56468 9304
rect 56716 8924 56756 9715
rect 57292 9428 57332 11647
rect 57772 11528 57812 11537
rect 57676 11488 57772 11528
rect 57580 10352 57620 10361
rect 57387 10268 57429 10277
rect 57387 10228 57388 10268
rect 57428 10228 57429 10268
rect 57387 10219 57429 10228
rect 57388 10134 57428 10219
rect 57580 10016 57620 10312
rect 57676 10184 57716 11488
rect 57772 11479 57812 11488
rect 57772 11024 57812 11033
rect 58060 11024 58100 12991
rect 58156 12713 58196 13084
rect 58155 12704 58197 12713
rect 58155 12664 58156 12704
rect 58196 12664 58197 12704
rect 58155 12655 58197 12664
rect 58156 12536 58196 12545
rect 58252 12536 58292 13579
rect 58635 13460 58677 13469
rect 58635 13420 58636 13460
rect 58676 13420 58677 13460
rect 58635 13411 58677 13420
rect 58444 13376 58484 13385
rect 58196 12496 58292 12536
rect 58348 13336 58444 13376
rect 58348 12536 58388 13336
rect 58444 13327 58484 13336
rect 58443 13208 58485 13217
rect 58443 13168 58444 13208
rect 58484 13168 58485 13208
rect 58443 13159 58485 13168
rect 58636 13208 58676 13411
rect 58636 13159 58676 13168
rect 58731 13208 58773 13217
rect 58731 13168 58732 13208
rect 58772 13168 58773 13208
rect 58731 13159 58773 13168
rect 58828 13208 58868 13663
rect 58924 13460 58964 13840
rect 58924 13411 58964 13420
rect 58924 13208 58964 13217
rect 58828 13168 58924 13208
rect 58156 12487 58196 12496
rect 58348 12487 58388 12496
rect 58252 12368 58292 12377
rect 58444 12368 58484 13159
rect 58539 13124 58581 13133
rect 58539 13084 58540 13124
rect 58580 13084 58581 13124
rect 58539 13075 58581 13084
rect 58292 12328 58484 12368
rect 58252 12319 58292 12328
rect 58251 12200 58293 12209
rect 58251 12160 58252 12200
rect 58292 12160 58293 12200
rect 58251 12151 58293 12160
rect 58252 11696 58292 12151
rect 58540 11705 58580 13075
rect 58732 13074 58772 13159
rect 57812 10984 58100 11024
rect 58156 11528 58196 11537
rect 57772 10975 57812 10984
rect 58059 10436 58101 10445
rect 58059 10396 58060 10436
rect 58100 10396 58101 10436
rect 58059 10387 58101 10396
rect 57867 10352 57909 10361
rect 57867 10312 57868 10352
rect 57908 10312 57909 10352
rect 57867 10303 57909 10312
rect 57772 10184 57812 10193
rect 57676 10144 57772 10184
rect 57772 10135 57812 10144
rect 57868 10184 57908 10303
rect 58060 10302 58100 10387
rect 57868 10135 57908 10144
rect 58060 10184 58100 10193
rect 58156 10184 58196 11488
rect 58252 11444 58292 11656
rect 58347 11696 58389 11705
rect 58347 11656 58348 11696
rect 58388 11656 58389 11696
rect 58347 11647 58389 11656
rect 58444 11696 58484 11705
rect 58348 11562 58388 11647
rect 58252 11404 58388 11444
rect 58348 10193 58388 11404
rect 58444 11201 58484 11656
rect 58539 11696 58581 11705
rect 58539 11656 58540 11696
rect 58580 11656 58581 11696
rect 58539 11647 58581 11656
rect 58828 11696 58868 13168
rect 58924 13159 58964 13168
rect 59019 12620 59061 12629
rect 59019 12580 59020 12620
rect 59060 12580 59061 12620
rect 59019 12571 59061 12580
rect 59020 12041 59060 12571
rect 59212 12545 59252 16192
rect 59308 16183 59348 16192
rect 59404 16064 59444 16073
rect 59596 16064 59636 17032
rect 59444 16024 59636 16064
rect 59692 16232 59732 16241
rect 59884 16232 59924 17116
rect 60055 17072 60095 17472
rect 60345 17072 60385 17472
rect 59732 16192 59924 16232
rect 59980 17032 60095 17072
rect 60268 17032 60385 17072
rect 60455 17072 60495 17472
rect 60745 17165 60785 17472
rect 60744 17156 60786 17165
rect 60744 17116 60745 17156
rect 60785 17116 60786 17156
rect 60744 17107 60786 17116
rect 60855 17072 60895 17472
rect 60939 17156 60981 17165
rect 61145 17156 61185 17472
rect 60939 17116 60940 17156
rect 60980 17116 60981 17156
rect 60939 17107 60981 17116
rect 61132 17116 61185 17156
rect 60455 17032 60500 17072
rect 59404 16015 59444 16024
rect 59499 15896 59541 15905
rect 59499 15856 59500 15896
rect 59540 15856 59541 15896
rect 59499 15847 59541 15856
rect 59500 15728 59540 15847
rect 59500 15679 59540 15688
rect 59500 15308 59540 15317
rect 59500 14729 59540 15268
rect 59499 14720 59541 14729
rect 59499 14680 59500 14720
rect 59540 14680 59541 14720
rect 59499 14671 59541 14680
rect 59403 14384 59445 14393
rect 59403 14344 59404 14384
rect 59444 14344 59445 14384
rect 59403 14335 59445 14344
rect 59404 14048 59444 14335
rect 59404 13999 59444 14008
rect 59307 13376 59349 13385
rect 59307 13336 59308 13376
rect 59348 13336 59349 13376
rect 59307 13327 59349 13336
rect 59211 12536 59253 12545
rect 59211 12496 59212 12536
rect 59252 12496 59253 12536
rect 59211 12487 59253 12496
rect 59308 12536 59348 13327
rect 59692 12629 59732 16192
rect 59788 16064 59828 16073
rect 59980 16064 60020 17032
rect 60268 16988 60308 17032
rect 59828 16024 60020 16064
rect 60076 16948 60308 16988
rect 60076 16232 60116 16948
rect 60460 16736 60500 17032
rect 60844 17032 60895 17072
rect 60844 16736 60884 17032
rect 60172 16696 60500 16736
rect 60556 16696 60884 16736
rect 60172 16484 60212 16696
rect 60172 16435 60212 16444
rect 60556 16484 60596 16696
rect 60940 16652 60980 17107
rect 60748 16612 60980 16652
rect 60748 16484 60788 16612
rect 60556 16435 60596 16444
rect 60652 16444 60788 16484
rect 60843 16484 60885 16493
rect 60843 16444 60844 16484
rect 60884 16444 60885 16484
rect 59788 16015 59828 16024
rect 59979 15392 60021 15401
rect 59979 15352 59980 15392
rect 60020 15352 60021 15392
rect 59979 15343 60021 15352
rect 59980 12980 60020 15343
rect 59884 12940 60020 12980
rect 59691 12620 59733 12629
rect 59691 12580 59692 12620
rect 59732 12580 59733 12620
rect 59691 12571 59733 12580
rect 59509 12549 59549 12558
rect 59549 12509 59636 12536
rect 59509 12496 59636 12509
rect 59308 12452 59348 12496
rect 59596 12452 59636 12496
rect 59308 12412 59540 12452
rect 59596 12412 59732 12452
rect 59500 12368 59540 12412
rect 59500 12328 59636 12368
rect 59404 12284 59444 12293
rect 59116 12244 59404 12284
rect 59019 12032 59061 12041
rect 59019 11992 59020 12032
rect 59060 11992 59061 12032
rect 59019 11983 59061 11992
rect 58828 11647 58868 11656
rect 59020 11696 59060 11705
rect 58923 11612 58965 11621
rect 58923 11572 58924 11612
rect 58964 11572 58965 11612
rect 58923 11563 58965 11572
rect 58924 11478 58964 11563
rect 58443 11192 58485 11201
rect 58923 11192 58965 11201
rect 58443 11152 58444 11192
rect 58484 11152 58580 11192
rect 58443 11143 58485 11152
rect 58100 10144 58196 10184
rect 58252 10184 58292 10193
rect 58060 10135 58100 10144
rect 58252 10016 58292 10144
rect 58347 10184 58389 10193
rect 58347 10144 58348 10184
rect 58388 10144 58389 10184
rect 58347 10135 58389 10144
rect 58444 10184 58484 10193
rect 57580 9976 58292 10016
rect 58348 10016 58388 10025
rect 58059 9680 58101 9689
rect 58059 9640 58060 9680
rect 58100 9640 58101 9680
rect 58059 9631 58101 9640
rect 57772 9512 57812 9521
rect 57676 9472 57772 9512
rect 57388 9428 57428 9437
rect 57292 9388 57388 9428
rect 57388 9379 57428 9388
rect 56716 8875 56756 8884
rect 57580 9260 57620 9269
rect 57580 8336 57620 9220
rect 57676 8672 57716 9472
rect 57772 9463 57812 9472
rect 57964 9512 58004 9521
rect 57772 9260 57812 9269
rect 57772 8849 57812 9220
rect 57964 8849 58004 9472
rect 58060 9512 58100 9631
rect 58060 9463 58100 9472
rect 58059 8924 58101 8933
rect 58059 8884 58060 8924
rect 58100 8884 58101 8924
rect 58059 8875 58101 8884
rect 57771 8840 57813 8849
rect 57771 8800 57772 8840
rect 57812 8800 57813 8840
rect 57771 8791 57813 8800
rect 57963 8840 58005 8849
rect 57963 8800 57964 8840
rect 58004 8800 58005 8840
rect 57963 8791 58005 8800
rect 57772 8672 57812 8681
rect 57676 8632 57772 8672
rect 57772 8623 57812 8632
rect 57868 8672 57908 8681
rect 57868 8513 57908 8632
rect 57964 8672 58004 8681
rect 57867 8504 57909 8513
rect 57867 8464 57868 8504
rect 57908 8464 57909 8504
rect 57867 8455 57909 8464
rect 57964 8336 58004 8632
rect 57580 8296 58004 8336
rect 56372 7960 56468 8000
rect 57196 8000 57236 8009
rect 56332 7951 56372 7960
rect 55563 7160 55605 7169
rect 55563 7120 55564 7160
rect 55604 7120 55605 7160
rect 55563 7111 55605 7120
rect 54988 6784 55316 6824
rect 54988 6488 55028 6784
rect 54988 6439 55028 6448
rect 55083 6488 55125 6497
rect 55083 6448 55084 6488
rect 55124 6448 55125 6488
rect 55083 6439 55125 6448
rect 54220 5514 54260 5599
rect 54700 5597 54740 5608
rect 54891 5648 54933 5657
rect 54891 5608 54892 5648
rect 54932 5608 54933 5648
rect 54891 5599 54933 5608
rect 54892 5514 54932 5599
rect 54027 4976 54069 4985
rect 54027 4936 54028 4976
rect 54068 4936 54069 4976
rect 54027 4927 54069 4936
rect 53835 4472 53877 4481
rect 53835 4432 53836 4472
rect 53876 4432 53877 4472
rect 53835 4423 53877 4432
rect 55084 4145 55124 6439
rect 55180 4304 55220 4313
rect 53259 4096 53260 4136
rect 53300 4096 53396 4136
rect 53643 4136 53685 4145
rect 53643 4096 53644 4136
rect 53684 4096 53685 4136
rect 53259 4087 53301 4096
rect 53643 4087 53685 4096
rect 55083 4136 55125 4145
rect 55083 4096 55084 4136
rect 55124 4096 55125 4136
rect 55083 4087 55125 4096
rect 53260 4068 53300 4087
rect 53644 4002 53684 4087
rect 52971 3968 53013 3977
rect 52971 3928 52972 3968
rect 53012 3928 53013 3968
rect 52971 3919 53013 3928
rect 54796 3968 54836 3979
rect 54796 3893 54836 3928
rect 52779 3884 52821 3893
rect 52779 3844 52780 3884
rect 52820 3844 52821 3884
rect 52779 3835 52821 3844
rect 54795 3884 54837 3893
rect 54795 3844 54796 3884
rect 54836 3844 54837 3884
rect 54795 3835 54837 3844
rect 52684 3499 52724 3508
rect 52780 3473 52820 3835
rect 53931 3632 53973 3641
rect 53931 3592 53932 3632
rect 53972 3592 53973 3632
rect 53931 3583 53973 3592
rect 53932 3498 53972 3583
rect 52588 3415 52628 3424
rect 52779 3464 52821 3473
rect 52779 3424 52780 3464
rect 52820 3424 52821 3464
rect 52779 3415 52821 3424
rect 55084 3464 55124 4087
rect 55180 3473 55220 4264
rect 55371 4220 55413 4229
rect 55371 4180 55372 4220
rect 55412 4180 55413 4220
rect 55371 4171 55413 4180
rect 55084 3415 55124 3424
rect 55179 3464 55221 3473
rect 55179 3424 55180 3464
rect 55220 3424 55221 3464
rect 55179 3415 55221 3424
rect 52780 3330 52820 3415
rect 52436 3256 52532 3296
rect 52396 3247 52436 3256
rect 54028 2792 54068 2801
rect 53932 2752 54028 2792
rect 8907 2708 8949 2717
rect 8907 2668 8908 2708
rect 8948 2668 8949 2708
rect 8907 2659 8949 2668
rect 52299 2708 52341 2717
rect 52299 2668 52300 2708
rect 52340 2668 52341 2708
rect 52299 2659 52341 2668
rect 3148 2573 3188 2584
rect 4299 2624 4341 2633
rect 4299 2584 4300 2624
rect 4340 2584 4341 2624
rect 4299 2575 4341 2584
rect 4779 2624 4821 2633
rect 4779 2584 4780 2624
rect 4820 2584 4821 2624
rect 4779 2575 4821 2584
rect 2956 2456 2996 2465
rect 2668 2416 2956 2456
rect 2956 2407 2996 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 53548 1952 53588 1961
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 53548 1373 53588 1912
rect 53932 1952 53972 2752
rect 54028 2743 54068 2752
rect 55372 2624 55412 4171
rect 55467 3968 55509 3977
rect 55467 3928 55468 3968
rect 55508 3928 55509 3968
rect 55467 3919 55509 3928
rect 55372 2575 55412 2584
rect 55468 2624 55508 3919
rect 55564 2900 55604 7111
rect 56908 7076 56948 7085
rect 55851 6488 55893 6497
rect 55851 6448 55852 6488
rect 55892 6448 55893 6488
rect 55851 6439 55893 6448
rect 55852 6354 55892 6439
rect 56908 6329 56948 7036
rect 57003 6824 57045 6833
rect 57003 6784 57004 6824
rect 57044 6784 57045 6824
rect 57003 6775 57045 6784
rect 57004 6656 57044 6775
rect 57004 6607 57044 6616
rect 57196 6488 57236 7960
rect 57292 7160 57332 7169
rect 57332 7120 57428 7160
rect 57292 7111 57332 7120
rect 57291 6488 57333 6497
rect 57196 6448 57292 6488
rect 57332 6448 57333 6488
rect 57291 6439 57333 6448
rect 56907 6320 56949 6329
rect 56907 6280 56908 6320
rect 56948 6280 56949 6320
rect 56907 6271 56949 6280
rect 57004 6236 57044 6245
rect 56620 5816 56660 5825
rect 56235 5648 56277 5657
rect 56235 5608 56236 5648
rect 56276 5608 56277 5648
rect 56235 5599 56277 5608
rect 56428 5648 56468 5657
rect 56236 5514 56276 5599
rect 56332 5564 56372 5573
rect 55756 5144 55796 5153
rect 55796 5104 56180 5144
rect 55756 5095 55796 5104
rect 56140 5060 56180 5104
rect 56140 5011 56180 5020
rect 56332 4985 56372 5524
rect 55659 4976 55701 4985
rect 55659 4936 55660 4976
rect 55700 4936 55701 4976
rect 55659 4927 55701 4936
rect 55852 4976 55892 4985
rect 55660 4817 55700 4927
rect 55659 4808 55701 4817
rect 55659 4768 55660 4808
rect 55700 4768 55701 4808
rect 55659 4759 55701 4768
rect 55852 4397 55892 4936
rect 55947 4976 55989 4985
rect 55947 4936 55948 4976
rect 55988 4936 55989 4976
rect 55947 4927 55989 4936
rect 56331 4976 56373 4985
rect 56331 4936 56332 4976
rect 56372 4936 56373 4976
rect 56331 4927 56373 4936
rect 55948 4842 55988 4927
rect 56139 4808 56181 4817
rect 56139 4768 56140 4808
rect 56180 4768 56181 4808
rect 56428 4808 56468 5608
rect 56524 4976 56564 4985
rect 56620 4976 56660 5776
rect 57004 5741 57044 6196
rect 57003 5732 57045 5741
rect 57003 5692 57004 5732
rect 57044 5692 57045 5732
rect 57003 5683 57045 5692
rect 56564 4936 56660 4976
rect 57292 4976 57332 6439
rect 57388 6320 57428 7120
rect 57964 6665 58004 8296
rect 58060 8672 58100 8875
rect 58060 8093 58100 8632
rect 58156 8429 58196 9976
rect 58251 9848 58293 9857
rect 58251 9808 58252 9848
rect 58292 9808 58293 9848
rect 58251 9799 58293 9808
rect 58252 8756 58292 9799
rect 58348 9689 58388 9976
rect 58347 9680 58389 9689
rect 58347 9640 58348 9680
rect 58388 9640 58389 9680
rect 58347 9631 58389 9640
rect 58348 9512 58388 9521
rect 58348 9101 58388 9472
rect 58347 9092 58389 9101
rect 58347 9052 58348 9092
rect 58388 9052 58389 9092
rect 58347 9043 58389 9052
rect 58252 8707 58292 8716
rect 58444 8672 58484 10144
rect 58540 10184 58580 11152
rect 58923 11152 58924 11192
rect 58964 11152 58965 11192
rect 58923 11143 58965 11152
rect 58924 11058 58964 11143
rect 59020 10940 59060 11656
rect 59116 11696 59156 12244
rect 59404 12235 59444 12244
rect 59499 12032 59541 12041
rect 59499 11992 59500 12032
rect 59540 11992 59541 12032
rect 59499 11983 59541 11992
rect 59116 11647 59156 11656
rect 59307 11612 59349 11621
rect 59307 11572 59308 11612
rect 59348 11572 59349 11612
rect 59307 11563 59349 11572
rect 59308 11478 59348 11563
rect 59307 11360 59349 11369
rect 59307 11320 59308 11360
rect 59348 11320 59349 11360
rect 59307 11311 59349 11320
rect 59020 10900 59252 10940
rect 59116 10772 59156 10781
rect 58732 10352 58772 10363
rect 58732 10277 58772 10312
rect 58731 10268 58773 10277
rect 58731 10228 58732 10268
rect 58772 10228 58773 10268
rect 58731 10219 58773 10228
rect 58923 10268 58965 10277
rect 58923 10228 58924 10268
rect 58964 10228 58965 10268
rect 58923 10219 58965 10228
rect 58540 10135 58580 10144
rect 58924 10134 58964 10219
rect 59116 10184 59156 10732
rect 59212 10361 59252 10900
rect 59211 10352 59253 10361
rect 59211 10312 59212 10352
rect 59252 10312 59253 10352
rect 59211 10303 59253 10312
rect 59116 10135 59156 10144
rect 59212 10100 59252 10303
rect 59308 10184 59348 11311
rect 59403 11192 59445 11201
rect 59403 11152 59404 11192
rect 59444 11152 59445 11192
rect 59403 11143 59445 11152
rect 59404 11108 59444 11143
rect 59404 11057 59444 11068
rect 59500 11024 59540 11983
rect 59500 10975 59540 10984
rect 59596 10856 59636 12328
rect 59692 12041 59732 12412
rect 59788 12368 59828 12377
rect 59691 12032 59733 12041
rect 59691 11992 59692 12032
rect 59732 11992 59733 12032
rect 59691 11983 59733 11992
rect 59692 11696 59732 11705
rect 59788 11696 59828 12328
rect 59732 11656 59828 11696
rect 59692 11647 59732 11656
rect 59788 11033 59828 11118
rect 59787 11024 59829 11033
rect 59787 10984 59788 11024
rect 59828 10984 59829 11024
rect 59787 10975 59829 10984
rect 59596 10816 59828 10856
rect 59691 10268 59733 10277
rect 59691 10228 59692 10268
rect 59732 10228 59733 10268
rect 59691 10219 59733 10228
rect 59500 10184 59540 10195
rect 59348 10144 59444 10184
rect 59308 10135 59348 10144
rect 59212 10051 59252 10060
rect 59307 9680 59349 9689
rect 59307 9640 59308 9680
rect 59348 9640 59349 9680
rect 59307 9631 59349 9640
rect 58635 9512 58677 9521
rect 58635 9472 58636 9512
rect 58676 9472 58677 9512
rect 58635 9463 58677 9472
rect 58732 9512 58772 9521
rect 58636 9378 58676 9463
rect 58732 8933 58772 9472
rect 59020 9260 59060 9269
rect 59212 9260 59252 9269
rect 58828 9220 59020 9260
rect 58731 8924 58773 8933
rect 58731 8884 58732 8924
rect 58772 8884 58773 8924
rect 58731 8875 58773 8884
rect 58731 8756 58773 8765
rect 58731 8716 58732 8756
rect 58772 8716 58773 8756
rect 58731 8707 58773 8716
rect 58635 8672 58677 8681
rect 58444 8632 58580 8672
rect 58443 8504 58485 8513
rect 58443 8464 58444 8504
rect 58484 8464 58485 8504
rect 58443 8455 58485 8464
rect 58155 8420 58197 8429
rect 58155 8380 58156 8420
rect 58196 8380 58197 8420
rect 58155 8371 58197 8380
rect 58059 8084 58101 8093
rect 58059 8044 58060 8084
rect 58100 8044 58101 8084
rect 58059 8035 58101 8044
rect 58060 7916 58100 8035
rect 58348 7916 58388 7925
rect 58060 7876 58348 7916
rect 58348 7867 58388 7876
rect 58444 7832 58484 8455
rect 58540 8252 58580 8632
rect 58635 8632 58636 8672
rect 58676 8632 58677 8672
rect 58635 8623 58677 8632
rect 58636 8538 58676 8623
rect 58732 8622 58772 8707
rect 58828 8672 58868 9220
rect 59020 9211 59060 9220
rect 59116 9220 59212 9260
rect 59019 9008 59061 9017
rect 59019 8968 59020 9008
rect 59060 8968 59061 9008
rect 59019 8959 59061 8968
rect 58828 8623 58868 8632
rect 59020 8672 59060 8959
rect 59116 8681 59156 9220
rect 59212 9211 59252 9220
rect 59211 8756 59253 8765
rect 59211 8716 59212 8756
rect 59252 8716 59253 8756
rect 59211 8707 59253 8716
rect 59020 8623 59060 8632
rect 59115 8672 59157 8681
rect 59115 8632 59116 8672
rect 59156 8632 59157 8672
rect 59115 8623 59157 8632
rect 59212 8672 59252 8707
rect 59212 8621 59252 8632
rect 59308 8672 59348 9631
rect 59404 9428 59444 10144
rect 59500 10109 59540 10144
rect 59692 10184 59732 10219
rect 59499 10100 59541 10109
rect 59499 10060 59500 10100
rect 59540 10060 59541 10100
rect 59499 10051 59541 10060
rect 59596 10100 59636 10109
rect 59404 9379 59444 9388
rect 59500 8924 59540 10051
rect 59596 9689 59636 10060
rect 59595 9680 59637 9689
rect 59595 9640 59596 9680
rect 59636 9640 59637 9680
rect 59595 9631 59637 9640
rect 59692 9521 59732 10144
rect 59500 8875 59540 8884
rect 59596 9512 59636 9521
rect 59596 8672 59636 9472
rect 59691 9512 59733 9521
rect 59691 9472 59692 9512
rect 59732 9472 59733 9512
rect 59691 9463 59733 9472
rect 59692 8756 59732 8765
rect 59788 8756 59828 10816
rect 59732 8716 59828 8756
rect 59692 8707 59732 8716
rect 59308 8623 59348 8632
rect 59404 8632 59636 8672
rect 59116 8504 59156 8513
rect 59404 8504 59444 8632
rect 59156 8464 59444 8504
rect 59499 8504 59541 8513
rect 59499 8464 59500 8504
rect 59540 8464 59541 8504
rect 59116 8455 59156 8464
rect 59499 8455 59541 8464
rect 58827 8420 58869 8429
rect 58827 8380 58828 8420
rect 58868 8380 58869 8420
rect 58827 8371 58869 8380
rect 58540 8212 58676 8252
rect 58539 8084 58581 8093
rect 58539 8044 58540 8084
rect 58580 8044 58581 8084
rect 58539 8035 58581 8044
rect 58540 8000 58580 8035
rect 58540 7949 58580 7960
rect 58636 8000 58676 8212
rect 58828 8000 58868 8371
rect 58676 7960 58772 8000
rect 58636 7951 58676 7960
rect 58444 7792 58676 7832
rect 58347 7748 58389 7757
rect 58347 7708 58348 7748
rect 58388 7708 58389 7748
rect 58347 7699 58389 7708
rect 58156 7160 58196 7169
rect 57963 6656 58005 6665
rect 57963 6616 57964 6656
rect 58004 6616 58005 6656
rect 57963 6607 58005 6616
rect 58059 6572 58101 6581
rect 58059 6532 58060 6572
rect 58100 6532 58101 6572
rect 58059 6523 58101 6532
rect 58060 6488 58100 6523
rect 58156 6497 58196 7120
rect 58060 6437 58100 6448
rect 58155 6488 58197 6497
rect 58155 6448 58156 6488
rect 58196 6448 58197 6488
rect 58155 6439 58197 6448
rect 58252 6488 58292 6497
rect 58252 6329 58292 6448
rect 58348 6488 58388 7699
rect 58539 6572 58581 6581
rect 58539 6532 58540 6572
rect 58580 6532 58581 6572
rect 58539 6523 58581 6532
rect 58348 6439 58388 6448
rect 58540 6438 58580 6523
rect 58636 6488 58676 7792
rect 58732 6824 58772 7960
rect 58828 7916 58868 7960
rect 58828 7876 59060 7916
rect 58827 7748 58869 7757
rect 58827 7708 58828 7748
rect 58868 7708 58869 7748
rect 58827 7699 58869 7708
rect 58828 7614 58868 7699
rect 58732 6784 58868 6824
rect 58731 6656 58773 6665
rect 58731 6616 58732 6656
rect 58772 6616 58773 6656
rect 58828 6656 58868 6784
rect 58828 6616 58964 6656
rect 58731 6607 58773 6616
rect 57388 6271 57428 6280
rect 58059 6320 58101 6329
rect 58059 6280 58060 6320
rect 58100 6280 58101 6320
rect 58059 6271 58101 6280
rect 58251 6320 58293 6329
rect 58251 6280 58252 6320
rect 58292 6280 58293 6320
rect 58251 6271 58293 6280
rect 58060 6186 58100 6271
rect 58059 6068 58101 6077
rect 58059 6028 58060 6068
rect 58100 6028 58101 6068
rect 58059 6019 58101 6028
rect 57388 4976 57428 4985
rect 57579 4976 57621 4985
rect 57292 4936 57388 4976
rect 57428 4936 57580 4976
rect 57620 4936 57621 4976
rect 56524 4927 56564 4936
rect 57388 4927 57428 4936
rect 57579 4927 57621 4936
rect 56715 4892 56757 4901
rect 56715 4852 56716 4892
rect 56756 4852 56757 4892
rect 56715 4843 56757 4852
rect 56523 4808 56565 4817
rect 56428 4768 56524 4808
rect 56564 4768 56565 4808
rect 56139 4759 56181 4768
rect 56523 4759 56565 4768
rect 55851 4388 55893 4397
rect 55851 4348 55852 4388
rect 55892 4348 55893 4388
rect 55851 4339 55893 4348
rect 55755 4220 55797 4229
rect 55755 4180 55756 4220
rect 55796 4180 55797 4220
rect 55755 4171 55797 4180
rect 55659 4136 55701 4145
rect 55659 4096 55660 4136
rect 55700 4096 55701 4136
rect 55659 4087 55701 4096
rect 55756 4136 55796 4171
rect 55660 4002 55700 4087
rect 55756 4085 55796 4096
rect 55852 4136 55892 4145
rect 55852 3977 55892 4096
rect 55948 4136 55988 4145
rect 55948 4061 55988 4096
rect 55947 4052 55989 4061
rect 55947 4012 55948 4052
rect 55988 4012 55989 4052
rect 55947 4003 55989 4012
rect 55851 3968 55893 3977
rect 55851 3928 55852 3968
rect 55892 3928 55893 3968
rect 55851 3919 55893 3928
rect 55948 3641 55988 4003
rect 55947 3632 55989 3641
rect 55947 3592 55948 3632
rect 55988 3592 56084 3632
rect 55947 3583 55989 3592
rect 55947 3464 55989 3473
rect 55947 3424 55948 3464
rect 55988 3424 55989 3464
rect 55947 3415 55989 3424
rect 55948 3330 55988 3415
rect 55564 2860 55700 2900
rect 55468 2575 55508 2584
rect 55564 2624 55604 2633
rect 55276 2456 55316 2465
rect 53932 1903 53972 1912
rect 54795 1952 54837 1961
rect 54795 1912 54796 1952
rect 54836 1912 54837 1952
rect 54795 1903 54837 1912
rect 54796 1818 54836 1903
rect 53547 1364 53589 1373
rect 53547 1324 53548 1364
rect 53588 1324 53589 1364
rect 53547 1315 53589 1324
rect 55276 1112 55316 2416
rect 55564 2129 55604 2584
rect 55563 2120 55605 2129
rect 55563 2080 55564 2120
rect 55604 2080 55605 2120
rect 55563 2071 55605 2080
rect 55660 1961 55700 2860
rect 55755 2708 55797 2717
rect 55755 2668 55756 2708
rect 55796 2668 55797 2708
rect 55755 2659 55797 2668
rect 55756 2624 55796 2659
rect 55756 2573 55796 2584
rect 55947 2624 55989 2633
rect 55947 2584 55948 2624
rect 55988 2584 55989 2624
rect 55947 2575 55989 2584
rect 56044 2624 56084 3592
rect 56140 3380 56180 4759
rect 56235 4472 56277 4481
rect 56235 4432 56236 4472
rect 56276 4432 56277 4472
rect 56235 4423 56277 4432
rect 56236 4136 56276 4423
rect 56236 4087 56276 4096
rect 56524 4136 56564 4759
rect 56524 4087 56564 4096
rect 56619 4052 56661 4061
rect 56619 4012 56620 4052
rect 56660 4012 56661 4052
rect 56619 4003 56661 4012
rect 56620 3918 56660 4003
rect 56331 3548 56373 3557
rect 56331 3508 56332 3548
rect 56372 3508 56373 3548
rect 56331 3499 56373 3508
rect 56332 3414 56372 3499
rect 56716 3464 56756 4843
rect 57003 4472 57045 4481
rect 57003 4432 57004 4472
rect 57044 4432 57045 4472
rect 57003 4423 57045 4432
rect 56811 4388 56853 4397
rect 56811 4348 56812 4388
rect 56852 4348 56853 4388
rect 56811 4339 56853 4348
rect 56812 3548 56852 4339
rect 56812 3499 56852 3508
rect 56908 4304 56948 4313
rect 56140 3340 56276 3380
rect 56139 3212 56181 3221
rect 56139 3172 56140 3212
rect 56180 3172 56181 3212
rect 56139 3163 56181 3172
rect 56044 2575 56084 2584
rect 55948 2490 55988 2575
rect 55852 2456 55892 2465
rect 55756 2416 55852 2456
rect 56140 2456 56180 3163
rect 56236 2624 56276 3340
rect 56716 3221 56756 3424
rect 56908 3464 56948 4264
rect 56908 3415 56948 3424
rect 56715 3212 56757 3221
rect 56715 3172 56716 3212
rect 56756 3172 56757 3212
rect 56715 3163 56757 3172
rect 56812 2792 56852 2801
rect 56524 2752 56812 2792
rect 56236 2575 56276 2584
rect 56428 2624 56468 2633
rect 56331 2456 56373 2465
rect 56140 2416 56276 2456
rect 55659 1952 55701 1961
rect 55659 1912 55660 1952
rect 55700 1912 55701 1952
rect 55659 1903 55701 1912
rect 55563 1448 55605 1457
rect 55563 1408 55564 1448
rect 55604 1408 55605 1448
rect 55563 1399 55605 1408
rect 55371 1364 55413 1373
rect 55371 1324 55372 1364
rect 55412 1324 55413 1364
rect 55371 1315 55413 1324
rect 55372 1230 55412 1315
rect 55372 1112 55412 1121
rect 55276 1072 55372 1112
rect 55372 1063 55412 1072
rect 55564 1112 55604 1399
rect 55564 1063 55604 1072
rect 55660 1112 55700 1121
rect 55756 1112 55796 2416
rect 55852 2407 55892 2416
rect 55947 2120 55989 2129
rect 55947 2080 55948 2120
rect 55988 2080 55989 2120
rect 55947 2071 55989 2080
rect 55948 1986 55988 2071
rect 56140 1952 56180 1961
rect 56236 1952 56276 2416
rect 56331 2416 56332 2456
rect 56372 2416 56373 2456
rect 56331 2407 56373 2416
rect 56332 2322 56372 2407
rect 56332 1952 56372 1961
rect 56236 1912 56332 1952
rect 55948 1700 55988 1709
rect 55852 1660 55948 1700
rect 55852 1121 55892 1660
rect 55948 1651 55988 1660
rect 55948 1364 55988 1373
rect 56140 1364 56180 1912
rect 56332 1903 56372 1912
rect 56236 1700 56276 1709
rect 56428 1700 56468 2584
rect 56524 2624 56564 2752
rect 56812 2743 56852 2752
rect 56524 2575 56564 2584
rect 56715 2624 56757 2633
rect 56908 2624 56948 2633
rect 56715 2584 56716 2624
rect 56756 2584 56757 2624
rect 56715 2575 56757 2584
rect 56812 2584 56908 2624
rect 56619 2540 56661 2549
rect 56619 2500 56620 2540
rect 56660 2500 56661 2540
rect 56619 2491 56661 2500
rect 56523 2456 56565 2465
rect 56523 2416 56524 2456
rect 56564 2416 56565 2456
rect 56523 2407 56565 2416
rect 56524 2036 56564 2407
rect 56524 1987 56564 1996
rect 56276 1660 56468 1700
rect 56236 1457 56276 1660
rect 56331 1532 56373 1541
rect 56331 1492 56332 1532
rect 56372 1492 56373 1532
rect 56331 1483 56373 1492
rect 56235 1448 56277 1457
rect 56235 1408 56236 1448
rect 56276 1408 56277 1448
rect 56235 1399 56277 1408
rect 55988 1324 56180 1364
rect 55948 1315 55988 1324
rect 55700 1072 55796 1112
rect 55851 1112 55893 1121
rect 55851 1072 55852 1112
rect 55892 1072 55893 1112
rect 55660 1063 55700 1072
rect 55851 1063 55893 1072
rect 56235 1112 56277 1121
rect 56235 1072 56236 1112
rect 56276 1072 56277 1112
rect 56235 1063 56277 1072
rect 56332 1112 56372 1483
rect 56332 1063 56372 1072
rect 56620 1112 56660 2491
rect 56716 2490 56756 2575
rect 56812 2129 56852 2584
rect 56908 2575 56948 2584
rect 57004 2549 57044 4423
rect 57291 4388 57333 4397
rect 57291 4348 57292 4388
rect 57332 4348 57333 4388
rect 57291 4339 57333 4348
rect 57099 4136 57141 4145
rect 57099 4096 57100 4136
rect 57140 4096 57141 4136
rect 57099 4087 57141 4096
rect 57292 4136 57332 4339
rect 57964 4313 58004 4398
rect 57387 4304 57429 4313
rect 57387 4264 57388 4304
rect 57428 4264 57429 4304
rect 57387 4255 57429 4264
rect 57963 4304 58005 4313
rect 57963 4264 57964 4304
rect 58004 4264 58005 4304
rect 57963 4255 58005 4264
rect 57292 4087 57332 4096
rect 57388 4136 57428 4255
rect 57388 4087 57428 4096
rect 57964 4136 58004 4145
rect 58060 4136 58100 6019
rect 58155 5648 58197 5657
rect 58155 5608 58156 5648
rect 58196 5608 58197 5648
rect 58155 5599 58197 5608
rect 58004 4096 58100 4136
rect 58156 4136 58196 5599
rect 58539 4808 58581 4817
rect 58539 4768 58540 4808
rect 58580 4768 58581 4808
rect 58539 4759 58581 4768
rect 58540 4674 58580 4759
rect 58636 4313 58676 6448
rect 58732 6488 58772 6607
rect 58635 4304 58677 4313
rect 58635 4264 58636 4304
rect 58676 4264 58677 4304
rect 58635 4255 58677 4264
rect 57964 4087 58004 4096
rect 57100 4002 57140 4087
rect 57196 3968 57236 3977
rect 57196 3557 57236 3928
rect 57195 3548 57237 3557
rect 57195 3508 57196 3548
rect 57236 3508 57237 3548
rect 57195 3499 57237 3508
rect 57100 2792 57140 2801
rect 57003 2540 57045 2549
rect 57003 2500 57004 2540
rect 57044 2500 57045 2540
rect 57003 2491 57045 2500
rect 56811 2120 56853 2129
rect 56811 2080 56812 2120
rect 56852 2080 56853 2120
rect 56811 2071 56853 2080
rect 56812 1541 56852 2071
rect 56908 1952 56948 1961
rect 57100 1952 57140 2752
rect 57387 2708 57429 2717
rect 57387 2668 57388 2708
rect 57428 2668 57429 2708
rect 57387 2659 57429 2668
rect 57291 2624 57333 2633
rect 57291 2584 57292 2624
rect 57332 2584 57333 2624
rect 57291 2575 57333 2584
rect 56948 1912 57140 1952
rect 56908 1903 56948 1912
rect 56811 1532 56853 1541
rect 56811 1492 56812 1532
rect 56852 1492 56853 1532
rect 56811 1483 56853 1492
rect 56620 1063 56660 1072
rect 57195 1112 57237 1121
rect 57195 1072 57196 1112
rect 57236 1072 57237 1112
rect 57195 1063 57237 1072
rect 57292 1112 57332 2575
rect 57388 1112 57428 2659
rect 58156 2633 58196 4096
rect 58251 4136 58293 4145
rect 58251 4096 58252 4136
rect 58292 4096 58293 4136
rect 58251 4087 58293 4096
rect 58252 4002 58292 4087
rect 58155 2624 58197 2633
rect 58155 2584 58156 2624
rect 58196 2584 58197 2624
rect 58155 2575 58197 2584
rect 57771 1952 57813 1961
rect 57771 1912 57772 1952
rect 57812 1912 57813 1952
rect 57771 1903 57813 1912
rect 57772 1818 57812 1903
rect 57484 1289 57524 1374
rect 57483 1280 57525 1289
rect 57483 1240 57484 1280
rect 57524 1240 57525 1280
rect 57483 1231 57525 1240
rect 57484 1112 57524 1121
rect 57388 1072 57484 1112
rect 57292 1063 57332 1072
rect 57484 1063 57524 1072
rect 58636 1112 58676 4255
rect 58732 4229 58772 6448
rect 58827 6488 58869 6497
rect 58827 6448 58828 6488
rect 58868 6448 58869 6488
rect 58827 6439 58869 6448
rect 58828 6354 58868 6439
rect 58924 5657 58964 6616
rect 59020 6581 59060 7876
rect 59307 6992 59349 7001
rect 59212 6952 59308 6992
rect 59348 6952 59349 6992
rect 59019 6572 59061 6581
rect 59019 6532 59020 6572
rect 59060 6532 59061 6572
rect 59019 6523 59061 6532
rect 59020 6077 59060 6523
rect 59212 6497 59252 6952
rect 59307 6943 59349 6952
rect 59308 6858 59348 6943
rect 59500 6749 59540 8455
rect 59595 8000 59637 8009
rect 59595 7960 59596 8000
rect 59636 7960 59637 8000
rect 59595 7951 59637 7960
rect 59499 6740 59541 6749
rect 59499 6700 59500 6740
rect 59540 6700 59541 6740
rect 59499 6691 59541 6700
rect 59307 6656 59349 6665
rect 59307 6616 59308 6656
rect 59348 6616 59349 6656
rect 59307 6607 59349 6616
rect 59211 6488 59253 6497
rect 59211 6448 59212 6488
rect 59252 6448 59253 6488
rect 59211 6439 59253 6448
rect 59308 6488 59348 6607
rect 59499 6572 59541 6581
rect 59499 6532 59500 6572
rect 59540 6532 59541 6572
rect 59499 6523 59541 6532
rect 59308 6439 59348 6448
rect 59500 6488 59540 6523
rect 59212 6354 59252 6439
rect 59500 6437 59540 6448
rect 59500 6236 59540 6245
rect 59019 6068 59061 6077
rect 59019 6028 59020 6068
rect 59060 6028 59061 6068
rect 59019 6019 59061 6028
rect 58923 5648 58965 5657
rect 58923 5608 58924 5648
rect 58964 5608 58965 5648
rect 58923 5599 58965 5608
rect 59212 5648 59252 5657
rect 58923 5480 58965 5489
rect 58923 5440 58924 5480
rect 58964 5440 58965 5480
rect 58923 5431 58965 5440
rect 58924 5060 58964 5431
rect 58924 5011 58964 5020
rect 59212 4808 59252 5608
rect 59403 5648 59445 5657
rect 59403 5608 59404 5648
rect 59444 5608 59445 5648
rect 59403 5599 59445 5608
rect 59500 5648 59540 6196
rect 59500 5599 59540 5608
rect 59404 5514 59444 5599
rect 59307 5480 59349 5489
rect 59307 5440 59308 5480
rect 59348 5440 59349 5480
rect 59307 5431 59349 5440
rect 59308 5346 59348 5431
rect 59403 5396 59445 5405
rect 59403 5356 59404 5396
rect 59444 5356 59445 5396
rect 59403 5347 59445 5356
rect 59307 5228 59349 5237
rect 59307 5188 59308 5228
rect 59348 5188 59349 5228
rect 59307 5179 59349 5188
rect 59308 4976 59348 5179
rect 59308 4927 59348 4936
rect 59212 4768 59348 4808
rect 59211 4304 59253 4313
rect 59211 4264 59212 4304
rect 59252 4264 59253 4304
rect 59211 4255 59253 4264
rect 58731 4220 58773 4229
rect 58731 4180 58732 4220
rect 58772 4180 58773 4220
rect 58731 4171 58773 4180
rect 59115 4220 59157 4229
rect 59115 4180 59116 4220
rect 59156 4180 59157 4220
rect 59115 4171 59157 4180
rect 58732 3137 58772 4171
rect 59019 4136 59061 4145
rect 59019 4096 59020 4136
rect 59060 4096 59061 4136
rect 59019 4087 59061 4096
rect 59116 4136 59156 4171
rect 59020 4002 59060 4087
rect 59116 4085 59156 4096
rect 59212 4136 59252 4255
rect 59212 4087 59252 4096
rect 59308 4136 59348 4768
rect 59308 4087 59348 4096
rect 59404 3884 59444 5347
rect 59020 3844 59444 3884
rect 58827 3212 58869 3221
rect 58827 3172 58828 3212
rect 58868 3172 58869 3212
rect 58827 3163 58869 3172
rect 58731 3128 58773 3137
rect 58731 3088 58732 3128
rect 58772 3088 58773 3128
rect 58731 3079 58773 3088
rect 58636 1063 58676 1072
rect 58732 1112 58772 3079
rect 58828 2624 58868 3163
rect 58828 2575 58868 2584
rect 58923 2624 58965 2633
rect 58923 2584 58924 2624
rect 58964 2584 58965 2624
rect 59020 2624 59060 3844
rect 59499 3716 59541 3725
rect 59499 3676 59500 3716
rect 59540 3676 59541 3716
rect 59499 3667 59541 3676
rect 59307 3464 59349 3473
rect 59307 3424 59308 3464
rect 59348 3424 59349 3464
rect 59307 3415 59349 3424
rect 59500 3464 59540 3667
rect 59500 3415 59540 3424
rect 59308 3330 59348 3415
rect 59403 3212 59445 3221
rect 59403 3172 59404 3212
rect 59444 3172 59445 3212
rect 59403 3163 59445 3172
rect 59404 3078 59444 3163
rect 59403 2960 59445 2969
rect 59403 2920 59404 2960
rect 59444 2920 59445 2960
rect 59403 2911 59445 2920
rect 59115 2876 59157 2885
rect 59115 2836 59116 2876
rect 59156 2836 59157 2876
rect 59115 2827 59157 2836
rect 59116 2742 59156 2827
rect 59116 2624 59156 2633
rect 59020 2584 59116 2624
rect 58923 2575 58965 2584
rect 59116 2575 59156 2584
rect 59211 2624 59253 2633
rect 59211 2584 59212 2624
rect 59252 2584 59253 2624
rect 59211 2575 59253 2584
rect 59404 2624 59444 2911
rect 59404 2575 59444 2584
rect 58924 2490 58964 2575
rect 58827 2456 58869 2465
rect 58827 2416 58828 2456
rect 58868 2416 58869 2456
rect 58827 2407 58869 2416
rect 58732 1063 58772 1072
rect 58828 1112 58868 2407
rect 58923 2120 58965 2129
rect 58923 2080 58924 2120
rect 58964 2080 58965 2120
rect 58923 2071 58965 2080
rect 58924 1986 58964 2071
rect 59116 1952 59156 1961
rect 58923 1700 58965 1709
rect 58923 1660 58924 1700
rect 58964 1660 58965 1700
rect 58923 1651 58965 1660
rect 58924 1566 58964 1651
rect 59020 1364 59060 1373
rect 59116 1364 59156 1912
rect 59060 1324 59156 1364
rect 59020 1315 59060 1324
rect 59020 1112 59060 1121
rect 58828 1063 58868 1072
rect 58924 1072 59020 1112
rect 56236 978 56276 1063
rect 57196 978 57236 1063
rect 58540 944 58580 953
rect 58924 944 58964 1072
rect 59020 1063 59060 1072
rect 59212 1112 59252 2575
rect 59500 1952 59540 1961
rect 59500 1289 59540 1912
rect 59307 1280 59349 1289
rect 59307 1240 59308 1280
rect 59348 1240 59349 1280
rect 59307 1231 59349 1240
rect 59499 1280 59541 1289
rect 59499 1240 59500 1280
rect 59540 1240 59541 1280
rect 59499 1231 59541 1240
rect 59212 1063 59252 1072
rect 59308 1112 59348 1231
rect 59308 1063 59348 1072
rect 59596 1112 59636 7951
rect 59884 7916 59924 12940
rect 60076 11117 60116 16192
rect 60460 16232 60500 16241
rect 60652 16232 60692 16444
rect 60843 16435 60885 16444
rect 60844 16350 60884 16435
rect 61036 16400 61076 16409
rect 60940 16360 61036 16400
rect 60500 16192 60692 16232
rect 60747 16232 60789 16241
rect 60747 16192 60748 16232
rect 60788 16192 60789 16232
rect 60363 15476 60405 15485
rect 60363 15436 60364 15476
rect 60404 15436 60405 15476
rect 60363 15427 60405 15436
rect 60171 15392 60213 15401
rect 60171 15352 60172 15392
rect 60212 15352 60213 15392
rect 60171 15343 60213 15352
rect 60172 15258 60212 15343
rect 60364 15342 60404 15427
rect 60363 15224 60405 15233
rect 60363 15184 60364 15224
rect 60404 15184 60405 15224
rect 60363 15175 60405 15184
rect 60171 14888 60213 14897
rect 60171 14848 60172 14888
rect 60212 14848 60213 14888
rect 60171 14839 60213 14848
rect 60172 12980 60212 14839
rect 60364 14804 60404 15175
rect 60364 14755 60404 14764
rect 60172 12940 60308 12980
rect 60075 11108 60117 11117
rect 60075 11068 60076 11108
rect 60116 11068 60117 11108
rect 60075 11059 60117 11068
rect 59980 9512 60020 9521
rect 60020 9472 60116 9512
rect 59980 9463 60020 9472
rect 60076 8840 60116 9472
rect 60076 8791 60116 8800
rect 59884 7867 59924 7876
rect 60268 7916 60308 12940
rect 60460 10529 60500 16192
rect 60747 16183 60789 16192
rect 60556 15560 60596 15569
rect 60748 15560 60788 16183
rect 60556 14972 60596 15520
rect 60556 14923 60596 14932
rect 60652 15520 60788 15560
rect 60940 15560 60980 16360
rect 61036 16351 61076 16360
rect 61132 16241 61172 17116
rect 61255 17072 61295 17472
rect 61545 17156 61585 17472
rect 61228 17032 61295 17072
rect 61420 17116 61585 17156
rect 61228 16493 61268 17032
rect 61227 16484 61269 16493
rect 61227 16444 61228 16484
rect 61268 16444 61269 16484
rect 61227 16435 61269 16444
rect 61131 16232 61173 16241
rect 61131 16192 61132 16232
rect 61172 16192 61173 16232
rect 61131 16183 61173 16192
rect 61420 16232 61460 17116
rect 61655 17072 61695 17472
rect 61516 17032 61695 17072
rect 61516 16484 61556 17032
rect 61945 16988 61985 17472
rect 62055 17072 62095 17472
rect 62345 17072 62385 17472
rect 62055 17032 62228 17072
rect 61945 16948 62132 16988
rect 61516 16435 61556 16444
rect 61707 16316 61749 16325
rect 61707 16276 61708 16316
rect 61748 16276 61749 16316
rect 61707 16267 61749 16276
rect 61420 15560 61460 16192
rect 61708 16182 61748 16267
rect 62092 16232 62132 16948
rect 62188 16484 62228 17032
rect 62188 16435 62228 16444
rect 62284 17032 62385 17072
rect 62455 17072 62495 17472
rect 62745 17156 62785 17472
rect 62668 17116 62785 17156
rect 62455 17032 62516 17072
rect 61900 16064 61940 16073
rect 61803 15560 61845 15569
rect 61420 15520 61748 15560
rect 60555 14804 60597 14813
rect 60555 14764 60556 14804
rect 60596 14764 60597 14804
rect 60555 14755 60597 14764
rect 60556 14720 60596 14755
rect 60556 14669 60596 14680
rect 60555 14300 60597 14309
rect 60555 14260 60556 14300
rect 60596 14260 60597 14300
rect 60555 14251 60597 14260
rect 60556 14216 60596 14251
rect 60556 14165 60596 14176
rect 60555 13040 60597 13049
rect 60555 13000 60556 13040
rect 60596 13000 60597 13040
rect 60555 12991 60597 13000
rect 60556 11696 60596 12991
rect 60652 12980 60692 15520
rect 60940 15511 60980 15520
rect 60939 15392 60981 15401
rect 60939 15352 60940 15392
rect 60980 15352 60981 15392
rect 60939 15343 60981 15352
rect 60748 14720 60788 14729
rect 60748 13712 60788 14680
rect 60843 14720 60885 14729
rect 60843 14680 60844 14720
rect 60884 14680 60885 14720
rect 60843 14671 60885 14680
rect 60844 14586 60884 14671
rect 60844 13964 60884 13973
rect 60940 13964 60980 15343
rect 61419 14804 61461 14813
rect 61419 14764 61420 14804
rect 61460 14764 61461 14804
rect 61419 14755 61461 14764
rect 61132 14720 61172 14731
rect 61132 14645 61172 14680
rect 61420 14720 61460 14755
rect 61420 14669 61460 14680
rect 61131 14636 61173 14645
rect 61131 14596 61132 14636
rect 61172 14596 61173 14636
rect 61131 14587 61173 14596
rect 61516 14636 61556 14645
rect 61036 14216 61076 14225
rect 61132 14216 61172 14587
rect 61076 14176 61172 14216
rect 61036 14167 61076 14176
rect 60884 13924 60980 13964
rect 61228 14048 61268 14057
rect 60844 13915 60884 13924
rect 61036 13796 61076 13805
rect 60748 13672 60980 13712
rect 60940 13469 60980 13672
rect 60939 13460 60981 13469
rect 60939 13420 60940 13460
rect 60980 13420 60981 13460
rect 60939 13411 60981 13420
rect 60844 13208 60884 13217
rect 60652 12940 60788 12980
rect 60556 11647 60596 11656
rect 60459 10520 60501 10529
rect 60459 10480 60460 10520
rect 60500 10480 60501 10520
rect 60459 10471 60501 10480
rect 60459 10100 60501 10109
rect 60459 10060 60460 10100
rect 60500 10060 60501 10100
rect 60459 10051 60501 10060
rect 60460 8672 60500 10051
rect 60268 7867 60308 7876
rect 60364 8632 60460 8672
rect 59692 7748 59732 7757
rect 59692 7160 59732 7708
rect 60076 7748 60116 7757
rect 60076 7328 60116 7708
rect 60364 7328 60404 8632
rect 60460 8623 60500 8632
rect 60651 8672 60693 8681
rect 60651 8632 60652 8672
rect 60692 8632 60693 8672
rect 60651 8623 60693 8632
rect 60556 8588 60596 8597
rect 59884 7288 60116 7328
rect 60172 7288 60404 7328
rect 60460 8000 60500 8009
rect 59732 7120 59828 7160
rect 59692 7111 59732 7120
rect 59692 5816 59732 5825
rect 59692 5237 59732 5776
rect 59691 5228 59733 5237
rect 59691 5188 59692 5228
rect 59732 5188 59733 5228
rect 59691 5179 59733 5188
rect 59788 4229 59828 7120
rect 59884 5405 59924 7288
rect 59979 7160 60021 7169
rect 59979 7120 59980 7160
rect 60020 7120 60021 7160
rect 59979 7111 60021 7120
rect 59980 7026 60020 7111
rect 60075 7076 60117 7085
rect 60075 7036 60076 7076
rect 60116 7036 60117 7076
rect 60075 7027 60117 7036
rect 60076 6942 60116 7027
rect 60075 6740 60117 6749
rect 60075 6700 60076 6740
rect 60116 6700 60117 6740
rect 60075 6691 60117 6700
rect 59979 6656 60021 6665
rect 59979 6616 59980 6656
rect 60020 6616 60021 6656
rect 59979 6607 60021 6616
rect 59883 5396 59925 5405
rect 59883 5356 59884 5396
rect 59924 5356 59925 5396
rect 59883 5347 59925 5356
rect 59787 4220 59829 4229
rect 59787 4180 59788 4220
rect 59828 4180 59829 4220
rect 59787 4171 59829 4180
rect 59787 3716 59829 3725
rect 59787 3676 59788 3716
rect 59828 3676 59829 3716
rect 59787 3667 59829 3676
rect 59692 3464 59732 3473
rect 59692 2885 59732 3424
rect 59691 2876 59733 2885
rect 59691 2836 59692 2876
rect 59732 2836 59733 2876
rect 59691 2827 59733 2836
rect 59788 2708 59828 3667
rect 59980 3473 60020 6607
rect 60076 6488 60116 6691
rect 60172 6665 60212 7288
rect 60267 7160 60309 7169
rect 60267 7120 60268 7160
rect 60308 7120 60309 7160
rect 60267 7111 60309 7120
rect 60171 6656 60213 6665
rect 60171 6616 60172 6656
rect 60212 6616 60213 6656
rect 60171 6607 60213 6616
rect 60172 6488 60212 6497
rect 60076 6448 60172 6488
rect 60172 5153 60212 6448
rect 60268 6329 60308 7111
rect 60460 6992 60500 7960
rect 60556 7160 60596 8548
rect 60652 8538 60692 8623
rect 60748 8177 60788 12940
rect 60844 12713 60884 13168
rect 60940 13208 60980 13411
rect 60940 13159 60980 13168
rect 60843 12704 60885 12713
rect 60843 12664 60844 12704
rect 60884 12664 60885 12704
rect 60843 12655 60885 12664
rect 60939 11696 60981 11705
rect 60939 11656 60940 11696
rect 60980 11656 60981 11696
rect 60939 11647 60981 11656
rect 60940 11192 60980 11647
rect 61036 11537 61076 13756
rect 61132 13460 61172 13469
rect 61228 13460 61268 14008
rect 61516 13973 61556 14596
rect 61611 14048 61653 14057
rect 61611 14008 61612 14048
rect 61652 14008 61653 14048
rect 61611 13999 61653 14008
rect 61515 13964 61557 13973
rect 61515 13924 61516 13964
rect 61556 13924 61557 13964
rect 61515 13915 61557 13924
rect 61516 13796 61556 13915
rect 61612 13914 61652 13999
rect 61516 13756 61652 13796
rect 61172 13420 61268 13460
rect 61132 13411 61172 13420
rect 61419 13292 61461 13301
rect 61419 13252 61420 13292
rect 61460 13252 61461 13292
rect 61419 13243 61461 13252
rect 61516 13245 61556 13254
rect 61132 13208 61172 13217
rect 61324 13208 61364 13217
rect 61172 13168 61324 13208
rect 61132 13159 61172 13168
rect 61324 13159 61364 13168
rect 61420 13208 61460 13243
rect 61420 13157 61460 13168
rect 61516 13133 61556 13205
rect 61612 13208 61652 13756
rect 61612 13159 61652 13168
rect 61515 13124 61557 13133
rect 61515 13084 61516 13124
rect 61556 13084 61557 13124
rect 61515 13075 61557 13084
rect 61708 12980 61748 15520
rect 61803 15520 61804 15560
rect 61844 15520 61845 15560
rect 61803 15511 61845 15520
rect 61804 15426 61844 15511
rect 61900 14981 61940 16024
rect 61899 14972 61941 14981
rect 61899 14932 61900 14972
rect 61940 14932 61941 14972
rect 61899 14923 61941 14932
rect 61804 14888 61844 14897
rect 61804 13208 61844 14848
rect 61996 14561 62036 14646
rect 61995 14552 62037 14561
rect 61995 14512 61996 14552
rect 62036 14512 62037 14552
rect 61995 14503 62037 14512
rect 61995 14384 62037 14393
rect 61995 14344 61996 14384
rect 62036 14344 62037 14384
rect 61995 14335 62037 14344
rect 61899 13460 61941 13469
rect 61899 13420 61900 13460
rect 61940 13420 61941 13460
rect 61899 13411 61941 13420
rect 61900 13326 61940 13411
rect 61996 13208 62036 14335
rect 62092 14225 62132 16192
rect 62284 16232 62324 17032
rect 62476 16484 62516 17032
rect 62476 16435 62516 16444
rect 62668 16241 62708 17116
rect 62855 17072 62895 17472
rect 63145 17156 63185 17472
rect 62764 17032 62895 17072
rect 62956 17116 63185 17156
rect 62764 16484 62804 17032
rect 62764 16435 62804 16444
rect 62380 16232 62420 16241
rect 62284 16192 62380 16232
rect 62187 14972 62229 14981
rect 62187 14932 62188 14972
rect 62228 14932 62229 14972
rect 62187 14923 62229 14932
rect 62188 14804 62228 14923
rect 62188 14755 62228 14764
rect 62091 14216 62133 14225
rect 62091 14176 62092 14216
rect 62132 14176 62133 14216
rect 62091 14167 62133 14176
rect 62187 14048 62229 14057
rect 62187 14008 62188 14048
rect 62228 14008 62229 14048
rect 62187 13999 62229 14008
rect 62188 13418 62228 13999
rect 62188 13369 62228 13378
rect 61804 13159 61844 13168
rect 61900 13168 61996 13208
rect 61708 12940 61844 12980
rect 61707 12032 61749 12041
rect 61707 11992 61708 12032
rect 61748 11992 61749 12032
rect 61707 11983 61749 11992
rect 61708 11948 61748 11983
rect 61708 11897 61748 11908
rect 61035 11528 61077 11537
rect 61035 11488 61036 11528
rect 61076 11488 61077 11528
rect 61035 11479 61077 11488
rect 60940 11143 60980 11152
rect 61036 11033 61076 11479
rect 61035 11024 61077 11033
rect 61035 10984 61036 11024
rect 61076 10984 61077 11024
rect 61035 10975 61077 10984
rect 60843 9512 60885 9521
rect 60843 9472 60844 9512
rect 60884 9472 60885 9512
rect 60843 9463 60885 9472
rect 60844 9378 60884 9463
rect 60747 8168 60789 8177
rect 60747 8128 60748 8168
rect 60788 8128 60789 8168
rect 60747 8119 60789 8128
rect 60844 8000 60884 8009
rect 60844 7328 60884 7960
rect 61708 8000 61748 8009
rect 61036 7328 61076 7337
rect 60844 7288 61036 7328
rect 61036 7279 61076 7288
rect 60652 7169 60692 7254
rect 60556 7111 60596 7120
rect 60651 7160 60693 7169
rect 60651 7120 60652 7160
rect 60692 7120 60693 7160
rect 60651 7111 60693 7120
rect 60844 7160 60884 7169
rect 60748 6992 60788 7001
rect 60364 6950 60404 6959
rect 60460 6952 60748 6992
rect 60748 6943 60788 6952
rect 60364 6488 60404 6910
rect 60364 6439 60404 6448
rect 60267 6320 60309 6329
rect 60267 6280 60268 6320
rect 60308 6280 60309 6320
rect 60267 6271 60309 6280
rect 60268 6186 60308 6271
rect 60844 5648 60884 7120
rect 61419 6656 61461 6665
rect 61419 6616 61420 6656
rect 61460 6616 61461 6656
rect 61419 6607 61461 6616
rect 61420 6488 61460 6607
rect 61420 6439 61460 6448
rect 61612 6488 61652 6497
rect 61516 6236 61556 6245
rect 61132 6196 61516 6236
rect 61036 5657 61076 5742
rect 60844 5405 60884 5608
rect 61035 5648 61077 5657
rect 61035 5608 61036 5648
rect 61076 5608 61077 5648
rect 61035 5599 61077 5608
rect 61132 5648 61172 6196
rect 61516 6187 61556 6196
rect 61515 5900 61557 5909
rect 61612 5900 61652 6448
rect 61515 5860 61516 5900
rect 61556 5860 61652 5900
rect 61515 5851 61557 5860
rect 61132 5599 61172 5608
rect 61324 5564 61364 5573
rect 60940 5480 60980 5489
rect 61324 5480 61364 5524
rect 60980 5440 61364 5480
rect 60940 5431 60980 5440
rect 60843 5396 60885 5405
rect 61516 5396 61556 5851
rect 61708 5816 61748 7960
rect 61804 6161 61844 12940
rect 61900 11369 61940 13168
rect 61996 13159 62036 13168
rect 62284 12980 62324 16192
rect 62380 16183 62420 16192
rect 62667 16232 62709 16241
rect 62956 16232 62996 17116
rect 63255 17072 63295 17472
rect 63545 17156 63585 17472
rect 63052 17032 63295 17072
rect 63340 17116 63585 17156
rect 63052 16484 63092 17032
rect 63340 16988 63380 17116
rect 63655 17072 63695 17472
rect 63945 17156 63985 17472
rect 63244 16948 63380 16988
rect 63436 17032 63695 17072
rect 63916 17116 63985 17156
rect 63244 16568 63284 16948
rect 63244 16528 63367 16568
rect 63052 16435 63092 16444
rect 62667 16192 62668 16232
rect 62708 16192 62709 16232
rect 62667 16183 62709 16192
rect 62860 16192 62956 16232
rect 62668 16098 62708 16183
rect 62571 15644 62613 15653
rect 62571 15604 62572 15644
rect 62612 15604 62613 15644
rect 62571 15595 62613 15604
rect 62572 14813 62612 15595
rect 62571 14804 62613 14813
rect 62571 14764 62572 14804
rect 62612 14764 62613 14804
rect 62571 14755 62613 14764
rect 62380 14720 62420 14729
rect 62380 14561 62420 14680
rect 62475 14720 62517 14729
rect 62475 14680 62476 14720
rect 62516 14680 62517 14720
rect 62475 14671 62517 14680
rect 62572 14720 62612 14755
rect 62476 14586 62516 14671
rect 62572 14670 62612 14680
rect 62764 14561 62804 14646
rect 62379 14552 62421 14561
rect 62379 14512 62380 14552
rect 62420 14512 62421 14552
rect 62379 14503 62421 14512
rect 62763 14552 62805 14561
rect 62763 14512 62764 14552
rect 62804 14512 62805 14552
rect 62763 14503 62805 14512
rect 62380 14057 62420 14503
rect 62860 14384 62900 16192
rect 62956 16183 62996 16192
rect 63051 16232 63093 16241
rect 63051 16192 63052 16232
rect 63092 16192 63093 16232
rect 63051 16183 63093 16192
rect 63327 16221 63367 16528
rect 63436 16484 63476 17032
rect 63436 16435 63476 16444
rect 63916 16316 63956 17116
rect 64055 17072 64095 17472
rect 64345 17156 64385 17472
rect 62956 15737 62996 15822
rect 62955 15728 62997 15737
rect 62955 15688 62956 15728
rect 62996 15688 62997 15728
rect 62955 15679 62997 15688
rect 62955 14888 62997 14897
rect 62955 14848 62956 14888
rect 62996 14848 62997 14888
rect 62955 14839 62997 14848
rect 62956 14804 62996 14839
rect 62956 14753 62996 14764
rect 62572 14344 62900 14384
rect 62379 14048 62421 14057
rect 62379 14008 62380 14048
rect 62420 14008 62421 14048
rect 62379 13999 62421 14008
rect 62476 14048 62516 14057
rect 62380 13385 62420 13999
rect 62379 13376 62421 13385
rect 62379 13336 62380 13376
rect 62420 13336 62421 13376
rect 62379 13327 62421 13336
rect 62476 13049 62516 14008
rect 62475 13040 62517 13049
rect 62475 13000 62476 13040
rect 62516 13000 62517 13040
rect 62475 12991 62517 13000
rect 62284 12940 62420 12980
rect 62091 12704 62133 12713
rect 62091 12664 62092 12704
rect 62132 12664 62133 12704
rect 61996 12629 62036 12660
rect 62091 12655 62133 12664
rect 61995 12620 62037 12629
rect 61995 12580 61996 12620
rect 62036 12580 62037 12620
rect 61995 12571 62037 12580
rect 61996 12536 62036 12571
rect 62092 12570 62132 12655
rect 61899 11360 61941 11369
rect 61899 11320 61900 11360
rect 61940 11320 61941 11360
rect 61899 11311 61941 11320
rect 61996 11108 62036 12496
rect 62188 12536 62228 12547
rect 62188 12461 62228 12496
rect 62283 12536 62325 12545
rect 62283 12496 62284 12536
rect 62324 12496 62325 12536
rect 62283 12487 62325 12496
rect 62187 12452 62229 12461
rect 62187 12412 62188 12452
rect 62228 12412 62229 12452
rect 62187 12403 62229 12412
rect 62284 12402 62324 12487
rect 62092 11864 62132 11873
rect 62132 11824 62228 11864
rect 62092 11815 62132 11824
rect 61900 11068 62036 11108
rect 61900 10193 61940 11068
rect 62188 11033 62228 11824
rect 62092 11024 62132 11033
rect 61995 10268 62037 10277
rect 61995 10228 61996 10268
rect 62036 10228 62037 10268
rect 61995 10219 62037 10228
rect 61899 10184 61941 10193
rect 61899 10144 61900 10184
rect 61940 10144 61941 10184
rect 61899 10135 61941 10144
rect 61996 9680 62036 10219
rect 61996 9631 62036 9640
rect 62092 9521 62132 10984
rect 62187 11024 62229 11033
rect 62187 10984 62188 11024
rect 62228 10984 62229 11024
rect 62187 10975 62229 10984
rect 62380 10520 62420 12940
rect 62475 12116 62517 12125
rect 62475 12076 62476 12116
rect 62516 12076 62517 12116
rect 62475 12067 62517 12076
rect 62284 10480 62420 10520
rect 62187 9596 62229 9605
rect 62187 9556 62188 9596
rect 62228 9556 62229 9596
rect 62187 9547 62229 9556
rect 62091 9512 62133 9521
rect 62091 9472 62092 9512
rect 62132 9472 62133 9512
rect 62091 9463 62133 9472
rect 62188 9462 62228 9547
rect 61899 8672 61941 8681
rect 61899 8632 61900 8672
rect 61940 8632 61941 8672
rect 61899 8623 61941 8632
rect 61900 7085 61940 8623
rect 62187 7748 62229 7757
rect 62187 7708 62188 7748
rect 62228 7708 62229 7748
rect 62187 7699 62229 7708
rect 62188 7160 62228 7699
rect 62188 7111 62228 7120
rect 61899 7076 61941 7085
rect 61899 7036 61900 7076
rect 61940 7036 61941 7076
rect 61899 7027 61941 7036
rect 62284 6833 62324 10480
rect 62380 10352 62420 10361
rect 62380 9512 62420 10312
rect 62476 9773 62516 12067
rect 62572 11285 62612 14344
rect 62667 14216 62709 14225
rect 62667 14176 62668 14216
rect 62708 14176 62709 14216
rect 62667 14167 62709 14176
rect 62571 11276 62613 11285
rect 62571 11236 62572 11276
rect 62612 11236 62613 11276
rect 62571 11227 62613 11236
rect 62475 9764 62517 9773
rect 62475 9724 62476 9764
rect 62516 9724 62517 9764
rect 62475 9715 62517 9724
rect 62572 9512 62612 9521
rect 62380 9472 62572 9512
rect 62572 9463 62612 9472
rect 62668 7328 62708 14167
rect 62955 13292 62997 13301
rect 62955 13252 62956 13292
rect 62996 13252 62997 13292
rect 62955 13243 62997 13252
rect 62859 13124 62901 13133
rect 62859 13084 62860 13124
rect 62900 13084 62901 13124
rect 62859 13075 62901 13084
rect 62763 12536 62805 12545
rect 62763 12496 62764 12536
rect 62804 12496 62805 12536
rect 62763 12487 62805 12496
rect 62764 11705 62804 12487
rect 62763 11696 62805 11705
rect 62763 11656 62764 11696
rect 62804 11656 62805 11696
rect 62763 11647 62805 11656
rect 62860 11696 62900 13075
rect 62764 11562 62804 11647
rect 62860 11192 62900 11656
rect 62956 11696 62996 13243
rect 63052 12125 63092 16183
rect 63327 15896 63367 16181
rect 63724 16276 63956 16316
rect 64012 17032 64095 17072
rect 64300 17116 64385 17156
rect 63724 16232 63764 16276
rect 64012 16232 64052 17032
rect 63724 16073 63764 16192
rect 63820 16192 64052 16232
rect 64108 16232 64148 16241
rect 64300 16232 64340 17116
rect 64455 17072 64495 17472
rect 64587 17156 64629 17165
rect 64745 17156 64785 17472
rect 64855 17165 64895 17472
rect 64587 17116 64588 17156
rect 64628 17116 64629 17156
rect 64587 17107 64629 17116
rect 64684 17116 64785 17156
rect 64854 17156 64896 17165
rect 65145 17156 65185 17472
rect 64854 17116 64855 17156
rect 64895 17116 64896 17156
rect 64148 16192 64340 16232
rect 64396 17032 64495 17072
rect 63820 16148 63860 16192
rect 63820 16099 63860 16108
rect 63723 16064 63765 16073
rect 63723 16024 63724 16064
rect 63764 16024 63765 16064
rect 63723 16015 63765 16024
rect 63244 15856 63367 15896
rect 63244 13553 63284 15856
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 64108 15065 64148 16192
rect 64204 16064 64244 16073
rect 64396 16064 64436 17032
rect 64588 16484 64628 17107
rect 64684 16913 64724 17116
rect 64854 17107 64896 17116
rect 64972 17116 65185 17156
rect 64683 16904 64725 16913
rect 64683 16864 64684 16904
rect 64724 16864 64725 16904
rect 64683 16855 64725 16864
rect 64588 16435 64628 16444
rect 64492 16232 64532 16241
rect 64684 16232 64724 16855
rect 64972 16241 65012 17116
rect 65255 17072 65295 17472
rect 65545 17156 65585 17472
rect 65068 17032 65295 17072
rect 65356 17116 65585 17156
rect 65068 16484 65108 17032
rect 65356 16997 65396 17116
rect 65655 17072 65695 17472
rect 65945 17156 65985 17472
rect 65452 17032 65695 17072
rect 65740 17116 65985 17156
rect 65355 16988 65397 16997
rect 65355 16948 65356 16988
rect 65396 16948 65397 16988
rect 65355 16939 65397 16948
rect 65068 16435 65108 16444
rect 64532 16192 64724 16232
rect 64971 16232 65013 16241
rect 64971 16192 64972 16232
rect 65012 16192 65013 16232
rect 64492 16183 64532 16192
rect 64971 16183 65013 16192
rect 65356 16232 65396 16939
rect 65452 16484 65492 17032
rect 65452 16435 65492 16444
rect 65740 16409 65780 17116
rect 66055 17072 66095 17472
rect 66345 17156 66385 17472
rect 65836 17032 66095 17072
rect 66316 17116 66385 17156
rect 65836 16484 65876 17032
rect 65836 16435 65876 16444
rect 65739 16400 65781 16409
rect 65739 16360 65740 16400
rect 65780 16360 65781 16400
rect 65739 16351 65781 16360
rect 65356 16183 65396 16192
rect 65740 16232 65780 16351
rect 65740 16183 65780 16192
rect 66124 16232 66164 16241
rect 66316 16232 66356 17116
rect 66455 17072 66495 17472
rect 66603 17156 66645 17165
rect 66745 17156 66785 17472
rect 66855 17165 66895 17472
rect 66603 17116 66604 17156
rect 66644 17116 66645 17156
rect 66603 17107 66645 17116
rect 66700 17116 66785 17156
rect 66854 17156 66896 17165
rect 67145 17156 67185 17472
rect 66854 17116 66855 17156
rect 66895 17116 66896 17156
rect 66164 16192 66356 16232
rect 66412 17032 66495 17072
rect 64972 16098 65012 16183
rect 64244 16024 64436 16064
rect 64204 16015 64244 16024
rect 66124 15905 66164 16192
rect 66220 16064 66260 16073
rect 66412 16064 66452 17032
rect 66604 16484 66644 17107
rect 66604 16435 66644 16444
rect 66260 16024 66452 16064
rect 66508 16232 66548 16241
rect 66700 16232 66740 17116
rect 66854 17107 66896 17116
rect 66988 17116 67185 17156
rect 66988 16232 67028 17116
rect 67255 17072 67295 17472
rect 67545 17072 67585 17472
rect 67084 17032 67295 17072
rect 67372 17032 67585 17072
rect 67655 17072 67695 17472
rect 67945 17156 67985 17472
rect 67756 17116 67985 17156
rect 67655 17032 67700 17072
rect 67084 16484 67124 17032
rect 67084 16435 67124 16444
rect 67372 16232 67412 17032
rect 67468 16484 67508 16493
rect 67660 16484 67700 17032
rect 67508 16444 67700 16484
rect 67468 16435 67508 16444
rect 66548 16192 66740 16232
rect 66796 16192 66988 16232
rect 66220 16015 66260 16024
rect 66123 15896 66165 15905
rect 66123 15856 66124 15896
rect 66164 15856 66165 15896
rect 66123 15847 66165 15856
rect 64875 15812 64917 15821
rect 64875 15772 64876 15812
rect 64916 15772 64917 15812
rect 64875 15763 64917 15772
rect 64876 15560 64916 15763
rect 64588 15520 64876 15560
rect 64107 15056 64149 15065
rect 64107 15016 64108 15056
rect 64148 15016 64149 15056
rect 64107 15007 64149 15016
rect 64204 14888 64244 14897
rect 64012 14848 64204 14888
rect 63435 14804 63477 14813
rect 63435 14764 63436 14804
rect 63476 14764 63477 14804
rect 63435 14755 63477 14764
rect 63723 14804 63765 14813
rect 63723 14764 63724 14804
rect 63764 14764 63765 14804
rect 63723 14755 63765 14764
rect 63915 14804 63957 14813
rect 63915 14764 63916 14804
rect 63956 14764 63957 14804
rect 63915 14755 63957 14764
rect 63243 13544 63285 13553
rect 63243 13504 63244 13544
rect 63284 13504 63285 13544
rect 63243 13495 63285 13504
rect 63436 12980 63476 14755
rect 63724 14561 63764 14755
rect 63820 14720 63860 14729
rect 63723 14552 63765 14561
rect 63723 14512 63724 14552
rect 63764 14512 63765 14552
rect 63723 14503 63765 14512
rect 63820 14477 63860 14680
rect 63916 14670 63956 14755
rect 64012 14720 64052 14848
rect 64204 14839 64244 14848
rect 64299 14804 64341 14813
rect 64299 14764 64300 14804
rect 64340 14764 64341 14804
rect 64299 14755 64341 14764
rect 64012 14671 64052 14680
rect 63819 14468 63861 14477
rect 63819 14428 63820 14468
rect 63860 14428 63861 14468
rect 63819 14419 63861 14428
rect 63820 14048 63860 14059
rect 63820 13973 63860 14008
rect 63915 14048 63957 14057
rect 64108 14048 64148 14057
rect 63915 14008 63916 14048
rect 63956 14008 63957 14048
rect 63915 13999 63957 14008
rect 64012 14008 64108 14048
rect 63627 13964 63669 13973
rect 63627 13924 63628 13964
rect 63668 13924 63669 13964
rect 63627 13915 63669 13924
rect 63819 13964 63861 13973
rect 63819 13924 63820 13964
rect 63860 13924 63861 13964
rect 63819 13915 63861 13924
rect 63628 13830 63668 13915
rect 63916 13914 63956 13999
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 63436 12940 63956 12980
rect 63627 12788 63669 12797
rect 63627 12748 63628 12788
rect 63668 12748 63669 12788
rect 63627 12739 63669 12748
rect 63296 12536 63336 12545
rect 63296 12200 63336 12496
rect 63628 12536 63668 12739
rect 63628 12487 63668 12496
rect 63723 12536 63765 12545
rect 63723 12496 63724 12536
rect 63764 12496 63765 12536
rect 63723 12487 63765 12496
rect 63724 12402 63764 12487
rect 63916 12452 63956 12940
rect 64012 12629 64052 14008
rect 64108 13999 64148 14008
rect 64108 13796 64148 13805
rect 64108 13208 64148 13756
rect 64204 13208 64244 13217
rect 64108 13168 64204 13208
rect 64204 13159 64244 13168
rect 64300 13208 64340 14755
rect 64588 14720 64628 15520
rect 64876 15511 64916 15520
rect 65068 15560 65108 15569
rect 65452 15560 65492 15569
rect 65108 15520 65300 15560
rect 65068 15511 65108 15520
rect 64972 15308 65012 15317
rect 65012 15268 65204 15308
rect 64972 15259 65012 15268
rect 64588 14671 64628 14680
rect 64875 14720 64917 14729
rect 64875 14680 64876 14720
rect 64916 14680 64917 14720
rect 64875 14671 64917 14680
rect 65164 14720 65204 15268
rect 65260 14981 65300 15520
rect 65259 14972 65301 14981
rect 65452 14972 65492 15520
rect 65739 15560 65781 15569
rect 65739 15520 65740 15560
rect 65780 15520 65781 15560
rect 65739 15511 65781 15520
rect 65836 15560 65876 15569
rect 65259 14932 65260 14972
rect 65300 14932 65396 14972
rect 65259 14923 65301 14932
rect 65259 14804 65301 14813
rect 65259 14764 65260 14804
rect 65300 14764 65301 14804
rect 65259 14755 65301 14764
rect 65164 14671 65204 14680
rect 65260 14720 65300 14755
rect 64492 14636 64532 14645
rect 64492 14477 64532 14596
rect 64876 14586 64916 14671
rect 65260 14669 65300 14680
rect 64491 14468 64533 14477
rect 64491 14428 64492 14468
rect 64532 14428 64533 14468
rect 64491 14419 64533 14428
rect 65259 14468 65301 14477
rect 65259 14428 65260 14468
rect 65300 14428 65301 14468
rect 65259 14419 65301 14428
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 64395 14048 64437 14057
rect 64395 14008 64396 14048
rect 64436 14008 64437 14048
rect 64395 13999 64437 14008
rect 64588 14048 64628 14057
rect 64300 13159 64340 13168
rect 64396 13040 64436 13999
rect 64492 13460 64532 13469
rect 64588 13460 64628 14008
rect 64532 13420 64628 13460
rect 64972 14048 65012 14057
rect 64492 13411 64532 13420
rect 64972 13376 65012 14008
rect 65164 13376 65204 13385
rect 64972 13336 65164 13376
rect 65164 13327 65204 13336
rect 64779 13292 64821 13301
rect 64779 13252 64780 13292
rect 64820 13252 64821 13292
rect 64779 13243 64821 13252
rect 64492 13208 64532 13217
rect 64684 13208 64724 13217
rect 64532 13168 64684 13208
rect 64492 13159 64532 13168
rect 64684 13159 64724 13168
rect 64780 13208 64820 13243
rect 64780 13157 64820 13168
rect 64875 13208 64917 13217
rect 64875 13168 64876 13208
rect 64916 13168 64917 13208
rect 64875 13159 64917 13168
rect 64972 13208 65012 13217
rect 65260 13208 65300 14419
rect 65356 14393 65396 14932
rect 65452 14923 65492 14932
rect 65452 14720 65492 14729
rect 65452 14561 65492 14680
rect 65451 14552 65493 14561
rect 65451 14512 65452 14552
rect 65492 14512 65493 14552
rect 65451 14503 65493 14512
rect 65355 14384 65397 14393
rect 65355 14344 65356 14384
rect 65396 14344 65397 14384
rect 65355 14335 65397 14344
rect 65740 14048 65780 15511
rect 65836 14888 65876 15520
rect 66219 15476 66261 15485
rect 66219 15436 66220 15476
rect 66260 15436 66261 15476
rect 66219 15427 66261 15436
rect 65932 14888 65972 14897
rect 65836 14848 65932 14888
rect 65932 14839 65972 14848
rect 65836 14048 65876 14057
rect 65740 14008 65836 14048
rect 65876 14008 66068 14048
rect 65836 13999 65876 14008
rect 65012 13168 65300 13208
rect 64972 13159 65012 13168
rect 64876 13074 64916 13159
rect 64396 13000 64628 13040
rect 64395 12788 64437 12797
rect 64395 12748 64396 12788
rect 64436 12748 64437 12788
rect 64395 12739 64437 12748
rect 64011 12620 64053 12629
rect 64011 12580 64012 12620
rect 64052 12580 64053 12620
rect 64011 12571 64053 12580
rect 64396 12536 64436 12739
rect 64588 12545 64628 13000
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 64396 12487 64436 12496
rect 64587 12536 64629 12545
rect 64587 12496 64588 12536
rect 64628 12496 64629 12536
rect 64587 12487 64629 12496
rect 64780 12536 64820 12545
rect 63916 12412 64148 12452
rect 63244 12160 63336 12200
rect 64012 12284 64052 12293
rect 63051 12116 63093 12125
rect 63051 12076 63052 12116
rect 63092 12076 63093 12116
rect 63051 12067 63093 12076
rect 63244 11948 63284 12160
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 63244 11908 63380 11948
rect 63340 11705 63380 11908
rect 62956 11453 62996 11656
rect 63052 11696 63092 11705
rect 63244 11696 63284 11705
rect 63092 11656 63244 11696
rect 63052 11647 63092 11656
rect 63244 11647 63284 11656
rect 63339 11696 63381 11705
rect 63339 11656 63340 11696
rect 63380 11656 63381 11696
rect 63339 11647 63381 11656
rect 63436 11696 63476 11707
rect 63436 11621 63476 11656
rect 63532 11696 63572 11705
rect 63435 11612 63477 11621
rect 63435 11572 63436 11612
rect 63476 11572 63477 11612
rect 63435 11563 63477 11572
rect 63340 11528 63380 11537
rect 62955 11444 62997 11453
rect 62955 11404 62956 11444
rect 62996 11404 62997 11444
rect 62955 11395 62997 11404
rect 62860 11152 63092 11192
rect 62955 11024 62997 11033
rect 62955 10984 62956 11024
rect 62996 10984 62997 11024
rect 62955 10975 62997 10984
rect 62956 10890 62996 10975
rect 62859 9176 62901 9185
rect 62859 9136 62860 9176
rect 62900 9136 62901 9176
rect 62859 9127 62901 9136
rect 62860 8681 62900 9127
rect 63052 8681 63092 11152
rect 63340 11108 63380 11488
rect 63340 11059 63380 11068
rect 63532 10856 63572 11656
rect 63820 11696 63860 11705
rect 63820 11369 63860 11656
rect 63915 11696 63957 11705
rect 63915 11656 63916 11696
rect 63956 11656 63957 11696
rect 63915 11647 63957 11656
rect 64012 11696 64052 12244
rect 64108 11696 64148 12412
rect 64588 12402 64628 12487
rect 64492 12284 64532 12293
rect 64203 11948 64245 11957
rect 64203 11908 64204 11948
rect 64244 11908 64245 11948
rect 64203 11899 64245 11908
rect 64204 11814 64244 11899
rect 64204 11696 64244 11705
rect 64108 11656 64204 11696
rect 64012 11647 64052 11656
rect 64204 11647 64244 11656
rect 64395 11696 64437 11705
rect 64395 11656 64396 11696
rect 64436 11656 64437 11696
rect 64395 11647 64437 11656
rect 64492 11696 64532 12244
rect 64780 11957 64820 12496
rect 65164 12536 65204 12545
rect 64779 11948 64821 11957
rect 64779 11908 64780 11948
rect 64820 11908 64821 11948
rect 64779 11899 64821 11908
rect 65164 11864 65204 12496
rect 65547 12536 65589 12545
rect 65547 12496 65548 12536
rect 65588 12496 65589 12536
rect 65547 12487 65589 12496
rect 66028 12536 66068 14008
rect 66028 12487 66068 12496
rect 65260 11864 65300 11873
rect 65164 11824 65260 11864
rect 65260 11815 65300 11824
rect 64492 11647 64532 11656
rect 63916 11562 63956 11647
rect 64396 11562 64436 11647
rect 64011 11444 64053 11453
rect 64011 11404 64012 11444
rect 64052 11404 64053 11444
rect 64011 11395 64053 11404
rect 63819 11360 63861 11369
rect 63819 11320 63820 11360
rect 63860 11320 63861 11360
rect 63819 11311 63861 11320
rect 63820 11033 63860 11311
rect 63819 11024 63861 11033
rect 63819 10984 63820 11024
rect 63860 10984 63861 11024
rect 63819 10975 63861 10984
rect 63436 10816 63572 10856
rect 63436 10436 63476 10816
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 63436 10387 63476 10396
rect 63435 10184 63477 10193
rect 63628 10184 63668 10193
rect 63435 10144 63436 10184
rect 63476 10144 63572 10184
rect 63435 10135 63477 10144
rect 63436 10050 63476 10135
rect 63435 9512 63477 9521
rect 63435 9472 63436 9512
rect 63476 9472 63477 9512
rect 63435 9463 63477 9472
rect 63436 9378 63476 9463
rect 63532 9353 63572 10144
rect 63628 10109 63668 10144
rect 63724 10184 63764 10193
rect 63627 10100 63669 10109
rect 63627 10060 63628 10100
rect 63668 10060 63669 10100
rect 63627 10051 63669 10060
rect 63531 9344 63573 9353
rect 63531 9304 63532 9344
rect 63572 9304 63573 9344
rect 63531 9295 63573 9304
rect 63628 9269 63668 10051
rect 63724 10025 63764 10144
rect 63723 10016 63765 10025
rect 63723 9976 63724 10016
rect 63764 9976 63765 10016
rect 63723 9967 63765 9976
rect 63627 9260 63669 9269
rect 63627 9220 63628 9260
rect 63668 9220 63669 9260
rect 63627 9211 63669 9220
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 63819 8924 63861 8933
rect 63819 8884 63820 8924
rect 63860 8884 63861 8924
rect 63819 8875 63861 8884
rect 62859 8672 62901 8681
rect 62859 8632 62860 8672
rect 62900 8632 62901 8672
rect 62859 8623 62901 8632
rect 63051 8672 63093 8681
rect 63051 8632 63052 8672
rect 63092 8632 63093 8672
rect 63051 8623 63093 8632
rect 63820 8672 63860 8875
rect 63820 8623 63860 8632
rect 63915 8672 63957 8681
rect 63915 8632 63916 8672
rect 63956 8632 63957 8672
rect 63915 8623 63957 8632
rect 64012 8672 64052 11395
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 64492 11024 64532 11033
rect 64204 10436 64244 10445
rect 64492 10436 64532 10984
rect 64683 11024 64725 11033
rect 64876 11024 64916 11033
rect 64683 10984 64684 11024
rect 64724 10984 64725 11024
rect 64683 10975 64725 10984
rect 64780 10984 64876 11024
rect 64587 10940 64629 10949
rect 64587 10900 64588 10940
rect 64628 10900 64629 10940
rect 64587 10891 64629 10900
rect 64588 10806 64628 10891
rect 64684 10890 64724 10975
rect 64244 10396 64532 10436
rect 64204 10387 64244 10396
rect 64780 10352 64820 10984
rect 64876 10975 64916 10984
rect 65068 11024 65108 11034
rect 65068 10949 65108 10984
rect 65164 11024 65204 11033
rect 65204 10984 65396 11024
rect 65164 10975 65204 10984
rect 65067 10940 65109 10949
rect 65067 10900 65068 10940
rect 65108 10900 65109 10940
rect 65067 10891 65109 10900
rect 64875 10772 64917 10781
rect 64875 10732 64876 10772
rect 64916 10732 64917 10772
rect 64875 10723 64917 10732
rect 64876 10638 64916 10723
rect 64780 10312 65012 10352
rect 64587 10184 64629 10193
rect 64876 10184 64916 10193
rect 64587 10144 64588 10184
rect 64628 10144 64629 10184
rect 64587 10135 64629 10144
rect 64780 10144 64876 10184
rect 64492 10100 64532 10109
rect 64492 10025 64532 10060
rect 64588 10050 64628 10135
rect 64491 10016 64533 10025
rect 64780 10016 64820 10144
rect 64876 10135 64916 10144
rect 64972 10025 65012 10312
rect 64491 9976 64492 10016
rect 64532 9976 64533 10016
rect 64491 9967 64533 9976
rect 64684 9976 64820 10016
rect 64971 10016 65013 10025
rect 64971 9976 64972 10016
rect 65012 9976 65013 10016
rect 65068 10016 65108 10891
rect 65259 10772 65301 10781
rect 65259 10732 65260 10772
rect 65300 10732 65301 10772
rect 65259 10723 65301 10732
rect 65260 10184 65300 10723
rect 65260 10135 65300 10144
rect 65068 9976 65300 10016
rect 64107 9680 64149 9689
rect 64107 9640 64108 9680
rect 64148 9640 64149 9680
rect 64492 9680 64532 9967
rect 64588 9680 64628 9689
rect 64492 9640 64588 9680
rect 64107 9631 64149 9640
rect 64588 9631 64628 9640
rect 64012 8623 64052 8632
rect 64108 8672 64148 9631
rect 64299 9344 64341 9353
rect 64299 9304 64300 9344
rect 64340 9304 64341 9344
rect 64299 9295 64341 9304
rect 64108 8623 64148 8632
rect 64300 8672 64340 9295
rect 64588 9260 64628 9269
rect 64588 8933 64628 9220
rect 64587 8924 64629 8933
rect 64587 8884 64588 8924
rect 64628 8884 64629 8924
rect 64587 8875 64629 8884
rect 64491 8840 64533 8849
rect 64491 8800 64492 8840
rect 64532 8800 64533 8840
rect 64491 8791 64533 8800
rect 64300 8623 64340 8632
rect 64395 8672 64437 8681
rect 64395 8632 64396 8672
rect 64436 8632 64437 8672
rect 64395 8623 64437 8632
rect 64492 8672 64532 8791
rect 64492 8623 64532 8632
rect 64588 8672 64628 8681
rect 62860 8168 62900 8623
rect 63916 8538 63956 8623
rect 64396 8588 64436 8623
rect 64396 8537 64436 8548
rect 64108 8168 64148 8177
rect 62860 8119 62900 8128
rect 63628 8128 64108 8168
rect 63628 8000 63668 8128
rect 64108 8119 64148 8128
rect 64588 8009 64628 8632
rect 63628 7951 63668 7960
rect 63819 8000 63861 8009
rect 63819 7960 63820 8000
rect 63860 7960 63861 8000
rect 63819 7951 63861 7960
rect 63916 8000 63956 8009
rect 64204 8000 64244 8009
rect 63956 7960 64052 8000
rect 63916 7951 63956 7960
rect 63820 7866 63860 7951
rect 62476 7288 62708 7328
rect 63052 7832 63092 7841
rect 62283 6824 62325 6833
rect 62283 6784 62284 6824
rect 62324 6784 62325 6824
rect 62283 6775 62325 6784
rect 61803 6152 61845 6161
rect 61803 6112 61804 6152
rect 61844 6112 61845 6152
rect 61803 6103 61845 6112
rect 61612 5776 61748 5816
rect 61612 5657 61652 5776
rect 61611 5648 61653 5657
rect 61611 5608 61612 5648
rect 61652 5608 61653 5648
rect 61611 5599 61653 5608
rect 61708 5648 61748 5657
rect 61748 5608 61844 5648
rect 61708 5599 61748 5608
rect 60843 5356 60844 5396
rect 60884 5356 60885 5396
rect 60843 5347 60885 5356
rect 61132 5356 61556 5396
rect 60171 5144 60213 5153
rect 60171 5104 60172 5144
rect 60212 5104 60213 5144
rect 60171 5095 60213 5104
rect 60459 5144 60501 5153
rect 60459 5104 60460 5144
rect 60500 5104 60501 5144
rect 60459 5095 60501 5104
rect 60171 4976 60213 4985
rect 60171 4936 60172 4976
rect 60212 4936 60213 4976
rect 60171 4927 60213 4936
rect 60172 4842 60212 4927
rect 60172 4304 60212 4313
rect 59979 3464 60021 3473
rect 59979 3424 59980 3464
rect 60020 3424 60021 3464
rect 59979 3415 60021 3424
rect 60076 3464 60116 3473
rect 60172 3464 60212 4264
rect 60116 3424 60212 3464
rect 60076 3415 60116 3424
rect 59692 2668 59828 2708
rect 60076 2792 60116 2801
rect 59692 2624 59732 2668
rect 60076 2624 60116 2752
rect 60268 2624 60308 2633
rect 60076 2584 60268 2624
rect 59692 2575 59732 2584
rect 60268 2575 60308 2584
rect 60363 2624 60405 2633
rect 60363 2584 60364 2624
rect 60404 2584 60405 2624
rect 60363 2575 60405 2584
rect 60460 2624 60500 5095
rect 60844 4481 60884 5347
rect 60939 4976 60981 4985
rect 60939 4936 60940 4976
rect 60980 4936 60981 4976
rect 60939 4927 60981 4936
rect 60843 4472 60885 4481
rect 60843 4432 60844 4472
rect 60884 4432 60885 4472
rect 60843 4423 60885 4432
rect 60843 4220 60885 4229
rect 60843 4180 60844 4220
rect 60884 4180 60885 4220
rect 60843 4171 60885 4180
rect 60844 4136 60884 4171
rect 60844 3053 60884 4096
rect 60940 3464 60980 4927
rect 61132 4136 61172 5356
rect 61612 4985 61652 5599
rect 61611 4976 61653 4985
rect 61611 4936 61612 4976
rect 61652 4936 61653 4976
rect 61611 4927 61653 4936
rect 61804 4808 61844 5608
rect 62283 5564 62325 5573
rect 62283 5524 62284 5564
rect 62324 5524 62325 5564
rect 62283 5515 62325 5524
rect 62284 5060 62324 5515
rect 62379 5144 62421 5153
rect 62379 5104 62380 5144
rect 62420 5104 62421 5144
rect 62379 5095 62421 5104
rect 62284 5011 62324 5020
rect 61804 4759 61844 4768
rect 62188 4976 62228 4985
rect 61324 4724 61364 4733
rect 61132 4087 61172 4096
rect 61227 4136 61269 4145
rect 61324 4136 61364 4684
rect 62188 4397 62228 4936
rect 62380 4976 62420 5095
rect 62380 4649 62420 4936
rect 62379 4640 62421 4649
rect 62379 4600 62380 4640
rect 62420 4600 62421 4640
rect 62379 4591 62421 4600
rect 61515 4388 61557 4397
rect 61515 4348 61516 4388
rect 61556 4348 61557 4388
rect 61515 4339 61557 4348
rect 62187 4388 62229 4397
rect 62187 4348 62188 4388
rect 62228 4348 62229 4388
rect 62187 4339 62229 4348
rect 61516 4254 61556 4339
rect 61227 4096 61228 4136
rect 61268 4096 61364 4136
rect 61227 4087 61269 4096
rect 61228 4002 61268 4087
rect 62476 3893 62516 7288
rect 62572 7160 62612 7169
rect 63052 7160 63092 7792
rect 63628 7757 63668 7842
rect 63627 7748 63669 7757
rect 63627 7708 63628 7748
rect 63668 7708 63669 7748
rect 63627 7699 63669 7708
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 62612 7120 63092 7160
rect 63436 7160 63476 7169
rect 62572 7111 62612 7120
rect 63339 6320 63381 6329
rect 63244 6280 63340 6320
rect 63380 6280 63381 6320
rect 62571 5648 62613 5657
rect 62571 5608 62572 5648
rect 62612 5608 62613 5648
rect 62571 5599 62613 5608
rect 62955 5648 62997 5657
rect 62955 5608 62956 5648
rect 62996 5608 62997 5648
rect 62955 5599 62997 5608
rect 62572 5514 62612 5599
rect 62763 4304 62805 4313
rect 62763 4264 62764 4304
rect 62804 4264 62805 4304
rect 62763 4255 62805 4264
rect 62475 3884 62517 3893
rect 62475 3844 62476 3884
rect 62516 3844 62517 3884
rect 62475 3835 62517 3844
rect 62091 3716 62133 3725
rect 62091 3676 62092 3716
rect 62132 3676 62133 3716
rect 62091 3667 62133 3676
rect 62092 3632 62132 3667
rect 62092 3581 62132 3592
rect 60843 3044 60885 3053
rect 60843 3004 60844 3044
rect 60884 3004 60885 3044
rect 60843 2995 60885 3004
rect 60940 2900 60980 3424
rect 61803 3464 61845 3473
rect 61803 3424 61804 3464
rect 61844 3424 61845 3464
rect 61803 3415 61845 3424
rect 60460 2575 60500 2584
rect 60556 2860 60980 2900
rect 59788 2540 59828 2551
rect 59788 2465 59828 2500
rect 60364 2490 60404 2575
rect 59787 2456 59829 2465
rect 60556 2456 60596 2860
rect 59787 2416 59788 2456
rect 59828 2416 59829 2456
rect 59787 2407 59829 2416
rect 60460 2416 60596 2456
rect 61515 2456 61557 2465
rect 61515 2416 61516 2456
rect 61556 2416 61557 2456
rect 60364 1952 60404 1961
rect 60460 1952 60500 2416
rect 61515 2407 61557 2416
rect 61516 2120 61556 2407
rect 61516 2071 61556 2080
rect 60404 1912 60500 1952
rect 60364 1903 60404 1912
rect 60460 1196 60500 1912
rect 61708 1952 61748 1961
rect 61516 1700 61556 1709
rect 60747 1280 60789 1289
rect 60747 1240 60748 1280
rect 60788 1240 60789 1280
rect 60747 1231 60789 1240
rect 60460 1147 60500 1156
rect 60748 1146 60788 1231
rect 61516 1112 61556 1660
rect 61708 1373 61748 1912
rect 61707 1364 61749 1373
rect 61707 1324 61708 1364
rect 61748 1324 61749 1364
rect 61707 1315 61749 1324
rect 61708 1112 61748 1121
rect 61516 1072 61708 1112
rect 59596 1063 59636 1072
rect 61708 1063 61748 1072
rect 61804 1112 61844 3415
rect 62764 2900 62804 4255
rect 62860 4052 62900 4061
rect 62860 3641 62900 4012
rect 62859 3632 62901 3641
rect 62859 3592 62860 3632
rect 62900 3592 62901 3632
rect 62859 3583 62901 3592
rect 62764 2860 62900 2900
rect 62188 2792 62228 2801
rect 62092 2752 62188 2792
rect 62092 1952 62132 2752
rect 62188 2743 62228 2752
rect 62092 1903 62132 1912
rect 62571 1364 62613 1373
rect 62571 1324 62572 1364
rect 62612 1324 62613 1364
rect 62571 1315 62613 1324
rect 61996 1280 62036 1289
rect 62379 1280 62421 1289
rect 62036 1240 62324 1280
rect 61996 1231 62036 1240
rect 61804 1063 61844 1072
rect 61996 1112 62036 1123
rect 61996 1037 62036 1072
rect 62284 1112 62324 1240
rect 62379 1240 62380 1280
rect 62420 1240 62421 1280
rect 62379 1231 62421 1240
rect 62284 1063 62324 1072
rect 62380 1112 62420 1231
rect 62572 1230 62612 1315
rect 62380 1063 62420 1072
rect 62572 1112 62612 1121
rect 62764 1112 62804 1121
rect 62612 1072 62764 1112
rect 62572 1063 62612 1072
rect 62764 1063 62804 1072
rect 62860 1112 62900 2860
rect 62956 1952 62996 5599
rect 63147 5060 63189 5069
rect 63147 5020 63148 5060
rect 63188 5020 63189 5060
rect 63147 5011 63189 5020
rect 63148 4926 63188 5011
rect 63244 4976 63284 6280
rect 63339 6271 63381 6280
rect 63340 6252 63380 6271
rect 63436 5657 63476 7120
rect 64012 7085 64052 7960
rect 64011 7076 64053 7085
rect 64011 7036 64012 7076
rect 64052 7036 64053 7076
rect 64011 7027 64053 7036
rect 64011 6908 64053 6917
rect 64011 6868 64012 6908
rect 64052 6868 64053 6908
rect 64011 6859 64053 6868
rect 64012 6581 64052 6859
rect 64011 6572 64053 6581
rect 64011 6532 64012 6572
rect 64052 6532 64053 6572
rect 64011 6523 64053 6532
rect 63627 6320 63669 6329
rect 63627 6280 63628 6320
rect 63668 6280 63669 6320
rect 63627 6271 63669 6280
rect 63628 6186 63668 6271
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 63723 5900 63765 5909
rect 63723 5860 63724 5900
rect 63764 5860 63765 5900
rect 63723 5851 63765 5860
rect 63724 5732 63764 5851
rect 63724 5683 63764 5692
rect 63435 5648 63477 5657
rect 63435 5608 63436 5648
rect 63476 5608 63477 5648
rect 63435 5599 63477 5608
rect 63532 4976 63572 4985
rect 63244 4936 63532 4976
rect 63532 4927 63572 4936
rect 64012 4817 64052 6523
rect 64204 5741 64244 7960
rect 64300 8000 64340 8009
rect 64203 5732 64245 5741
rect 64203 5692 64204 5732
rect 64244 5692 64245 5732
rect 64203 5683 64245 5692
rect 64300 5237 64340 7960
rect 64395 8000 64437 8009
rect 64395 7960 64396 8000
rect 64436 7960 64437 8000
rect 64395 7951 64437 7960
rect 64587 8000 64629 8009
rect 64587 7960 64588 8000
rect 64628 7960 64629 8000
rect 64587 7951 64629 7960
rect 64684 8000 64724 9976
rect 64971 9967 65013 9976
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 64779 9680 64821 9689
rect 65260 9680 65300 9976
rect 64779 9640 64780 9680
rect 64820 9640 64821 9680
rect 64779 9631 64821 9640
rect 64972 9640 65300 9680
rect 64780 9512 64820 9631
rect 64875 9596 64917 9605
rect 64875 9556 64876 9596
rect 64916 9556 64917 9596
rect 64875 9547 64917 9556
rect 64780 9463 64820 9472
rect 64876 9462 64916 9547
rect 64972 9512 65012 9640
rect 65356 9596 65396 10984
rect 65451 10688 65493 10697
rect 65451 10648 65452 10688
rect 65492 10648 65493 10688
rect 65451 10639 65493 10648
rect 65452 10193 65492 10639
rect 65451 10184 65493 10193
rect 65451 10144 65452 10184
rect 65492 10144 65493 10184
rect 65451 10135 65493 10144
rect 65356 9547 65396 9556
rect 64972 9463 65012 9472
rect 65068 9512 65108 9521
rect 64779 9260 64821 9269
rect 64779 9220 64780 9260
rect 64820 9220 64821 9260
rect 64779 9211 64821 9220
rect 64780 8756 64820 9211
rect 64971 8840 65013 8849
rect 64971 8800 64972 8840
rect 65012 8800 65013 8840
rect 64971 8791 65013 8800
rect 64780 8707 64820 8716
rect 64972 8706 65012 8791
rect 65068 8681 65108 9472
rect 65260 9512 65300 9521
rect 65260 9344 65300 9472
rect 65452 9512 65492 10135
rect 65452 9463 65492 9472
rect 65548 9344 65588 12487
rect 66220 11873 66260 15427
rect 66508 14309 66548 16192
rect 66699 15560 66741 15569
rect 66699 15520 66700 15560
rect 66740 15520 66741 15560
rect 66699 15511 66741 15520
rect 66700 15426 66740 15511
rect 66507 14300 66549 14309
rect 66507 14260 66508 14300
rect 66548 14260 66549 14300
rect 66507 14251 66549 14260
rect 66796 12041 66836 16192
rect 66988 16183 67028 16192
rect 67084 16192 67372 16232
rect 66891 15980 66933 15989
rect 66891 15940 66892 15980
rect 66932 15940 66933 15980
rect 66891 15931 66933 15940
rect 66892 12980 66932 15931
rect 66987 14468 67029 14477
rect 66987 14428 66988 14468
rect 67028 14428 67029 14468
rect 66987 14419 67029 14428
rect 66988 14216 67028 14419
rect 66988 14167 67028 14176
rect 66892 12940 67028 12980
rect 66795 12032 66837 12041
rect 66795 11992 66796 12032
rect 66836 11992 66837 12032
rect 66795 11983 66837 11992
rect 66219 11864 66261 11873
rect 66219 11824 66220 11864
rect 66260 11824 66261 11864
rect 66219 11815 66261 11824
rect 65740 10856 65780 10865
rect 65644 10816 65740 10856
rect 65644 10184 65684 10816
rect 65740 10807 65780 10816
rect 65644 10135 65684 10144
rect 66508 10184 66548 10193
rect 65643 10016 65685 10025
rect 65643 9976 65644 10016
rect 65684 9976 65685 10016
rect 65643 9967 65685 9976
rect 65260 9304 65588 9344
rect 65067 8672 65109 8681
rect 65644 8672 65684 9967
rect 66508 9521 66548 10144
rect 66891 10100 66933 10109
rect 66891 10060 66892 10100
rect 66932 10060 66933 10100
rect 66891 10051 66933 10060
rect 66892 9596 66932 10051
rect 66892 9547 66932 9556
rect 66507 9512 66549 9521
rect 66507 9472 66508 9512
rect 66548 9472 66549 9512
rect 66507 9463 66549 9472
rect 66123 8840 66165 8849
rect 66123 8800 66124 8840
rect 66164 8800 66165 8840
rect 66123 8791 66165 8800
rect 65067 8632 65068 8672
rect 65108 8632 65109 8672
rect 65067 8623 65109 8632
rect 65548 8632 65684 8672
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 64971 8168 65013 8177
rect 64971 8128 64972 8168
rect 65012 8128 65013 8168
rect 64971 8119 65013 8128
rect 64396 7412 64436 7951
rect 64588 7412 64628 7421
rect 64396 7372 64588 7412
rect 64588 7363 64628 7372
rect 64684 7253 64724 7960
rect 64972 8000 65012 8119
rect 65259 8084 65301 8093
rect 65259 8044 65260 8084
rect 65300 8044 65301 8084
rect 65259 8035 65301 8044
rect 64972 7951 65012 7960
rect 65067 8000 65109 8009
rect 65067 7960 65068 8000
rect 65108 7960 65109 8000
rect 65067 7951 65109 7960
rect 65068 7866 65108 7951
rect 65260 7412 65300 8035
rect 65548 8000 65588 8632
rect 66028 8588 66068 8597
rect 65644 8548 66028 8588
rect 65644 8168 65684 8548
rect 66028 8539 66068 8548
rect 65644 8119 65684 8128
rect 65739 8084 65781 8093
rect 65739 8044 65740 8084
rect 65780 8044 65781 8084
rect 65739 8035 65781 8044
rect 65356 7748 65396 7757
rect 65396 7708 65492 7748
rect 65356 7699 65396 7708
rect 65356 7412 65396 7421
rect 65260 7372 65356 7412
rect 65356 7363 65396 7372
rect 64683 7244 64725 7253
rect 64683 7204 64684 7244
rect 64724 7204 64725 7244
rect 64683 7195 64725 7204
rect 64780 7160 64820 7169
rect 64780 7001 64820 7120
rect 64876 7085 64916 7170
rect 64972 7160 65012 7169
rect 64875 7076 64917 7085
rect 64875 7036 64876 7076
rect 64916 7036 64917 7076
rect 64875 7027 64917 7036
rect 64972 7001 65012 7120
rect 65067 7160 65109 7169
rect 65067 7120 65068 7160
rect 65108 7120 65109 7160
rect 65067 7111 65109 7120
rect 65260 7160 65300 7169
rect 64779 6992 64821 7001
rect 64779 6952 64780 6992
rect 64820 6952 64821 6992
rect 64779 6943 64821 6952
rect 64971 6992 65013 7001
rect 64971 6952 64972 6992
rect 65012 6952 65013 6992
rect 65068 6992 65108 7111
rect 65260 7076 65300 7120
rect 65452 7160 65492 7708
rect 65452 7111 65492 7120
rect 65355 7076 65397 7085
rect 65260 7036 65356 7076
rect 65396 7036 65397 7076
rect 65355 7027 65397 7036
rect 65068 6952 65300 6992
rect 64971 6943 65013 6952
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 65260 5984 65300 6952
rect 65260 5944 65396 5984
rect 64587 5816 64629 5825
rect 64587 5776 64588 5816
rect 64628 5776 64629 5816
rect 64587 5767 64629 5776
rect 65067 5816 65109 5825
rect 65067 5776 65068 5816
rect 65108 5776 65109 5816
rect 65067 5767 65109 5776
rect 64491 5732 64533 5741
rect 64491 5692 64492 5732
rect 64532 5692 64533 5732
rect 64491 5683 64533 5692
rect 64395 5648 64437 5657
rect 64395 5608 64396 5648
rect 64436 5608 64437 5648
rect 64395 5599 64437 5608
rect 64299 5228 64341 5237
rect 64299 5188 64300 5228
rect 64340 5188 64341 5228
rect 64299 5179 64341 5188
rect 64396 4976 64436 5599
rect 64108 4936 64396 4976
rect 64011 4808 64053 4817
rect 64011 4768 64012 4808
rect 64052 4768 64053 4808
rect 64011 4759 64053 4768
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 63435 4220 63477 4229
rect 63435 4180 63436 4220
rect 63476 4180 63477 4220
rect 63435 4171 63477 4180
rect 63244 4136 63284 4145
rect 63244 3716 63284 4096
rect 63244 3676 63380 3716
rect 63340 3338 63380 3676
rect 63340 3289 63380 3298
rect 63051 3128 63093 3137
rect 63051 3088 63052 3128
rect 63092 3088 63093 3128
rect 63051 3079 63093 3088
rect 62956 1903 62996 1912
rect 63052 1784 63092 3079
rect 62860 1063 62900 1072
rect 62956 1744 63092 1784
rect 62956 1112 62996 1744
rect 62956 1063 62996 1072
rect 63051 1112 63093 1121
rect 63051 1072 63052 1112
rect 63092 1072 63093 1112
rect 63436 1112 63476 4171
rect 64108 4136 64148 4936
rect 64396 4927 64436 4936
rect 64203 4808 64245 4817
rect 64492 4808 64532 5683
rect 64588 5648 64628 5767
rect 64588 5599 64628 5608
rect 64779 5648 64821 5657
rect 64779 5608 64780 5648
rect 64820 5608 64821 5648
rect 64779 5599 64821 5608
rect 64876 5648 64916 5657
rect 64780 5514 64820 5599
rect 64876 5489 64916 5608
rect 65068 5648 65108 5767
rect 65163 5732 65205 5741
rect 65163 5692 65164 5732
rect 65204 5692 65205 5732
rect 65163 5683 65205 5692
rect 65068 5599 65108 5608
rect 65164 5648 65204 5683
rect 65164 5597 65204 5608
rect 65260 5648 65300 5657
rect 64684 5480 64724 5489
rect 64684 5069 64724 5440
rect 64875 5480 64917 5489
rect 64875 5440 64876 5480
rect 64916 5440 64917 5480
rect 64875 5431 64917 5440
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 65260 5237 65300 5608
rect 65356 5648 65396 5944
rect 65548 5741 65588 7960
rect 65740 8000 65780 8035
rect 65740 7949 65780 7960
rect 65836 8000 65876 8009
rect 66028 8000 66068 8009
rect 66124 8000 66164 8791
rect 66508 8681 66548 9463
rect 66412 8672 66452 8681
rect 65836 7841 65876 7960
rect 65932 7960 66028 8000
rect 66068 7960 66164 8000
rect 66219 8000 66261 8009
rect 66219 7960 66220 8000
rect 66260 7960 66261 8000
rect 65835 7832 65877 7841
rect 65835 7792 65836 7832
rect 65876 7792 65877 7832
rect 65835 7783 65877 7792
rect 65739 7244 65781 7253
rect 65739 7204 65740 7244
rect 65780 7204 65781 7244
rect 65739 7195 65781 7204
rect 65740 6488 65780 7195
rect 65932 7001 65972 7960
rect 66028 7951 66068 7960
rect 66219 7951 66261 7960
rect 66220 7866 66260 7951
rect 66123 7832 66165 7841
rect 66123 7792 66124 7832
rect 66164 7792 66165 7832
rect 66412 7832 66452 8632
rect 66507 8672 66549 8681
rect 66507 8632 66508 8672
rect 66548 8632 66549 8672
rect 66507 8623 66549 8632
rect 66508 7832 66548 7841
rect 66412 7792 66508 7832
rect 66123 7783 66165 7792
rect 66508 7783 66548 7792
rect 66124 7698 66164 7783
rect 66123 7160 66165 7169
rect 66123 7120 66124 7160
rect 66164 7120 66165 7160
rect 66123 7111 66165 7120
rect 66220 7160 66260 7169
rect 65931 6992 65973 7001
rect 65931 6952 65932 6992
rect 65972 6952 65973 6992
rect 65931 6943 65973 6952
rect 65644 6448 65740 6488
rect 65547 5732 65589 5741
rect 65547 5692 65548 5732
rect 65588 5692 65589 5732
rect 65547 5683 65589 5692
rect 65259 5228 65301 5237
rect 65259 5188 65260 5228
rect 65300 5188 65301 5228
rect 65259 5179 65301 5188
rect 64683 5060 64725 5069
rect 64683 5020 64684 5060
rect 64724 5020 64725 5060
rect 64683 5011 64725 5020
rect 64203 4768 64204 4808
rect 64244 4768 64245 4808
rect 64203 4759 64245 4768
rect 64396 4768 64532 4808
rect 64108 4087 64148 4096
rect 64011 3632 64053 3641
rect 64011 3592 64012 3632
rect 64052 3592 64053 3632
rect 64011 3583 64053 3592
rect 64012 3498 64052 3583
rect 64108 3473 64148 3558
rect 63820 3464 63860 3473
rect 63820 3212 63860 3424
rect 63915 3464 63957 3473
rect 63915 3424 63916 3464
rect 63956 3424 63957 3464
rect 63915 3415 63957 3424
rect 64107 3464 64149 3473
rect 64107 3424 64108 3464
rect 64148 3424 64149 3464
rect 64107 3415 64149 3424
rect 63916 3330 63956 3415
rect 64204 3296 64244 4759
rect 64396 4313 64436 4768
rect 65260 4649 65300 5179
rect 65356 5144 65396 5608
rect 65548 5144 65588 5153
rect 65356 5104 65548 5144
rect 65548 5095 65588 5104
rect 64491 4640 64533 4649
rect 64491 4600 64492 4640
rect 64532 4600 64533 4640
rect 64491 4591 64533 4600
rect 65259 4640 65301 4649
rect 65259 4600 65260 4640
rect 65300 4600 65301 4640
rect 65259 4591 65301 4600
rect 64395 4304 64437 4313
rect 64395 4264 64396 4304
rect 64436 4264 64437 4304
rect 64395 4255 64437 4264
rect 64299 3464 64341 3473
rect 64299 3424 64300 3464
rect 64340 3424 64341 3464
rect 64299 3415 64341 3424
rect 64396 3464 64436 4255
rect 64396 3415 64436 3424
rect 64492 3464 64532 4591
rect 64683 4556 64725 4565
rect 64683 4516 64684 4556
rect 64724 4516 64725 4556
rect 64683 4507 64725 4516
rect 64300 3330 64340 3415
rect 64108 3256 64244 3296
rect 63820 3172 64052 3212
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 64012 2876 64052 3172
rect 64012 2827 64052 2836
rect 63724 2624 63764 2633
rect 63724 2120 63764 2584
rect 63819 2624 63861 2633
rect 63819 2584 63820 2624
rect 63860 2584 63861 2624
rect 63819 2575 63861 2584
rect 64012 2624 64052 2633
rect 64108 2624 64148 3256
rect 64492 3137 64532 3424
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 64588 3330 64628 3415
rect 64491 3128 64533 3137
rect 64491 3088 64492 3128
rect 64532 3088 64533 3128
rect 64491 3079 64533 3088
rect 64684 3053 64724 4507
rect 65644 4229 65684 6448
rect 65740 6439 65780 6448
rect 65835 5480 65877 5489
rect 65835 5440 65836 5480
rect 65876 5440 65877 5480
rect 65835 5431 65877 5440
rect 65836 5144 65876 5431
rect 65836 5095 65876 5104
rect 65932 4985 65972 6943
rect 66124 6572 66164 7111
rect 66220 7085 66260 7120
rect 66412 7160 66452 7169
rect 66219 7076 66261 7085
rect 66219 7036 66220 7076
rect 66260 7036 66261 7076
rect 66219 7027 66261 7036
rect 66316 7076 66356 7085
rect 66124 6523 66164 6532
rect 66027 6488 66069 6497
rect 66027 6448 66028 6488
rect 66068 6448 66069 6488
rect 66027 6439 66069 6448
rect 66028 6354 66068 6439
rect 66123 5732 66165 5741
rect 66123 5692 66124 5732
rect 66164 5692 66165 5732
rect 66123 5683 66165 5692
rect 65740 4976 65780 4985
rect 65740 4817 65780 4936
rect 65931 4976 65973 4985
rect 65931 4936 65932 4976
rect 65972 4936 65973 4976
rect 65931 4927 65973 4936
rect 66028 4976 66068 4985
rect 65932 4842 65972 4927
rect 65739 4808 65781 4817
rect 65739 4768 65740 4808
rect 65780 4768 65781 4808
rect 65739 4759 65781 4768
rect 65835 4304 65877 4313
rect 65835 4264 65836 4304
rect 65876 4264 65877 4304
rect 65835 4255 65877 4264
rect 65643 4220 65685 4229
rect 65643 4180 65644 4220
rect 65684 4180 65685 4220
rect 65643 4171 65685 4180
rect 65548 4136 65588 4145
rect 65260 4061 65300 4092
rect 65259 4052 65301 4061
rect 65259 4012 65260 4052
rect 65300 4012 65301 4052
rect 65548 4052 65588 4096
rect 65644 4052 65684 4171
rect 65836 4136 65876 4255
rect 65836 4087 65876 4096
rect 65548 4012 65684 4052
rect 65931 4052 65973 4061
rect 66028 4052 66068 4936
rect 66124 4481 66164 5683
rect 66220 4976 66260 7027
rect 66316 5657 66356 7036
rect 66412 6320 66452 7120
rect 66700 7160 66740 7169
rect 66700 7001 66740 7120
rect 66892 7160 66932 7171
rect 66892 7085 66932 7120
rect 66796 7076 66836 7085
rect 66699 6992 66741 7001
rect 66699 6952 66700 6992
rect 66740 6952 66741 6992
rect 66699 6943 66741 6952
rect 66700 6488 66740 6497
rect 66412 6271 66452 6280
rect 66508 6448 66700 6488
rect 66412 5900 66452 5909
rect 66508 5900 66548 6448
rect 66700 6439 66740 6448
rect 66452 5860 66548 5900
rect 66412 5851 66452 5860
rect 66411 5732 66453 5741
rect 66411 5692 66412 5732
rect 66452 5692 66453 5732
rect 66411 5683 66453 5692
rect 66315 5648 66357 5657
rect 66315 5608 66316 5648
rect 66356 5608 66357 5648
rect 66315 5599 66357 5608
rect 66412 5648 66452 5683
rect 66412 5597 66452 5608
rect 66603 5648 66645 5657
rect 66603 5608 66604 5648
rect 66644 5608 66645 5648
rect 66603 5599 66645 5608
rect 66700 5648 66740 5657
rect 66796 5648 66836 7036
rect 66891 7076 66933 7085
rect 66891 7036 66892 7076
rect 66932 7036 66933 7076
rect 66891 7027 66933 7036
rect 66892 6497 66932 7027
rect 66891 6488 66933 6497
rect 66891 6448 66892 6488
rect 66932 6448 66933 6488
rect 66891 6439 66933 6448
rect 66740 5608 66836 5648
rect 66700 5599 66740 5608
rect 66604 5514 66644 5599
rect 66316 5104 66548 5144
rect 66316 5060 66356 5104
rect 66316 5011 66356 5020
rect 66220 4565 66260 4936
rect 66412 4976 66452 4985
rect 66219 4556 66261 4565
rect 66219 4516 66220 4556
rect 66260 4516 66261 4556
rect 66219 4507 66261 4516
rect 66123 4472 66165 4481
rect 66123 4432 66124 4472
rect 66164 4432 66165 4472
rect 66123 4423 66165 4432
rect 65931 4012 65932 4052
rect 65972 4012 66068 4052
rect 65259 4003 65301 4012
rect 65931 4003 65973 4012
rect 65260 3968 65300 4003
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 65260 3473 65300 3928
rect 65932 3918 65972 4003
rect 65259 3464 65301 3473
rect 65259 3424 65260 3464
rect 65300 3424 65301 3464
rect 65259 3415 65301 3424
rect 66124 3464 66164 4423
rect 66220 4388 66260 4397
rect 66412 4388 66452 4936
rect 66260 4348 66452 4388
rect 66220 4339 66260 4348
rect 66412 4052 66452 4061
rect 66220 4012 66412 4052
rect 66220 3632 66260 4012
rect 66412 4003 66452 4012
rect 66220 3583 66260 3592
rect 66508 3557 66548 5104
rect 66603 4976 66645 4985
rect 66603 4936 66604 4976
rect 66644 4936 66645 4976
rect 66603 4927 66645 4936
rect 66315 3548 66357 3557
rect 66315 3508 66316 3548
rect 66356 3508 66357 3548
rect 66315 3499 66357 3508
rect 66507 3548 66549 3557
rect 66507 3508 66508 3548
rect 66548 3508 66549 3548
rect 66507 3499 66549 3508
rect 64779 3380 64821 3389
rect 64779 3340 64780 3380
rect 64820 3340 64821 3380
rect 64779 3331 64821 3340
rect 64683 3044 64725 3053
rect 64683 3004 64684 3044
rect 64724 3004 64725 3044
rect 64683 2995 64725 3004
rect 64203 2960 64245 2969
rect 64203 2920 64204 2960
rect 64244 2920 64245 2960
rect 64203 2911 64245 2920
rect 64052 2584 64148 2624
rect 64204 2624 64244 2911
rect 64780 2900 64820 3331
rect 66124 2969 66164 3424
rect 66316 3464 66356 3499
rect 66604 3473 66644 4927
rect 66892 4808 66932 4817
rect 66796 4768 66892 4808
rect 66796 4136 66836 4768
rect 66892 4759 66932 4768
rect 66891 4304 66933 4313
rect 66891 4264 66892 4304
rect 66932 4264 66933 4304
rect 66891 4255 66933 4264
rect 66796 4087 66836 4096
rect 66316 3413 66356 3424
rect 66412 3464 66452 3473
rect 66412 3296 66452 3424
rect 66603 3464 66645 3473
rect 66603 3424 66604 3464
rect 66644 3424 66645 3464
rect 66603 3415 66645 3424
rect 66796 3464 66836 3473
rect 66892 3464 66932 4255
rect 66988 3725 67028 12940
rect 67084 10277 67124 16192
rect 67372 16183 67412 16192
rect 67756 16232 67796 17116
rect 68055 17072 68095 17472
rect 68345 17156 68385 17472
rect 67852 17032 68095 17072
rect 68140 17116 68385 17156
rect 67852 16484 67892 17032
rect 67852 16435 67892 16444
rect 67659 16148 67701 16157
rect 67659 16108 67660 16148
rect 67700 16108 67701 16148
rect 67659 16099 67701 16108
rect 67179 14804 67221 14813
rect 67179 14764 67180 14804
rect 67220 14764 67221 14804
rect 67179 14755 67221 14764
rect 67180 14670 67220 14755
rect 67564 14636 67604 14645
rect 67372 14552 67412 14561
rect 67412 14512 67508 14552
rect 67372 14503 67412 14512
rect 67275 14468 67317 14477
rect 67275 14428 67276 14468
rect 67316 14428 67317 14468
rect 67275 14419 67317 14428
rect 67276 14048 67316 14419
rect 67468 14300 67508 14512
rect 67564 14477 67604 14596
rect 67563 14468 67605 14477
rect 67563 14428 67564 14468
rect 67604 14428 67605 14468
rect 67563 14419 67605 14428
rect 67468 14260 67604 14300
rect 67467 14132 67509 14141
rect 67467 14092 67468 14132
rect 67508 14092 67509 14132
rect 67467 14083 67509 14092
rect 67276 13999 67316 14008
rect 67371 14048 67413 14057
rect 67371 14008 67372 14048
rect 67412 14008 67413 14048
rect 67371 13999 67413 14008
rect 67372 13914 67412 13999
rect 67468 13998 67508 14083
rect 67564 14048 67604 14260
rect 67275 13796 67317 13805
rect 67275 13756 67276 13796
rect 67316 13756 67317 13796
rect 67275 13747 67317 13756
rect 67179 12788 67221 12797
rect 67179 12748 67180 12788
rect 67220 12748 67221 12788
rect 67179 12739 67221 12748
rect 67180 12704 67220 12739
rect 67180 12653 67220 12664
rect 67276 10520 67316 13747
rect 67564 13301 67604 14008
rect 67660 13805 67700 16099
rect 67659 13796 67701 13805
rect 67659 13756 67660 13796
rect 67700 13756 67701 13796
rect 67659 13747 67701 13756
rect 67563 13292 67605 13301
rect 67563 13252 67564 13292
rect 67604 13252 67605 13292
rect 67563 13243 67605 13252
rect 67756 12980 67796 16192
rect 68140 16232 68180 17116
rect 68455 17072 68495 17472
rect 68745 17156 68785 17472
rect 68236 17032 68495 17072
rect 68716 17116 68785 17156
rect 68236 16484 68276 17032
rect 68236 16435 68276 16444
rect 67947 15896 67989 15905
rect 67947 15856 67948 15896
rect 67988 15856 67989 15896
rect 67947 15847 67989 15856
rect 67851 15812 67893 15821
rect 67851 15772 67852 15812
rect 67892 15772 67893 15812
rect 67851 15763 67893 15772
rect 67852 15728 67892 15763
rect 67852 15677 67892 15688
rect 67948 15140 67988 15847
rect 67852 15100 67988 15140
rect 68044 15392 68084 15401
rect 67852 13721 67892 15100
rect 67948 14720 67988 14729
rect 68044 14720 68084 15352
rect 67988 14680 68084 14720
rect 67948 14671 67988 14680
rect 68140 14552 68180 16192
rect 68235 16232 68277 16241
rect 68235 16192 68236 16232
rect 68276 16192 68277 16232
rect 68235 16183 68277 16192
rect 68524 16232 68564 16241
rect 68716 16232 68756 17116
rect 68855 17072 68895 17472
rect 69145 17240 69185 17472
rect 69255 17324 69295 17472
rect 69255 17284 69332 17324
rect 68564 16192 68756 16232
rect 68812 17032 68895 17072
rect 69004 17200 69185 17240
rect 67948 14512 68180 14552
rect 67851 13712 67893 13721
rect 67851 13672 67852 13712
rect 67892 13672 67893 13712
rect 67851 13663 67893 13672
rect 67756 12940 67892 12980
rect 67372 12536 67412 12545
rect 67756 12536 67796 12545
rect 67372 11957 67412 12496
rect 67468 12496 67756 12536
rect 67371 11948 67413 11957
rect 67371 11908 67372 11948
rect 67412 11908 67413 11948
rect 67371 11899 67413 11908
rect 67468 11864 67508 12496
rect 67756 12487 67796 12496
rect 67468 11815 67508 11824
rect 67852 10772 67892 12940
rect 67756 10732 67892 10772
rect 67659 10688 67701 10697
rect 67659 10648 67660 10688
rect 67700 10648 67701 10688
rect 67659 10639 67701 10648
rect 67276 10480 67412 10520
rect 67275 10352 67317 10361
rect 67275 10312 67276 10352
rect 67316 10312 67317 10352
rect 67275 10303 67317 10312
rect 67083 10268 67125 10277
rect 67083 10228 67084 10268
rect 67124 10228 67125 10268
rect 67083 10219 67125 10228
rect 67276 9512 67316 10303
rect 67276 9463 67316 9472
rect 67275 8672 67317 8681
rect 67275 8632 67276 8672
rect 67316 8632 67317 8672
rect 67275 8623 67317 8632
rect 67276 8538 67316 8623
rect 67084 6488 67124 6497
rect 67084 5816 67124 6448
rect 67180 5816 67220 5825
rect 67084 5776 67180 5816
rect 67180 5767 67220 5776
rect 66987 3716 67029 3725
rect 66987 3676 66988 3716
rect 67028 3676 67029 3716
rect 66987 3667 67029 3676
rect 66836 3424 66932 3464
rect 66796 3415 66836 3424
rect 66700 3296 66740 3305
rect 66412 3256 66700 3296
rect 66700 3247 66740 3256
rect 66123 2960 66165 2969
rect 66123 2920 66124 2960
rect 66164 2920 66165 2960
rect 66123 2911 66165 2920
rect 63820 2490 63860 2575
rect 64012 2288 64052 2584
rect 64204 2575 64244 2584
rect 64396 2836 64628 2876
rect 64396 2624 64436 2836
rect 64491 2708 64533 2717
rect 64491 2668 64492 2708
rect 64532 2668 64533 2708
rect 64491 2659 64533 2668
rect 64396 2575 64436 2584
rect 64492 2624 64532 2659
rect 64492 2573 64532 2584
rect 64300 2456 64340 2465
rect 64340 2416 64436 2456
rect 64300 2407 64340 2416
rect 64012 2248 64244 2288
rect 64108 2120 64148 2129
rect 63724 2080 64108 2120
rect 64108 2071 64148 2080
rect 64108 1700 64148 1709
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 64011 1364 64053 1373
rect 64011 1324 64012 1364
rect 64052 1324 64053 1364
rect 64011 1315 64053 1324
rect 63724 1112 63764 1121
rect 63436 1072 63724 1112
rect 63051 1063 63093 1072
rect 63724 1063 63764 1072
rect 64012 1112 64052 1315
rect 64108 1121 64148 1660
rect 64012 1063 64052 1072
rect 64107 1112 64149 1121
rect 64107 1072 64108 1112
rect 64148 1072 64149 1112
rect 64107 1063 64149 1072
rect 61995 1028 62037 1037
rect 61995 988 61996 1028
rect 62036 988 62037 1028
rect 61995 979 62037 988
rect 63052 978 63092 1063
rect 64108 978 64148 1063
rect 64204 1037 64244 2248
rect 64396 1952 64436 2416
rect 64492 1952 64532 1961
rect 64396 1912 64492 1952
rect 64588 1952 64628 2836
rect 64684 2860 64820 2900
rect 67372 2900 67412 10480
rect 67660 10436 67700 10639
rect 67660 10387 67700 10396
rect 67659 10268 67701 10277
rect 67659 10228 67660 10268
rect 67700 10228 67701 10268
rect 67659 10219 67701 10228
rect 67660 4901 67700 10219
rect 67756 9185 67796 10732
rect 67851 10352 67893 10361
rect 67851 10312 67852 10352
rect 67892 10312 67893 10352
rect 67851 10303 67893 10312
rect 67852 10218 67892 10303
rect 67755 9176 67797 9185
rect 67755 9136 67756 9176
rect 67796 9136 67797 9176
rect 67755 9127 67797 9136
rect 67948 7328 67988 14512
rect 68139 14216 68181 14225
rect 68139 14176 68140 14216
rect 68180 14176 68181 14216
rect 68139 14167 68181 14176
rect 68043 14132 68085 14141
rect 68043 14092 68044 14132
rect 68084 14092 68085 14132
rect 68043 14083 68085 14092
rect 68044 14048 68084 14083
rect 68044 13997 68084 14008
rect 68140 14048 68180 14167
rect 68140 13999 68180 14008
rect 68236 13880 68276 16183
rect 68524 16073 68564 16192
rect 68523 16064 68565 16073
rect 68523 16024 68524 16064
rect 68564 16024 68565 16064
rect 68523 16015 68565 16024
rect 68620 16064 68660 16073
rect 68812 16064 68852 17032
rect 69004 16988 69044 17200
rect 68908 16948 69044 16988
rect 68908 16241 68948 16948
rect 69292 16736 69332 17284
rect 69545 17156 69585 17472
rect 69004 16696 69332 16736
rect 69388 17116 69585 17156
rect 69004 16484 69044 16696
rect 69004 16435 69044 16444
rect 68907 16232 68949 16241
rect 69388 16232 69428 17116
rect 69655 17072 69695 17472
rect 69945 17156 69985 17472
rect 69484 17032 69695 17072
rect 69772 17116 69985 17156
rect 69484 16484 69524 17032
rect 69484 16435 69524 16444
rect 68907 16192 68908 16232
rect 68948 16192 68949 16232
rect 68907 16183 68949 16192
rect 69292 16192 69388 16232
rect 68908 16098 68948 16183
rect 68660 16024 68852 16064
rect 68620 16015 68660 16024
rect 69292 15989 69332 16192
rect 69388 16183 69428 16192
rect 69772 16232 69812 17116
rect 70055 17072 70095 17472
rect 70345 17156 70385 17472
rect 69868 17032 70095 17072
rect 70156 17116 70385 17156
rect 69868 16484 69908 17032
rect 69868 16435 69908 16444
rect 70156 16241 70196 17116
rect 70455 17072 70495 17472
rect 70745 17156 70785 17472
rect 70252 17032 70495 17072
rect 70540 17116 70785 17156
rect 70252 16484 70292 17032
rect 70252 16435 70292 16444
rect 69772 16157 69812 16192
rect 70155 16232 70197 16241
rect 70155 16192 70156 16232
rect 70196 16192 70197 16232
rect 70155 16183 70197 16192
rect 70540 16232 70580 17116
rect 70855 17072 70895 17472
rect 71145 17156 71185 17472
rect 70636 17032 70895 17072
rect 70937 17116 71185 17156
rect 70636 16484 70676 17032
rect 70937 16988 70977 17116
rect 71255 17072 71295 17472
rect 71403 17156 71445 17165
rect 71545 17156 71585 17472
rect 71655 17165 71695 17472
rect 71403 17116 71404 17156
rect 71444 17116 71445 17156
rect 71403 17107 71445 17116
rect 71500 17116 71585 17156
rect 71654 17156 71696 17165
rect 71945 17156 71985 17472
rect 71654 17116 71655 17156
rect 71695 17116 71696 17156
rect 70636 16435 70676 16444
rect 70924 16948 70977 16988
rect 71020 17032 71295 17072
rect 69771 16148 69813 16157
rect 69771 16108 69772 16148
rect 69812 16108 69813 16148
rect 69771 16099 69813 16108
rect 70156 16098 70196 16183
rect 70540 16073 70580 16192
rect 70924 16232 70964 16948
rect 71020 16484 71060 17032
rect 71020 16435 71060 16444
rect 71404 16484 71444 17107
rect 71404 16435 71444 16444
rect 69387 16064 69429 16073
rect 69387 16024 69388 16064
rect 69428 16024 69429 16064
rect 69387 16015 69429 16024
rect 70539 16064 70581 16073
rect 70539 16024 70540 16064
rect 70580 16024 70581 16064
rect 70539 16015 70581 16024
rect 69291 15980 69333 15989
rect 69291 15940 69292 15980
rect 69332 15940 69333 15980
rect 69291 15931 69333 15940
rect 68716 15485 68756 15570
rect 68811 15560 68853 15569
rect 68811 15520 68812 15560
rect 68852 15520 68853 15560
rect 68811 15511 68853 15520
rect 68715 15476 68757 15485
rect 68715 15436 68716 15476
rect 68756 15436 68757 15476
rect 68715 15427 68757 15436
rect 68715 15308 68757 15317
rect 68715 15268 68716 15308
rect 68756 15268 68757 15308
rect 68715 15259 68757 15268
rect 68332 14048 68372 14057
rect 68524 14048 68564 14057
rect 68372 14008 68524 14048
rect 68332 13999 68372 14008
rect 68524 13999 68564 14008
rect 68619 14048 68661 14057
rect 68619 14008 68620 14048
rect 68660 14008 68661 14048
rect 68619 13999 68661 14008
rect 68716 14048 68756 15259
rect 68812 14720 68852 15511
rect 68907 15308 68949 15317
rect 68907 15268 68908 15308
rect 68948 15268 68949 15308
rect 68907 15259 68949 15268
rect 68908 15174 68948 15259
rect 68907 14720 68949 14729
rect 68852 14680 68908 14720
rect 68948 14680 68949 14720
rect 68812 14671 68852 14680
rect 68907 14671 68949 14680
rect 68811 14132 68853 14141
rect 68811 14092 68812 14132
rect 68852 14092 68853 14132
rect 68811 14083 68853 14092
rect 67852 7288 67988 7328
rect 68044 13840 68276 13880
rect 67852 5909 67892 7288
rect 67947 7160 67989 7169
rect 67947 7120 67948 7160
rect 67988 7120 67989 7160
rect 67947 7111 67989 7120
rect 67948 6488 67988 7111
rect 67948 6439 67988 6448
rect 67851 5900 67893 5909
rect 67851 5860 67852 5900
rect 67892 5860 67893 5900
rect 67851 5851 67893 5860
rect 67659 4892 67701 4901
rect 67659 4852 67660 4892
rect 67700 4852 67701 4892
rect 67659 4843 67701 4852
rect 67755 4724 67797 4733
rect 67755 4684 67756 4724
rect 67796 4684 67797 4724
rect 67755 4675 67797 4684
rect 67660 4136 67700 4145
rect 67660 3044 67700 4096
rect 67564 3004 67700 3044
rect 67372 2860 67508 2900
rect 64684 2633 64724 2860
rect 66508 2792 66548 2801
rect 64779 2708 64821 2717
rect 64779 2668 64780 2708
rect 64820 2668 64821 2708
rect 64779 2659 64821 2668
rect 64683 2624 64725 2633
rect 64683 2584 64684 2624
rect 64724 2584 64725 2624
rect 64683 2575 64725 2584
rect 64780 2574 64820 2659
rect 64875 2624 64917 2633
rect 64875 2584 64876 2624
rect 64916 2584 64917 2624
rect 64875 2575 64917 2584
rect 65259 2624 65301 2633
rect 65259 2584 65260 2624
rect 65300 2584 65301 2624
rect 65259 2575 65301 2584
rect 64876 2490 64916 2575
rect 64683 2456 64725 2465
rect 64683 2416 64684 2456
rect 64724 2416 64725 2456
rect 64683 2407 64725 2416
rect 64684 2036 64724 2407
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 65260 2129 65300 2575
rect 65259 2120 65301 2129
rect 65259 2080 65260 2120
rect 65300 2080 65301 2120
rect 65259 2071 65301 2080
rect 64684 1996 64820 2036
rect 64588 1912 64724 1952
rect 64492 1903 64532 1912
rect 64684 1289 64724 1912
rect 64396 1280 64436 1289
rect 64683 1280 64725 1289
rect 64436 1240 64628 1280
rect 64396 1231 64436 1240
rect 64588 1112 64628 1240
rect 64683 1240 64684 1280
rect 64724 1240 64725 1280
rect 64683 1231 64725 1240
rect 64684 1146 64724 1231
rect 64588 1063 64628 1072
rect 64780 1112 64820 1996
rect 64876 1952 64916 1961
rect 64916 1912 65012 1952
rect 64876 1903 64916 1912
rect 64972 1280 65012 1912
rect 65260 1373 65300 2071
rect 65739 1952 65781 1961
rect 65739 1912 65740 1952
rect 65780 1912 65781 1952
rect 65739 1903 65781 1912
rect 65740 1818 65780 1903
rect 65259 1364 65301 1373
rect 65259 1324 65260 1364
rect 65300 1324 65301 1364
rect 65259 1315 65301 1324
rect 64972 1231 65012 1240
rect 64780 1063 64820 1072
rect 66027 1112 66069 1121
rect 66027 1072 66028 1112
rect 66068 1072 66069 1112
rect 66027 1063 66069 1072
rect 66412 1112 66452 1121
rect 66508 1112 66548 2752
rect 67468 2549 67508 2860
rect 66891 2540 66933 2549
rect 66891 2500 66892 2540
rect 66932 2500 66933 2540
rect 66891 2491 66933 2500
rect 67467 2540 67509 2549
rect 67467 2500 67468 2540
rect 67508 2500 67509 2540
rect 67467 2491 67509 2500
rect 66892 2129 66932 2491
rect 67371 2456 67413 2465
rect 67371 2416 67372 2456
rect 67412 2416 67413 2456
rect 67371 2407 67413 2416
rect 66891 2120 66933 2129
rect 66891 2080 66892 2120
rect 66932 2080 66933 2120
rect 66891 2071 66933 2080
rect 66892 1986 66932 2071
rect 67275 1952 67317 1961
rect 67275 1912 67276 1952
rect 67316 1912 67317 1952
rect 67275 1903 67317 1912
rect 67372 1952 67412 2407
rect 67564 2288 67604 3004
rect 67756 2900 67796 4675
rect 67468 2248 67604 2288
rect 67660 2860 67796 2900
rect 67468 1961 67508 2248
rect 67563 2036 67605 2045
rect 67563 1996 67564 2036
rect 67604 1996 67605 2036
rect 67563 1987 67605 1996
rect 67372 1903 67412 1912
rect 67467 1952 67509 1961
rect 67467 1912 67468 1952
rect 67508 1912 67509 1952
rect 67467 1903 67509 1912
rect 67564 1952 67604 1987
rect 66452 1072 66548 1112
rect 67276 1112 67316 1903
rect 67564 1901 67604 1912
rect 67660 1952 67700 2860
rect 67947 2624 67989 2633
rect 67947 2584 67948 2624
rect 67988 2584 67989 2624
rect 67947 2575 67989 2584
rect 67660 1903 67700 1912
rect 67948 1952 67988 2575
rect 67948 1903 67988 1912
rect 68044 1709 68084 13840
rect 68331 13796 68373 13805
rect 68331 13756 68332 13796
rect 68372 13756 68373 13796
rect 68331 13747 68373 13756
rect 68139 13712 68181 13721
rect 68139 13672 68140 13712
rect 68180 13672 68181 13712
rect 68139 13663 68181 13672
rect 68140 9680 68180 13663
rect 68332 13662 68372 13747
rect 68620 13208 68660 13999
rect 68620 13049 68660 13168
rect 68716 13208 68756 14008
rect 68812 14048 68852 14083
rect 68812 13997 68852 14008
rect 68812 13217 68852 13302
rect 68524 13040 68564 13049
rect 68427 12872 68469 12881
rect 68427 12832 68428 12872
rect 68468 12832 68469 12872
rect 68427 12823 68469 12832
rect 68428 10613 68468 12823
rect 68524 11696 68564 13000
rect 68619 13040 68661 13049
rect 68619 13000 68620 13040
rect 68660 13000 68661 13040
rect 68619 12991 68661 13000
rect 68716 12713 68756 13168
rect 68811 13208 68853 13217
rect 68811 13168 68812 13208
rect 68852 13168 68853 13208
rect 68811 13159 68853 13168
rect 68811 13040 68853 13049
rect 68811 13000 68812 13040
rect 68852 13000 68853 13040
rect 68811 12991 68853 13000
rect 68812 12881 68852 12991
rect 68811 12872 68853 12881
rect 68811 12832 68812 12872
rect 68852 12832 68853 12872
rect 68811 12823 68853 12832
rect 68715 12704 68757 12713
rect 68715 12664 68716 12704
rect 68756 12664 68757 12704
rect 68715 12655 68757 12664
rect 68620 12536 68660 12545
rect 68908 12536 68948 14671
rect 69195 14384 69237 14393
rect 69195 14344 69196 14384
rect 69236 14344 69237 14384
rect 69195 14335 69237 14344
rect 69004 14216 69044 14225
rect 69004 14057 69044 14176
rect 69099 14132 69141 14141
rect 69099 14092 69100 14132
rect 69140 14092 69141 14132
rect 69099 14083 69141 14092
rect 69003 14048 69045 14057
rect 69003 14008 69004 14048
rect 69044 14008 69045 14048
rect 69003 13999 69045 14008
rect 69100 13880 69140 14083
rect 69196 13973 69236 14335
rect 69195 13964 69237 13973
rect 69195 13924 69196 13964
rect 69236 13924 69237 13964
rect 69195 13915 69237 13924
rect 69004 13840 69140 13880
rect 69004 13208 69044 13840
rect 69196 13830 69236 13915
rect 69291 13292 69333 13301
rect 69291 13252 69292 13292
rect 69332 13252 69333 13292
rect 69291 13243 69333 13252
rect 69004 13159 69044 13168
rect 69100 13208 69140 13219
rect 69100 13133 69140 13168
rect 69292 13208 69332 13243
rect 69099 13124 69141 13133
rect 69099 13084 69100 13124
rect 69140 13084 69141 13124
rect 69099 13075 69141 13084
rect 69196 13040 69236 13049
rect 69003 12704 69045 12713
rect 69003 12664 69004 12704
rect 69044 12664 69045 12704
rect 69003 12655 69045 12664
rect 68660 12496 68948 12536
rect 68620 12487 68660 12496
rect 68907 11948 68949 11957
rect 68907 11908 68908 11948
rect 68948 11908 68949 11948
rect 68907 11899 68949 11908
rect 68908 11814 68948 11899
rect 68908 11696 68948 11705
rect 68524 11656 68908 11696
rect 68908 11647 68948 11656
rect 68907 11528 68949 11537
rect 68907 11488 68908 11528
rect 68948 11488 68949 11528
rect 68907 11479 68949 11488
rect 68908 11024 68948 11479
rect 68812 10984 68908 11024
rect 68427 10604 68469 10613
rect 68427 10564 68428 10604
rect 68468 10564 68469 10604
rect 68427 10555 68469 10564
rect 68427 10436 68469 10445
rect 68427 10396 68428 10436
rect 68468 10396 68469 10436
rect 68427 10387 68469 10396
rect 68331 10184 68373 10193
rect 68331 10144 68332 10184
rect 68372 10144 68373 10184
rect 68331 10135 68373 10144
rect 68428 10184 68468 10387
rect 68812 10277 68852 10984
rect 68908 10975 68948 10984
rect 69004 10949 69044 12655
rect 69099 12368 69141 12377
rect 69099 12328 69100 12368
rect 69140 12328 69141 12368
rect 69099 12319 69141 12328
rect 69100 11696 69140 12319
rect 69100 11647 69140 11656
rect 69196 11696 69236 13000
rect 69292 12989 69332 13168
rect 69291 12980 69333 12989
rect 69291 12940 69292 12980
rect 69332 12940 69333 12980
rect 69291 12931 69333 12940
rect 69388 12872 69428 16015
rect 70924 15905 70964 16192
rect 71308 16232 71348 16241
rect 71500 16232 71540 17116
rect 71654 17107 71696 17116
rect 71788 17116 71985 17156
rect 71348 16192 71540 16232
rect 71788 16232 71828 17116
rect 72055 17072 72095 17472
rect 72345 17156 72385 17472
rect 71884 17032 72095 17072
rect 72172 17116 72385 17156
rect 71884 16484 71924 17032
rect 71884 16435 71924 16444
rect 71308 16183 71348 16192
rect 70923 15896 70965 15905
rect 70923 15856 70924 15896
rect 70964 15856 70965 15896
rect 70923 15847 70965 15856
rect 71115 15644 71157 15653
rect 71115 15604 71116 15644
rect 71156 15604 71157 15644
rect 71115 15595 71157 15604
rect 70059 15560 70101 15569
rect 70059 15520 70060 15560
rect 70100 15520 70101 15560
rect 70059 15511 70101 15520
rect 70156 15560 70196 15569
rect 70348 15560 70388 15569
rect 70196 15520 70292 15560
rect 70156 15511 70196 15520
rect 69868 15476 69908 15487
rect 69868 15401 69908 15436
rect 70060 15426 70100 15511
rect 69867 15392 69909 15401
rect 69867 15352 69868 15392
rect 69908 15352 69909 15392
rect 69867 15343 69909 15352
rect 69676 15308 69716 15317
rect 69676 14048 69716 15268
rect 69964 14552 70004 14561
rect 70004 14512 70100 14552
rect 69964 14503 70004 14512
rect 70060 14141 70100 14512
rect 70252 14225 70292 15520
rect 70348 15476 70388 15520
rect 70924 15560 70964 15569
rect 70731 15476 70773 15485
rect 70348 15436 70676 15476
rect 70348 15308 70388 15317
rect 70540 15308 70580 15317
rect 70348 14720 70388 15268
rect 70348 14671 70388 14680
rect 70444 15268 70540 15308
rect 70251 14216 70293 14225
rect 70251 14176 70252 14216
rect 70292 14176 70293 14216
rect 70251 14167 70293 14176
rect 70059 14132 70101 14141
rect 70059 14092 70060 14132
rect 70100 14092 70101 14132
rect 70059 14083 70101 14092
rect 69484 14008 69676 14048
rect 69484 13301 69524 14008
rect 69676 13999 69716 14008
rect 69963 14048 70005 14057
rect 69963 14008 69964 14048
rect 70004 14008 70005 14048
rect 69963 13999 70005 14008
rect 69964 13914 70004 13999
rect 70060 13998 70100 14083
rect 69675 13544 69717 13553
rect 69675 13504 69676 13544
rect 69716 13504 69717 13544
rect 69675 13495 69717 13504
rect 70059 13544 70101 13553
rect 70059 13504 70060 13544
rect 70100 13504 70101 13544
rect 70059 13495 70101 13504
rect 69483 13292 69525 13301
rect 69483 13252 69484 13292
rect 69524 13252 69525 13292
rect 69483 13243 69525 13252
rect 69196 11647 69236 11656
rect 69292 12832 69428 12872
rect 69195 11528 69237 11537
rect 69195 11488 69196 11528
rect 69236 11488 69237 11528
rect 69195 11479 69237 11488
rect 69099 11024 69141 11033
rect 69099 10984 69100 11024
rect 69140 10984 69141 11024
rect 69099 10975 69141 10984
rect 69196 11024 69236 11479
rect 69292 11444 69332 12832
rect 69484 11696 69524 13243
rect 69579 13208 69621 13217
rect 69579 13168 69580 13208
rect 69620 13168 69621 13208
rect 69579 13159 69621 13168
rect 69676 13208 69716 13495
rect 69676 13159 69716 13168
rect 69868 13208 69908 13217
rect 69580 12293 69620 13159
rect 69772 13124 69812 13133
rect 69675 12956 69717 12965
rect 69675 12916 69676 12956
rect 69716 12916 69717 12956
rect 69675 12907 69717 12916
rect 69579 12284 69621 12293
rect 69579 12244 69580 12284
rect 69620 12244 69621 12284
rect 69579 12235 69621 12244
rect 69676 11873 69716 12907
rect 69772 12881 69812 13084
rect 69771 12872 69813 12881
rect 69771 12832 69772 12872
rect 69812 12832 69813 12872
rect 69771 12823 69813 12832
rect 69771 12284 69813 12293
rect 69771 12244 69772 12284
rect 69812 12244 69813 12284
rect 69771 12235 69813 12244
rect 69675 11864 69717 11873
rect 69675 11824 69676 11864
rect 69716 11824 69717 11864
rect 69772 11864 69812 12235
rect 69868 11948 69908 13168
rect 70060 13208 70100 13495
rect 70156 13460 70196 13469
rect 70252 13460 70292 14167
rect 70196 13420 70292 13460
rect 70348 13796 70388 13805
rect 70156 13411 70196 13420
rect 70060 13159 70100 13168
rect 70252 13208 70292 13217
rect 70348 13208 70388 13756
rect 70444 13553 70484 15268
rect 70540 15259 70580 15268
rect 70636 15140 70676 15436
rect 70731 15436 70732 15476
rect 70772 15436 70773 15476
rect 70731 15427 70773 15436
rect 70540 15100 70676 15140
rect 70540 14216 70580 15100
rect 70732 14897 70772 15427
rect 70827 15224 70869 15233
rect 70827 15184 70828 15224
rect 70868 15184 70869 15224
rect 70827 15175 70869 15184
rect 70731 14888 70773 14897
rect 70731 14848 70732 14888
rect 70772 14848 70773 14888
rect 70731 14839 70773 14848
rect 70732 14720 70772 14729
rect 70828 14720 70868 15175
rect 70772 14680 70868 14720
rect 70732 14671 70772 14680
rect 70924 14636 70964 15520
rect 71019 15560 71061 15569
rect 71019 15520 71020 15560
rect 71060 15520 71061 15560
rect 71019 15511 71061 15520
rect 71116 15560 71156 15595
rect 71020 15426 71060 15511
rect 71116 15509 71156 15520
rect 71308 15392 71348 15401
rect 71308 15233 71348 15352
rect 71307 15224 71349 15233
rect 71307 15184 71308 15224
rect 71348 15184 71349 15224
rect 71307 15175 71349 15184
rect 70924 14596 71156 14636
rect 70827 14468 70869 14477
rect 70827 14428 70828 14468
rect 70868 14428 70869 14468
rect 70827 14419 70869 14428
rect 70732 14216 70772 14225
rect 70540 14176 70732 14216
rect 70732 14167 70772 14176
rect 70540 13964 70580 13973
rect 70828 13964 70868 14419
rect 70923 14300 70965 14309
rect 70923 14260 70924 14300
rect 70964 14260 70965 14300
rect 70923 14251 70965 14260
rect 70580 13924 70868 13964
rect 70924 13964 70964 14251
rect 71116 14216 71156 14596
rect 71116 14167 71156 14176
rect 70540 13915 70580 13924
rect 70732 13796 70772 13805
rect 70443 13544 70485 13553
rect 70443 13504 70444 13544
rect 70484 13504 70485 13544
rect 70443 13495 70485 13504
rect 70732 13385 70772 13756
rect 70924 13721 70964 13924
rect 71116 13796 71156 13805
rect 70923 13712 70965 13721
rect 70923 13672 70924 13712
rect 70964 13672 70965 13712
rect 70923 13663 70965 13672
rect 70924 13544 70964 13663
rect 70828 13504 70964 13544
rect 70443 13376 70485 13385
rect 70443 13336 70444 13376
rect 70484 13336 70485 13376
rect 70443 13327 70485 13336
rect 70731 13376 70773 13385
rect 70731 13336 70732 13376
rect 70772 13336 70773 13376
rect 70731 13327 70773 13336
rect 70292 13168 70388 13208
rect 70252 13159 70292 13168
rect 70444 12980 70484 13327
rect 70539 13208 70581 13217
rect 70539 13168 70540 13208
rect 70580 13168 70581 13208
rect 70539 13159 70581 13168
rect 70252 12940 70484 12980
rect 70059 12872 70101 12881
rect 70059 12832 70060 12872
rect 70100 12832 70101 12872
rect 70059 12823 70101 12832
rect 69963 12536 70005 12545
rect 69963 12496 69964 12536
rect 70004 12496 70005 12536
rect 69963 12487 70005 12496
rect 70060 12536 70100 12823
rect 70252 12620 70292 12940
rect 70540 12704 70580 13159
rect 70828 13124 70868 13504
rect 70732 13084 70868 13124
rect 70924 13376 70964 13385
rect 69964 12402 70004 12487
rect 70060 12377 70100 12496
rect 70156 12580 70292 12620
rect 70059 12368 70101 12377
rect 70059 12328 70060 12368
rect 70100 12328 70101 12368
rect 70059 12319 70101 12328
rect 70156 12200 70196 12580
rect 70252 12578 70292 12580
rect 70252 12529 70292 12538
rect 70348 12664 70580 12704
rect 70635 12704 70677 12713
rect 70635 12664 70636 12704
rect 70676 12664 70677 12704
rect 70252 12377 70292 12462
rect 70251 12368 70293 12377
rect 70251 12328 70252 12368
rect 70292 12328 70293 12368
rect 70251 12319 70293 12328
rect 70348 12284 70388 12664
rect 70635 12655 70677 12664
rect 70444 12536 70484 12547
rect 70444 12461 70484 12496
rect 70539 12536 70581 12545
rect 70539 12496 70540 12536
rect 70580 12496 70581 12536
rect 70539 12487 70581 12496
rect 70443 12452 70485 12461
rect 70443 12412 70444 12452
rect 70484 12412 70485 12452
rect 70443 12403 70485 12412
rect 70348 12244 70484 12284
rect 70156 12160 70292 12200
rect 70156 11948 70196 11957
rect 69868 11908 70156 11948
rect 70156 11899 70196 11908
rect 69772 11824 69908 11864
rect 69675 11815 69717 11824
rect 69771 11696 69813 11705
rect 69524 11656 69716 11696
rect 69484 11647 69524 11656
rect 69292 11404 69428 11444
rect 69196 10975 69236 10984
rect 69003 10940 69045 10949
rect 69003 10900 69004 10940
rect 69044 10900 69045 10940
rect 69003 10891 69045 10900
rect 69100 10890 69140 10975
rect 69388 10940 69428 11404
rect 69292 10900 69428 10940
rect 69579 10940 69621 10949
rect 69579 10900 69580 10940
rect 69620 10900 69621 10940
rect 69676 10940 69716 11656
rect 69771 11656 69772 11696
rect 69812 11656 69813 11696
rect 69771 11647 69813 11656
rect 69772 11562 69812 11647
rect 69868 11612 69908 11824
rect 69868 11537 69908 11572
rect 69867 11528 69909 11537
rect 69867 11488 69868 11528
rect 69908 11488 69909 11528
rect 69867 11479 69909 11488
rect 69964 10940 70004 10949
rect 69676 10900 69964 10940
rect 70252 10940 70292 12160
rect 70444 11696 70484 12244
rect 70540 11948 70580 12487
rect 70540 11899 70580 11908
rect 70636 11705 70676 12655
rect 70444 11033 70484 11656
rect 70635 11696 70677 11705
rect 70635 11656 70636 11696
rect 70676 11656 70677 11696
rect 70635 11647 70677 11656
rect 70636 11562 70676 11647
rect 70443 11024 70485 11033
rect 70443 10984 70444 11024
rect 70484 10984 70485 11024
rect 70443 10975 70485 10984
rect 70348 10940 70388 10949
rect 70252 10900 70348 10940
rect 68908 10772 68948 10781
rect 68948 10732 69044 10772
rect 68908 10723 68948 10732
rect 68811 10268 68853 10277
rect 68811 10228 68812 10268
rect 68852 10228 68853 10268
rect 68811 10219 68853 10228
rect 68236 10100 68276 10111
rect 68236 10025 68276 10060
rect 68332 10050 68372 10135
rect 68235 10016 68277 10025
rect 68235 9976 68236 10016
rect 68276 9976 68277 10016
rect 68235 9967 68277 9976
rect 68428 9932 68468 10144
rect 68523 10184 68565 10193
rect 68523 10144 68524 10184
rect 68564 10144 68565 10184
rect 68523 10135 68565 10144
rect 68716 10184 68756 10193
rect 68524 10050 68564 10135
rect 68716 10025 68756 10144
rect 68908 10184 68948 10193
rect 68908 10109 68948 10144
rect 69004 10184 69044 10732
rect 69292 10352 69332 10900
rect 69579 10891 69621 10900
rect 69964 10891 70004 10900
rect 70348 10891 70388 10900
rect 70540 10940 70580 10949
rect 70732 10940 70772 13084
rect 70924 12980 70964 13336
rect 71116 13217 71156 13756
rect 71115 13208 71157 13217
rect 71115 13168 71116 13208
rect 71156 13168 71157 13208
rect 71115 13159 71157 13168
rect 70828 12940 70964 12980
rect 70828 12536 70868 12940
rect 70828 12487 70868 12496
rect 71211 12536 71253 12545
rect 71211 12496 71212 12536
rect 71252 12496 71253 12536
rect 71211 12487 71253 12496
rect 71116 10940 71156 10949
rect 70580 10900 70772 10940
rect 70828 10900 71116 10940
rect 70540 10891 70580 10900
rect 69580 10806 69620 10891
rect 69388 10772 69428 10781
rect 69388 10529 69428 10732
rect 69772 10772 69812 10781
rect 70156 10772 70196 10781
rect 69387 10520 69429 10529
rect 69387 10480 69388 10520
rect 69428 10480 69429 10520
rect 69387 10471 69429 10480
rect 69579 10436 69621 10445
rect 69579 10396 69580 10436
rect 69620 10396 69621 10436
rect 69579 10387 69621 10396
rect 69196 10312 69332 10352
rect 69387 10352 69429 10361
rect 69387 10312 69388 10352
rect 69428 10312 69429 10352
rect 69099 10268 69141 10277
rect 69099 10228 69100 10268
rect 69140 10228 69141 10268
rect 69099 10219 69141 10228
rect 69004 10135 69044 10144
rect 68811 10100 68853 10109
rect 68811 10060 68812 10100
rect 68852 10060 68853 10100
rect 68908 10100 68960 10109
rect 68908 10060 68919 10100
rect 68959 10060 68960 10100
rect 68811 10051 68853 10060
rect 68918 10051 68960 10060
rect 68715 10016 68757 10025
rect 68715 9976 68716 10016
rect 68756 9976 68757 10016
rect 68715 9967 68757 9976
rect 68812 9966 68852 10051
rect 68428 9892 68564 9932
rect 68140 9640 68468 9680
rect 68140 9512 68180 9521
rect 68140 8681 68180 9472
rect 68428 8924 68468 9640
rect 68428 8875 68468 8884
rect 68139 8672 68181 8681
rect 68139 8632 68140 8672
rect 68180 8632 68181 8672
rect 68139 8623 68181 8632
rect 68428 8504 68468 8513
rect 68331 8084 68373 8093
rect 68331 8044 68332 8084
rect 68372 8044 68373 8084
rect 68331 8035 68373 8044
rect 68332 7950 68372 8035
rect 68428 8009 68468 8464
rect 68427 8000 68469 8009
rect 68427 7960 68428 8000
rect 68468 7960 68469 8000
rect 68427 7951 68469 7960
rect 68524 6329 68564 9892
rect 68715 8840 68757 8849
rect 68715 8800 68716 8840
rect 68756 8800 68757 8840
rect 68715 8791 68757 8800
rect 68716 8000 68756 8791
rect 68908 8756 68948 8765
rect 69100 8756 69140 10219
rect 68948 8716 69140 8756
rect 68908 8707 68948 8716
rect 68716 7951 68756 7960
rect 69100 8504 69140 8513
rect 69100 7001 69140 8464
rect 69196 7085 69236 10312
rect 69387 10303 69429 10312
rect 69292 10184 69332 10193
rect 69388 10184 69428 10303
rect 69332 10144 69428 10184
rect 69483 10184 69525 10193
rect 69483 10144 69484 10184
rect 69524 10144 69525 10184
rect 69292 10135 69332 10144
rect 69483 10135 69525 10144
rect 69580 10184 69620 10387
rect 69772 10361 69812 10732
rect 69868 10732 70156 10772
rect 69771 10352 69813 10361
rect 69771 10312 69772 10352
rect 69812 10312 69813 10352
rect 69771 10303 69813 10312
rect 69676 10193 69716 10278
rect 69580 10135 69620 10144
rect 69675 10184 69717 10193
rect 69675 10144 69676 10184
rect 69716 10144 69717 10184
rect 69868 10184 69908 10732
rect 70156 10723 70196 10732
rect 70732 10772 70772 10781
rect 70828 10772 70868 10900
rect 70772 10732 70868 10772
rect 70924 10772 70964 10781
rect 70732 10723 70772 10732
rect 70924 10688 70964 10732
rect 70828 10648 70964 10688
rect 70155 10604 70197 10613
rect 70155 10564 70156 10604
rect 70196 10564 70197 10604
rect 70155 10555 70197 10564
rect 69964 10352 70004 10361
rect 70004 10312 70100 10352
rect 69964 10303 70004 10312
rect 69868 10144 70004 10184
rect 69675 10135 69717 10144
rect 69292 9680 69332 9689
rect 69484 9680 69524 10135
rect 69867 10016 69909 10025
rect 69867 9976 69868 10016
rect 69908 9976 69909 10016
rect 69867 9967 69909 9976
rect 69675 9932 69717 9941
rect 69675 9892 69676 9932
rect 69716 9892 69717 9932
rect 69675 9883 69717 9892
rect 69332 9640 69524 9680
rect 69292 9631 69332 9640
rect 69484 9512 69524 9640
rect 69579 9596 69621 9605
rect 69579 9556 69580 9596
rect 69620 9556 69621 9596
rect 69579 9547 69621 9556
rect 69484 9463 69524 9472
rect 69580 9512 69620 9547
rect 69580 9461 69620 9472
rect 69579 9260 69621 9269
rect 69579 9220 69580 9260
rect 69620 9220 69621 9260
rect 69579 9211 69621 9220
rect 69483 8756 69525 8765
rect 69483 8716 69484 8756
rect 69524 8716 69525 8756
rect 69483 8707 69525 8716
rect 69292 8672 69332 8681
rect 69292 7580 69332 8632
rect 69484 8672 69524 8707
rect 69484 8621 69524 8632
rect 69580 8672 69620 9211
rect 69676 8681 69716 9883
rect 69772 9512 69812 9523
rect 69772 9437 69812 9472
rect 69771 9428 69813 9437
rect 69771 9388 69772 9428
rect 69812 9388 69813 9428
rect 69771 9379 69813 9388
rect 69771 9260 69813 9269
rect 69771 9220 69772 9260
rect 69812 9220 69813 9260
rect 69771 9211 69813 9220
rect 69772 9126 69812 9211
rect 69868 8924 69908 9967
rect 69964 9521 70004 10144
rect 69963 9512 70005 9521
rect 69963 9472 69964 9512
rect 70004 9472 70005 9512
rect 69963 9463 70005 9472
rect 69963 9344 70005 9353
rect 69963 9304 69964 9344
rect 70004 9304 70005 9344
rect 69963 9295 70005 9304
rect 69964 9210 70004 9295
rect 69868 8875 69908 8884
rect 69580 8623 69620 8632
rect 69675 8672 69717 8681
rect 69675 8632 69676 8672
rect 69716 8632 69717 8672
rect 69675 8623 69717 8632
rect 69772 8672 69812 8681
rect 69867 8672 69909 8681
rect 69812 8632 69868 8672
rect 69908 8632 69909 8672
rect 69772 8623 69812 8632
rect 69867 8623 69909 8632
rect 69964 8672 70004 8681
rect 70060 8672 70100 10312
rect 70156 10268 70196 10555
rect 70348 10352 70388 10363
rect 70348 10277 70388 10312
rect 70731 10352 70773 10361
rect 70731 10312 70732 10352
rect 70772 10312 70773 10352
rect 70731 10303 70773 10312
rect 70156 10219 70196 10228
rect 70347 10268 70389 10277
rect 70347 10228 70348 10268
rect 70388 10228 70389 10268
rect 70347 10219 70389 10228
rect 70155 10100 70197 10109
rect 70155 10060 70156 10100
rect 70196 10060 70197 10100
rect 70155 10051 70197 10060
rect 70443 10100 70485 10109
rect 70443 10060 70444 10100
rect 70484 10060 70485 10100
rect 70443 10051 70485 10060
rect 70540 10100 70580 10109
rect 70156 9512 70196 10051
rect 70347 9596 70389 9605
rect 70347 9556 70348 9596
rect 70388 9556 70389 9596
rect 70347 9547 70389 9556
rect 70156 9463 70196 9472
rect 70251 9512 70293 9521
rect 70251 9472 70252 9512
rect 70292 9472 70293 9512
rect 70251 9463 70293 9472
rect 70252 9378 70292 9463
rect 70251 9260 70293 9269
rect 70251 9220 70252 9260
rect 70292 9220 70293 9260
rect 70251 9211 70293 9220
rect 70155 8840 70197 8849
rect 70155 8800 70156 8840
rect 70196 8800 70197 8840
rect 70155 8791 70197 8800
rect 70156 8706 70196 8791
rect 70004 8632 70100 8672
rect 69964 8623 70004 8632
rect 69388 8504 69428 8513
rect 69388 8093 69428 8464
rect 69387 8084 69429 8093
rect 69387 8044 69388 8084
rect 69428 8044 69429 8084
rect 69387 8035 69429 8044
rect 69580 8000 69620 8009
rect 69676 8000 69716 8623
rect 70252 8588 70292 9211
rect 70156 8548 70292 8588
rect 69771 8504 69813 8513
rect 69771 8464 69772 8504
rect 69812 8464 69813 8504
rect 69771 8455 69813 8464
rect 69620 7960 69716 8000
rect 69292 7540 69524 7580
rect 69388 7328 69428 7337
rect 69195 7076 69237 7085
rect 69195 7036 69196 7076
rect 69236 7036 69237 7076
rect 69195 7027 69237 7036
rect 69099 6992 69141 7001
rect 69099 6952 69100 6992
rect 69140 6952 69141 6992
rect 69099 6943 69141 6952
rect 69100 6656 69140 6665
rect 69196 6656 69236 7027
rect 69140 6616 69236 6656
rect 69100 6607 69140 6616
rect 69388 6497 69428 7288
rect 69484 6992 69524 7540
rect 69580 7169 69620 7960
rect 69772 7328 69812 8455
rect 69867 7748 69909 7757
rect 69867 7708 69868 7748
rect 69908 7708 69909 7748
rect 69867 7699 69909 7708
rect 69676 7288 69812 7328
rect 69579 7160 69621 7169
rect 69579 7120 69580 7160
rect 69620 7120 69621 7160
rect 69579 7111 69621 7120
rect 69676 7160 69716 7288
rect 69580 6992 69620 7001
rect 69484 6952 69580 6992
rect 69580 6943 69620 6952
rect 69676 6656 69716 7120
rect 69484 6616 69716 6656
rect 69772 7160 69812 7169
rect 69292 6488 69332 6497
rect 68523 6320 68565 6329
rect 68523 6280 68524 6320
rect 68564 6280 68565 6320
rect 68523 6271 68565 6280
rect 69292 5909 69332 6448
rect 69387 6488 69429 6497
rect 69387 6448 69388 6488
rect 69428 6448 69429 6488
rect 69387 6439 69429 6448
rect 69387 6320 69429 6329
rect 69387 6280 69388 6320
rect 69428 6280 69429 6320
rect 69387 6271 69429 6280
rect 69291 5900 69333 5909
rect 69291 5860 69292 5900
rect 69332 5860 69333 5900
rect 69291 5851 69333 5860
rect 69291 5732 69333 5741
rect 69291 5692 69292 5732
rect 69332 5692 69333 5732
rect 69291 5683 69333 5692
rect 69292 5648 69332 5683
rect 68715 4976 68757 4985
rect 68715 4936 68716 4976
rect 68756 4936 68757 4976
rect 68715 4927 68757 4936
rect 68908 4976 68948 4985
rect 69099 4976 69141 4985
rect 68948 4936 69044 4976
rect 68908 4927 68948 4936
rect 68235 3464 68277 3473
rect 68235 3424 68236 3464
rect 68276 3424 68277 3464
rect 68235 3415 68277 3424
rect 68620 3464 68660 3473
rect 68236 2624 68276 3415
rect 68331 3212 68373 3221
rect 68331 3172 68332 3212
rect 68372 3172 68373 3212
rect 68331 3163 68373 3172
rect 68236 2575 68276 2584
rect 68332 2624 68372 3163
rect 68620 2900 68660 3424
rect 68716 3464 68756 4927
rect 68907 4724 68949 4733
rect 68907 4684 68908 4724
rect 68948 4684 68949 4724
rect 68907 4675 68949 4684
rect 68908 4590 68948 4675
rect 69004 4565 69044 4936
rect 69099 4936 69100 4976
rect 69140 4936 69141 4976
rect 69099 4927 69141 4936
rect 69196 4976 69236 4985
rect 69292 4976 69332 5608
rect 69388 5648 69428 6271
rect 69388 5396 69428 5608
rect 69484 5648 69524 6616
rect 69675 6488 69717 6497
rect 69675 6448 69676 6488
rect 69716 6448 69717 6488
rect 69675 6439 69717 6448
rect 69676 6354 69716 6439
rect 69772 6329 69812 7120
rect 69868 7160 69908 7699
rect 69868 7111 69908 7120
rect 70060 7160 70100 7169
rect 70156 7160 70196 8548
rect 70348 7916 70388 9547
rect 70444 9428 70484 10051
rect 70444 9379 70484 9388
rect 70540 9353 70580 10060
rect 70635 9680 70677 9689
rect 70635 9640 70636 9680
rect 70676 9640 70677 9680
rect 70635 9631 70677 9640
rect 70636 9546 70676 9631
rect 70539 9344 70581 9353
rect 70539 9304 70540 9344
rect 70580 9304 70581 9344
rect 70539 9295 70581 9304
rect 70636 9260 70676 9269
rect 70636 8681 70676 9220
rect 70732 8756 70772 10303
rect 70828 9605 70868 10648
rect 71019 10436 71061 10445
rect 71019 10396 71020 10436
rect 71060 10396 71061 10436
rect 71019 10387 71061 10396
rect 70923 10184 70965 10193
rect 70923 10144 70924 10184
rect 70964 10144 70965 10184
rect 70923 10135 70965 10144
rect 70924 10050 70964 10135
rect 70827 9596 70869 9605
rect 70827 9556 70828 9596
rect 70868 9556 70869 9596
rect 70827 9547 70869 9556
rect 70828 9512 70868 9547
rect 70828 9462 70868 9472
rect 70923 9512 70965 9521
rect 70923 9472 70924 9512
rect 70964 9472 70965 9512
rect 70923 9463 70965 9472
rect 71020 9512 71060 10387
rect 71116 9689 71156 10900
rect 71115 9680 71157 9689
rect 71115 9640 71116 9680
rect 71156 9640 71157 9680
rect 71115 9631 71157 9640
rect 71020 9463 71060 9472
rect 70924 9378 70964 9463
rect 71212 9344 71252 12487
rect 71308 10856 71348 10865
rect 71308 10193 71348 10816
rect 71404 10697 71444 16192
rect 71499 15644 71541 15653
rect 71499 15604 71500 15644
rect 71540 15604 71541 15644
rect 71499 15595 71541 15604
rect 71500 14057 71540 15595
rect 71595 14720 71637 14729
rect 71595 14680 71596 14720
rect 71636 14680 71637 14720
rect 71595 14671 71637 14680
rect 71499 14048 71541 14057
rect 71499 14008 71500 14048
rect 71540 14008 71541 14048
rect 71499 13999 71541 14008
rect 71596 12980 71636 14671
rect 71596 12965 71732 12980
rect 71596 12956 71733 12965
rect 71596 12940 71692 12956
rect 71691 12916 71692 12940
rect 71732 12916 71733 12956
rect 71691 12907 71733 12916
rect 71692 12545 71732 12907
rect 71788 12797 71828 16192
rect 72172 16232 72212 17116
rect 72455 17072 72495 17472
rect 72745 17156 72785 17472
rect 72268 17032 72495 17072
rect 72556 17116 72785 17156
rect 72268 16484 72308 17032
rect 72268 16435 72308 16444
rect 72172 15737 72212 16192
rect 72556 16232 72596 17116
rect 72855 17072 72895 17472
rect 73145 17156 73185 17472
rect 72652 17032 72895 17072
rect 72940 17116 73185 17156
rect 72652 16484 72692 17032
rect 72652 16435 72692 16444
rect 72940 16232 72980 17116
rect 73255 17072 73295 17472
rect 73545 17240 73585 17472
rect 73036 17032 73295 17072
rect 73420 17200 73585 17240
rect 73036 16484 73076 17032
rect 73420 16988 73460 17200
rect 73655 17072 73695 17472
rect 73945 17156 73985 17472
rect 73036 16435 73076 16444
rect 73324 16948 73460 16988
rect 73516 17032 73695 17072
rect 73900 17116 73985 17156
rect 72556 15821 72596 16192
rect 72748 16192 72940 16232
rect 72555 15812 72597 15821
rect 72555 15772 72556 15812
rect 72596 15772 72597 15812
rect 72555 15763 72597 15772
rect 72171 15728 72213 15737
rect 72171 15688 72172 15728
rect 72212 15688 72213 15728
rect 72171 15679 72213 15688
rect 72748 15653 72788 16192
rect 72940 16183 72980 16192
rect 73131 16232 73173 16241
rect 73131 16192 73132 16232
rect 73172 16192 73173 16232
rect 73131 16183 73173 16192
rect 73324 16232 73364 16948
rect 73420 16484 73460 16493
rect 73516 16484 73556 17032
rect 73460 16444 73556 16484
rect 73420 16416 73460 16444
rect 73708 16232 73748 16241
rect 73900 16232 73940 17116
rect 74055 17072 74095 17472
rect 74345 17156 74385 17472
rect 72747 15644 72789 15653
rect 72747 15604 72748 15644
rect 72788 15604 72789 15644
rect 72747 15595 72789 15604
rect 72652 15392 72692 15401
rect 72171 14552 72213 14561
rect 72171 14512 72172 14552
rect 72212 14512 72213 14552
rect 72171 14503 72213 14512
rect 72172 14132 72212 14503
rect 72172 14083 72212 14092
rect 72556 14048 72596 14057
rect 72652 14048 72692 15352
rect 72748 14972 72788 15595
rect 72748 14923 72788 14932
rect 72596 14008 72692 14048
rect 72556 13999 72596 14008
rect 72076 13376 72116 13385
rect 72116 13336 72692 13376
rect 72076 13327 72116 13336
rect 72652 13208 72692 13336
rect 72652 13159 72692 13168
rect 72267 13124 72309 13133
rect 72267 13084 72268 13124
rect 72308 13084 72309 13124
rect 72267 13075 72309 13084
rect 72268 12990 72308 13075
rect 71787 12788 71829 12797
rect 71787 12748 71788 12788
rect 71828 12748 71829 12788
rect 71787 12739 71829 12748
rect 72843 12704 72885 12713
rect 72843 12664 72844 12704
rect 72884 12664 72885 12704
rect 72843 12655 72885 12664
rect 72844 12570 72884 12655
rect 71691 12536 71733 12545
rect 71691 12496 71692 12536
rect 71732 12496 71733 12536
rect 71691 12487 71733 12496
rect 71692 12402 71732 12487
rect 72940 11696 72980 11705
rect 72556 11612 72596 11621
rect 72556 11201 72596 11572
rect 72555 11192 72597 11201
rect 72555 11152 72556 11192
rect 72596 11152 72597 11192
rect 72555 11143 72597 11152
rect 72940 10856 72980 11656
rect 73036 10856 73076 10865
rect 72940 10816 73036 10856
rect 73036 10807 73076 10816
rect 71403 10688 71445 10697
rect 71403 10648 71404 10688
rect 71444 10648 71445 10688
rect 71403 10639 71445 10648
rect 72939 10436 72981 10445
rect 72939 10396 72940 10436
rect 72980 10396 72981 10436
rect 72939 10387 72981 10396
rect 72940 10302 72980 10387
rect 71307 10184 71349 10193
rect 71307 10144 71308 10184
rect 71348 10144 71349 10184
rect 71307 10135 71349 10144
rect 71788 10184 71828 10193
rect 71788 10109 71828 10144
rect 71787 10100 71829 10109
rect 71787 10060 71788 10100
rect 71828 10060 71829 10100
rect 71787 10051 71829 10060
rect 72843 10100 72885 10109
rect 72843 10060 72844 10100
rect 72884 10060 72885 10100
rect 72843 10051 72885 10060
rect 71788 9941 71828 10051
rect 71787 9932 71829 9941
rect 71787 9892 71788 9932
rect 71828 9892 71829 9932
rect 71787 9883 71829 9892
rect 71979 9680 72021 9689
rect 71979 9640 71980 9680
rect 72020 9640 72021 9680
rect 71979 9631 72021 9640
rect 71307 9596 71349 9605
rect 71307 9556 71308 9596
rect 71348 9556 71349 9596
rect 71307 9547 71349 9556
rect 71308 9512 71348 9547
rect 71308 9461 71348 9472
rect 71500 9512 71540 9521
rect 71020 9304 71252 9344
rect 71307 9344 71349 9353
rect 71307 9304 71308 9344
rect 71348 9304 71349 9344
rect 70732 8716 70868 8756
rect 70635 8672 70677 8681
rect 70635 8632 70636 8672
rect 70676 8632 70677 8672
rect 70635 8623 70677 8632
rect 70828 8672 70868 8716
rect 70731 8588 70773 8597
rect 70731 8548 70732 8588
rect 70772 8548 70773 8588
rect 70731 8539 70773 8548
rect 70732 8168 70772 8539
rect 70732 8119 70772 8128
rect 70100 7120 70196 7160
rect 70252 7876 70388 7916
rect 70252 7160 70292 7876
rect 70347 7748 70389 7757
rect 70347 7708 70348 7748
rect 70388 7708 70389 7748
rect 70347 7699 70389 7708
rect 70731 7748 70773 7757
rect 70731 7708 70732 7748
rect 70772 7708 70773 7748
rect 70731 7699 70773 7708
rect 70348 7179 70388 7699
rect 70732 7614 70772 7699
rect 70348 7130 70388 7139
rect 70443 7160 70485 7169
rect 69963 7076 70005 7085
rect 69963 7036 69964 7076
rect 70004 7036 70005 7076
rect 69963 7027 70005 7036
rect 69771 6320 69813 6329
rect 69771 6280 69772 6320
rect 69812 6280 69813 6320
rect 69771 6271 69813 6280
rect 69771 5900 69813 5909
rect 69771 5860 69772 5900
rect 69812 5860 69813 5900
rect 69771 5851 69813 5860
rect 69772 5766 69812 5851
rect 69484 5480 69524 5608
rect 69580 5648 69620 5657
rect 69772 5648 69812 5657
rect 69620 5608 69772 5648
rect 69580 5599 69620 5608
rect 69772 5599 69812 5608
rect 69964 5648 70004 7027
rect 70060 6917 70100 7120
rect 70252 7076 70292 7120
rect 70443 7120 70444 7160
rect 70484 7120 70485 7160
rect 70443 7111 70485 7120
rect 70252 7036 70388 7076
rect 70156 6992 70196 7001
rect 70059 6908 70101 6917
rect 70059 6868 70060 6908
rect 70100 6868 70101 6908
rect 70059 6859 70101 6868
rect 69964 5599 70004 5608
rect 70060 5648 70100 5657
rect 70156 5648 70196 6952
rect 70251 6908 70293 6917
rect 70251 6868 70252 6908
rect 70292 6868 70293 6908
rect 70251 6859 70293 6868
rect 70100 5608 70196 5648
rect 70060 5599 70100 5608
rect 69484 5440 69908 5480
rect 69388 5356 69524 5396
rect 69236 4936 69332 4976
rect 69196 4927 69236 4936
rect 69100 4842 69140 4927
rect 69388 4808 69428 4817
rect 69003 4556 69045 4565
rect 69003 4516 69004 4556
rect 69044 4516 69045 4556
rect 69003 4507 69045 4516
rect 68907 4472 68949 4481
rect 68907 4432 68908 4472
rect 68948 4432 68949 4472
rect 68907 4423 68949 4432
rect 68811 4304 68853 4313
rect 68811 4264 68812 4304
rect 68852 4264 68853 4304
rect 68811 4255 68853 4264
rect 68812 4170 68852 4255
rect 68716 3053 68756 3424
rect 68908 3464 68948 4423
rect 69388 4136 69428 4768
rect 69484 4229 69524 5356
rect 69483 4220 69525 4229
rect 69483 4180 69484 4220
rect 69524 4180 69525 4220
rect 69483 4171 69525 4180
rect 69388 4087 69428 4096
rect 69004 4052 69044 4061
rect 69004 3641 69044 4012
rect 69291 4052 69333 4061
rect 69291 4012 69292 4052
rect 69332 4012 69333 4052
rect 69291 4003 69333 4012
rect 69003 3632 69045 3641
rect 69003 3592 69004 3632
rect 69044 3592 69045 3632
rect 69003 3583 69045 3592
rect 68908 3415 68948 3424
rect 69196 3464 69236 3473
rect 68908 3296 68948 3305
rect 69196 3296 69236 3424
rect 69292 3464 69332 4003
rect 69387 3632 69429 3641
rect 69387 3592 69388 3632
rect 69428 3592 69429 3632
rect 69387 3583 69429 3592
rect 69388 3498 69428 3583
rect 69868 3473 69908 5440
rect 70252 4565 70292 6859
rect 70348 4985 70388 7036
rect 70444 6488 70484 7111
rect 70540 6488 70580 6497
rect 70444 6448 70540 6488
rect 70347 4976 70389 4985
rect 70347 4936 70348 4976
rect 70388 4936 70389 4976
rect 70347 4927 70389 4936
rect 70251 4556 70293 4565
rect 70251 4516 70252 4556
rect 70292 4516 70293 4556
rect 70251 4507 70293 4516
rect 69963 4220 70005 4229
rect 69963 4180 69964 4220
rect 70004 4180 70005 4220
rect 69963 4171 70005 4180
rect 69292 3415 69332 3424
rect 69484 3464 69524 3473
rect 69772 3464 69812 3473
rect 69524 3424 69772 3464
rect 69484 3415 69524 3424
rect 69772 3415 69812 3424
rect 69867 3464 69909 3473
rect 69867 3424 69868 3464
rect 69908 3424 69909 3464
rect 69867 3415 69909 3424
rect 69964 3464 70004 4171
rect 70252 4136 70292 4145
rect 68948 3256 69236 3296
rect 68908 3247 68948 3256
rect 68907 3128 68949 3137
rect 68907 3088 68908 3128
rect 68948 3088 68949 3128
rect 68907 3079 68949 3088
rect 68715 3044 68757 3053
rect 68715 3004 68716 3044
rect 68756 3004 68757 3044
rect 68715 2995 68757 3004
rect 68908 2900 68948 3079
rect 69868 3053 69908 3415
rect 69964 3221 70004 3424
rect 70059 3464 70101 3473
rect 70059 3424 70060 3464
rect 70100 3424 70101 3464
rect 70059 3415 70101 3424
rect 70060 3330 70100 3415
rect 69963 3212 70005 3221
rect 69963 3172 69964 3212
rect 70004 3172 70005 3212
rect 69963 3163 70005 3172
rect 69003 3044 69045 3053
rect 69003 3004 69004 3044
rect 69044 3004 69045 3044
rect 69003 2995 69045 3004
rect 69867 3044 69909 3053
rect 69867 3004 69868 3044
rect 69908 3004 69909 3044
rect 69867 2995 69909 3004
rect 68332 2575 68372 2584
rect 68428 2860 68660 2900
rect 68812 2860 68948 2900
rect 68428 2624 68468 2860
rect 68716 2792 68756 2801
rect 68139 2456 68181 2465
rect 68139 2416 68140 2456
rect 68180 2416 68181 2456
rect 68139 2407 68181 2416
rect 68140 2322 68180 2407
rect 68235 2120 68277 2129
rect 68235 2080 68236 2120
rect 68276 2080 68277 2120
rect 68235 2071 68277 2080
rect 68236 1952 68276 2071
rect 68236 1903 68276 1912
rect 68332 1952 68372 1961
rect 68428 1952 68468 2584
rect 68524 2752 68716 2792
rect 68524 2045 68564 2752
rect 68716 2743 68756 2752
rect 68620 2624 68660 2633
rect 68523 2036 68565 2045
rect 68523 1996 68524 2036
rect 68564 1996 68565 2036
rect 68523 1987 68565 1996
rect 68372 1912 68468 1952
rect 68332 1903 68372 1912
rect 67372 1700 67412 1709
rect 67372 1121 67412 1660
rect 68043 1700 68085 1709
rect 68043 1660 68044 1700
rect 68084 1660 68085 1700
rect 68043 1651 68085 1660
rect 68428 1364 68468 1912
rect 68428 1315 68468 1324
rect 66412 1063 66452 1072
rect 67276 1063 67316 1072
rect 67371 1112 67413 1121
rect 67371 1072 67372 1112
rect 67412 1072 67413 1112
rect 67371 1063 67413 1072
rect 64203 1028 64245 1037
rect 64203 988 64204 1028
rect 64244 988 64245 1028
rect 64203 979 64245 988
rect 66028 978 66068 1063
rect 58580 904 58964 944
rect 68524 944 68564 1987
rect 68620 1784 68660 2584
rect 68812 2624 68852 2860
rect 68812 2575 68852 2584
rect 69004 2624 69044 2995
rect 69004 2575 69044 2584
rect 69196 2624 69236 2633
rect 69100 2540 69140 2549
rect 69100 2120 69140 2500
rect 69196 2129 69236 2584
rect 68620 1735 68660 1744
rect 68716 2080 69140 2120
rect 69195 2120 69237 2129
rect 69195 2080 69196 2120
rect 69236 2080 69237 2120
rect 68716 1616 68756 2080
rect 69195 2071 69237 2080
rect 70252 1961 70292 4096
rect 68620 1576 68756 1616
rect 68812 1952 68852 1961
rect 68620 1112 68660 1576
rect 68812 1364 68852 1912
rect 69196 1952 69236 1961
rect 70059 1952 70101 1961
rect 69236 1912 69332 1952
rect 69196 1903 69236 1912
rect 69003 1868 69045 1877
rect 69003 1828 69004 1868
rect 69044 1828 69045 1868
rect 69003 1819 69045 1828
rect 68908 1364 68948 1373
rect 68812 1324 68908 1364
rect 68908 1315 68948 1324
rect 68620 1063 68660 1072
rect 68716 1112 68756 1121
rect 68716 944 68756 1072
rect 68908 1112 68948 1121
rect 69004 1112 69044 1819
rect 69292 1280 69332 1912
rect 70059 1912 70060 1952
rect 70100 1912 70101 1952
rect 70059 1903 70101 1912
rect 70251 1952 70293 1961
rect 70251 1912 70252 1952
rect 70292 1912 70293 1952
rect 70251 1903 70293 1912
rect 70060 1818 70100 1903
rect 70444 1364 70484 6448
rect 70540 6439 70580 6448
rect 70828 5825 70868 8632
rect 70923 8672 70965 8681
rect 70923 8632 70924 8672
rect 70964 8632 70965 8672
rect 70923 8623 70965 8632
rect 70924 7169 70964 8623
rect 70923 7160 70965 7169
rect 70923 7120 70924 7160
rect 70964 7120 70965 7160
rect 70923 7111 70965 7120
rect 70827 5816 70869 5825
rect 70827 5776 70828 5816
rect 70868 5776 70869 5816
rect 70827 5767 70869 5776
rect 70828 3557 70868 5767
rect 70827 3548 70869 3557
rect 70827 3508 70828 3548
rect 70868 3508 70869 3548
rect 70827 3499 70869 3508
rect 70444 1315 70484 1324
rect 69292 1231 69332 1240
rect 70923 1280 70965 1289
rect 70923 1240 70924 1280
rect 70964 1240 70965 1280
rect 70923 1231 70965 1240
rect 68948 1072 69044 1112
rect 69771 1112 69813 1121
rect 69771 1072 69772 1112
rect 69812 1072 69813 1112
rect 68908 1063 68948 1072
rect 69771 1063 69813 1072
rect 70924 1112 70964 1231
rect 71020 1121 71060 9304
rect 71307 9295 71349 9304
rect 71115 8672 71157 8681
rect 71115 8632 71116 8672
rect 71156 8632 71157 8672
rect 71115 8623 71157 8632
rect 71116 8538 71156 8623
rect 71211 8588 71253 8597
rect 71211 8548 71212 8588
rect 71252 8548 71253 8588
rect 71211 8539 71253 8548
rect 71212 8454 71252 8539
rect 71308 8000 71348 9295
rect 71404 9260 71444 9269
rect 71404 8765 71444 9220
rect 71500 8924 71540 9472
rect 71692 9512 71732 9523
rect 71692 9437 71732 9472
rect 71883 9512 71925 9521
rect 71883 9472 71884 9512
rect 71924 9472 71925 9512
rect 71883 9463 71925 9472
rect 71691 9428 71733 9437
rect 71691 9388 71692 9428
rect 71732 9388 71733 9428
rect 71691 9379 71733 9388
rect 71500 8875 71540 8884
rect 71788 9260 71828 9269
rect 71403 8756 71445 8765
rect 71403 8716 71404 8756
rect 71444 8716 71445 8756
rect 71403 8707 71445 8716
rect 71404 8177 71444 8707
rect 71692 8588 71732 8597
rect 71500 8548 71692 8588
rect 71403 8168 71445 8177
rect 71403 8128 71404 8168
rect 71444 8128 71445 8168
rect 71403 8119 71445 8128
rect 71500 8168 71540 8548
rect 71692 8539 71732 8548
rect 71500 8119 71540 8128
rect 71404 8000 71444 8009
rect 71595 8000 71637 8009
rect 71308 7960 71404 8000
rect 71444 7960 71540 8000
rect 71404 7951 71444 7960
rect 71212 7160 71252 7169
rect 71116 5900 71156 5909
rect 71212 5900 71252 7120
rect 71403 7160 71445 7169
rect 71403 7120 71404 7160
rect 71444 7120 71445 7160
rect 71500 7160 71540 7960
rect 71595 7960 71596 8000
rect 71636 7960 71637 8000
rect 71595 7951 71637 7960
rect 71692 8000 71732 8009
rect 71788 8000 71828 9220
rect 71884 8681 71924 9463
rect 71980 9437 72020 9631
rect 71979 9428 72021 9437
rect 71979 9388 71980 9428
rect 72020 9388 72021 9428
rect 71979 9379 72021 9388
rect 71883 8672 71925 8681
rect 71883 8632 71884 8672
rect 71924 8632 71925 8672
rect 71883 8623 71925 8632
rect 71732 7960 71828 8000
rect 71692 7951 71732 7960
rect 71596 7866 71636 7951
rect 71596 7160 71636 7169
rect 71500 7120 71596 7160
rect 71403 7111 71445 7120
rect 71307 7076 71349 7085
rect 71307 7036 71308 7076
rect 71348 7036 71349 7076
rect 71307 7027 71349 7036
rect 71308 6942 71348 7027
rect 71404 6404 71444 7111
rect 71156 5860 71252 5900
rect 71308 6364 71444 6404
rect 71116 5851 71156 5860
rect 71115 4976 71157 4985
rect 71115 4936 71116 4976
rect 71156 4936 71157 4976
rect 71115 4927 71157 4936
rect 71116 1877 71156 4927
rect 71308 4724 71348 6364
rect 71403 5732 71445 5741
rect 71403 5692 71404 5732
rect 71444 5692 71445 5732
rect 71403 5683 71445 5692
rect 71404 5648 71444 5683
rect 71404 5597 71444 5608
rect 71499 5648 71541 5657
rect 71499 5608 71500 5648
rect 71540 5608 71541 5648
rect 71499 5599 71541 5608
rect 71500 5514 71540 5599
rect 71596 4985 71636 7120
rect 71788 7160 71828 7171
rect 71788 7085 71828 7120
rect 71883 7160 71925 7169
rect 71883 7120 71884 7160
rect 71924 7120 71925 7160
rect 71883 7111 71925 7120
rect 71787 7076 71829 7085
rect 71787 7036 71788 7076
rect 71828 7036 71829 7076
rect 71787 7027 71829 7036
rect 71884 7026 71924 7111
rect 71692 6992 71732 7001
rect 71692 6572 71732 6952
rect 71884 6572 71924 6581
rect 71692 6532 71884 6572
rect 71884 6523 71924 6532
rect 71692 6236 71732 6245
rect 71692 5741 71732 6196
rect 71787 5816 71829 5825
rect 71787 5776 71788 5816
rect 71828 5776 71829 5816
rect 71787 5767 71829 5776
rect 71691 5732 71733 5741
rect 71691 5692 71692 5732
rect 71732 5692 71733 5732
rect 71691 5683 71733 5692
rect 71788 5648 71828 5767
rect 71980 5648 72020 9379
rect 72172 9344 72212 9353
rect 72076 8672 72116 8681
rect 72172 8672 72212 9304
rect 72116 8632 72212 8672
rect 72844 8672 72884 10051
rect 72940 8672 72980 8681
rect 72844 8632 72940 8672
rect 72076 8623 72116 8632
rect 72940 8623 72980 8632
rect 73132 8084 73172 16183
rect 73324 12713 73364 16192
rect 73516 16192 73708 16232
rect 73748 16192 73940 16232
rect 73996 17032 74095 17072
rect 74188 17116 74385 17156
rect 73516 14300 73556 16192
rect 73708 16183 73748 16192
rect 73804 16064 73844 16073
rect 73996 16064 74036 17032
rect 74188 16232 74228 17116
rect 74455 17072 74495 17472
rect 74745 17072 74785 17472
rect 74284 17032 74495 17072
rect 74572 17032 74785 17072
rect 74855 17072 74895 17472
rect 75145 17156 75185 17472
rect 74956 17116 75185 17156
rect 74855 17032 74900 17072
rect 74284 16484 74324 17032
rect 74284 16435 74324 16444
rect 74572 16232 74612 17032
rect 74668 16484 74708 16493
rect 74860 16484 74900 17032
rect 74708 16444 74900 16484
rect 74668 16435 74708 16444
rect 74956 16241 74996 17116
rect 75255 17072 75295 17472
rect 75545 17156 75585 17472
rect 75052 17032 75295 17072
rect 75340 17116 75585 17156
rect 75052 16484 75092 17032
rect 75052 16435 75092 16444
rect 74228 16192 74516 16232
rect 74188 16183 74228 16192
rect 73844 16024 74036 16064
rect 73804 16015 73844 16024
rect 74283 15392 74325 15401
rect 74283 15352 74284 15392
rect 74324 15352 74325 15392
rect 74283 15343 74325 15352
rect 73612 14848 74132 14888
rect 73612 14720 73652 14848
rect 73612 14671 73652 14680
rect 73803 14720 73845 14729
rect 73803 14680 73804 14720
rect 73844 14680 73845 14720
rect 73803 14671 73845 14680
rect 73900 14720 73940 14729
rect 73804 14586 73844 14671
rect 73900 14561 73940 14680
rect 74092 14720 74132 14848
rect 74092 14671 74132 14680
rect 74188 14720 74228 14729
rect 73707 14552 73749 14561
rect 73707 14512 73708 14552
rect 73748 14512 73749 14552
rect 73707 14503 73749 14512
rect 73899 14552 73941 14561
rect 73899 14512 73900 14552
rect 73940 14512 73941 14552
rect 73899 14503 73941 14512
rect 73708 14418 73748 14503
rect 74188 14393 74228 14680
rect 74284 14720 74324 15343
rect 74284 14671 74324 14680
rect 74380 14720 74420 14729
rect 74380 14645 74420 14680
rect 74379 14636 74421 14645
rect 74379 14596 74380 14636
rect 74420 14596 74421 14636
rect 74379 14587 74421 14596
rect 74380 14393 74420 14587
rect 74187 14384 74229 14393
rect 74187 14344 74188 14384
rect 74228 14344 74229 14384
rect 74187 14335 74229 14344
rect 74379 14384 74421 14393
rect 74379 14344 74380 14384
rect 74420 14344 74421 14384
rect 74379 14335 74421 14344
rect 73516 14260 73748 14300
rect 73445 14048 73485 14057
rect 73445 13292 73485 14008
rect 73611 13628 73653 13637
rect 73611 13588 73612 13628
rect 73652 13588 73653 13628
rect 73611 13579 73653 13588
rect 73445 13252 73523 13292
rect 73483 13217 73523 13252
rect 73483 13208 73556 13217
rect 73483 13168 73516 13208
rect 73516 12965 73556 13168
rect 73515 12956 73557 12965
rect 73515 12916 73516 12956
rect 73556 12916 73557 12956
rect 73515 12907 73557 12916
rect 73323 12704 73365 12713
rect 73323 12664 73324 12704
rect 73364 12664 73365 12704
rect 73323 12655 73365 12664
rect 73516 11696 73556 12907
rect 73612 11864 73652 13579
rect 73708 12980 73748 14260
rect 74476 14132 74516 16192
rect 74092 14092 74516 14132
rect 73708 12940 74036 12980
rect 73612 11824 73940 11864
rect 73804 11696 73844 11705
rect 73516 11656 73804 11696
rect 73804 11647 73844 11656
rect 73900 10352 73940 11824
rect 73996 10445 74036 12940
rect 73995 10436 74037 10445
rect 73995 10396 73996 10436
rect 74036 10396 74037 10436
rect 73995 10387 74037 10396
rect 73708 10312 73940 10352
rect 73516 10100 73556 10109
rect 73516 9185 73556 10060
rect 73515 9176 73557 9185
rect 73515 9136 73516 9176
rect 73556 9136 73557 9176
rect 73515 9127 73557 9136
rect 72940 8044 73172 8084
rect 73611 8084 73653 8093
rect 73611 8044 73612 8084
rect 73652 8044 73653 8084
rect 72364 7328 72404 7337
rect 72171 7160 72213 7169
rect 72171 7120 72172 7160
rect 72212 7120 72213 7160
rect 72171 7111 72213 7120
rect 72172 5732 72212 7111
rect 72268 6488 72308 6497
rect 72364 6488 72404 7288
rect 72308 6448 72404 6488
rect 72268 6439 72308 6448
rect 72172 5683 72212 5692
rect 72076 5648 72116 5657
rect 71980 5608 72076 5648
rect 71788 5599 71828 5608
rect 72076 5599 72116 5608
rect 72267 5648 72309 5657
rect 72267 5608 72268 5648
rect 72308 5608 72309 5648
rect 72267 5599 72309 5608
rect 72268 5514 72308 5599
rect 71692 5144 71732 5153
rect 71732 5104 72020 5144
rect 71692 5095 71732 5104
rect 71595 4976 71637 4985
rect 71788 4976 71828 4985
rect 71595 4936 71596 4976
rect 71636 4936 71637 4976
rect 71595 4927 71637 4936
rect 71692 4936 71788 4976
rect 71596 4842 71636 4927
rect 71308 4684 71636 4724
rect 71499 4304 71541 4313
rect 71499 4264 71500 4304
rect 71540 4264 71541 4304
rect 71499 4255 71541 4264
rect 71404 3968 71444 3977
rect 71211 3548 71253 3557
rect 71211 3508 71212 3548
rect 71252 3508 71253 3548
rect 71211 3499 71253 3508
rect 71212 3464 71252 3499
rect 71404 3473 71444 3928
rect 71212 2633 71252 3424
rect 71403 3464 71445 3473
rect 71403 3424 71404 3464
rect 71444 3424 71445 3464
rect 71403 3415 71445 3424
rect 71500 3464 71540 4255
rect 71596 4136 71636 4684
rect 71596 3800 71636 4096
rect 71692 4061 71732 4936
rect 71788 4927 71828 4936
rect 71883 4976 71925 4985
rect 71883 4936 71884 4976
rect 71924 4936 71925 4976
rect 71883 4927 71925 4936
rect 71884 4842 71924 4927
rect 71788 4136 71828 4145
rect 71691 4052 71733 4061
rect 71691 4012 71692 4052
rect 71732 4012 71733 4052
rect 71691 4003 71733 4012
rect 71692 3918 71732 4003
rect 71596 3760 71732 3800
rect 71500 3415 71540 3424
rect 71595 3464 71637 3473
rect 71595 3424 71596 3464
rect 71636 3424 71637 3464
rect 71595 3415 71637 3424
rect 71596 3330 71636 3415
rect 71692 3137 71732 3760
rect 71788 3296 71828 4096
rect 71980 4136 72020 5104
rect 72075 5060 72117 5069
rect 72075 5020 72076 5060
rect 72116 5020 72117 5060
rect 72075 5011 72117 5020
rect 72076 4976 72116 5011
rect 72076 4724 72116 4936
rect 72171 4976 72213 4985
rect 72171 4936 72172 4976
rect 72212 4936 72213 4976
rect 72171 4927 72213 4936
rect 72268 4976 72308 4985
rect 72172 4842 72212 4927
rect 72076 4684 72212 4724
rect 71980 4087 72020 4096
rect 72075 3464 72117 3473
rect 72075 3424 72076 3464
rect 72116 3424 72117 3464
rect 72075 3415 72117 3424
rect 72172 3464 72212 4684
rect 72268 4397 72308 4936
rect 72460 4808 72500 4817
rect 72364 4768 72460 4808
rect 72267 4388 72309 4397
rect 72267 4348 72268 4388
rect 72308 4348 72309 4388
rect 72267 4339 72309 4348
rect 72364 4136 72404 4768
rect 72460 4759 72500 4768
rect 72459 4556 72501 4565
rect 72459 4516 72460 4556
rect 72500 4516 72501 4556
rect 72459 4507 72501 4516
rect 72460 4397 72500 4507
rect 72459 4388 72501 4397
rect 72459 4348 72460 4388
rect 72500 4348 72501 4388
rect 72459 4339 72501 4348
rect 72364 4087 72404 4096
rect 72172 3415 72212 3424
rect 72364 3464 72404 3473
rect 72460 3464 72500 4339
rect 72404 3424 72500 3464
rect 72364 3415 72404 3424
rect 72076 3330 72116 3415
rect 71884 3296 71924 3305
rect 71788 3256 71884 3296
rect 71884 3247 71924 3256
rect 71979 3212 72021 3221
rect 71979 3172 71980 3212
rect 72020 3172 72021 3212
rect 71979 3163 72021 3172
rect 72364 3212 72404 3221
rect 71691 3128 71733 3137
rect 71691 3088 71692 3128
rect 71732 3088 71733 3128
rect 71691 3079 71733 3088
rect 71787 3044 71829 3053
rect 71787 3004 71788 3044
rect 71828 3004 71829 3044
rect 71787 2995 71829 3004
rect 71500 2792 71540 2801
rect 71211 2624 71253 2633
rect 71211 2584 71212 2624
rect 71252 2584 71253 2624
rect 71211 2575 71253 2584
rect 71211 2120 71253 2129
rect 71211 2080 71212 2120
rect 71252 2080 71253 2120
rect 71211 2071 71253 2080
rect 71212 1986 71252 2071
rect 71404 1952 71444 1961
rect 71500 1952 71540 2752
rect 71788 2624 71828 2995
rect 71980 2900 72020 3163
rect 71788 2575 71828 2584
rect 71884 2860 72020 2900
rect 72364 2900 72404 3172
rect 72940 2900 72980 8044
rect 73611 8035 73653 8044
rect 73612 7950 73652 8035
rect 73035 7916 73077 7925
rect 73035 7876 73036 7916
rect 73076 7876 73077 7916
rect 73035 7867 73077 7876
rect 73036 6320 73076 7867
rect 73132 6488 73172 6497
rect 73172 6448 73268 6488
rect 73132 6439 73172 6448
rect 73036 6280 73172 6320
rect 73132 2900 73172 6280
rect 73228 4136 73268 6448
rect 73611 5564 73653 5573
rect 73611 5524 73612 5564
rect 73652 5524 73653 5564
rect 73611 5515 73653 5524
rect 73612 5430 73652 5515
rect 73268 4096 73364 4136
rect 73228 4087 73268 4096
rect 72267 2876 72309 2885
rect 71884 2624 71924 2860
rect 72267 2836 72268 2876
rect 72308 2836 72309 2876
rect 72364 2860 72788 2900
rect 72940 2860 73076 2900
rect 73132 2860 73268 2900
rect 72267 2827 72309 2836
rect 71884 2575 71924 2584
rect 71979 2624 72021 2633
rect 71979 2584 71980 2624
rect 72020 2584 72021 2624
rect 71979 2575 72021 2584
rect 72268 2624 72308 2827
rect 71980 2490 72020 2575
rect 72268 2549 72308 2584
rect 72556 2624 72596 2633
rect 72267 2540 72309 2549
rect 72267 2500 72268 2540
rect 72308 2500 72309 2540
rect 72267 2491 72309 2500
rect 71692 2456 71732 2465
rect 71732 2416 71924 2456
rect 71692 2407 71732 2416
rect 71788 1952 71828 1961
rect 71500 1912 71788 1952
rect 71115 1868 71157 1877
rect 71115 1828 71116 1868
rect 71156 1828 71157 1868
rect 71115 1819 71157 1828
rect 71404 1373 71444 1912
rect 71788 1903 71828 1912
rect 71403 1364 71445 1373
rect 71403 1324 71404 1364
rect 71444 1324 71445 1364
rect 71403 1315 71445 1324
rect 71884 1121 71924 2416
rect 72556 2213 72596 2584
rect 72651 2624 72693 2633
rect 72651 2584 72652 2624
rect 72692 2584 72693 2624
rect 72651 2575 72693 2584
rect 72652 2490 72692 2575
rect 72555 2204 72597 2213
rect 72555 2164 72556 2204
rect 72596 2164 72597 2204
rect 72555 2155 72597 2164
rect 72651 1952 72693 1961
rect 72651 1912 72652 1952
rect 72692 1912 72693 1952
rect 72651 1903 72693 1912
rect 72652 1818 72692 1903
rect 72459 1364 72501 1373
rect 72459 1324 72460 1364
rect 72500 1324 72501 1364
rect 72459 1315 72501 1324
rect 72075 1280 72117 1289
rect 72075 1240 72076 1280
rect 72116 1240 72117 1280
rect 72075 1231 72117 1240
rect 70924 1063 70964 1072
rect 71019 1112 71061 1121
rect 71019 1072 71020 1112
rect 71060 1072 71061 1112
rect 71019 1063 71061 1072
rect 71211 1112 71253 1121
rect 71211 1072 71212 1112
rect 71252 1072 71253 1112
rect 71211 1063 71253 1072
rect 71883 1112 71925 1121
rect 71883 1072 71884 1112
rect 71924 1072 71925 1112
rect 71883 1063 71925 1072
rect 72076 1112 72116 1231
rect 72460 1230 72500 1315
rect 72076 1063 72116 1072
rect 72459 1112 72501 1121
rect 72459 1072 72460 1112
rect 72500 1072 72501 1112
rect 72459 1063 72501 1072
rect 72651 1112 72693 1121
rect 72651 1072 72652 1112
rect 72692 1072 72693 1112
rect 72651 1063 72693 1072
rect 72748 1112 72788 2860
rect 72939 2792 72981 2801
rect 72939 2752 72940 2792
rect 72980 2752 72981 2792
rect 72939 2743 72981 2752
rect 72940 2658 72980 2743
rect 73036 2129 73076 2860
rect 73131 2708 73173 2717
rect 73131 2668 73132 2708
rect 73172 2668 73173 2708
rect 73131 2659 73173 2668
rect 73132 2213 73172 2659
rect 73228 2624 73268 2860
rect 73131 2204 73173 2213
rect 73131 2164 73132 2204
rect 73172 2164 73173 2204
rect 73131 2155 73173 2164
rect 73035 2120 73077 2129
rect 73035 2080 73036 2120
rect 73076 2080 73077 2120
rect 73035 2071 73077 2080
rect 72748 1063 72788 1072
rect 69772 978 69812 1063
rect 71212 978 71252 1063
rect 72460 978 72500 1063
rect 72652 978 72692 1063
rect 68524 904 68756 944
rect 73132 944 73172 2155
rect 73228 1289 73268 2584
rect 73324 2876 73364 4096
rect 73708 2900 73748 10312
rect 73900 10184 73940 10193
rect 73940 10144 74036 10184
rect 73900 10135 73940 10144
rect 73996 9344 74036 10144
rect 74092 9521 74132 14092
rect 74572 13964 74612 16192
rect 74955 16232 74997 16241
rect 74955 16192 74956 16232
rect 74996 16192 74997 16232
rect 74955 16183 74997 16192
rect 75340 16232 75380 17116
rect 75655 17072 75695 17472
rect 75945 17240 75985 17472
rect 75436 17032 75695 17072
rect 75820 17200 75985 17240
rect 75436 16484 75476 17032
rect 75436 16435 75476 16444
rect 75724 16232 75764 16241
rect 75820 16232 75860 17200
rect 76055 17072 76095 17472
rect 76345 17072 76385 17472
rect 75380 16192 75476 16232
rect 75340 16183 75380 16192
rect 74956 16098 74996 16183
rect 75147 15560 75189 15569
rect 75147 15520 75148 15560
rect 75188 15520 75189 15560
rect 75147 15511 75189 15520
rect 75340 15560 75380 15569
rect 75148 15426 75188 15511
rect 74667 15308 74709 15317
rect 74667 15268 74668 15308
rect 74708 15268 74709 15308
rect 74667 15259 74709 15268
rect 75244 15308 75284 15317
rect 74668 14720 74708 15259
rect 74763 14804 74805 14813
rect 74763 14764 74764 14804
rect 74804 14764 74805 14804
rect 74763 14755 74805 14764
rect 74668 14671 74708 14680
rect 74667 14552 74709 14561
rect 74667 14512 74668 14552
rect 74708 14512 74709 14552
rect 74667 14503 74709 14512
rect 74188 13924 74612 13964
rect 74091 9512 74133 9521
rect 74091 9472 74092 9512
rect 74132 9472 74133 9512
rect 74091 9463 74133 9472
rect 73996 9295 74036 9304
rect 74092 8924 74132 9463
rect 74188 9008 74228 13924
rect 74668 13880 74708 14503
rect 74764 14048 74804 14755
rect 75244 14729 75284 15268
rect 75340 14972 75380 15520
rect 75340 14923 75380 14932
rect 75436 14804 75476 16192
rect 75628 16192 75724 16232
rect 75764 16192 75860 16232
rect 76012 17032 76095 17072
rect 76300 17032 76385 17072
rect 76455 17072 76495 17472
rect 76455 17032 76532 17072
rect 75532 14897 75572 14982
rect 75531 14888 75573 14897
rect 75531 14848 75532 14888
rect 75572 14848 75573 14888
rect 75531 14839 75573 14848
rect 75340 14764 75476 14804
rect 74956 14720 74996 14729
rect 74956 14561 74996 14680
rect 75243 14720 75285 14729
rect 75243 14680 75244 14720
rect 75284 14680 75285 14720
rect 75243 14671 75285 14680
rect 75051 14636 75093 14645
rect 75051 14596 75052 14636
rect 75092 14596 75093 14636
rect 75051 14587 75093 14596
rect 74955 14552 74997 14561
rect 74955 14512 74956 14552
rect 74996 14512 74997 14552
rect 74955 14503 74997 14512
rect 75052 14502 75092 14587
rect 74764 13999 74804 14008
rect 74955 14048 74997 14057
rect 74955 14008 74956 14048
rect 74996 14008 74997 14048
rect 74955 13999 74997 14008
rect 75052 14048 75092 14057
rect 75243 14048 75285 14057
rect 75092 14008 75188 14048
rect 75052 13999 75092 14008
rect 74956 13914 74996 13999
rect 74764 13880 74804 13889
rect 74668 13840 74764 13880
rect 74764 13831 74804 13840
rect 74571 13796 74613 13805
rect 74571 13756 74572 13796
rect 74612 13756 74613 13796
rect 74571 13747 74613 13756
rect 74572 13662 74612 13747
rect 74668 13292 74708 13303
rect 74668 13217 74708 13252
rect 74764 13252 74996 13292
rect 74667 13208 74709 13217
rect 74667 13168 74668 13208
rect 74708 13168 74709 13208
rect 74667 13159 74709 13168
rect 74379 13124 74421 13133
rect 74379 13084 74380 13124
rect 74420 13084 74421 13124
rect 74379 13075 74421 13084
rect 74283 13040 74325 13049
rect 74283 13000 74284 13040
rect 74324 13000 74325 13040
rect 74283 12991 74325 13000
rect 74284 12536 74324 12991
rect 74380 12704 74420 13075
rect 74764 12980 74804 13252
rect 74956 13208 74996 13252
rect 75148 13217 75188 14008
rect 75243 14008 75244 14048
rect 75284 14008 75285 14048
rect 75243 13999 75285 14008
rect 74956 13159 74996 13168
rect 75052 13208 75092 13217
rect 74860 13049 74900 13134
rect 74859 13040 74901 13049
rect 74963 13040 75005 13049
rect 74859 13000 74860 13040
rect 74900 13000 74901 13040
rect 74859 12991 74901 13000
rect 74956 13000 74964 13040
rect 75004 13000 75005 13040
rect 74956 12991 75005 13000
rect 74668 12940 74804 12980
rect 74380 12655 74420 12664
rect 74475 12704 74517 12713
rect 74475 12664 74476 12704
rect 74516 12664 74517 12704
rect 74475 12655 74517 12664
rect 74284 12487 74324 12496
rect 74476 12536 74516 12655
rect 74476 12487 74516 12496
rect 74572 12536 74612 12545
rect 74572 12377 74612 12496
rect 74571 12368 74613 12377
rect 74571 12328 74572 12368
rect 74612 12328 74613 12368
rect 74571 12319 74613 12328
rect 74668 11192 74708 12940
rect 74763 12620 74805 12629
rect 74763 12580 74764 12620
rect 74804 12580 74805 12620
rect 74763 12571 74805 12580
rect 74764 12536 74804 12571
rect 74764 12485 74804 12496
rect 74956 12536 74996 12991
rect 75052 12797 75092 13168
rect 75147 13208 75189 13217
rect 75147 13168 75148 13208
rect 75188 13168 75189 13208
rect 75147 13159 75189 13168
rect 75148 13074 75188 13159
rect 75244 13133 75284 13999
rect 75243 13124 75285 13133
rect 75243 13084 75244 13124
rect 75284 13084 75285 13124
rect 75243 13075 75285 13084
rect 75340 12980 75380 14764
rect 75532 14678 75572 14687
rect 75532 14477 75572 14638
rect 75531 14468 75573 14477
rect 75531 14428 75532 14468
rect 75572 14428 75573 14468
rect 75531 14419 75573 14428
rect 75628 13637 75668 16192
rect 75724 16183 75764 16192
rect 75820 16064 75860 16073
rect 76012 16064 76052 17032
rect 75860 16024 76052 16064
rect 76300 16232 76340 17032
rect 76492 16484 76532 17032
rect 76745 16988 76785 17472
rect 76855 17072 76895 17472
rect 77145 17072 77185 17472
rect 77255 17072 77295 17472
rect 77545 17072 77585 17472
rect 77655 17072 77695 17472
rect 77945 17072 77985 17472
rect 78055 17072 78095 17472
rect 78345 17156 78385 17472
rect 76855 17032 76916 17072
rect 77145 17032 77204 17072
rect 77255 17032 77300 17072
rect 77545 17032 77588 17072
rect 76745 16948 76820 16988
rect 76492 16435 76532 16444
rect 76588 16232 76628 16241
rect 76300 16192 76588 16232
rect 76780 16232 76820 16948
rect 76876 16484 76916 17032
rect 76876 16435 76916 16444
rect 76971 16232 77013 16241
rect 76780 16192 76972 16232
rect 77012 16192 77013 16232
rect 75820 16015 75860 16024
rect 76203 14888 76245 14897
rect 76203 14848 76204 14888
rect 76244 14848 76245 14888
rect 76203 14839 76245 14848
rect 75724 14729 75764 14814
rect 75723 14720 75765 14729
rect 75723 14680 75724 14720
rect 75764 14680 75765 14720
rect 75723 14671 75765 14680
rect 75820 14720 75860 14729
rect 75820 14216 75860 14680
rect 76204 14720 76244 14839
rect 76204 14671 76244 14680
rect 76011 14384 76053 14393
rect 76011 14344 76012 14384
rect 76052 14344 76053 14384
rect 76011 14335 76053 14344
rect 75820 14176 75956 14216
rect 75916 14132 75956 14176
rect 75916 14083 75956 14092
rect 75820 14048 75860 14057
rect 75820 13721 75860 14008
rect 76012 14048 76052 14335
rect 76012 13999 76052 14008
rect 75819 13712 75861 13721
rect 75819 13672 75820 13712
rect 75860 13672 75861 13712
rect 75819 13663 75861 13672
rect 75627 13628 75669 13637
rect 75627 13588 75628 13628
rect 75668 13588 75669 13628
rect 75627 13579 75669 13588
rect 76108 13376 76148 13385
rect 75435 13292 75477 13301
rect 75435 13252 75436 13292
rect 75476 13252 75477 13292
rect 75435 13243 75477 13252
rect 75723 13292 75765 13301
rect 75723 13252 75724 13292
rect 75764 13252 75765 13292
rect 75723 13243 75765 13252
rect 75148 12940 75380 12980
rect 75436 13208 75476 13243
rect 75051 12788 75093 12797
rect 75051 12748 75052 12788
rect 75092 12748 75093 12788
rect 75051 12739 75093 12748
rect 74956 12487 74996 12496
rect 75052 12536 75092 12545
rect 74763 12368 74805 12377
rect 74763 12328 74764 12368
rect 74804 12328 74805 12368
rect 74763 12319 74805 12328
rect 74764 12234 74804 12319
rect 75052 11957 75092 12496
rect 74956 11948 74996 11957
rect 75051 11948 75093 11957
rect 74996 11908 75052 11948
rect 75092 11908 75093 11948
rect 74956 11899 74996 11908
rect 75051 11899 75093 11908
rect 75052 11814 75092 11899
rect 74956 11528 74996 11537
rect 74859 11360 74901 11369
rect 74859 11320 74860 11360
rect 74900 11320 74901 11360
rect 74859 11311 74901 11320
rect 74668 11152 74804 11192
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 74764 11024 74804 11152
rect 74668 10890 74708 10975
rect 74764 10865 74804 10984
rect 74860 11024 74900 11311
rect 74860 10949 74900 10984
rect 74956 11024 74996 11488
rect 75148 11192 75188 12940
rect 75243 12788 75285 12797
rect 75243 12748 75244 12788
rect 75284 12748 75285 12788
rect 75243 12739 75285 12748
rect 75244 11369 75284 12739
rect 75436 11864 75476 13168
rect 75724 13208 75764 13243
rect 75724 13157 75764 13168
rect 75819 13208 75861 13217
rect 75819 13168 75820 13208
rect 75860 13168 75861 13208
rect 75819 13159 75861 13168
rect 75820 13074 75860 13159
rect 76108 12980 76148 13336
rect 76108 12940 76244 12980
rect 76107 12704 76149 12713
rect 76107 12664 76108 12704
rect 76148 12664 76149 12704
rect 76107 12655 76149 12664
rect 75531 12620 75573 12629
rect 75531 12580 75532 12620
rect 75572 12580 75573 12620
rect 75531 12571 75573 12580
rect 76108 12620 76148 12655
rect 75340 11824 75476 11864
rect 75340 11696 75380 11824
rect 75340 11537 75380 11656
rect 75435 11696 75477 11705
rect 75435 11656 75436 11696
rect 75476 11656 75477 11696
rect 75435 11647 75477 11656
rect 75339 11528 75381 11537
rect 75339 11488 75340 11528
rect 75380 11488 75381 11528
rect 75339 11479 75381 11488
rect 75243 11360 75285 11369
rect 75243 11320 75244 11360
rect 75284 11320 75285 11360
rect 75243 11311 75285 11320
rect 74956 10975 74996 10984
rect 75052 11152 75188 11192
rect 75243 11192 75285 11201
rect 75436 11192 75476 11647
rect 75243 11152 75244 11192
rect 75284 11152 75285 11192
rect 74859 10940 74901 10949
rect 74859 10900 74860 10940
rect 74900 10900 74901 10940
rect 74859 10891 74901 10900
rect 74763 10856 74805 10865
rect 74763 10816 74764 10856
rect 74804 10816 74805 10856
rect 74763 10807 74805 10816
rect 74764 10529 74804 10807
rect 74763 10520 74805 10529
rect 74763 10480 74764 10520
rect 74804 10480 74805 10520
rect 74763 10471 74805 10480
rect 74763 10184 74805 10193
rect 74763 10144 74764 10184
rect 74804 10144 74900 10184
rect 74763 10135 74805 10144
rect 74764 10050 74804 10135
rect 74188 8968 74420 9008
rect 74092 8875 74132 8884
rect 74284 8840 74324 8849
rect 73996 8000 74036 8009
rect 74284 8000 74324 8800
rect 74036 7960 74324 8000
rect 73996 7951 74036 7960
rect 74284 6656 74324 6665
rect 74380 6656 74420 8968
rect 74860 8000 74900 10144
rect 74860 7951 74900 7960
rect 74324 6616 74420 6656
rect 74284 6607 74324 6616
rect 74476 6320 74516 6329
rect 74284 6236 74324 6245
rect 74284 5825 74324 6196
rect 74283 5816 74325 5825
rect 74283 5776 74284 5816
rect 74324 5776 74325 5816
rect 74283 5767 74325 5776
rect 73996 5648 74036 5657
rect 74476 5648 74516 6280
rect 75052 5732 75092 11152
rect 75243 11143 75285 11152
rect 75340 11152 75476 11192
rect 75244 11058 75284 11143
rect 75147 11024 75189 11033
rect 75147 10984 75148 11024
rect 75188 10984 75189 11024
rect 75147 10975 75189 10984
rect 75340 11024 75380 11152
rect 75340 10975 75380 10984
rect 75436 11024 75476 11033
rect 75532 11024 75572 12571
rect 76108 12569 76148 12580
rect 76012 12536 76052 12545
rect 75916 12496 76012 12536
rect 75723 11948 75765 11957
rect 75723 11908 75724 11948
rect 75764 11908 75765 11948
rect 75723 11899 75765 11908
rect 75628 11696 75668 11705
rect 75628 11621 75668 11656
rect 75724 11696 75764 11899
rect 75724 11647 75764 11656
rect 75628 11612 75670 11621
rect 75628 11572 75629 11612
rect 75669 11572 75670 11612
rect 75628 11563 75670 11572
rect 75916 11453 75956 12496
rect 76012 12487 76052 12496
rect 76204 12536 76244 12940
rect 76204 12487 76244 12496
rect 76012 11864 76052 11873
rect 76052 11824 76148 11864
rect 76012 11815 76052 11824
rect 76011 11528 76053 11537
rect 76011 11488 76012 11528
rect 76052 11488 76053 11528
rect 76011 11479 76053 11488
rect 75915 11444 75957 11453
rect 75915 11404 75916 11444
rect 75956 11404 75957 11444
rect 75915 11395 75957 11404
rect 75628 11024 75668 11033
rect 75820 11024 75860 11033
rect 75532 10984 75628 11024
rect 75668 10984 75764 11024
rect 75148 10890 75188 10975
rect 75243 10940 75285 10949
rect 75243 10900 75244 10940
rect 75284 10900 75285 10940
rect 75243 10891 75285 10900
rect 75244 9521 75284 10891
rect 75339 10856 75381 10865
rect 75339 10816 75340 10856
rect 75380 10816 75381 10856
rect 75436 10856 75476 10984
rect 75628 10975 75668 10984
rect 75628 10856 75668 10865
rect 75436 10816 75628 10856
rect 75339 10807 75381 10816
rect 75628 10807 75668 10816
rect 75243 9512 75285 9521
rect 75243 9472 75244 9512
rect 75284 9472 75285 9512
rect 75243 9463 75285 9472
rect 75244 7169 75284 9463
rect 75340 8756 75380 10807
rect 75724 10184 75764 10984
rect 75820 10781 75860 10984
rect 75916 11024 75956 11033
rect 75819 10772 75861 10781
rect 75819 10732 75820 10772
rect 75860 10732 75861 10772
rect 75819 10723 75861 10732
rect 75916 10445 75956 10984
rect 76012 10856 76052 11479
rect 76108 11024 76148 11824
rect 76203 11696 76245 11705
rect 76203 11656 76204 11696
rect 76244 11656 76245 11696
rect 76203 11647 76245 11656
rect 76204 11108 76244 11647
rect 76300 11285 76340 16192
rect 76588 16183 76628 16192
rect 76971 16183 77013 16192
rect 77164 16232 77204 17032
rect 77260 16484 77300 17032
rect 77260 16435 77300 16444
rect 76972 16098 77012 16183
rect 77164 15560 77204 16192
rect 76396 15520 77204 15560
rect 77548 16232 77588 17032
rect 77644 17032 77695 17072
rect 77932 17032 77985 17072
rect 78028 17032 78095 17072
rect 78220 17116 78385 17156
rect 77644 16484 77684 17032
rect 77644 16435 77684 16444
rect 76396 12797 76436 15520
rect 76684 15392 76724 15401
rect 76588 14720 76628 14729
rect 76684 14720 76724 15352
rect 76628 14680 76724 14720
rect 77452 14720 77492 14729
rect 76588 14671 76628 14680
rect 77163 14216 77205 14225
rect 77163 14176 77164 14216
rect 77204 14176 77205 14216
rect 77163 14167 77205 14176
rect 76972 14048 77012 14057
rect 76492 14008 76972 14048
rect 76492 13460 76532 14008
rect 76972 13999 77012 14008
rect 76492 13411 76532 13420
rect 76587 13376 76629 13385
rect 77068 13376 77108 13385
rect 76587 13336 76588 13376
rect 76628 13336 76629 13376
rect 76587 13327 76629 13336
rect 76780 13336 77068 13376
rect 76492 13208 76532 13236
rect 76588 13208 76628 13327
rect 76532 13168 76628 13208
rect 76492 13159 76532 13168
rect 76395 12788 76437 12797
rect 76395 12748 76396 12788
rect 76436 12748 76437 12788
rect 76395 12739 76437 12748
rect 76588 12620 76628 13168
rect 76684 13208 76724 13217
rect 76684 12713 76724 13168
rect 76780 13208 76820 13336
rect 77068 13327 77108 13336
rect 77164 13301 77204 14167
rect 77356 14048 77396 14057
rect 77260 14008 77356 14048
rect 77260 13385 77300 14008
rect 77356 13999 77396 14008
rect 77452 13880 77492 14680
rect 77356 13840 77492 13880
rect 77259 13376 77301 13385
rect 77259 13336 77260 13376
rect 77300 13336 77301 13376
rect 77259 13327 77301 13336
rect 77163 13292 77205 13301
rect 77163 13252 77164 13292
rect 77204 13252 77205 13292
rect 77163 13243 77205 13252
rect 76780 13159 76820 13168
rect 76972 13208 77012 13219
rect 76972 13133 77012 13168
rect 77164 13208 77204 13243
rect 77164 13158 77204 13168
rect 76971 13124 77013 13133
rect 76971 13084 76972 13124
rect 77012 13084 77013 13124
rect 76971 13075 77013 13084
rect 76683 12704 76725 12713
rect 76683 12664 76684 12704
rect 76724 12664 76725 12704
rect 76683 12655 76725 12664
rect 76396 12580 76628 12620
rect 76396 11696 76436 12580
rect 76876 12536 76916 12545
rect 76492 12496 76876 12536
rect 76492 11948 76532 12496
rect 76876 12487 76916 12496
rect 76492 11899 76532 11908
rect 76492 11696 76532 11705
rect 76396 11656 76492 11696
rect 76395 11444 76437 11453
rect 76395 11404 76396 11444
rect 76436 11404 76437 11444
rect 76492 11444 76532 11656
rect 76683 11696 76725 11705
rect 76683 11656 76684 11696
rect 76724 11656 76725 11696
rect 76683 11647 76725 11656
rect 76780 11696 76820 11705
rect 76972 11696 77012 13075
rect 77356 12965 77396 13840
rect 77451 13376 77493 13385
rect 77451 13336 77452 13376
rect 77492 13336 77493 13376
rect 77451 13327 77493 13336
rect 77452 13242 77492 13327
rect 77548 12980 77588 16192
rect 77739 16232 77781 16241
rect 77739 16192 77740 16232
rect 77780 16192 77781 16232
rect 77739 16183 77781 16192
rect 77932 16232 77972 17032
rect 78028 16484 78068 17032
rect 78028 16435 78068 16444
rect 77355 12956 77397 12965
rect 77355 12916 77356 12956
rect 77396 12916 77397 12956
rect 77355 12907 77397 12916
rect 77452 12940 77588 12980
rect 77260 12536 77300 12545
rect 77300 12496 77396 12536
rect 77260 12487 77300 12496
rect 77356 11864 77396 12496
rect 77356 11815 77396 11824
rect 76820 11656 76916 11696
rect 76780 11647 76820 11656
rect 76684 11562 76724 11647
rect 76876 11528 76916 11656
rect 76972 11647 77012 11656
rect 77164 11696 77204 11707
rect 77164 11621 77204 11656
rect 77068 11612 77108 11621
rect 77068 11528 77108 11572
rect 77163 11612 77205 11621
rect 77163 11572 77164 11612
rect 77204 11572 77205 11612
rect 77163 11563 77205 11572
rect 76876 11488 77108 11528
rect 77259 11444 77301 11453
rect 76492 11404 76820 11444
rect 76395 11395 76437 11404
rect 76299 11276 76341 11285
rect 76299 11236 76300 11276
rect 76340 11236 76341 11276
rect 76299 11227 76341 11236
rect 76204 11059 76244 11068
rect 76108 10975 76148 10984
rect 76311 11024 76351 11032
rect 76396 11024 76436 11395
rect 76587 11276 76629 11285
rect 76587 11236 76588 11276
rect 76628 11236 76629 11276
rect 76587 11227 76629 11236
rect 76311 11023 76436 11024
rect 76351 10984 76436 11023
rect 76311 10974 76351 10983
rect 76492 10929 76532 10938
rect 76299 10856 76341 10865
rect 76012 10816 76244 10856
rect 75915 10436 75957 10445
rect 75915 10396 75916 10436
rect 75956 10396 75957 10436
rect 75915 10387 75957 10396
rect 75916 10302 75956 10387
rect 75436 10144 75764 10184
rect 76204 10184 76244 10816
rect 76299 10816 76300 10856
rect 76340 10816 76341 10856
rect 76299 10807 76341 10816
rect 75436 9017 75476 10144
rect 76204 10100 76244 10144
rect 76108 10060 76244 10100
rect 75531 10016 75573 10025
rect 75531 9976 75532 10016
rect 75572 9976 75573 10016
rect 75531 9967 75573 9976
rect 75916 10016 75956 10025
rect 75532 9680 75572 9967
rect 75916 9764 75956 9976
rect 76011 10016 76053 10025
rect 76011 9976 76012 10016
rect 76052 9976 76053 10016
rect 76011 9967 76053 9976
rect 75916 9724 75965 9764
rect 75925 9680 75965 9724
rect 75532 9631 75572 9640
rect 75916 9640 75965 9680
rect 75628 9512 75668 9521
rect 75532 9472 75628 9512
rect 75435 9008 75477 9017
rect 75435 8968 75436 9008
rect 75476 8968 75477 9008
rect 75435 8959 75477 8968
rect 75532 8756 75572 9472
rect 75628 9463 75668 9472
rect 75723 9512 75765 9521
rect 75723 9472 75724 9512
rect 75764 9472 75765 9512
rect 75723 9463 75765 9472
rect 75820 9512 75860 9521
rect 75916 9512 75956 9640
rect 75860 9472 75956 9512
rect 76012 9512 76052 9967
rect 75820 9463 75860 9472
rect 76012 9463 76052 9472
rect 75724 9378 75764 9463
rect 75723 9260 75765 9269
rect 75723 9220 75724 9260
rect 75764 9220 75765 9260
rect 75723 9211 75765 9220
rect 76012 9260 76052 9271
rect 75340 8716 75572 8756
rect 75435 7748 75477 7757
rect 75435 7708 75436 7748
rect 75476 7708 75477 7748
rect 75435 7699 75477 7708
rect 75243 7160 75285 7169
rect 75243 7120 75244 7160
rect 75284 7120 75285 7160
rect 75243 7111 75285 7120
rect 75436 7160 75476 7699
rect 75532 7580 75572 8716
rect 75628 8672 75668 8681
rect 75628 8597 75668 8632
rect 75724 8672 75764 9211
rect 76012 9185 76052 9220
rect 76011 9176 76053 9185
rect 76011 9136 76012 9176
rect 76052 9136 76053 9176
rect 76011 9127 76053 9136
rect 75819 9008 75861 9017
rect 75819 8968 75820 9008
rect 75860 8968 75861 9008
rect 75819 8959 75861 8968
rect 75820 8672 75860 8959
rect 75915 8924 75957 8933
rect 75915 8884 75916 8924
rect 75956 8884 75957 8924
rect 75915 8875 75957 8884
rect 75916 8790 75956 8875
rect 75916 8672 75956 8681
rect 75820 8632 75916 8672
rect 75627 8588 75669 8597
rect 75627 8548 75628 8588
rect 75668 8548 75669 8588
rect 75627 8539 75669 8548
rect 75628 7757 75668 8539
rect 75724 8084 75764 8632
rect 75724 8044 75860 8084
rect 75723 7916 75765 7925
rect 75723 7876 75724 7916
rect 75764 7876 75765 7916
rect 75723 7867 75765 7876
rect 75627 7748 75669 7757
rect 75627 7708 75628 7748
rect 75668 7708 75669 7748
rect 75627 7699 75669 7708
rect 75532 7540 75668 7580
rect 75436 7111 75476 7120
rect 75531 7160 75573 7169
rect 75531 7120 75532 7160
rect 75572 7120 75573 7160
rect 75531 7111 75573 7120
rect 75628 7160 75668 7540
rect 75532 7026 75572 7111
rect 75628 6992 75668 7120
rect 75724 7160 75764 7867
rect 75820 7673 75860 8044
rect 75819 7664 75861 7673
rect 75819 7624 75820 7664
rect 75860 7624 75861 7664
rect 75819 7615 75861 7624
rect 75724 7111 75764 7120
rect 75819 7160 75861 7169
rect 75819 7120 75820 7160
rect 75860 7120 75861 7160
rect 75819 7111 75861 7120
rect 75916 7160 75956 8632
rect 76108 8672 76148 10060
rect 76300 9680 76340 10807
rect 76492 10436 76532 10889
rect 76588 10604 76628 11227
rect 76684 10781 76724 10866
rect 76683 10772 76725 10781
rect 76683 10732 76684 10772
rect 76724 10732 76725 10772
rect 76683 10723 76725 10732
rect 76588 10564 76724 10604
rect 76396 10396 76532 10436
rect 76587 10436 76629 10445
rect 76587 10396 76588 10436
rect 76628 10396 76629 10436
rect 76396 10016 76436 10396
rect 76587 10387 76629 10396
rect 76491 10268 76533 10277
rect 76491 10228 76492 10268
rect 76532 10228 76533 10268
rect 76491 10219 76533 10228
rect 76492 10184 76532 10219
rect 76492 10133 76532 10144
rect 76588 10184 76628 10387
rect 76588 10135 76628 10144
rect 76684 10016 76724 10564
rect 76396 9976 76532 10016
rect 76492 9689 76532 9976
rect 76588 9976 76724 10016
rect 76491 9680 76533 9689
rect 76300 9640 76436 9680
rect 76300 9512 76340 9521
rect 76204 9498 76244 9507
rect 76204 9437 76244 9458
rect 76202 9428 76244 9437
rect 76202 9388 76203 9428
rect 76243 9388 76244 9428
rect 76202 9379 76244 9388
rect 76203 9364 76243 9379
rect 76300 8933 76340 9472
rect 76299 8924 76341 8933
rect 76299 8884 76300 8924
rect 76340 8884 76341 8924
rect 76299 8875 76341 8884
rect 76204 8672 76244 8681
rect 76108 8632 76204 8672
rect 76108 7832 76148 8632
rect 76204 8623 76244 8632
rect 76396 8168 76436 9640
rect 76491 9640 76492 9680
rect 76532 9640 76533 9680
rect 76491 9631 76533 9640
rect 76492 9428 76532 9631
rect 76492 9379 76532 9388
rect 76491 9260 76533 9269
rect 76491 9220 76492 9260
rect 76532 9220 76533 9260
rect 76491 9211 76533 9220
rect 76492 8672 76532 9211
rect 76588 9092 76628 9976
rect 76780 9521 76820 11404
rect 77259 11404 77260 11444
rect 77300 11404 77301 11444
rect 77259 11395 77301 11404
rect 77068 11024 77108 11033
rect 76876 10984 77068 11024
rect 76876 10436 76916 10984
rect 77068 10975 77108 10984
rect 77260 11024 77300 11395
rect 77260 10949 77300 10984
rect 77259 10940 77301 10949
rect 77259 10900 77260 10940
rect 77300 10900 77301 10940
rect 77259 10891 77301 10900
rect 76971 10856 77013 10865
rect 77260 10860 77300 10891
rect 76971 10816 76972 10856
rect 77012 10816 77013 10856
rect 76971 10807 77013 10816
rect 76876 10387 76916 10396
rect 76779 9512 76821 9521
rect 76779 9472 76780 9512
rect 76820 9472 76821 9512
rect 76779 9463 76821 9472
rect 76683 9344 76725 9353
rect 76683 9304 76684 9344
rect 76724 9304 76725 9344
rect 76683 9295 76725 9304
rect 76684 9210 76724 9295
rect 76588 9052 76724 9092
rect 76492 8623 76532 8632
rect 76587 8588 76629 8597
rect 76587 8548 76588 8588
rect 76628 8548 76629 8588
rect 76587 8539 76629 8548
rect 76588 8454 76628 8539
rect 76396 8128 76628 8168
rect 76204 8009 76244 8094
rect 76299 8084 76341 8093
rect 76299 8044 76300 8084
rect 76340 8044 76341 8084
rect 76299 8035 76341 8044
rect 76203 8000 76245 8009
rect 76203 7960 76204 8000
rect 76244 7960 76245 8000
rect 76203 7951 76245 7960
rect 76300 7950 76340 8035
rect 76395 8000 76437 8009
rect 76395 7960 76396 8000
rect 76436 7960 76437 8000
rect 76395 7951 76437 7960
rect 76492 8000 76532 8009
rect 76396 7866 76436 7951
rect 76108 7792 76340 7832
rect 76011 7748 76053 7757
rect 76011 7708 76012 7748
rect 76052 7708 76053 7748
rect 76011 7699 76053 7708
rect 76012 7614 76052 7699
rect 76107 7664 76149 7673
rect 76107 7624 76108 7664
rect 76148 7624 76149 7664
rect 76107 7615 76149 7624
rect 76011 7244 76053 7253
rect 76011 7204 76012 7244
rect 76052 7204 76053 7244
rect 76011 7195 76053 7204
rect 75916 7111 75956 7120
rect 75628 6952 75764 6992
rect 75628 6488 75668 6497
rect 75052 5692 75188 5732
rect 74036 5608 74516 5648
rect 74860 5648 74900 5657
rect 74900 5608 75092 5648
rect 73996 5599 74036 5608
rect 74860 5599 74900 5608
rect 74284 4808 74324 4817
rect 74188 4768 74284 4808
rect 73803 3548 73845 3557
rect 73803 3508 73804 3548
rect 73844 3508 73845 3548
rect 73803 3499 73845 3508
rect 73804 3414 73844 3499
rect 74188 3464 74228 4768
rect 74284 4759 74324 4768
rect 74379 4472 74421 4481
rect 74379 4432 74380 4472
rect 74420 4432 74421 4472
rect 74379 4423 74421 4432
rect 74380 4304 74420 4423
rect 74859 4388 74901 4397
rect 74859 4348 74860 4388
rect 74900 4348 74901 4388
rect 74859 4339 74901 4348
rect 74380 4255 74420 4264
rect 74860 3473 74900 4339
rect 74188 3415 74228 3424
rect 74859 3464 74901 3473
rect 74859 3424 74860 3464
rect 74900 3424 74901 3464
rect 74859 3415 74901 3424
rect 75052 3464 75092 5608
rect 75148 4481 75188 5692
rect 75628 5657 75668 6448
rect 75724 6488 75764 6952
rect 75724 6439 75764 6448
rect 75820 6488 75860 7111
rect 76012 7076 76052 7195
rect 76012 7027 76052 7036
rect 76108 7160 76148 7615
rect 76011 6908 76053 6917
rect 76011 6868 76012 6908
rect 76052 6868 76053 6908
rect 76011 6859 76053 6868
rect 76012 6488 76052 6859
rect 76108 6740 76148 7120
rect 76204 7160 76244 7169
rect 76204 6917 76244 7120
rect 76203 6908 76245 6917
rect 76203 6868 76204 6908
rect 76244 6868 76245 6908
rect 76203 6859 76245 6868
rect 76107 6700 76148 6740
rect 76107 6656 76147 6700
rect 76107 6616 76148 6656
rect 75917 6480 76052 6488
rect 75820 6439 75860 6448
rect 75916 6451 76052 6480
rect 75956 6448 76052 6451
rect 75956 6440 75957 6448
rect 75916 6402 75956 6411
rect 76011 5900 76053 5909
rect 76011 5860 76012 5900
rect 76052 5860 76053 5900
rect 76011 5851 76053 5860
rect 76012 5766 76052 5851
rect 75627 5648 75669 5657
rect 75627 5608 75628 5648
rect 75668 5608 75669 5648
rect 75627 5599 75669 5608
rect 76108 5564 76148 6616
rect 76204 6488 76244 6497
rect 76300 6488 76340 7792
rect 76492 7253 76532 7960
rect 76491 7244 76533 7253
rect 76491 7204 76492 7244
rect 76532 7204 76533 7244
rect 76491 7195 76533 7204
rect 76588 7076 76628 8128
rect 76244 6448 76340 6488
rect 76492 7036 76628 7076
rect 76492 6488 76532 7036
rect 76587 6908 76629 6917
rect 76587 6868 76588 6908
rect 76628 6868 76629 6908
rect 76587 6859 76629 6868
rect 76204 6439 76244 6448
rect 76492 5825 76532 6448
rect 76588 6488 76628 6859
rect 76588 5909 76628 6448
rect 76587 5900 76629 5909
rect 76587 5860 76588 5900
rect 76628 5860 76629 5900
rect 76587 5851 76629 5860
rect 76491 5816 76533 5825
rect 76491 5776 76492 5816
rect 76532 5776 76533 5816
rect 76491 5767 76533 5776
rect 76203 5648 76245 5657
rect 76203 5608 76204 5648
rect 76244 5608 76245 5648
rect 76203 5599 76245 5608
rect 76395 5648 76437 5657
rect 76395 5608 76396 5648
rect 76436 5608 76437 5648
rect 76395 5599 76437 5608
rect 76492 5648 76532 5657
rect 76012 5524 76148 5564
rect 75916 4976 75956 4985
rect 75147 4472 75189 4481
rect 75147 4432 75148 4472
rect 75188 4432 75189 4472
rect 75147 4423 75189 4432
rect 75148 4264 75668 4304
rect 75148 4136 75188 4264
rect 75148 4087 75188 4096
rect 75340 4136 75380 4147
rect 75340 4061 75380 4096
rect 75436 4136 75476 4145
rect 75339 4052 75381 4061
rect 75339 4012 75340 4052
rect 75380 4012 75381 4052
rect 75339 4003 75381 4012
rect 75244 3968 75284 3977
rect 75244 3557 75284 3928
rect 75436 3641 75476 4096
rect 75628 4136 75668 4264
rect 75916 4145 75956 4936
rect 76012 4976 76052 5524
rect 76204 5514 76244 5599
rect 76299 5564 76341 5573
rect 76299 5524 76300 5564
rect 76340 5524 76341 5564
rect 76299 5515 76341 5524
rect 76300 5430 76340 5515
rect 76396 5514 76436 5599
rect 76492 5153 76532 5608
rect 76107 5144 76149 5153
rect 76107 5104 76108 5144
rect 76148 5104 76149 5144
rect 76107 5095 76149 5104
rect 76491 5144 76533 5153
rect 76491 5104 76492 5144
rect 76532 5104 76533 5144
rect 76491 5095 76533 5104
rect 76108 5010 76148 5095
rect 76012 4313 76052 4936
rect 76204 4976 76244 4985
rect 76011 4304 76053 4313
rect 76011 4264 76012 4304
rect 76052 4264 76053 4304
rect 76204 4304 76244 4936
rect 76204 4264 76436 4304
rect 76011 4255 76053 4264
rect 75628 4087 75668 4096
rect 75724 4136 75764 4145
rect 75435 3632 75477 3641
rect 75435 3592 75436 3632
rect 75476 3592 75477 3632
rect 75435 3583 75477 3592
rect 75243 3548 75285 3557
rect 75243 3508 75244 3548
rect 75284 3508 75285 3548
rect 75243 3499 75285 3508
rect 74667 3380 74709 3389
rect 74667 3340 74668 3380
rect 74708 3340 74709 3380
rect 74667 3331 74709 3340
rect 73516 2876 73556 2885
rect 73324 2836 73516 2876
rect 73324 1961 73364 2836
rect 73516 2827 73556 2836
rect 73612 2860 73748 2900
rect 73612 2717 73652 2860
rect 73611 2708 73653 2717
rect 73611 2668 73612 2708
rect 73652 2668 73653 2708
rect 73611 2659 73653 2668
rect 74379 2708 74421 2717
rect 74379 2668 74380 2708
rect 74420 2668 74421 2708
rect 74379 2659 74421 2668
rect 73803 2624 73845 2633
rect 73803 2584 73804 2624
rect 73844 2584 73845 2624
rect 73803 2575 73845 2584
rect 74187 2624 74229 2633
rect 74187 2584 74188 2624
rect 74228 2584 74229 2624
rect 74187 2575 74229 2584
rect 74380 2624 74420 2659
rect 73804 2120 73844 2575
rect 74091 2540 74133 2549
rect 74091 2500 74092 2540
rect 74132 2500 74133 2540
rect 74091 2491 74133 2500
rect 73804 1961 73844 2080
rect 73323 1952 73365 1961
rect 73323 1912 73324 1952
rect 73364 1912 73365 1952
rect 73323 1903 73365 1912
rect 73803 1952 73845 1961
rect 73803 1912 73804 1952
rect 73844 1912 73845 1952
rect 73803 1903 73845 1912
rect 73996 1952 74036 1963
rect 73996 1877 74036 1912
rect 74092 1952 74132 2491
rect 74188 2129 74228 2575
rect 74380 2573 74420 2584
rect 74572 2624 74612 2633
rect 74668 2624 74708 3331
rect 74612 2584 74708 2624
rect 74572 2575 74612 2584
rect 74476 2540 74516 2549
rect 74476 2204 74516 2500
rect 74284 2164 74516 2204
rect 74187 2120 74229 2129
rect 74187 2080 74188 2120
rect 74228 2080 74229 2120
rect 74187 2071 74229 2080
rect 74188 1952 74228 1961
rect 74092 1912 74188 1952
rect 73995 1868 74037 1877
rect 73995 1828 73996 1868
rect 74036 1828 74037 1868
rect 73995 1819 74037 1828
rect 73996 1700 74036 1709
rect 73227 1280 73269 1289
rect 73227 1240 73228 1280
rect 73268 1240 73269 1280
rect 73227 1231 73269 1240
rect 73996 1121 74036 1660
rect 74092 1205 74132 1912
rect 74188 1903 74228 1912
rect 74284 1952 74324 2164
rect 74379 2036 74421 2045
rect 74379 1996 74380 2036
rect 74420 1996 74421 2036
rect 74379 1987 74421 1996
rect 74284 1903 74324 1912
rect 74091 1196 74133 1205
rect 74091 1156 74092 1196
rect 74132 1156 74133 1196
rect 74091 1147 74133 1156
rect 73995 1112 74037 1121
rect 73995 1072 73996 1112
rect 74036 1072 74037 1112
rect 73995 1063 74037 1072
rect 74380 1112 74420 1987
rect 74571 1952 74613 1961
rect 74571 1912 74572 1952
rect 74612 1912 74613 1952
rect 74571 1903 74613 1912
rect 74668 1952 74708 2584
rect 74668 1903 74708 1912
rect 74860 1952 74900 3415
rect 74956 2792 74996 2801
rect 74956 2120 74996 2752
rect 75052 2633 75092 3424
rect 75339 3128 75381 3137
rect 75339 3088 75340 3128
rect 75380 3088 75381 3128
rect 75339 3079 75381 3088
rect 75147 2792 75189 2801
rect 75147 2752 75148 2792
rect 75188 2752 75189 2792
rect 75147 2743 75189 2752
rect 75051 2624 75093 2633
rect 75051 2584 75052 2624
rect 75092 2584 75093 2624
rect 75051 2575 75093 2584
rect 75148 2624 75188 2743
rect 75148 2575 75188 2584
rect 75340 2624 75380 3079
rect 75724 3053 75764 4096
rect 75820 4136 75860 4145
rect 75820 3221 75860 4096
rect 75915 4136 75957 4145
rect 76204 4136 76244 4145
rect 75915 4096 75916 4136
rect 75956 4096 75957 4136
rect 75915 4087 75957 4096
rect 76012 4096 76204 4136
rect 75916 4002 75956 4087
rect 75819 3212 75861 3221
rect 75819 3172 75820 3212
rect 75860 3172 75861 3212
rect 75819 3163 75861 3172
rect 75723 3044 75765 3053
rect 75723 3004 75724 3044
rect 75764 3004 75765 3044
rect 75723 2995 75765 3004
rect 75340 2575 75380 2584
rect 75243 2540 75285 2549
rect 75243 2500 75244 2540
rect 75284 2500 75285 2540
rect 75243 2491 75285 2500
rect 75244 2406 75284 2491
rect 74956 2080 75380 2120
rect 74860 1903 74900 1912
rect 75148 1952 75188 1961
rect 74572 1818 74612 1903
rect 74860 1784 74900 1793
rect 75148 1784 75188 1912
rect 75243 1952 75285 1961
rect 75243 1912 75244 1952
rect 75284 1912 75285 1952
rect 75243 1903 75285 1912
rect 75244 1818 75284 1903
rect 74900 1744 75188 1784
rect 74860 1735 74900 1744
rect 74380 1063 74420 1072
rect 75244 1112 75284 1121
rect 75340 1112 75380 2080
rect 75436 1961 75476 2046
rect 75435 1952 75477 1961
rect 75435 1912 75436 1952
rect 75476 1912 75477 1952
rect 75435 1903 75477 1912
rect 75628 1952 75668 1961
rect 75436 1784 75476 1793
rect 75628 1784 75668 1912
rect 75476 1744 75668 1784
rect 75436 1735 75476 1744
rect 75284 1072 75380 1112
rect 75627 1112 75669 1121
rect 75627 1072 75628 1112
rect 75668 1072 75669 1112
rect 75244 1063 75284 1072
rect 75627 1063 75669 1072
rect 75628 978 75668 1063
rect 73228 944 73268 953
rect 73132 904 73228 944
rect 75724 944 75764 2995
rect 75820 1121 75860 3163
rect 76012 2885 76052 4096
rect 76204 4087 76244 4096
rect 76299 4136 76341 4145
rect 76299 4096 76300 4136
rect 76340 4096 76341 4136
rect 76299 4087 76341 4096
rect 76204 3632 76244 3641
rect 76300 3632 76340 4087
rect 76244 3592 76340 3632
rect 76204 3583 76244 3592
rect 76396 3473 76436 4264
rect 76491 4220 76533 4229
rect 76491 4180 76492 4220
rect 76532 4180 76533 4220
rect 76684 4220 76724 9052
rect 76780 8000 76820 9463
rect 76875 8840 76917 8849
rect 76875 8800 76876 8840
rect 76916 8800 76917 8840
rect 76875 8791 76917 8800
rect 76876 8706 76916 8791
rect 76972 8177 77012 10807
rect 77164 10772 77204 10781
rect 77204 10732 77300 10772
rect 77164 10723 77204 10732
rect 77068 10100 77108 10109
rect 77068 9680 77108 10060
rect 77164 9680 77204 9689
rect 77068 9640 77164 9680
rect 77164 9631 77204 9640
rect 77067 9512 77109 9521
rect 77067 9472 77068 9512
rect 77108 9472 77109 9512
rect 77067 9463 77109 9472
rect 77260 9512 77300 10732
rect 77452 10352 77492 12940
rect 77740 10940 77780 16183
rect 77932 12980 77972 16192
rect 78220 16232 78260 17116
rect 78455 17072 78495 17472
rect 78745 17156 78785 17472
rect 78316 17032 78495 17072
rect 78604 17116 78785 17156
rect 78316 16484 78356 17032
rect 78316 16435 78356 16444
rect 78604 16232 78644 17116
rect 78855 17072 78895 17472
rect 78987 17156 79029 17165
rect 78987 17116 78988 17156
rect 79028 17116 79029 17156
rect 78987 17107 79029 17116
rect 78700 17032 78895 17072
rect 78700 16484 78740 17032
rect 78700 16435 78740 16444
rect 78988 16484 79028 17107
rect 79145 17072 79185 17472
rect 79255 17156 79295 17472
rect 79371 17156 79413 17165
rect 79255 17116 79316 17156
rect 79145 17032 79220 17072
rect 78988 16435 79028 16444
rect 78260 16192 78356 16232
rect 78220 16183 78260 16192
rect 78220 14048 78260 14057
rect 78220 12980 78260 14008
rect 77932 12940 78068 12980
rect 78124 12965 78260 12980
rect 77740 10900 77972 10940
rect 77356 10312 77492 10352
rect 77644 10856 77684 10865
rect 77356 9689 77396 10312
rect 77452 10184 77492 10193
rect 77644 10184 77684 10816
rect 77739 10772 77781 10781
rect 77739 10732 77740 10772
rect 77780 10732 77781 10772
rect 77739 10723 77781 10732
rect 77492 10144 77684 10184
rect 77452 10135 77492 10144
rect 77740 10100 77780 10723
rect 77835 10268 77877 10277
rect 77835 10228 77836 10268
rect 77876 10228 77877 10268
rect 77835 10219 77877 10228
rect 77836 10109 77876 10219
rect 77548 10060 77780 10100
rect 77835 10100 77877 10109
rect 77835 10060 77836 10100
rect 77876 10060 77877 10100
rect 77355 9680 77397 9689
rect 77355 9640 77356 9680
rect 77396 9640 77397 9680
rect 77355 9631 77397 9640
rect 77068 9378 77108 9463
rect 77260 9437 77300 9472
rect 77356 9512 77396 9521
rect 77451 9512 77493 9521
rect 77396 9472 77452 9512
rect 77492 9472 77493 9512
rect 77356 9463 77396 9472
rect 77451 9463 77493 9472
rect 77548 9512 77588 10060
rect 77835 10051 77877 10060
rect 77259 9428 77301 9437
rect 77259 9388 77260 9428
rect 77300 9388 77301 9428
rect 77259 9379 77301 9388
rect 77548 9260 77588 9472
rect 77643 9512 77685 9521
rect 77643 9472 77644 9512
rect 77684 9472 77685 9512
rect 77643 9463 77685 9472
rect 77740 9512 77780 9521
rect 77836 9512 77876 10051
rect 77780 9472 77876 9512
rect 77740 9463 77780 9472
rect 77644 9378 77684 9463
rect 77356 9220 77588 9260
rect 77739 9260 77781 9269
rect 77739 9220 77740 9260
rect 77780 9220 77781 9260
rect 77068 8588 77108 8597
rect 76971 8168 77013 8177
rect 76971 8128 76972 8168
rect 77012 8128 77013 8168
rect 76971 8119 77013 8128
rect 77068 8168 77108 8548
rect 77068 8119 77108 8128
rect 76972 8000 77012 8009
rect 76780 7960 76972 8000
rect 76780 5648 76820 7960
rect 76972 7951 77012 7960
rect 77163 8000 77205 8009
rect 77163 7960 77164 8000
rect 77204 7960 77205 8000
rect 77163 7951 77205 7960
rect 77260 8000 77300 8009
rect 77164 7866 77204 7951
rect 77067 7580 77109 7589
rect 77067 7540 77068 7580
rect 77108 7540 77109 7580
rect 77067 7531 77109 7540
rect 76876 7160 76916 7169
rect 76876 6320 76916 7120
rect 77068 7160 77108 7531
rect 77260 7421 77300 7960
rect 77259 7412 77301 7421
rect 77259 7372 77260 7412
rect 77300 7372 77301 7412
rect 77259 7363 77301 7372
rect 77068 7111 77108 7120
rect 77356 7160 77396 9220
rect 77739 9211 77781 9220
rect 77740 8933 77780 9211
rect 77739 8924 77781 8933
rect 77739 8884 77740 8924
rect 77780 8884 77781 8924
rect 77739 8875 77781 8884
rect 77643 8840 77685 8849
rect 77643 8800 77644 8840
rect 77684 8800 77685 8840
rect 77643 8791 77685 8800
rect 77451 8672 77493 8681
rect 77451 8632 77452 8672
rect 77492 8632 77493 8672
rect 77451 8623 77493 8632
rect 77452 8538 77492 8623
rect 77451 8168 77493 8177
rect 77451 8128 77452 8168
rect 77492 8128 77493 8168
rect 77451 8119 77493 8128
rect 77452 8000 77492 8119
rect 77452 7589 77492 7960
rect 77547 8000 77589 8009
rect 77547 7960 77548 8000
rect 77588 7960 77589 8000
rect 77547 7951 77589 7960
rect 77644 8000 77684 8791
rect 77644 7951 77684 7960
rect 77548 7866 77588 7951
rect 77451 7580 77493 7589
rect 77451 7540 77452 7580
rect 77492 7540 77493 7580
rect 77451 7531 77493 7540
rect 77451 7412 77493 7421
rect 77451 7372 77452 7412
rect 77492 7372 77493 7412
rect 77451 7363 77493 7372
rect 77452 7278 77492 7363
rect 76972 7076 77012 7085
rect 76972 6656 77012 7036
rect 76972 6616 77300 6656
rect 76876 6271 76916 6280
rect 77068 6488 77108 6497
rect 77068 5900 77108 6448
rect 77068 5851 77108 5860
rect 77260 5657 77300 6616
rect 77356 6320 77396 7120
rect 77451 7160 77493 7169
rect 77451 7120 77452 7160
rect 77492 7120 77493 7160
rect 77451 7111 77493 7120
rect 77548 7160 77588 7169
rect 77740 7160 77780 8875
rect 77835 8672 77877 8681
rect 77835 8632 77836 8672
rect 77876 8632 77877 8672
rect 77835 8623 77877 8632
rect 77836 7832 77876 8623
rect 77836 7783 77876 7792
rect 77836 7328 77876 7339
rect 77836 7253 77876 7288
rect 77835 7244 77877 7253
rect 77835 7204 77836 7244
rect 77876 7204 77877 7244
rect 77835 7195 77877 7204
rect 77588 7120 77780 7160
rect 77548 7111 77588 7120
rect 77452 6488 77492 7111
rect 77932 7076 77972 10900
rect 78028 10109 78068 12940
rect 78123 12956 78260 12965
rect 78123 12916 78124 12956
rect 78164 12940 78260 12956
rect 78164 12916 78165 12940
rect 78123 12907 78165 12916
rect 78124 12536 78164 12907
rect 78124 12487 78164 12496
rect 78316 12293 78356 16192
rect 78604 14720 78644 16192
rect 78891 16232 78933 16241
rect 78891 16192 78892 16232
rect 78932 16192 78933 16232
rect 78891 16183 78933 16192
rect 79180 16232 79220 17032
rect 79276 16484 79316 17116
rect 79371 17116 79372 17156
rect 79412 17116 79413 17156
rect 79371 17107 79413 17116
rect 79276 16435 79316 16444
rect 78892 16098 78932 16183
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 78604 14680 78740 14720
rect 78603 14552 78645 14561
rect 78603 14512 78604 14552
rect 78644 14512 78645 14552
rect 78603 14503 78645 14512
rect 78604 14418 78644 14503
rect 78700 14225 78740 14680
rect 79180 14561 79220 16192
rect 79372 15560 79412 17107
rect 79545 17072 79585 17472
rect 79655 17165 79695 17472
rect 79654 17156 79696 17165
rect 79654 17116 79655 17156
rect 79695 17116 79696 17156
rect 79654 17107 79696 17116
rect 79468 17032 79585 17072
rect 79468 15728 79508 17032
rect 79468 15679 79508 15688
rect 79372 15511 79412 15520
rect 79179 14552 79221 14561
rect 79179 14512 79180 14552
rect 79220 14512 79221 14552
rect 79179 14503 79221 14512
rect 78699 14216 78741 14225
rect 78699 14176 78700 14216
rect 78740 14176 78741 14216
rect 78699 14167 78741 14176
rect 79371 14216 79413 14225
rect 79371 14176 79372 14216
rect 79412 14176 79413 14216
rect 79371 14167 79413 14176
rect 79372 14082 79412 14167
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 78315 12284 78357 12293
rect 78315 12244 78316 12284
rect 78356 12244 78357 12284
rect 78315 12235 78357 12244
rect 79275 12284 79317 12293
rect 79275 12244 79276 12284
rect 79316 12244 79317 12284
rect 79275 12235 79317 12244
rect 78316 11621 78356 12235
rect 79276 12150 79316 12235
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 78315 11612 78357 11621
rect 78315 11572 78316 11612
rect 78356 11572 78357 11612
rect 78315 11563 78357 11572
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 79468 10268 79508 10277
rect 78315 10184 78357 10193
rect 78315 10144 78316 10184
rect 78356 10144 78357 10184
rect 78315 10135 78357 10144
rect 78027 10100 78069 10109
rect 78027 10060 78028 10100
rect 78068 10060 78069 10100
rect 78027 10051 78069 10060
rect 78316 8672 78356 10135
rect 79468 10109 79508 10228
rect 79467 10100 79509 10109
rect 79467 10060 79468 10100
rect 79508 10060 79509 10100
rect 79467 10051 79509 10060
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 79467 8924 79509 8933
rect 79467 8884 79468 8924
rect 79508 8884 79509 8924
rect 79467 8875 79509 8884
rect 79468 8790 79508 8875
rect 78316 8623 78356 8632
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 77452 6439 77492 6448
rect 77740 7036 77972 7076
rect 77356 6280 77492 6320
rect 77068 5648 77108 5657
rect 76780 5608 77068 5648
rect 77068 5599 77108 5608
rect 77259 5648 77301 5657
rect 77259 5608 77260 5648
rect 77300 5608 77301 5648
rect 77259 5599 77301 5608
rect 77356 5648 77396 5657
rect 77452 5648 77492 6280
rect 77740 5984 77780 7036
rect 78316 6488 78356 6497
rect 77740 5944 77876 5984
rect 77739 5816 77781 5825
rect 77739 5776 77740 5816
rect 77780 5776 77781 5816
rect 77739 5767 77781 5776
rect 77548 5648 77588 5657
rect 77452 5608 77548 5648
rect 77260 5514 77300 5599
rect 77356 5480 77396 5608
rect 77548 5599 77588 5608
rect 77740 5648 77780 5767
rect 77740 5599 77780 5608
rect 77644 5564 77684 5573
rect 77644 5480 77684 5524
rect 77836 5480 77876 5944
rect 77356 5440 77684 5480
rect 77740 5440 77876 5480
rect 77740 5396 77780 5440
rect 77644 5356 77780 5396
rect 77644 5144 77684 5356
rect 77260 5104 77684 5144
rect 76963 4989 77003 4998
rect 76876 4949 76963 4976
rect 76876 4936 77003 4949
rect 77164 4976 77204 4985
rect 76876 4388 76916 4936
rect 77164 4892 77204 4936
rect 76876 4339 76916 4348
rect 76972 4852 77204 4892
rect 76684 4180 76916 4220
rect 76491 4171 76533 4180
rect 76492 4136 76532 4171
rect 76492 4085 76532 4096
rect 76587 4136 76629 4145
rect 76587 4096 76588 4136
rect 76628 4096 76629 4136
rect 76587 4087 76629 4096
rect 76588 4002 76628 4087
rect 76491 3632 76533 3641
rect 76491 3592 76492 3632
rect 76532 3592 76533 3632
rect 76491 3583 76533 3592
rect 76492 3498 76532 3583
rect 76395 3464 76437 3473
rect 76395 3424 76396 3464
rect 76436 3424 76437 3464
rect 76395 3415 76437 3424
rect 76587 3464 76629 3473
rect 76587 3424 76588 3464
rect 76628 3424 76629 3464
rect 76587 3415 76629 3424
rect 76684 3464 76724 3473
rect 76396 3330 76436 3415
rect 76588 3330 76628 3415
rect 76011 2876 76053 2885
rect 76011 2836 76012 2876
rect 76052 2836 76053 2876
rect 76011 2827 76053 2836
rect 76108 2792 76148 2801
rect 75915 1952 75957 1961
rect 75915 1912 75916 1952
rect 75956 1912 75957 1952
rect 75915 1903 75957 1912
rect 76012 1952 76052 1961
rect 76108 1952 76148 2752
rect 76684 2549 76724 3424
rect 76876 2900 76916 4180
rect 76972 3137 77012 4852
rect 77068 4724 77108 4733
rect 77108 4684 77204 4724
rect 77068 4675 77108 4684
rect 77164 4061 77204 4684
rect 77260 4229 77300 5104
rect 77644 4989 77684 5104
rect 77452 4976 77492 4985
rect 77492 4936 77588 4976
rect 77644 4940 77684 4949
rect 77452 4927 77492 4936
rect 77548 4892 77588 4936
rect 77548 4852 77677 4892
rect 77451 4808 77493 4817
rect 77451 4768 77452 4808
rect 77492 4768 77493 4808
rect 77637 4808 77677 4852
rect 77835 4808 77877 4817
rect 77637 4768 77684 4808
rect 77451 4759 77493 4768
rect 77259 4220 77301 4229
rect 77259 4180 77260 4220
rect 77300 4180 77301 4220
rect 77259 4171 77301 4180
rect 77452 4136 77492 4759
rect 77452 4087 77492 4096
rect 77548 4724 77588 4733
rect 77068 4052 77108 4061
rect 77068 3632 77108 4012
rect 77163 4052 77205 4061
rect 77163 4012 77164 4052
rect 77204 4012 77396 4052
rect 77163 4003 77205 4012
rect 77164 3918 77204 4003
rect 77260 3632 77300 3641
rect 77068 3592 77260 3632
rect 77260 3583 77300 3592
rect 77164 3464 77204 3473
rect 77356 3464 77396 4012
rect 77204 3424 77300 3464
rect 77164 3415 77204 3424
rect 76971 3128 77013 3137
rect 76971 3088 76972 3128
rect 77012 3088 77013 3128
rect 76971 3079 77013 3088
rect 76779 2876 76821 2885
rect 76779 2836 76780 2876
rect 76820 2836 76821 2876
rect 76876 2860 77012 2900
rect 77260 2885 77300 3424
rect 77356 3415 77396 3424
rect 77452 3464 77492 3473
rect 77548 3464 77588 4684
rect 77644 4313 77684 4768
rect 77835 4768 77836 4808
rect 77876 4768 77877 4808
rect 77835 4759 77877 4768
rect 77836 4674 77876 4759
rect 77643 4304 77685 4313
rect 77643 4264 77644 4304
rect 77684 4264 77685 4304
rect 77643 4255 77685 4264
rect 77644 3473 77684 4255
rect 78316 4136 78356 6448
rect 79468 6236 79508 6245
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 79468 5825 79508 6196
rect 79467 5816 79509 5825
rect 79467 5776 79468 5816
rect 79508 5776 79509 5816
rect 79467 5767 79509 5776
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 79467 4220 79509 4229
rect 79467 4180 79468 4220
rect 79508 4180 79509 4220
rect 79467 4171 79509 4180
rect 77492 3424 77588 3464
rect 77643 3464 77685 3473
rect 77643 3424 77644 3464
rect 77684 3424 77685 3464
rect 77452 3415 77492 3424
rect 77643 3415 77685 3424
rect 77835 3128 77877 3137
rect 77835 3088 77836 3128
rect 77876 3088 77877 3128
rect 77835 3079 77877 3088
rect 76779 2827 76821 2836
rect 76780 2624 76820 2827
rect 76780 2575 76820 2584
rect 76875 2624 76917 2633
rect 76875 2584 76876 2624
rect 76916 2584 76917 2624
rect 76972 2624 77012 2860
rect 77259 2876 77301 2885
rect 77259 2836 77260 2876
rect 77300 2836 77301 2876
rect 77259 2827 77301 2836
rect 77068 2624 77108 2633
rect 76972 2584 77068 2624
rect 76875 2575 76917 2584
rect 76203 2540 76245 2549
rect 76203 2500 76204 2540
rect 76244 2500 76245 2540
rect 76203 2491 76245 2500
rect 76683 2540 76725 2549
rect 76683 2500 76684 2540
rect 76724 2500 76725 2540
rect 76683 2491 76725 2500
rect 76052 1912 76148 1952
rect 76012 1903 76052 1912
rect 75819 1112 75861 1121
rect 75819 1072 75820 1112
rect 75860 1072 75861 1112
rect 75819 1063 75861 1072
rect 75916 1112 75956 1903
rect 75916 1063 75956 1072
rect 76012 1112 76052 1121
rect 76012 944 76052 1072
rect 76107 1112 76149 1121
rect 76107 1072 76108 1112
rect 76148 1072 76149 1112
rect 76107 1063 76149 1072
rect 76204 1112 76244 2491
rect 76876 1961 76916 2575
rect 77068 2045 77108 2584
rect 77163 2540 77205 2549
rect 77163 2500 77164 2540
rect 77204 2500 77205 2540
rect 77163 2491 77205 2500
rect 77164 2406 77204 2491
rect 77067 2036 77109 2045
rect 77067 1996 77068 2036
rect 77108 1996 77109 2036
rect 77067 1987 77109 1996
rect 76875 1952 76917 1961
rect 76875 1912 76876 1952
rect 76916 1912 76917 1952
rect 76875 1903 76917 1912
rect 76876 1818 76916 1903
rect 77068 1364 77108 1987
rect 77260 1877 77300 2827
rect 77452 2792 77492 2801
rect 77452 2624 77492 2752
rect 77644 2624 77684 2633
rect 77452 2584 77644 2624
rect 77644 2575 77684 2584
rect 77836 2624 77876 3079
rect 78123 2876 78165 2885
rect 78123 2836 78124 2876
rect 78164 2836 78165 2876
rect 78123 2827 78165 2836
rect 77836 2575 77876 2584
rect 77740 2540 77780 2549
rect 77740 2381 77780 2500
rect 78027 2540 78069 2549
rect 78027 2500 78028 2540
rect 78068 2500 78069 2540
rect 78027 2491 78069 2500
rect 77739 2372 77781 2381
rect 77739 2332 77740 2372
rect 77780 2332 77781 2372
rect 77739 2323 77781 2332
rect 77740 2129 77780 2323
rect 77739 2120 77781 2129
rect 77739 2080 77740 2120
rect 77780 2080 77781 2120
rect 77739 2071 77781 2080
rect 78028 2120 78068 2491
rect 78028 2071 78068 2080
rect 78124 1952 78164 2827
rect 78219 2792 78261 2801
rect 78219 2752 78220 2792
rect 78260 2752 78261 2792
rect 78219 2743 78261 2752
rect 78220 2658 78260 2743
rect 78316 1961 78356 4096
rect 79468 4086 79508 4171
rect 78603 3464 78645 3473
rect 78603 3424 78604 3464
rect 78644 3424 78645 3464
rect 78603 3415 78645 3424
rect 78411 2372 78453 2381
rect 78411 2332 78412 2372
rect 78452 2332 78453 2372
rect 78411 2323 78453 2332
rect 78220 1952 78260 1961
rect 78124 1912 78220 1952
rect 78220 1903 78260 1912
rect 78315 1952 78357 1961
rect 78315 1912 78316 1952
rect 78356 1912 78357 1952
rect 78315 1903 78357 1912
rect 78412 1952 78452 2323
rect 78412 1903 78452 1912
rect 78508 1952 78548 1961
rect 78604 1952 78644 3415
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 79179 2792 79221 2801
rect 79179 2752 79180 2792
rect 79220 2752 79221 2792
rect 79179 2743 79221 2752
rect 78700 1952 78740 1961
rect 78604 1912 78700 1952
rect 77259 1868 77301 1877
rect 77259 1828 77260 1868
rect 77300 1828 77301 1868
rect 77259 1819 77301 1828
rect 77068 1315 77108 1324
rect 78220 1700 78260 1709
rect 78220 1289 78260 1660
rect 78219 1280 78261 1289
rect 78219 1240 78220 1280
rect 78260 1240 78261 1280
rect 78219 1231 78261 1240
rect 76204 1063 76244 1072
rect 78220 1112 78260 1121
rect 78316 1112 78356 1903
rect 78508 1784 78548 1912
rect 78700 1903 78740 1912
rect 78891 1952 78933 1961
rect 78891 1912 78892 1952
rect 78932 1912 78933 1952
rect 78891 1903 78933 1912
rect 78892 1818 78932 1903
rect 78796 1784 78836 1793
rect 78508 1744 78796 1784
rect 78796 1735 78836 1744
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 78260 1072 78356 1112
rect 79084 1112 79124 1121
rect 79180 1112 79220 2743
rect 79467 1280 79509 1289
rect 79467 1240 79468 1280
rect 79508 1240 79509 1280
rect 79467 1231 79509 1240
rect 79124 1072 79220 1112
rect 79468 1112 79508 1231
rect 78220 1063 78260 1072
rect 79084 1063 79124 1072
rect 79468 1063 79508 1072
rect 76108 978 76148 1063
rect 75724 904 76052 944
rect 58540 895 58580 904
rect 73228 895 73268 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 56908 38032 56948 38072
rect 58252 38032 58292 38072
rect 652 37528 692 37568
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 844 25936 884 25976
rect 652 25768 692 25808
rect 844 25096 884 25136
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 844 23836 884 23876
rect 844 23584 884 23624
rect 652 23248 692 23288
rect 556 22408 596 22448
rect 652 21568 692 21608
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 54700 36772 54740 36812
rect 55660 37360 55700 37400
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 49228 36016 49268 36056
rect 50572 36016 50612 36056
rect 50380 35932 50420 35972
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 49708 35176 49748 35216
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 46156 34504 46196 34544
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 42220 32908 42260 32948
rect 42700 32908 42740 32948
rect 42124 32656 42164 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 41452 31312 41492 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 41068 31060 41108 31100
rect 40204 30808 40244 30848
rect 40204 30640 40244 30680
rect 40876 30556 40916 30596
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 39724 30220 39764 30260
rect 40204 30220 40244 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 37708 27700 37748 27740
rect 38380 28204 38420 28244
rect 38668 27868 38708 27908
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 33004 26944 33044 26984
rect 34252 26944 34292 26984
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 3916 25096 3956 25136
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 1996 23836 2036 23876
rect 1420 23584 1460 23624
rect 1804 23584 1844 23624
rect 2188 23584 2228 23624
rect 1516 23164 1556 23204
rect 1420 23080 1460 23120
rect 1900 23080 1940 23120
rect 2092 23080 2132 23120
rect 1708 22828 1748 22868
rect 2764 22828 2804 22868
rect 1900 21484 1940 21524
rect 940 20812 980 20852
rect 652 20728 692 20768
rect 844 20728 884 20768
rect 2668 20056 2708 20096
rect 1996 19972 2036 20012
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 1708 18460 1748 18500
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 844 14932 884 14972
rect 652 14848 692 14888
rect 1516 14932 1556 14972
rect 652 14008 692 14048
rect 652 13168 692 13208
rect 1324 14680 1364 14720
rect 1516 14176 1556 14216
rect 1228 13252 1268 13292
rect 652 12328 692 12368
rect 556 12244 596 12284
rect 1132 11740 1172 11780
rect 652 11488 692 11528
rect 1420 12664 1460 12704
rect 1324 12412 1364 12452
rect 1516 12244 1556 12284
rect 1036 10732 1076 10772
rect 652 9808 692 9848
rect 844 10060 884 10100
rect 652 8968 692 9008
rect 652 8128 692 8168
rect 652 7288 692 7328
rect 556 7204 596 7244
rect 652 6448 692 6488
rect 844 9388 884 9428
rect 844 9136 884 9176
rect 1036 8548 1076 8588
rect 2380 17116 2420 17156
rect 2188 16864 2228 16904
rect 2572 16528 2612 16568
rect 1804 15520 1844 15560
rect 1996 14848 2036 14888
rect 2188 14764 2228 14804
rect 1708 14596 1748 14636
rect 2188 14344 2228 14384
rect 1708 14008 1748 14048
rect 2092 14008 2132 14048
rect 2380 14680 2420 14720
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3052 21484 3092 21524
rect 3244 21400 3284 21440
rect 3628 21400 3668 21440
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 3628 21064 3668 21104
rect 3532 20728 3572 20768
rect 3820 21064 3860 21104
rect 3724 20560 3764 20600
rect 3628 20476 3668 20516
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4108 23080 4148 23120
rect 4012 21484 4052 21524
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 32236 25936 32276 25976
rect 33196 25936 33236 25976
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 35020 26860 35060 26900
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 34924 26272 34964 26312
rect 34444 26104 34484 26144
rect 34444 25936 34484 25976
rect 33388 25852 33428 25892
rect 33868 25852 33908 25892
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 31756 25348 31796 25388
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 29740 24760 29780 24800
rect 7468 24676 7508 24716
rect 4780 23080 4820 23120
rect 6988 21988 7028 22028
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4396 21484 4436 21524
rect 5068 20812 5108 20852
rect 4396 20644 4436 20684
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 5356 20476 5396 20516
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4108 18376 4148 18416
rect 3340 17116 3380 17156
rect 2956 16864 2996 16904
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4876 19804 4916 19844
rect 4876 18544 4916 18584
rect 4204 17032 4244 17072
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 3340 16444 3380 16484
rect 2572 14848 2612 14888
rect 2476 14344 2516 14384
rect 1996 13924 2036 13964
rect 1900 11152 1940 11192
rect 1804 11068 1844 11108
rect 1324 10984 1364 11024
rect 1516 10060 1556 10100
rect 1708 10396 1748 10436
rect 2284 13924 2324 13964
rect 2956 15688 2996 15728
rect 2860 15604 2900 15644
rect 3148 15520 3188 15560
rect 4012 16612 4052 16652
rect 3820 16276 3860 16316
rect 3628 16024 3668 16064
rect 3916 16024 3956 16064
rect 3820 15688 3860 15728
rect 3532 15604 3572 15644
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 2956 14428 2996 14468
rect 2668 14008 2708 14048
rect 3340 14680 3380 14720
rect 3244 14596 3284 14636
rect 3244 14428 3284 14468
rect 2572 13924 2612 13964
rect 4012 15772 4052 15812
rect 3532 14176 3572 14216
rect 2476 12832 2516 12872
rect 2380 12664 2420 12704
rect 2764 13168 2804 13208
rect 3628 14008 3668 14048
rect 3820 14008 3860 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 3532 13252 3572 13292
rect 2956 13168 2996 13208
rect 2668 12748 2708 12788
rect 2572 12328 2612 12368
rect 2764 12328 2804 12368
rect 2188 11152 2228 11192
rect 1612 9136 1652 9176
rect 1708 8716 1748 8756
rect 2284 10816 2324 10856
rect 2476 10984 2516 11024
rect 2476 10396 2516 10436
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4396 16444 4436 16484
rect 4204 16276 4244 16316
rect 4588 17032 4628 17072
rect 5068 19720 5108 19760
rect 5356 18544 5396 18584
rect 5164 17032 5204 17072
rect 5068 16612 5108 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4204 15772 4244 15812
rect 4396 15688 4436 15728
rect 4588 15520 4628 15560
rect 4780 15520 4820 15560
rect 4012 14596 4052 14636
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4204 14176 4244 14216
rect 5068 15520 5108 15560
rect 4876 14764 4916 14804
rect 4396 13168 4436 13208
rect 4108 12832 4148 12872
rect 4492 13000 4532 13040
rect 6988 16444 7028 16484
rect 7372 15268 7412 15308
rect 7276 14176 7316 14216
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 5164 13168 5204 13208
rect 4972 12748 5012 12788
rect 2956 11488 2996 11528
rect 3532 11488 3572 11528
rect 3436 11152 3476 11192
rect 3532 11068 3572 11108
rect 3724 11488 3764 11528
rect 4780 12496 4820 12536
rect 4012 11488 4052 11528
rect 4012 10984 4052 11024
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 2860 10312 2900 10352
rect 3052 10312 3092 10352
rect 3244 10228 3284 10268
rect 2572 8968 2612 9008
rect 2380 8632 2420 8672
rect 2284 8548 2324 8588
rect 940 7708 980 7748
rect 844 7204 884 7244
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 1036 7624 1076 7664
rect 1516 7708 1556 7748
rect 1996 7624 2036 7664
rect 1324 6280 1364 6320
rect 1804 5692 1844 5732
rect 1228 5104 1268 5144
rect 2870 9808 2910 9848
rect 2764 9304 2804 9344
rect 2764 8884 2804 8924
rect 3436 9808 3476 9848
rect 3532 9304 3572 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3340 8884 3380 8924
rect 3724 9472 3764 9512
rect 4684 11488 4724 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 5068 10984 5108 11024
rect 5452 12496 5492 12536
rect 5356 12328 5396 12368
rect 4876 10228 4916 10268
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3052 8800 3092 8840
rect 2956 8716 2996 8756
rect 3148 8716 3188 8756
rect 2668 8464 2708 8504
rect 2764 8044 2804 8084
rect 2572 7960 2612 8000
rect 2380 7036 2420 7076
rect 2188 6280 2228 6320
rect 2476 6280 2516 6320
rect 2668 6448 2708 6488
rect 2878 7960 2918 8000
rect 3724 8632 3764 8672
rect 2878 7624 2918 7664
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2860 6700 2900 6740
rect 3724 7960 3764 8000
rect 3628 7708 3668 7748
rect 4108 9304 4148 9344
rect 4588 9472 4628 9512
rect 5068 9976 5108 10016
rect 5068 8800 5108 8840
rect 4108 8464 4148 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4300 7960 4340 8000
rect 4108 7036 4148 7076
rect 4972 7708 5012 7748
rect 4492 7036 4532 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3532 6532 3572 6572
rect 2668 6280 2708 6320
rect 2668 6028 2708 6068
rect 2476 5608 2516 5648
rect 2284 5104 2324 5144
rect 2476 5104 2516 5144
rect 1804 4852 1844 4892
rect 2188 4852 2228 4892
rect 1900 4600 1940 4640
rect 1036 3928 1076 3968
rect 1228 3340 1268 3380
rect 652 3172 692 3212
rect 844 2752 884 2792
rect 2092 4096 2132 4136
rect 2380 4768 2420 4808
rect 2476 4684 2516 4724
rect 2284 4600 2324 4640
rect 2092 3340 2132 3380
rect 1516 2752 1556 2792
rect 1708 2668 1748 2708
rect 3052 6448 3092 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 2956 5692 2996 5732
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 2878 4096 2918 4136
rect 3628 5692 3668 5732
rect 4876 6700 4916 6740
rect 4492 6532 4532 6572
rect 4204 6448 4244 6488
rect 5836 12328 5876 12368
rect 5644 11656 5684 11696
rect 6220 11656 6260 11696
rect 7372 10984 7412 11024
rect 7180 9976 7220 10016
rect 30988 25264 31028 25304
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 28396 23080 28436 23120
rect 29548 23920 29588 23960
rect 30892 23920 30932 23960
rect 31660 25096 31700 25136
rect 31084 23668 31124 23708
rect 32812 25264 32852 25304
rect 33004 25180 33044 25220
rect 32140 25096 32180 25136
rect 31852 24844 31892 24884
rect 31660 23752 31700 23792
rect 31468 23668 31508 23708
rect 28972 23164 29012 23204
rect 29548 23164 29588 23204
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 28300 22492 28340 22532
rect 27628 22408 27668 22448
rect 27916 22408 27956 22448
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 23212 21652 23252 21692
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 22828 20560 22868 20600
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 10828 19972 10868 20012
rect 11116 20056 11156 20096
rect 9580 19552 9620 19592
rect 10924 19552 10964 19592
rect 10060 19216 10100 19256
rect 11692 20056 11732 20096
rect 8908 18712 8948 18752
rect 11020 18712 11060 18752
rect 8620 15184 8660 15224
rect 8620 14176 8660 14216
rect 7468 8464 7508 8504
rect 7180 7708 7220 7748
rect 5068 6448 5108 6488
rect 7372 6448 7412 6488
rect 4108 5776 4148 5816
rect 4108 5608 4148 5648
rect 3820 4768 3860 4808
rect 3916 4096 3956 4136
rect 3820 4012 3860 4052
rect 2572 2584 2612 2624
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 4780 4768 4820 4808
rect 4012 3592 4052 3632
rect 2956 3424 2996 3464
rect 4588 4096 4628 4136
rect 6220 5608 6260 5648
rect 7372 5440 7412 5480
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 5260 4012 5300 4052
rect 4396 3592 4436 3632
rect 4588 3256 4628 3296
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 3148 2668 3188 2708
rect 1420 2500 1460 2540
rect 2476 2500 2516 2540
rect 5068 3424 5108 3464
rect 5260 3424 5300 3464
rect 7468 3424 7508 3464
rect 10924 18460 10964 18500
rect 10636 16528 10676 16568
rect 21772 19804 21812 19844
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 14668 19468 14708 19508
rect 21772 19300 21812 19340
rect 11884 19132 11924 19172
rect 12076 18628 12116 18668
rect 13516 19216 13556 19256
rect 12268 19132 12308 19172
rect 22348 19132 22388 19172
rect 21964 18964 22004 19004
rect 22252 18964 22292 19004
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 22540 19048 22580 19088
rect 22444 18712 22484 18752
rect 22156 18544 22196 18584
rect 12268 18460 12308 18500
rect 14668 18460 14708 18500
rect 22348 18460 22388 18500
rect 21964 18292 22004 18332
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 26188 20896 26228 20936
rect 25900 20812 25940 20852
rect 25516 20140 25556 20180
rect 23500 19804 23540 19844
rect 23692 19804 23732 19844
rect 23020 18712 23060 18752
rect 22924 18292 22964 18332
rect 22732 17704 22772 17744
rect 22924 17704 22964 17744
rect 23404 18544 23444 18584
rect 23212 17620 23252 17660
rect 23116 17536 23156 17576
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 21964 17368 22004 17408
rect 26380 20812 26420 20852
rect 23692 18460 23732 18500
rect 24460 18880 24500 18920
rect 23980 18292 24020 18332
rect 25036 18712 25076 18752
rect 24844 18628 24884 18668
rect 24268 18208 24308 18248
rect 23884 18124 23924 18164
rect 24076 18124 24116 18164
rect 24268 17788 24308 17828
rect 23692 17704 23732 17744
rect 23596 17536 23636 17576
rect 23500 17116 23540 17156
rect 23788 17452 23828 17492
rect 23404 16948 23444 16988
rect 11788 16612 11828 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 24844 18460 24884 18500
rect 24748 18292 24788 18332
rect 25420 19048 25460 19088
rect 25900 19132 25940 19172
rect 25804 18964 25844 19004
rect 25996 18796 26036 18836
rect 25708 18712 25748 18752
rect 26668 20560 26708 20600
rect 26572 20056 26612 20096
rect 26764 20140 26804 20180
rect 26380 19888 26420 19928
rect 26572 19888 26612 19928
rect 26956 21484 26996 21524
rect 27148 21400 27188 21440
rect 27532 20896 27572 20936
rect 27148 20812 27188 20852
rect 27724 22324 27764 22364
rect 28204 22324 28244 22364
rect 27340 20728 27380 20768
rect 27628 20728 27668 20768
rect 26956 20560 26996 20600
rect 27340 20560 27380 20600
rect 26956 19888 26996 19928
rect 28492 22240 28532 22280
rect 28204 21652 28244 21692
rect 27820 21568 27860 21608
rect 28012 21148 28052 21188
rect 27916 20728 27956 20768
rect 28684 22072 28724 22112
rect 28300 21148 28340 21188
rect 28588 21568 28628 21608
rect 28492 21400 28532 21440
rect 28492 20728 28532 20768
rect 28876 21568 28916 21608
rect 29068 21736 29108 21776
rect 29452 21568 29492 21608
rect 28972 20812 29012 20852
rect 28876 20728 28916 20768
rect 27820 20140 27860 20180
rect 28972 19804 29012 19844
rect 29068 19384 29108 19424
rect 29260 19384 29300 19424
rect 27724 19300 27764 19340
rect 26188 18712 26228 18752
rect 26476 19048 26516 19088
rect 26380 18544 26420 18584
rect 27244 18796 27284 18836
rect 26860 18628 26900 18668
rect 26764 18544 26804 18584
rect 26092 18460 26132 18500
rect 25516 18376 25556 18416
rect 24556 18040 24596 18080
rect 28588 18796 28628 18836
rect 27820 18544 27860 18584
rect 27436 18292 27476 18332
rect 29068 19132 29108 19172
rect 28972 18712 29012 18752
rect 28396 18292 28436 18332
rect 27916 18208 27956 18248
rect 26668 17620 26708 17660
rect 25804 17536 25844 17576
rect 25324 17452 25364 17492
rect 27244 17452 27284 17492
rect 27436 17536 27476 17576
rect 24556 16948 24596 16988
rect 28972 18460 29012 18500
rect 29836 22240 29876 22280
rect 29644 22072 29684 22112
rect 30796 22492 30836 22532
rect 30700 22408 30740 22448
rect 30604 22240 30644 22280
rect 30028 22072 30068 22112
rect 30028 21904 30068 21944
rect 30316 20980 30356 21020
rect 29548 20056 29588 20096
rect 29548 19804 29588 19844
rect 29932 19132 29972 19172
rect 30220 19300 30260 19340
rect 30124 19048 30164 19088
rect 29452 18964 29492 19004
rect 30028 18964 30068 19004
rect 29356 18040 29396 18080
rect 28780 17452 28820 17492
rect 24460 16276 24500 16316
rect 11692 16024 11732 16064
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 29740 18712 29780 18752
rect 30988 22912 31028 22952
rect 30796 20476 30836 20516
rect 31180 23416 31220 23456
rect 31180 23080 31220 23120
rect 31372 23416 31412 23456
rect 31180 22324 31220 22364
rect 32236 24760 32276 24800
rect 32428 24592 32468 24632
rect 33868 25264 33908 25304
rect 34540 25264 34580 25304
rect 33484 25180 33524 25220
rect 33100 25012 33140 25052
rect 33292 25096 33332 25136
rect 33484 24844 33524 24884
rect 32716 24256 32756 24296
rect 32140 23836 32180 23876
rect 32236 23752 32276 23792
rect 31564 22408 31604 22448
rect 32140 23164 32180 23204
rect 31852 23080 31892 23120
rect 31756 22996 31796 23036
rect 31660 22324 31700 22364
rect 32236 23080 32276 23120
rect 32716 23836 32756 23876
rect 32620 23248 32660 23288
rect 32140 22996 32180 23036
rect 31564 22240 31604 22280
rect 31756 22240 31796 22280
rect 31468 21652 31508 21692
rect 31756 21400 31796 21440
rect 31372 20560 31412 20600
rect 31660 19300 31700 19340
rect 30316 18880 30356 18920
rect 29644 18208 29684 18248
rect 29836 17704 29876 17744
rect 29932 17620 29972 17660
rect 29548 17536 29588 17576
rect 30316 17620 30356 17660
rect 30220 17452 30260 17492
rect 30124 17116 30164 17156
rect 31084 19216 31124 19256
rect 30700 18628 30740 18668
rect 31180 18544 31220 18584
rect 31660 18544 31700 18584
rect 30508 18292 30548 18332
rect 31564 18292 31604 18332
rect 30412 17284 30452 17324
rect 30604 17284 30644 17324
rect 30508 17116 30548 17156
rect 31372 17704 31412 17744
rect 31564 17704 31604 17744
rect 31276 17368 31316 17408
rect 31084 15856 31124 15896
rect 29452 15520 29492 15560
rect 30220 15352 30260 15392
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 30220 14008 30260 14048
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 31564 15352 31604 15392
rect 31852 19300 31892 19340
rect 32332 22240 32372 22280
rect 32236 22156 32276 22196
rect 32332 21652 32372 21692
rect 32716 23080 32756 23120
rect 33196 24592 33236 24632
rect 34636 25180 34676 25220
rect 35596 26860 35636 26900
rect 35212 26776 35252 26816
rect 35308 26104 35348 26144
rect 35212 25936 35252 25976
rect 35692 26776 35732 26816
rect 39628 28540 39668 28580
rect 40780 30388 40820 30428
rect 40012 29800 40052 29840
rect 40012 28708 40052 28748
rect 40684 29800 40724 29840
rect 40780 29128 40820 29168
rect 40396 28624 40436 28664
rect 40396 28456 40436 28496
rect 35788 26272 35828 26312
rect 37036 26356 37076 26396
rect 35116 25852 35156 25892
rect 35596 25264 35636 25304
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 35020 24844 35060 24884
rect 33868 24508 33908 24548
rect 34156 24424 34196 24464
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 33004 23668 33044 23708
rect 32908 23248 32948 23288
rect 32908 22408 32948 22448
rect 32812 22156 32852 22196
rect 32908 21820 32948 21860
rect 32140 21568 32180 21608
rect 32620 21568 32660 21608
rect 32716 20476 32756 20516
rect 32524 20224 32564 20264
rect 32044 19384 32084 19424
rect 31948 19048 31988 19088
rect 31852 18964 31892 19004
rect 31852 18124 31892 18164
rect 31756 17452 31796 17492
rect 31852 15604 31892 15644
rect 31468 14680 31508 14720
rect 31276 14092 31316 14132
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 33004 20140 33044 20180
rect 32908 19888 32948 19928
rect 33004 19552 33044 19592
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 32908 19384 32948 19424
rect 33292 19384 33332 19424
rect 32236 18712 32276 18752
rect 32620 18712 32660 18752
rect 32140 18460 32180 18500
rect 32332 18460 32372 18500
rect 33004 18628 33044 18668
rect 33196 18628 33236 18668
rect 32428 18376 32468 18416
rect 32812 18208 32852 18248
rect 32716 17956 32756 17996
rect 32428 17788 32468 17828
rect 32332 17704 32372 17744
rect 32140 17620 32180 17660
rect 32716 17284 32756 17324
rect 32908 17284 32948 17324
rect 32140 15604 32180 15644
rect 31756 14932 31796 14972
rect 31756 14428 31796 14468
rect 31564 14008 31604 14048
rect 32044 14764 32084 14804
rect 32428 15520 32468 15560
rect 32236 14512 32276 14552
rect 32716 14932 32756 14972
rect 32620 14512 32660 14552
rect 32428 14428 32468 14468
rect 31852 14176 31892 14216
rect 32236 14092 32276 14132
rect 31948 13924 31988 13964
rect 32620 13924 32660 13964
rect 32620 13252 32660 13292
rect 31660 13168 31700 13208
rect 33868 18712 33908 18752
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 33388 17956 33428 17996
rect 33196 17704 33236 17744
rect 33484 17704 33524 17744
rect 35692 25012 35732 25052
rect 35596 24928 35636 24968
rect 35212 24256 35252 24296
rect 35116 23920 35156 23960
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 35692 24088 35732 24128
rect 36268 26104 36308 26144
rect 36460 26104 36500 26144
rect 35980 25852 36020 25892
rect 36172 25852 36212 25892
rect 35884 25432 35924 25472
rect 35884 24760 35924 24800
rect 36076 25180 36116 25220
rect 36460 25936 36500 25976
rect 36556 24844 36596 24884
rect 36268 24760 36308 24800
rect 36172 24592 36212 24632
rect 36172 23920 36212 23960
rect 36076 23752 36116 23792
rect 35788 23164 35828 23204
rect 35212 22492 35252 22532
rect 35692 22156 35732 22196
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 35212 21652 35252 21692
rect 36940 24592 36980 24632
rect 36652 23752 36692 23792
rect 36268 23584 36308 23624
rect 36268 23332 36308 23372
rect 36460 22576 36500 22616
rect 36268 22156 36308 22196
rect 36172 21904 36212 21944
rect 36844 23248 36884 23288
rect 38380 26104 38420 26144
rect 38092 26020 38132 26060
rect 37228 25852 37268 25892
rect 38092 25432 38132 25472
rect 37228 25264 37268 25304
rect 37036 24424 37076 24464
rect 38476 25852 38516 25892
rect 38476 25180 38516 25220
rect 38380 25096 38420 25136
rect 38860 26860 38900 26900
rect 39628 27196 39668 27236
rect 39052 26860 39092 26900
rect 39820 27616 39860 27656
rect 40396 28288 40436 28328
rect 41644 30724 41684 30764
rect 41740 30640 41780 30680
rect 41452 30556 41492 30596
rect 42124 30556 42164 30596
rect 41644 30472 41684 30512
rect 41068 28960 41108 29000
rect 40972 28372 41012 28412
rect 41356 29716 41396 29756
rect 41548 29632 41588 29672
rect 41260 28960 41300 29000
rect 41260 28372 41300 28412
rect 40972 28204 41012 28244
rect 40396 27700 40436 27740
rect 40300 27616 40340 27656
rect 40972 27616 41012 27656
rect 40492 27364 40532 27404
rect 41068 27364 41108 27404
rect 40492 27112 40532 27152
rect 39724 26692 39764 26732
rect 39916 26692 39956 26732
rect 39628 26608 39668 26648
rect 39244 26188 39284 26228
rect 40108 26776 40148 26816
rect 39820 26188 39860 26228
rect 38956 26020 38996 26060
rect 38860 25852 38900 25892
rect 39148 25600 39188 25640
rect 39532 25684 39572 25724
rect 39532 25516 39572 25556
rect 39436 25348 39476 25388
rect 39340 25264 39380 25304
rect 39628 25264 39668 25304
rect 39820 25264 39860 25304
rect 40204 26692 40244 26732
rect 40012 25516 40052 25556
rect 40108 25348 40148 25388
rect 39148 25012 39188 25052
rect 37996 24760 38036 24800
rect 37516 24088 37556 24128
rect 37324 23752 37364 23792
rect 37036 23332 37076 23372
rect 37324 23164 37364 23204
rect 37900 23248 37940 23288
rect 36748 22576 36788 22616
rect 37132 22912 37172 22952
rect 37228 22576 37268 22616
rect 36556 21736 36596 21776
rect 35788 21568 35828 21608
rect 36076 21568 36116 21608
rect 36268 21568 36308 21608
rect 36172 21484 36212 21524
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 36076 20476 36116 20516
rect 34444 19888 34484 19928
rect 34828 19888 34868 19928
rect 35020 19804 35060 19844
rect 34924 19636 34964 19676
rect 36460 21568 36500 21608
rect 36748 21652 36788 21692
rect 36268 19888 36308 19928
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 35308 18628 35348 18668
rect 34252 18544 34292 18584
rect 34156 18460 34196 18500
rect 35500 18460 35540 18500
rect 34348 17788 34388 17828
rect 33964 17284 34004 17324
rect 34348 17536 34388 17576
rect 34060 17116 34100 17156
rect 33004 16276 33044 16316
rect 33580 17032 33620 17072
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 34060 16696 34100 16736
rect 33868 16444 33908 16484
rect 33772 16276 33812 16316
rect 34252 16444 34292 16484
rect 33196 15688 33236 15728
rect 33964 15856 34004 15896
rect 33484 15772 33524 15812
rect 32908 14932 32948 14972
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 35116 17284 35156 17324
rect 35788 18628 35828 18668
rect 35692 18544 35732 18584
rect 36172 18628 36212 18668
rect 35692 18376 35732 18416
rect 38092 23752 38132 23792
rect 37612 23020 37652 23060
rect 37996 22912 38036 22952
rect 38092 22156 38132 22196
rect 38092 21652 38132 21692
rect 39244 24088 39284 24128
rect 38860 23920 38900 23960
rect 38764 23752 38804 23792
rect 39724 25180 39764 25220
rect 38956 23584 38996 23624
rect 38476 23080 38516 23120
rect 39148 23080 39188 23120
rect 39244 22240 39284 22280
rect 39628 24424 39668 24464
rect 40396 26692 40436 26732
rect 40300 26188 40340 26228
rect 40012 25180 40052 25220
rect 40204 25180 40244 25220
rect 40876 27028 40916 27068
rect 41452 29128 41492 29168
rect 41548 28624 41588 28664
rect 41452 28540 41492 28580
rect 41452 28288 41492 28328
rect 41356 27784 41396 27824
rect 41260 27196 41300 27236
rect 40780 26776 40820 26816
rect 40684 26356 40724 26396
rect 41548 28204 41588 28244
rect 41548 27364 41588 27404
rect 41452 26944 41492 26984
rect 42892 32656 42932 32696
rect 42412 32488 42452 32528
rect 42316 31144 42356 31184
rect 42316 30556 42356 30596
rect 42220 30304 42260 30344
rect 42124 29968 42164 30008
rect 41836 29716 41876 29756
rect 41740 29632 41780 29672
rect 41740 28792 41780 28832
rect 42028 28960 42068 29000
rect 41932 28540 41972 28580
rect 42220 28876 42260 28916
rect 42604 31144 42644 31184
rect 42508 30976 42548 31016
rect 42604 30640 42644 30680
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 49228 34504 49268 34544
rect 47020 34168 47060 34208
rect 46828 33160 46868 33200
rect 46060 32908 46100 32948
rect 46252 32908 46292 32948
rect 44716 32488 44756 32528
rect 44620 32152 44660 32192
rect 42892 31228 42932 31268
rect 42796 30808 42836 30848
rect 43084 31144 43124 31184
rect 43468 31228 43508 31268
rect 43468 31060 43508 31100
rect 43852 31144 43892 31184
rect 43180 30892 43220 30932
rect 42988 30472 43028 30512
rect 42508 30388 42548 30428
rect 42796 30304 42836 30344
rect 42412 29800 42452 29840
rect 42316 28708 42356 28748
rect 41740 27028 41780 27068
rect 42604 28204 42644 28244
rect 41644 26860 41684 26900
rect 41452 26356 41492 26396
rect 41260 26104 41300 26144
rect 40780 25684 40820 25724
rect 40396 25516 40436 25556
rect 39916 25012 39956 25052
rect 39916 24592 39956 24632
rect 40012 24424 40052 24464
rect 38380 21064 38420 21104
rect 38380 20896 38420 20936
rect 37612 20224 37652 20264
rect 38284 20224 38324 20264
rect 37708 19888 37748 19928
rect 37516 19804 37556 19844
rect 38092 19888 38132 19928
rect 37900 19636 37940 19676
rect 36460 18460 36500 18500
rect 36364 18208 36404 18248
rect 36652 18208 36692 18248
rect 36460 17872 36500 17912
rect 35596 17284 35636 17324
rect 34732 16444 34772 16484
rect 36652 16780 36692 16820
rect 37420 18460 37460 18500
rect 37036 17956 37076 17996
rect 36844 17788 36884 17828
rect 36844 17452 36884 17492
rect 36844 16276 36884 16316
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 35596 15772 35636 15812
rect 37132 16864 37172 16904
rect 37036 16192 37076 16232
rect 38092 17116 38132 17156
rect 37324 16444 37364 16484
rect 37996 16444 38036 16484
rect 37516 16360 37556 16400
rect 37708 16192 37748 16232
rect 36364 15772 36404 15812
rect 34828 15688 34868 15728
rect 35212 15688 35252 15728
rect 33580 15436 33620 15476
rect 34348 15520 34388 15560
rect 34156 15352 34196 15392
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 33100 14848 33140 14888
rect 33388 14764 33428 14804
rect 32812 13504 32852 13544
rect 33100 13504 33140 13544
rect 35116 15604 35156 15644
rect 34924 15520 34964 15560
rect 34924 15352 34964 15392
rect 34348 14848 34388 14888
rect 35404 15436 35444 15476
rect 35212 14848 35252 14888
rect 35116 14764 35156 14804
rect 34348 14680 34388 14720
rect 33772 14176 33812 14216
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 34924 13252 34964 13292
rect 32812 13168 32852 13208
rect 35020 13168 35060 13208
rect 35308 14680 35348 14720
rect 35212 13084 35252 13124
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 29932 12496 29972 12536
rect 31372 12496 31412 12536
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 33868 11908 33908 11948
rect 34828 11908 34868 11948
rect 35020 11824 35060 11864
rect 34828 11656 34868 11696
rect 35308 11656 35348 11696
rect 35500 13252 35540 13292
rect 36268 15688 36308 15728
rect 35980 15520 36020 15560
rect 35692 15100 35732 15140
rect 36460 15436 36500 15476
rect 37228 15688 37268 15728
rect 36940 15604 36980 15644
rect 37804 15604 37844 15644
rect 36556 15352 36596 15392
rect 36844 15352 36884 15392
rect 35980 14680 36020 14720
rect 36844 15100 36884 15140
rect 36748 14680 36788 14720
rect 37228 14680 37268 14720
rect 37516 15520 37556 15560
rect 37324 14428 37364 14468
rect 37420 14344 37460 14384
rect 37132 14092 37172 14132
rect 36748 13336 36788 13376
rect 35980 13084 36020 13124
rect 35596 12328 35636 12368
rect 35500 11572 35540 11612
rect 35404 11488 35444 11528
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 36556 12664 36596 12704
rect 36268 12328 36308 12368
rect 36748 12328 36788 12368
rect 36172 11908 36212 11948
rect 36268 11824 36308 11864
rect 36652 11824 36692 11864
rect 37324 14008 37364 14048
rect 36844 11656 36884 11696
rect 35980 10984 36020 11024
rect 36556 11068 36596 11108
rect 36748 10984 36788 11024
rect 37036 10984 37076 11024
rect 38092 14680 38132 14720
rect 38284 19888 38324 19928
rect 38476 20728 38516 20768
rect 39148 21568 39188 21608
rect 39052 20896 39092 20936
rect 38956 20728 38996 20768
rect 39148 20728 39188 20768
rect 39436 20728 39476 20768
rect 39436 20560 39476 20600
rect 39340 20140 39380 20180
rect 38668 19888 38708 19928
rect 38476 19804 38516 19844
rect 38380 18628 38420 18668
rect 39148 20056 39188 20096
rect 39052 19804 39092 19844
rect 38956 19216 38996 19256
rect 40492 24928 40532 24968
rect 40588 24844 40628 24884
rect 40876 24928 40916 24968
rect 40204 24508 40244 24548
rect 40684 24508 40724 24548
rect 41164 24844 41204 24884
rect 40876 24508 40916 24548
rect 40108 24340 40148 24380
rect 41164 24592 41204 24632
rect 41068 24508 41108 24548
rect 41740 26692 41780 26732
rect 40876 23920 40916 23960
rect 40492 23836 40532 23876
rect 40684 23836 40724 23876
rect 40108 23416 40148 23456
rect 40204 22072 40244 22112
rect 39532 19636 39572 19676
rect 39436 19384 39476 19424
rect 40780 23752 40820 23792
rect 40876 23248 40916 23288
rect 41644 24340 41684 24380
rect 41452 23920 41492 23960
rect 41260 23836 41300 23876
rect 40780 22240 40820 22280
rect 40684 21652 40724 21692
rect 41356 23248 41396 23288
rect 42124 25264 42164 25304
rect 42316 24592 42356 24632
rect 42220 23836 42260 23876
rect 41740 23668 41780 23708
rect 41644 23164 41684 23204
rect 41548 22912 41588 22952
rect 41356 21904 41396 21944
rect 41260 21652 41300 21692
rect 40492 20980 40532 21020
rect 40972 20140 41012 20180
rect 40780 19888 40820 19928
rect 40396 19636 40436 19676
rect 40780 19552 40820 19592
rect 40396 19300 40436 19340
rect 39436 19216 39476 19256
rect 39436 18712 39476 18752
rect 38668 18544 38708 18584
rect 38572 18460 38612 18500
rect 38572 18208 38612 18248
rect 38284 17956 38324 17996
rect 38284 17284 38324 17324
rect 38956 17788 38996 17828
rect 38476 16360 38516 16400
rect 38380 15604 38420 15644
rect 38572 15520 38612 15560
rect 38572 14428 38612 14468
rect 38092 11908 38132 11948
rect 37996 11656 38036 11696
rect 37612 11572 37652 11612
rect 38092 11572 38132 11612
rect 37516 11488 37556 11528
rect 37708 10984 37748 11024
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 36460 10144 36500 10184
rect 37228 10144 37268 10184
rect 38572 14008 38612 14048
rect 38476 13084 38516 13124
rect 38764 14008 38804 14048
rect 38668 13168 38708 13208
rect 38860 11992 38900 12032
rect 38860 11656 38900 11696
rect 38860 11320 38900 11360
rect 39244 16444 39284 16484
rect 39148 15520 39188 15560
rect 39436 14680 39476 14720
rect 39340 14596 39380 14636
rect 39148 14344 39188 14384
rect 39340 14260 39380 14300
rect 39148 14008 39188 14048
rect 43372 30724 43412 30764
rect 43756 30640 43796 30680
rect 43756 30472 43796 30512
rect 43948 30640 43988 30680
rect 43852 29968 43892 30008
rect 45004 32152 45044 32192
rect 44812 31648 44852 31688
rect 45004 31312 45044 31352
rect 44812 30976 44852 31016
rect 44716 30220 44756 30260
rect 44620 30052 44660 30092
rect 43084 29716 43124 29756
rect 43468 29296 43508 29336
rect 45772 30892 45812 30932
rect 46444 32572 46484 32612
rect 46348 31732 46388 31772
rect 46156 31564 46196 31604
rect 45004 30220 45044 30260
rect 45964 30220 46004 30260
rect 46060 30136 46100 30176
rect 45868 30052 45908 30092
rect 45004 29296 45044 29336
rect 45100 29128 45140 29168
rect 46348 30304 46388 30344
rect 46252 30136 46292 30176
rect 46156 29212 46196 29252
rect 46348 30052 46388 30092
rect 47020 33160 47060 33200
rect 47116 32824 47156 32864
rect 47788 32908 47828 32948
rect 47308 32572 47348 32612
rect 46924 32488 46964 32528
rect 47308 32152 47348 32192
rect 46828 31900 46868 31940
rect 46732 31564 46772 31604
rect 46636 31312 46676 31352
rect 47212 31312 47252 31352
rect 47212 30640 47252 30680
rect 46444 29716 46484 29756
rect 46060 29128 46100 29168
rect 44140 27784 44180 27824
rect 43564 27700 43604 27740
rect 43276 27616 43316 27656
rect 43084 27364 43124 27404
rect 45004 27784 45044 27824
rect 43372 27112 43412 27152
rect 43276 26776 43316 26816
rect 43180 26188 43220 26228
rect 42988 25264 43028 25304
rect 43276 24760 43316 24800
rect 44716 26860 44756 26900
rect 44044 26356 44084 26396
rect 43660 26104 43700 26144
rect 43660 25852 43700 25892
rect 43660 25264 43700 25304
rect 44044 25180 44084 25220
rect 43372 23500 43412 23540
rect 42028 22912 42068 22952
rect 42412 22240 42452 22280
rect 42412 21652 42452 21692
rect 42508 21568 42548 21608
rect 41260 19384 41300 19424
rect 41548 20980 41588 21020
rect 42412 20896 42452 20936
rect 42508 20728 42548 20768
rect 41644 19552 41684 19592
rect 41452 19132 41492 19172
rect 40972 19048 41012 19088
rect 40204 18628 40244 18668
rect 40012 18544 40052 18584
rect 39820 17704 39860 17744
rect 40396 18460 40436 18500
rect 39724 16864 39764 16904
rect 40108 16276 40148 16316
rect 39820 16024 39860 16064
rect 39916 15856 39956 15896
rect 40204 15940 40244 15980
rect 40300 15856 40340 15896
rect 40204 15520 40244 15560
rect 40012 15436 40052 15476
rect 40012 14680 40052 14720
rect 39724 14512 39764 14552
rect 41164 18712 41204 18752
rect 41068 18544 41108 18584
rect 41548 18376 41588 18416
rect 41932 19384 41972 19424
rect 42892 20560 42932 20600
rect 42796 20476 42836 20516
rect 42604 19972 42644 20012
rect 42508 19636 42548 19676
rect 42316 19216 42356 19256
rect 42124 19132 42164 19172
rect 42028 18712 42068 18752
rect 41644 18124 41684 18164
rect 41740 17956 41780 17996
rect 42124 18544 42164 18584
rect 42028 18376 42068 18416
rect 41164 17284 41204 17324
rect 41932 17704 41972 17744
rect 41932 17116 41972 17156
rect 41068 17032 41108 17072
rect 41452 16948 41492 16988
rect 40492 15940 40532 15980
rect 41836 17032 41876 17072
rect 40588 15688 40628 15728
rect 40492 15520 40532 15560
rect 40876 15520 40916 15560
rect 39820 14176 39860 14216
rect 39628 14092 39668 14132
rect 41164 14176 41204 14216
rect 39244 13924 39284 13964
rect 40108 13840 40148 13880
rect 39340 13336 39380 13376
rect 40396 14008 40436 14048
rect 40300 13084 40340 13124
rect 41356 14260 41396 14300
rect 41260 13924 41300 13964
rect 39532 12328 39572 12368
rect 39148 11992 39188 12032
rect 38956 10984 38996 11024
rect 40684 12496 40724 12536
rect 39436 11572 39476 11612
rect 39340 11068 39380 11108
rect 39532 11320 39572 11360
rect 39148 10900 39188 10940
rect 39532 10900 39572 10940
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 39340 10060 39380 10100
rect 40972 10060 41012 10100
rect 40684 9640 40724 9680
rect 40876 9556 40916 9596
rect 40108 9472 40148 9512
rect 40780 9472 40820 9512
rect 41260 9556 41300 9596
rect 41836 15940 41876 15980
rect 42220 18292 42260 18332
rect 42124 18124 42164 18164
rect 42220 17200 42260 17240
rect 42700 19804 42740 19844
rect 42604 18628 42644 18668
rect 42796 19216 42836 19256
rect 42796 18544 42836 18584
rect 42508 18376 42548 18416
rect 42412 18292 42452 18332
rect 42604 17788 42644 17828
rect 43564 22492 43604 22532
rect 44140 25012 44180 25052
rect 44908 27028 44948 27068
rect 45100 27028 45140 27068
rect 45292 26944 45332 26984
rect 45004 26608 45044 26648
rect 44908 25936 44948 25976
rect 44908 25348 44948 25388
rect 45100 26104 45140 26144
rect 45196 25432 45236 25472
rect 45676 28288 45716 28328
rect 45580 27700 45620 27740
rect 46348 28288 46388 28328
rect 45964 27784 46004 27824
rect 46444 27784 46484 27824
rect 46540 27700 46580 27740
rect 47116 30304 47156 30344
rect 46924 30220 46964 30260
rect 46348 27532 46388 27572
rect 45676 26944 45716 26984
rect 46060 26944 46100 26984
rect 45676 26608 45716 26648
rect 45772 25936 45812 25976
rect 45580 25852 45620 25892
rect 45484 25432 45524 25472
rect 45388 25180 45428 25220
rect 44428 24592 44468 24632
rect 44236 24256 44276 24296
rect 43948 23584 43988 23624
rect 43660 22240 43700 22280
rect 43564 21904 43604 21944
rect 44044 21568 44084 21608
rect 43948 20896 43988 20936
rect 43084 20812 43124 20852
rect 43084 20560 43124 20600
rect 43276 20560 43316 20600
rect 43084 20140 43124 20180
rect 43276 20140 43316 20180
rect 43084 19972 43124 20012
rect 42988 19804 43028 19844
rect 42892 18460 42932 18500
rect 42892 18292 42932 18332
rect 42892 18124 42932 18164
rect 42796 17704 42836 17744
rect 42700 17620 42740 17660
rect 42604 17116 42644 17156
rect 42028 15940 42068 15980
rect 41548 14008 41588 14048
rect 41644 13168 41684 13208
rect 42028 15520 42068 15560
rect 41932 13840 41972 13880
rect 41548 13084 41588 13124
rect 41548 12328 41588 12368
rect 41548 11656 41588 11696
rect 42220 14680 42260 14720
rect 41932 12496 41972 12536
rect 42412 16444 42452 16484
rect 42508 16276 42548 16316
rect 42604 16024 42644 16064
rect 42508 15520 42548 15560
rect 42412 13588 42452 13628
rect 43276 19720 43316 19760
rect 43084 18880 43124 18920
rect 43180 18628 43220 18668
rect 43084 18460 43124 18500
rect 43084 18040 43124 18080
rect 43084 17620 43124 17660
rect 42988 17200 43028 17240
rect 42892 17032 42932 17072
rect 42796 16360 42836 16400
rect 43084 16864 43124 16904
rect 43660 20812 43700 20852
rect 44716 24256 44756 24296
rect 44620 23752 44660 23792
rect 44428 23584 44468 23624
rect 44524 23500 44564 23540
rect 44620 23164 44660 23204
rect 45580 25264 45620 25304
rect 45484 25012 45524 25052
rect 44908 24424 44948 24464
rect 45004 23920 45044 23960
rect 45004 23668 45044 23708
rect 45004 23416 45044 23456
rect 44908 23248 44948 23288
rect 47596 29800 47636 29840
rect 47212 29716 47252 29756
rect 47212 28876 47252 28916
rect 47212 27784 47252 27824
rect 46636 26944 46676 26984
rect 46444 26776 46484 26816
rect 46636 26776 46676 26816
rect 46060 25852 46100 25892
rect 46060 25432 46100 25472
rect 45868 24424 45908 24464
rect 45196 24256 45236 24296
rect 45388 24256 45428 24296
rect 45196 23920 45236 23960
rect 45100 22996 45140 23036
rect 45964 23752 46004 23792
rect 46636 25600 46676 25640
rect 46444 25432 46484 25472
rect 46540 25264 46580 25304
rect 46444 25012 46484 25052
rect 47404 27616 47444 27656
rect 47308 27532 47348 27572
rect 47212 26776 47252 26816
rect 47884 32824 47924 32864
rect 48940 34336 48980 34376
rect 49228 34252 49268 34292
rect 49036 34168 49076 34208
rect 49036 33664 49076 33704
rect 48364 33412 48404 33452
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 48748 32992 48788 33032
rect 48652 32908 48692 32948
rect 47980 32152 48020 32192
rect 48364 32152 48404 32192
rect 49036 32908 49076 32948
rect 49228 33664 49268 33704
rect 49228 33412 49268 33452
rect 49516 34336 49556 34376
rect 48844 32572 48884 32612
rect 48940 32068 48980 32108
rect 48748 31984 48788 32024
rect 49324 32572 49364 32612
rect 49228 32320 49268 32360
rect 49132 32152 49172 32192
rect 48460 31900 48500 31940
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 49228 31816 49268 31856
rect 49036 31564 49076 31604
rect 49036 31312 49076 31352
rect 49228 31312 49268 31352
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 48364 29800 48404 29840
rect 49036 29800 49076 29840
rect 49420 32320 49460 32360
rect 50284 34252 50324 34292
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 50092 32152 50132 32192
rect 49996 32068 50036 32108
rect 49612 31900 49652 31940
rect 49516 31816 49556 31856
rect 49516 31144 49556 31184
rect 49324 30640 49364 30680
rect 49132 29632 49172 29672
rect 47788 28960 47828 29000
rect 48748 28876 48788 28916
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 48844 28120 48884 28160
rect 47692 27784 47732 27824
rect 47788 27700 47828 27740
rect 47692 27616 47732 27656
rect 47788 27532 47828 27572
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 47596 26860 47636 26900
rect 48268 26776 48308 26816
rect 47980 26608 48020 26648
rect 47116 26020 47156 26060
rect 47020 25936 47060 25976
rect 46924 25600 46964 25640
rect 46732 25348 46772 25388
rect 46828 24844 46868 24884
rect 47020 24844 47060 24884
rect 46636 24004 46676 24044
rect 46156 23920 46196 23960
rect 45292 23080 45332 23120
rect 45484 23080 45524 23120
rect 46060 23416 46100 23456
rect 46156 23332 46196 23372
rect 46636 23332 46676 23372
rect 46636 23164 46676 23204
rect 45580 22996 45620 23036
rect 44812 21568 44852 21608
rect 44140 20728 44180 20768
rect 45004 20896 45044 20936
rect 44908 20728 44948 20768
rect 45292 21736 45332 21776
rect 45484 22240 45524 22280
rect 45292 21568 45332 21608
rect 45388 21484 45428 21524
rect 45676 21736 45716 21776
rect 45388 21232 45428 21272
rect 45484 20728 45524 20768
rect 45868 21484 45908 21524
rect 44236 20056 44276 20096
rect 43852 19972 43892 20012
rect 44332 19972 44372 20012
rect 45004 20560 45044 20600
rect 46252 22240 46292 22280
rect 48076 26020 48116 26060
rect 47980 25600 48020 25640
rect 47596 23752 47636 23792
rect 46732 22240 46772 22280
rect 46060 20728 46100 20768
rect 46540 21316 46580 21356
rect 44908 20140 44948 20180
rect 44044 19888 44084 19928
rect 43852 18880 43892 18920
rect 43660 18712 43700 18752
rect 43756 16864 43796 16904
rect 44716 19888 44756 19928
rect 44524 19552 44564 19592
rect 44620 19048 44660 19088
rect 44332 18880 44372 18920
rect 44140 18712 44180 18752
rect 43948 18544 43988 18584
rect 44428 18628 44468 18668
rect 44620 18628 44660 18668
rect 43948 17788 43988 17828
rect 44044 17704 44084 17744
rect 44908 17536 44948 17576
rect 44332 17200 44372 17240
rect 43948 17032 43988 17072
rect 44716 17032 44756 17072
rect 44140 16864 44180 16904
rect 43372 16696 43412 16736
rect 43084 16612 43124 16652
rect 43084 16360 43124 16400
rect 43173 16276 43213 16316
rect 43372 15856 43412 15896
rect 42988 15520 43028 15560
rect 43180 15520 43220 15560
rect 42700 14680 42740 14720
rect 42700 14176 42740 14216
rect 42604 14092 42644 14132
rect 42988 14680 43028 14720
rect 43276 14680 43316 14720
rect 42892 14092 42932 14132
rect 43180 14092 43220 14132
rect 42700 13588 42740 13628
rect 42316 12916 42356 12956
rect 42028 12412 42068 12452
rect 41836 11656 41876 11696
rect 42796 13168 42836 13208
rect 43468 13840 43508 13880
rect 43276 13504 43316 13544
rect 43660 14008 43700 14048
rect 43852 13840 43892 13880
rect 43660 13252 43700 13292
rect 42508 12496 42548 12536
rect 42028 10480 42068 10520
rect 41644 10228 41684 10268
rect 41932 10228 41972 10268
rect 42988 12412 43028 12452
rect 42604 11992 42644 12032
rect 42604 11656 42644 11696
rect 42604 11152 42644 11192
rect 42316 10900 42356 10940
rect 42220 10228 42260 10268
rect 41836 10144 41876 10184
rect 41740 10060 41780 10100
rect 41356 9472 41396 9512
rect 43276 12916 43316 12956
rect 43564 12916 43604 12956
rect 44524 16696 44564 16736
rect 44140 16444 44180 16484
rect 44620 14008 44660 14048
rect 45676 20056 45716 20096
rect 45292 19972 45332 20012
rect 45292 19300 45332 19340
rect 45196 18628 45236 18668
rect 45100 16948 45140 16988
rect 45100 16360 45140 16400
rect 45004 15268 45044 15308
rect 45484 18544 45524 18584
rect 46060 18628 46100 18668
rect 46252 18376 46292 18416
rect 46828 18544 46868 18584
rect 46828 18292 46868 18332
rect 46828 18040 46868 18080
rect 46444 17788 46484 17828
rect 45580 17620 45620 17660
rect 45580 17452 45620 17492
rect 45484 17368 45524 17408
rect 45388 17032 45428 17072
rect 45292 16276 45332 16316
rect 45292 16108 45332 16148
rect 45484 16024 45524 16064
rect 45964 17704 46004 17744
rect 45772 17116 45812 17156
rect 45676 16948 45716 16988
rect 46252 17704 46292 17744
rect 46156 17116 46196 17156
rect 46060 16780 46100 16820
rect 46252 16276 46292 16316
rect 46060 16192 46100 16232
rect 45772 16024 45812 16064
rect 46060 15856 46100 15896
rect 45196 13756 45236 13796
rect 44332 13252 44372 13292
rect 44716 13252 44756 13292
rect 45484 13504 45524 13544
rect 45580 13252 45620 13292
rect 43276 11572 43316 11612
rect 42316 10144 42356 10184
rect 41548 9304 41588 9344
rect 41932 9304 41972 9344
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 41548 8716 41588 8756
rect 42316 9220 42356 9260
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 42700 9640 42740 9680
rect 42988 9724 43028 9764
rect 43084 9640 43124 9680
rect 43660 9640 43700 9680
rect 42508 8716 42548 8756
rect 42988 9556 43028 9596
rect 42892 9472 42932 9512
rect 42988 9304 43028 9344
rect 45388 12916 45428 12956
rect 44812 11992 44852 12032
rect 45292 11908 45332 11948
rect 43948 11068 43988 11108
rect 43852 10228 43892 10268
rect 44140 10900 44180 10940
rect 44332 10564 44372 10604
rect 44140 10228 44180 10268
rect 43852 9640 43892 9680
rect 44236 9808 44276 9848
rect 44044 9220 44084 9260
rect 44236 9388 44276 9428
rect 44140 8716 44180 8756
rect 42796 8632 42836 8672
rect 42412 8044 42452 8084
rect 44140 8128 44180 8168
rect 45676 13168 45716 13208
rect 46540 17704 46580 17744
rect 46444 15436 46484 15476
rect 46156 14680 46196 14720
rect 46540 14680 46580 14720
rect 48748 26608 48788 26648
rect 48268 25936 48308 25976
rect 48556 25936 48596 25976
rect 49132 25936 49172 25976
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 49420 29632 49460 29672
rect 50956 35932 50996 35972
rect 51052 35764 51092 35804
rect 50476 34336 50516 34376
rect 50476 33412 50516 33452
rect 50380 32656 50420 32696
rect 55948 37360 55988 37400
rect 55852 36772 55892 36812
rect 55948 36688 55988 36728
rect 56236 37192 56276 37232
rect 57580 37192 57620 37232
rect 57580 36772 57620 36812
rect 56428 36688 56468 36728
rect 56044 36520 56084 36560
rect 51436 35764 51476 35804
rect 51532 35260 51572 35300
rect 51244 34504 51284 34544
rect 51436 34336 51476 34376
rect 51628 33748 51668 33788
rect 52300 35764 52340 35804
rect 51820 35092 51860 35132
rect 52780 35260 52820 35300
rect 52108 35008 52148 35048
rect 54508 35260 54548 35300
rect 55660 35848 55700 35888
rect 56332 36436 56372 36476
rect 55852 35680 55892 35720
rect 55468 35512 55508 35552
rect 53356 35176 53396 35216
rect 53740 35092 53780 35132
rect 52204 34504 52244 34544
rect 52204 34336 52244 34376
rect 51724 33412 51764 33452
rect 50764 32992 50804 33032
rect 50572 32824 50612 32864
rect 50764 32740 50804 32780
rect 50476 32320 50516 32360
rect 49996 31732 50036 31772
rect 49708 31312 49748 31352
rect 50668 32572 50708 32612
rect 50476 31732 50516 31772
rect 50092 31312 50132 31352
rect 50380 31312 50420 31352
rect 50188 31228 50228 31268
rect 49708 31144 49748 31184
rect 49900 31144 49940 31184
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 49516 29296 49556 29336
rect 49804 30640 49844 30680
rect 51052 32572 51092 32612
rect 51244 32740 51284 32780
rect 50956 32320 50996 32360
rect 50860 31732 50900 31772
rect 50860 31312 50900 31352
rect 50476 31144 50516 31184
rect 50764 31144 50804 31184
rect 52492 33496 52532 33536
rect 53452 33496 53492 33536
rect 52204 32740 52244 32780
rect 51820 32152 51860 32192
rect 53740 33328 53780 33368
rect 53644 32992 53684 33032
rect 50572 30808 50612 30848
rect 50476 30640 50516 30680
rect 51532 30808 51572 30848
rect 50380 30388 50420 30428
rect 50188 30304 50228 30344
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 49804 29296 49844 29336
rect 50092 29296 50132 29336
rect 50380 29884 50420 29924
rect 50284 29464 50324 29504
rect 50668 30220 50708 30260
rect 51244 30640 51284 30680
rect 50572 29632 50612 29672
rect 49708 29128 49748 29168
rect 50380 29044 50420 29084
rect 49516 28960 49556 29000
rect 50284 28960 50324 29000
rect 49612 28792 49652 28832
rect 49996 28288 50036 28328
rect 50092 28120 50132 28160
rect 50188 28036 50228 28076
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 49420 27532 49460 27572
rect 49612 27196 49652 27236
rect 50092 27196 50132 27236
rect 50956 30220 50996 30260
rect 51532 30136 51572 30176
rect 51436 30052 51476 30092
rect 51052 29968 51092 30008
rect 51052 29716 51092 29756
rect 51340 29968 51380 30008
rect 50956 29464 50996 29504
rect 51244 29464 51284 29504
rect 51052 29212 51092 29252
rect 50860 29128 50900 29168
rect 51436 29716 51476 29756
rect 50572 28792 50612 28832
rect 50956 28792 50996 28832
rect 50476 28708 50516 28748
rect 50956 28624 50996 28664
rect 50572 28120 50612 28160
rect 50380 28036 50420 28076
rect 50380 27868 50420 27908
rect 50284 26944 50324 26984
rect 49612 26776 49652 26816
rect 50284 26776 50324 26816
rect 50668 27868 50708 27908
rect 49516 26692 49556 26732
rect 49420 26272 49460 26312
rect 49324 25516 49364 25556
rect 48172 25012 48212 25052
rect 49420 25012 49460 25052
rect 48268 23752 48308 23792
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 48748 24004 48788 24044
rect 48076 23668 48116 23708
rect 49324 23752 49364 23792
rect 49036 23248 49076 23288
rect 48748 23080 48788 23120
rect 48940 23080 48980 23120
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 47980 22492 48020 22532
rect 47692 21316 47732 21356
rect 48556 22240 48596 22280
rect 50188 26692 50228 26732
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 50188 26440 50228 26480
rect 50188 26272 50228 26312
rect 49612 26104 49652 26144
rect 49996 26104 50036 26144
rect 50572 26692 50612 26732
rect 50764 26608 50804 26648
rect 49612 25516 49652 25556
rect 49996 25264 50036 25304
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 50668 26272 50708 26312
rect 50668 25264 50708 25304
rect 50380 24928 50420 24968
rect 50572 24928 50612 24968
rect 49708 24592 49748 24632
rect 50380 24592 50420 24632
rect 51052 28204 51092 28244
rect 51340 29044 51380 29084
rect 51724 29884 51764 29924
rect 51436 28624 51476 28664
rect 51244 28120 51284 28160
rect 51244 27868 51284 27908
rect 51244 26944 51284 26984
rect 52396 31312 52436 31352
rect 52492 29800 52532 29840
rect 51820 29128 51860 29168
rect 52492 29044 52532 29084
rect 51724 28960 51764 29000
rect 51724 28372 51764 28412
rect 51820 28288 51860 28328
rect 51724 27868 51764 27908
rect 51724 27700 51764 27740
rect 51916 27616 51956 27656
rect 51820 27364 51860 27404
rect 51628 26944 51668 26984
rect 51532 26776 51572 26816
rect 51436 26104 51476 26144
rect 50668 24844 50708 24884
rect 49612 24508 49652 24548
rect 49996 24508 50036 24548
rect 50476 24424 50516 24464
rect 50092 24004 50132 24044
rect 50188 23836 50228 23876
rect 50092 23584 50132 23624
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 49996 23248 50036 23288
rect 50100 23248 50132 23288
rect 50132 23248 50140 23288
rect 49900 23080 49940 23120
rect 49804 23035 49844 23036
rect 49804 22996 49844 23035
rect 49036 21568 49076 21608
rect 50380 23836 50420 23876
rect 51148 24844 51188 24884
rect 50860 24508 50900 24548
rect 50764 24004 50804 24044
rect 50572 23920 50612 23960
rect 50860 23920 50900 23960
rect 50476 23164 50516 23204
rect 50284 23080 50324 23120
rect 50956 23836 50996 23876
rect 50764 23668 50804 23708
rect 50668 23332 50708 23372
rect 50860 23332 50900 23372
rect 51724 26104 51764 26144
rect 52108 28288 52148 28328
rect 52108 27700 52148 27740
rect 52396 28120 52436 28160
rect 52300 27952 52340 27992
rect 52204 27616 52244 27656
rect 52108 27364 52148 27404
rect 52588 28288 52628 28328
rect 52396 27532 52436 27572
rect 52300 26776 52340 26816
rect 52300 26608 52340 26648
rect 52108 26272 52148 26312
rect 52300 26272 52340 26312
rect 52588 26272 52628 26312
rect 51820 25852 51860 25892
rect 51340 24592 51380 24632
rect 51244 23920 51284 23960
rect 51148 23752 51188 23792
rect 51436 24508 51476 24548
rect 51724 24844 51764 24884
rect 51916 24844 51956 24884
rect 51820 24508 51860 24548
rect 51532 24424 51572 24464
rect 51820 24172 51860 24212
rect 51532 23752 51572 23792
rect 51436 23584 51476 23624
rect 50764 23164 50804 23204
rect 50668 23080 50708 23120
rect 50380 22492 50420 22532
rect 50092 22240 50132 22280
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 49420 21484 49460 21524
rect 49612 21568 49652 21608
rect 49516 21400 49556 21440
rect 48844 21316 48884 21356
rect 48364 21232 48404 21272
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 50380 21820 50420 21860
rect 50380 21652 50420 21692
rect 50284 20980 50324 21020
rect 50764 22912 50804 22952
rect 50572 21820 50612 21860
rect 51340 23164 51380 23204
rect 51436 23080 51476 23120
rect 51244 22996 51284 23036
rect 51148 22492 51188 22532
rect 50668 21484 50708 21524
rect 51052 21652 51092 21692
rect 50956 21568 50996 21608
rect 50860 21484 50900 21524
rect 50764 21064 50804 21104
rect 52492 26020 52532 26060
rect 53548 32824 53588 32864
rect 54028 33832 54068 33872
rect 53932 33748 53972 33788
rect 54028 33664 54068 33704
rect 54028 33496 54068 33536
rect 54028 33328 54068 33368
rect 53548 32572 53588 32612
rect 53932 32152 53972 32192
rect 53548 31816 53588 31856
rect 52876 30472 52916 30512
rect 53644 29212 53684 29252
rect 52972 28456 53012 28496
rect 52108 25264 52148 25304
rect 52108 24592 52148 24632
rect 52108 23752 52148 23792
rect 51820 23416 51860 23456
rect 51820 22576 51860 22616
rect 51532 21232 51572 21272
rect 52012 23164 52052 23204
rect 52588 25180 52628 25220
rect 52876 24592 52916 24632
rect 53356 27196 53396 27236
rect 54412 33832 54452 33872
rect 54316 33328 54356 33368
rect 54796 35092 54836 35132
rect 54508 33328 54548 33368
rect 54220 32152 54260 32192
rect 54124 31312 54164 31352
rect 54028 30388 54068 30428
rect 54508 32824 54548 32864
rect 54700 33664 54740 33704
rect 54988 34840 55028 34880
rect 54892 33748 54932 33788
rect 54412 32740 54452 32780
rect 54604 32656 54644 32696
rect 54796 32824 54836 32864
rect 55276 33664 55316 33704
rect 56140 35512 56180 35552
rect 56044 35176 56084 35216
rect 55852 35008 55892 35048
rect 55180 33412 55220 33452
rect 56140 34840 56180 34880
rect 54508 32152 54548 32192
rect 54412 32068 54452 32108
rect 54412 31900 54452 31940
rect 54700 32320 54740 32360
rect 54892 32236 54932 32276
rect 54988 32152 55028 32192
rect 54988 31900 55028 31940
rect 54796 30808 54836 30848
rect 54796 30640 54836 30680
rect 54604 30472 54644 30512
rect 54700 30220 54740 30260
rect 54988 30220 55028 30260
rect 55372 32236 55412 32276
rect 55276 32152 55316 32192
rect 55660 32152 55700 32192
rect 56044 34336 56084 34376
rect 57100 36436 57140 36476
rect 56620 35848 56660 35888
rect 56332 34588 56372 34628
rect 56236 34252 56276 34292
rect 56332 32236 56372 32276
rect 55948 31732 55988 31772
rect 55276 31144 55316 31184
rect 55564 31144 55604 31184
rect 55180 30388 55220 30428
rect 55084 30136 55124 30176
rect 55468 30304 55508 30344
rect 55756 31144 55796 31184
rect 55948 30976 55988 31016
rect 57100 35932 57140 35972
rect 56908 35512 56948 35552
rect 57388 36688 57428 36728
rect 57292 36520 57332 36560
rect 57196 35176 57236 35216
rect 58540 38116 58580 38156
rect 59308 38116 59348 38156
rect 58924 37948 58964 37988
rect 59116 37948 59156 37988
rect 58636 37276 58676 37316
rect 58924 36940 58964 36980
rect 58828 36856 58868 36896
rect 58444 36772 58484 36812
rect 58828 36688 58868 36728
rect 59500 37360 59540 37400
rect 59404 37276 59444 37316
rect 59308 37192 59348 37232
rect 59020 36184 59060 36224
rect 58636 36016 58676 36056
rect 58636 35848 58676 35888
rect 58252 35680 58292 35720
rect 57772 35176 57812 35216
rect 57484 35092 57524 35132
rect 57964 35092 58004 35132
rect 57580 34840 57620 34880
rect 58060 34504 58100 34544
rect 58060 34336 58100 34376
rect 57772 34000 57812 34040
rect 57580 32824 57620 32864
rect 58252 34336 58292 34376
rect 59116 35848 59156 35888
rect 59596 37276 59636 37316
rect 59500 36184 59540 36224
rect 59596 36016 59636 36056
rect 59500 35932 59540 35972
rect 59308 35848 59348 35888
rect 59212 35764 59252 35804
rect 58924 35680 58964 35720
rect 58828 35092 58868 35132
rect 58732 34588 58772 34628
rect 58636 34168 58676 34208
rect 58348 34000 58388 34040
rect 58444 33916 58484 33956
rect 58540 33748 58580 33788
rect 58348 33412 58388 33452
rect 58156 33076 58196 33116
rect 58252 32824 58292 32864
rect 59500 35764 59540 35804
rect 59596 35680 59636 35720
rect 59404 34588 59444 34628
rect 58924 33412 58964 33452
rect 58924 33244 58964 33284
rect 58636 32992 58676 33032
rect 58156 32740 58196 32780
rect 57676 32656 57716 32696
rect 56812 32152 56852 32192
rect 57196 31564 57236 31604
rect 56140 31144 56180 31184
rect 56140 30976 56180 31016
rect 55852 30640 55892 30680
rect 55564 29968 55604 30008
rect 54796 29884 54836 29924
rect 54700 29800 54740 29840
rect 55084 29800 55124 29840
rect 54028 29212 54068 29252
rect 54316 29212 54356 29252
rect 53932 28960 53972 29000
rect 53260 26860 53300 26900
rect 53260 26692 53300 26732
rect 52684 24004 52724 24044
rect 52588 23752 52628 23792
rect 52780 23248 52820 23288
rect 52492 23080 52532 23120
rect 52684 23080 52724 23120
rect 52204 22996 52244 23036
rect 52300 22912 52340 22952
rect 52396 22744 52436 22784
rect 52684 22828 52724 22868
rect 52108 22156 52148 22196
rect 51916 20980 51956 21020
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 51628 20476 51668 20516
rect 47212 20140 47252 20180
rect 47596 20140 47636 20180
rect 48940 20140 48980 20180
rect 50860 20140 50900 20180
rect 51532 20140 51572 20180
rect 47500 19384 47540 19424
rect 47500 18460 47540 18500
rect 47020 18376 47060 18416
rect 47500 17452 47540 17492
rect 47692 18544 47732 18584
rect 47788 18460 47828 18500
rect 47596 17368 47636 17408
rect 47500 17200 47540 17240
rect 47020 17032 47060 17072
rect 47308 16864 47348 16904
rect 47116 16780 47156 16820
rect 47212 16192 47252 16232
rect 47404 16276 47444 16316
rect 47308 15856 47348 15896
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 48940 19636 48980 19676
rect 47884 16528 47924 16568
rect 49036 19216 49076 19256
rect 48652 18712 48692 18752
rect 49036 18880 49076 18920
rect 49036 18712 49076 18752
rect 49228 18880 49268 18920
rect 49612 19636 49652 19676
rect 51532 19552 51572 19592
rect 49132 18628 49172 18668
rect 49324 18628 49364 18668
rect 48844 18544 48884 18584
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 49612 18880 49652 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 49804 18460 49844 18500
rect 50572 18460 50612 18500
rect 49516 18040 49556 18080
rect 48940 17788 48980 17828
rect 49516 17788 49556 17828
rect 48748 17704 48788 17744
rect 48364 17032 48404 17072
rect 49804 17788 49844 17828
rect 49612 17704 49652 17744
rect 50092 17704 50132 17744
rect 50476 18292 50516 18332
rect 50380 17704 50420 17744
rect 49420 17284 49460 17324
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 49612 17200 49652 17240
rect 49228 17116 49268 17156
rect 48652 16948 48692 16988
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 49612 16528 49652 16568
rect 48268 16276 48308 16316
rect 48652 16276 48692 16316
rect 49420 16276 49460 16316
rect 47500 16192 47540 16232
rect 47500 15856 47540 15896
rect 48268 15856 48308 15896
rect 47308 15016 47348 15056
rect 46924 14260 46964 14300
rect 45964 14176 46004 14216
rect 45868 13336 45908 13376
rect 45772 13000 45812 13040
rect 46156 14008 46196 14048
rect 46348 14008 46388 14048
rect 46156 13168 46196 13208
rect 46540 13252 46580 13292
rect 46444 13084 46484 13124
rect 45868 12916 45908 12956
rect 47020 14176 47060 14216
rect 47404 14176 47444 14216
rect 47884 15520 47924 15560
rect 47788 14008 47828 14048
rect 48172 15520 48212 15560
rect 48076 15016 48116 15056
rect 48076 14680 48116 14720
rect 47596 13420 47636 13460
rect 47404 13252 47444 13292
rect 45868 11656 45908 11696
rect 47500 12748 47540 12788
rect 46828 11152 46868 11192
rect 46732 11068 46772 11108
rect 46252 10900 46292 10940
rect 44812 10144 44852 10184
rect 45484 9472 45524 9512
rect 44524 9220 44564 9260
rect 45388 8632 45428 8672
rect 44812 8548 44852 8588
rect 44428 8044 44468 8084
rect 44908 8128 44948 8168
rect 45580 9304 45620 9344
rect 45388 7708 45428 7748
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 46924 10900 46964 10940
rect 46828 10648 46868 10688
rect 46348 10144 46388 10184
rect 47116 10480 47156 10520
rect 46348 9220 46388 9260
rect 46732 9472 46772 9512
rect 46732 9220 46772 9260
rect 46636 8632 46676 8672
rect 46252 8128 46292 8168
rect 45676 7960 45716 8000
rect 46540 7960 46580 8000
rect 47116 9472 47156 9512
rect 47020 9388 47060 9428
rect 46924 8716 46964 8756
rect 46828 8548 46868 8588
rect 48076 13168 48116 13208
rect 49996 17032 50036 17072
rect 50476 17536 50516 17576
rect 50380 17200 50420 17240
rect 49900 16864 49940 16904
rect 50188 16864 50228 16904
rect 50476 16780 50516 16820
rect 49900 16192 49940 16232
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 50380 15436 50420 15476
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 48844 13420 48884 13460
rect 47980 13084 48020 13124
rect 48076 13000 48116 13040
rect 47788 12748 47828 12788
rect 47692 12664 47732 12704
rect 48172 12664 48212 12704
rect 48268 12580 48308 12620
rect 48652 12496 48692 12536
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 49228 13252 49268 13292
rect 49324 13084 49364 13124
rect 49036 12496 49076 12536
rect 47884 11656 47924 11696
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 48268 11908 48308 11948
rect 48556 11824 48596 11864
rect 48460 11656 48500 11696
rect 48364 11572 48404 11612
rect 49708 13168 49748 13208
rect 49516 12664 49556 12704
rect 49132 12412 49172 12452
rect 49228 11824 49268 11864
rect 49036 11656 49076 11696
rect 49228 11656 49268 11696
rect 49516 12496 49556 12536
rect 49420 12412 49460 12452
rect 49516 11572 49556 11612
rect 48940 10984 48980 11024
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 49708 12664 49748 12704
rect 50092 11656 50132 11696
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 50380 15016 50420 15056
rect 51532 18460 51572 18500
rect 51340 18292 51380 18332
rect 51244 17956 51284 17996
rect 51148 17620 51188 17660
rect 50668 17284 50708 17324
rect 50764 17032 50804 17072
rect 50668 16864 50708 16904
rect 50572 16360 50612 16400
rect 50572 15520 50612 15560
rect 50572 14092 50612 14132
rect 50476 13588 50516 13628
rect 50476 13168 50516 13208
rect 50284 11656 50324 11696
rect 50188 11152 50228 11192
rect 50188 10984 50228 11024
rect 49420 10648 49460 10688
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 49228 10480 49268 10520
rect 47980 9388 48020 9428
rect 46828 8128 46868 8168
rect 47020 8128 47060 8168
rect 47500 8128 47540 8168
rect 47692 8128 47732 8168
rect 46732 7960 46772 8000
rect 46636 7120 46676 7160
rect 47308 7960 47348 8000
rect 47116 7120 47156 7160
rect 46828 6532 46868 6572
rect 45580 6448 45620 6488
rect 45484 6364 45524 6404
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 45868 5020 45908 5060
rect 47500 7708 47540 7748
rect 47500 7372 47540 7412
rect 47404 6448 47444 6488
rect 48940 10144 48980 10184
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 48460 8716 48500 8756
rect 48076 8632 48116 8672
rect 48268 8128 48308 8168
rect 47788 7372 47828 7412
rect 47980 7372 48020 7412
rect 47884 6448 47924 6488
rect 47308 6364 47348 6404
rect 47404 5776 47444 5816
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 47308 5608 47348 5648
rect 47308 5020 47348 5060
rect 47596 5776 47636 5816
rect 47500 5440 47540 5480
rect 47404 4768 47444 4808
rect 48268 7708 48308 7748
rect 48556 8548 48596 8588
rect 48556 7960 48596 8000
rect 49036 8548 49076 8588
rect 48844 8128 48884 8168
rect 49036 8212 49076 8252
rect 48940 7960 48980 8000
rect 48460 7708 48500 7748
rect 48748 7708 48788 7748
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 48364 7372 48404 7412
rect 49036 7372 49076 7412
rect 48748 7204 48788 7244
rect 48364 7120 48404 7160
rect 49516 10396 49556 10436
rect 49420 7960 49460 8000
rect 49804 10144 49844 10184
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 51052 17032 51092 17072
rect 51244 16780 51284 16820
rect 51244 16192 51284 16232
rect 51052 15520 51092 15560
rect 50764 13672 50804 13712
rect 51436 17200 51476 17240
rect 51436 16276 51476 16316
rect 52012 19048 52052 19088
rect 52300 21988 52340 22028
rect 52300 21568 52340 21608
rect 52684 22240 52724 22280
rect 52588 22156 52628 22196
rect 52588 21568 52628 21608
rect 52972 22912 53012 22952
rect 53548 24592 53588 24632
rect 54220 29128 54260 29168
rect 54700 28792 54740 28832
rect 54508 27952 54548 27992
rect 54796 28456 54836 28496
rect 55180 29128 55220 29168
rect 55372 29128 55412 29168
rect 55084 28960 55124 29000
rect 55276 28540 55316 28580
rect 55660 29632 55700 29672
rect 56620 31312 56660 31352
rect 56236 30304 56276 30344
rect 56044 29968 56084 30008
rect 55852 29884 55892 29924
rect 56044 29632 56084 29672
rect 55948 29212 55988 29252
rect 55660 28876 55700 28916
rect 55564 28792 55604 28832
rect 55468 28540 55508 28580
rect 55180 27700 55220 27740
rect 54220 27028 54260 27068
rect 55660 28288 55700 28328
rect 55852 29128 55892 29168
rect 55948 28708 55988 28748
rect 55756 28120 55796 28160
rect 55372 27532 55412 27572
rect 55948 27616 55988 27656
rect 55660 27028 55700 27068
rect 55468 26608 55508 26648
rect 55468 26104 55508 26144
rect 54892 25936 54932 25976
rect 54700 25852 54740 25892
rect 54700 25348 54740 25388
rect 55276 25264 55316 25304
rect 55468 25264 55508 25304
rect 54700 25096 54740 25136
rect 54028 24256 54068 24296
rect 55468 25096 55508 25136
rect 55180 24676 55220 24716
rect 54700 23752 54740 23792
rect 54124 23584 54164 23624
rect 54316 23248 54356 23288
rect 53644 23164 53684 23204
rect 55564 24004 55604 24044
rect 56236 29800 56276 29840
rect 56332 29212 56372 29252
rect 56428 28624 56468 28664
rect 56428 28288 56468 28328
rect 57100 28120 57140 28160
rect 56812 27700 56852 27740
rect 56332 27616 56372 27656
rect 56044 26608 56084 26648
rect 55756 26104 55796 26144
rect 56236 25936 56276 25976
rect 57004 26272 57044 26312
rect 56236 25264 56276 25304
rect 55756 25096 55796 25136
rect 56140 24592 56180 24632
rect 57100 25096 57140 25136
rect 56332 24508 56372 24548
rect 57388 31312 57428 31352
rect 57580 31312 57620 31352
rect 58540 32740 58580 32780
rect 58252 31984 58292 32024
rect 59212 33244 59252 33284
rect 59020 33076 59060 33116
rect 59116 32152 59156 32192
rect 59308 32152 59348 32192
rect 60268 37276 60308 37316
rect 62572 37948 62612 37988
rect 62380 37360 62420 37400
rect 60364 36856 60404 36896
rect 59788 34504 59828 34544
rect 59596 34168 59636 34208
rect 59500 34084 59540 34124
rect 58348 31732 58388 31772
rect 59308 31984 59348 32024
rect 59308 31732 59348 31772
rect 59116 31312 59156 31352
rect 57964 30808 58004 30848
rect 57676 30724 57716 30764
rect 59020 30892 59060 30932
rect 58636 30640 58676 30680
rect 58540 30304 58580 30344
rect 58828 29884 58868 29924
rect 58732 28624 58772 28664
rect 58540 28036 58580 28076
rect 58444 27784 58484 27824
rect 57964 27280 58004 27320
rect 57676 26944 57716 26984
rect 57484 26776 57524 26816
rect 57292 26104 57332 26144
rect 57676 26020 57716 26060
rect 57388 25936 57428 25976
rect 57196 24424 57236 24464
rect 55756 24004 55796 24044
rect 57676 24340 57716 24380
rect 55852 23920 55892 23960
rect 57292 23920 57332 23960
rect 54796 23164 54836 23204
rect 54604 23080 54644 23120
rect 55276 23164 55316 23204
rect 53545 22828 53585 22868
rect 52876 22156 52916 22196
rect 52300 20560 52340 20600
rect 52684 20980 52724 21020
rect 52588 20476 52628 20516
rect 51628 17200 51668 17240
rect 51724 17116 51764 17156
rect 51628 17032 51668 17072
rect 51916 17704 51956 17744
rect 51628 16528 51668 16568
rect 51532 16192 51572 16232
rect 51724 16360 51764 16400
rect 51916 16696 51956 16736
rect 51820 16192 51860 16232
rect 51340 15856 51380 15896
rect 51244 15352 51284 15392
rect 51244 14176 51284 14216
rect 51820 15856 51860 15896
rect 51724 14260 51764 14300
rect 51436 13672 51476 13712
rect 50956 13588 50996 13628
rect 50860 13252 50900 13292
rect 51628 13420 51668 13460
rect 51244 12916 51284 12956
rect 51628 12580 51668 12620
rect 52300 17452 52340 17492
rect 52300 17116 52340 17156
rect 52492 17368 52532 17408
rect 52396 17032 52436 17072
rect 52684 17368 52724 17408
rect 52588 17284 52628 17324
rect 52780 17200 52820 17240
rect 52588 17116 52628 17156
rect 54055 22996 54095 23036
rect 53945 22744 53985 22784
rect 54455 22912 54495 22952
rect 54855 22744 54895 22784
rect 56044 23332 56084 23372
rect 56620 23416 56660 23456
rect 56428 23248 56468 23288
rect 56812 23416 56852 23456
rect 56908 23164 56948 23204
rect 57292 23500 57332 23540
rect 57196 23164 57236 23204
rect 57580 23500 57620 23540
rect 57676 23416 57716 23456
rect 58156 27028 58196 27068
rect 58060 25096 58100 25136
rect 58060 24676 58100 24716
rect 58252 26944 58292 26984
rect 58444 27028 58484 27068
rect 58828 26776 58868 26816
rect 58348 25936 58388 25976
rect 58540 26104 58580 26144
rect 59692 33664 59732 33704
rect 59788 32236 59828 32276
rect 59404 31564 59444 31604
rect 60364 34168 60404 34208
rect 59980 34084 60020 34124
rect 60268 33748 60308 33788
rect 59980 33496 60020 33536
rect 59884 31900 59924 31940
rect 59788 31732 59828 31772
rect 59788 31312 59828 31352
rect 59884 31144 59924 31184
rect 59692 31060 59732 31100
rect 61132 37276 61172 37316
rect 62284 37276 62324 37316
rect 61804 36940 61844 36980
rect 61132 36856 61172 36896
rect 60556 36688 60596 36728
rect 61708 36688 61748 36728
rect 62380 36856 62420 36896
rect 61516 35680 61556 35720
rect 62380 36688 62420 36728
rect 61900 35932 61940 35972
rect 61612 35008 61652 35048
rect 61516 34336 61556 34376
rect 61900 35008 61940 35048
rect 61804 34924 61844 34964
rect 61996 34924 62036 34964
rect 61708 34672 61748 34712
rect 61612 33916 61652 33956
rect 60460 33664 60500 33704
rect 61708 33748 61748 33788
rect 62284 34924 62324 34964
rect 61996 34504 62036 34544
rect 61996 34336 62036 34376
rect 62188 34336 62228 34376
rect 62188 34084 62228 34124
rect 61996 34000 62036 34040
rect 61900 33664 61940 33704
rect 62380 34000 62420 34040
rect 62380 33664 62420 33704
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 63340 36772 63380 36812
rect 63916 36772 63956 36812
rect 67468 38200 67508 38240
rect 67084 38116 67124 38156
rect 66316 37948 66356 37988
rect 64972 37360 65012 37400
rect 65644 37360 65684 37400
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 62956 36604 62996 36644
rect 63148 36604 63188 36644
rect 62860 35176 62900 35216
rect 64012 36688 64052 36728
rect 63244 36436 63284 36476
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 62764 34924 62804 34964
rect 63148 34588 63188 34628
rect 62860 34336 62900 34376
rect 62764 34252 62804 34292
rect 63148 34252 63188 34292
rect 62668 33832 62708 33872
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 64012 34588 64052 34628
rect 60940 33076 60980 33116
rect 60940 32404 60980 32444
rect 60076 31480 60116 31520
rect 61324 32740 61364 32780
rect 60748 31900 60788 31940
rect 60652 31396 60692 31436
rect 60364 31228 60404 31268
rect 60556 31144 60596 31184
rect 60268 31060 60308 31100
rect 59596 30808 59636 30848
rect 60076 30808 60116 30848
rect 59596 30556 59636 30596
rect 59404 29464 59444 29504
rect 59116 29212 59156 29252
rect 59692 29884 59732 29924
rect 59980 30640 60020 30680
rect 59980 30052 60020 30092
rect 60268 30556 60308 30596
rect 60268 30388 60308 30428
rect 59020 28540 59060 28580
rect 59884 29296 59924 29336
rect 60172 29464 60212 29504
rect 59404 28540 59444 28580
rect 59308 28120 59348 28160
rect 60364 29968 60404 30008
rect 60364 29128 60404 29168
rect 60556 29044 60596 29084
rect 59884 28288 59924 28328
rect 59212 27784 59252 27824
rect 59308 27616 59348 27656
rect 59116 26860 59156 26900
rect 59692 27784 59732 27824
rect 59884 27784 59924 27824
rect 59788 27532 59828 27572
rect 59500 27364 59540 27404
rect 59116 26608 59156 26648
rect 58924 26440 58964 26480
rect 59020 26272 59060 26312
rect 59308 26356 59348 26396
rect 58924 25768 58964 25808
rect 58732 25600 58772 25640
rect 58636 25264 58676 25304
rect 58444 25096 58484 25136
rect 58636 24592 58676 24632
rect 59212 25180 59252 25220
rect 59020 24592 59060 24632
rect 59788 27196 59828 27236
rect 59980 27364 60020 27404
rect 59884 27028 59924 27068
rect 60364 28288 60404 28328
rect 60844 31564 60884 31604
rect 61036 31144 61076 31184
rect 61036 30640 61076 30680
rect 60940 30220 60980 30260
rect 60748 29968 60788 30008
rect 60844 29128 60884 29168
rect 61132 30388 61172 30428
rect 61228 30052 61268 30092
rect 61996 33328 62036 33368
rect 61900 32824 61940 32864
rect 61612 32152 61652 32192
rect 61804 32152 61844 32192
rect 61420 30220 61460 30260
rect 61996 32572 62036 32612
rect 61996 31480 62036 31520
rect 61900 31312 61940 31352
rect 61132 29044 61172 29084
rect 61036 28792 61076 28832
rect 60652 28456 60692 28496
rect 60268 27532 60308 27572
rect 59980 26860 60020 26900
rect 59500 26608 59540 26648
rect 59692 26608 59732 26648
rect 59692 26440 59732 26480
rect 59500 26104 59540 26144
rect 59404 25936 59444 25976
rect 59884 26104 59924 26144
rect 59500 25180 59540 25220
rect 59692 25180 59732 25220
rect 59308 24760 59348 24800
rect 58060 23752 58100 23792
rect 58348 23752 58388 23792
rect 57964 23500 58004 23540
rect 58060 23416 58100 23456
rect 59596 24760 59636 24800
rect 59500 24676 59540 24716
rect 59884 24928 59924 24968
rect 59788 24676 59828 24716
rect 59692 24592 59732 24632
rect 59884 24592 59924 24632
rect 60076 26440 60116 26480
rect 60460 27448 60500 27488
rect 60364 27112 60404 27152
rect 60268 26272 60308 26312
rect 60076 26104 60116 26144
rect 60652 28288 60692 28328
rect 60940 27868 60980 27908
rect 60844 27616 60884 27656
rect 60940 27280 60980 27320
rect 60748 27196 60788 27236
rect 60844 26860 60884 26900
rect 60556 26692 60596 26732
rect 60460 26272 60500 26312
rect 60460 26104 60500 26144
rect 60364 25096 60404 25136
rect 60460 25012 60500 25052
rect 60268 24928 60308 24968
rect 60172 24676 60212 24716
rect 60364 24760 60404 24800
rect 60460 24592 60500 24632
rect 59980 24340 60020 24380
rect 60364 24340 60404 24380
rect 60652 26188 60692 26228
rect 61132 27616 61172 27656
rect 61708 28288 61748 28328
rect 61900 27784 61940 27824
rect 61324 27448 61364 27488
rect 61228 27280 61268 27320
rect 61996 27028 62036 27068
rect 61324 26524 61364 26564
rect 61228 26272 61268 26312
rect 60748 25852 60788 25892
rect 60652 25096 60692 25136
rect 60844 25768 60884 25808
rect 61036 26020 61076 26060
rect 61228 26020 61268 26060
rect 61132 25936 61172 25976
rect 60940 25096 60980 25136
rect 60748 24676 60788 24716
rect 58444 23668 58484 23708
rect 58855 22828 58895 22868
rect 61132 24592 61172 24632
rect 61612 26188 61652 26228
rect 61516 25264 61556 25304
rect 61708 24928 61748 24968
rect 62476 32824 62516 32864
rect 62284 31816 62324 31856
rect 63244 33664 63284 33704
rect 63148 33580 63188 33620
rect 63052 33496 63092 33536
rect 62572 32572 62612 32612
rect 62572 32236 62612 32276
rect 62764 32068 62804 32108
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 63244 32908 63284 32948
rect 62956 32656 62996 32696
rect 62956 32236 62996 32276
rect 63148 32824 63188 32864
rect 65356 36688 65396 36728
rect 64396 36604 64436 36644
rect 64492 36016 64532 36056
rect 64396 35848 64436 35888
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 63340 32572 63380 32612
rect 63244 32320 63284 32360
rect 63436 32236 63476 32276
rect 63244 32068 63284 32108
rect 63916 32740 63956 32780
rect 64108 32656 64148 32696
rect 64012 32320 64052 32360
rect 64300 32236 64340 32276
rect 64588 32572 64628 32612
rect 64492 32152 64532 32192
rect 63148 31816 63188 31856
rect 63052 31648 63092 31688
rect 62572 31228 62612 31268
rect 63148 31312 63188 31352
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 63051 31228 63091 31268
rect 62476 30724 62516 30764
rect 62284 27028 62324 27068
rect 62284 26860 62324 26900
rect 62284 24424 62324 24464
rect 62188 24088 62228 24128
rect 62860 30388 62900 30428
rect 63052 30220 63092 30260
rect 62956 30052 62996 30092
rect 63244 31144 63284 31184
rect 63436 30220 63476 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 63340 30136 63380 30176
rect 62956 28960 62996 29000
rect 64108 31816 64148 31856
rect 64012 29884 64052 29924
rect 63628 29800 63668 29840
rect 63820 29800 63860 29840
rect 63148 29716 63188 29756
rect 63340 29632 63380 29672
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 65260 32152 65300 32192
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 63532 29128 63572 29168
rect 63436 29044 63476 29084
rect 63148 28288 63188 28328
rect 62860 27196 62900 27236
rect 63916 29128 63956 29168
rect 64012 29044 64052 29084
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 63724 28456 63764 28496
rect 63532 27952 63572 27992
rect 63436 27532 63476 27572
rect 64012 28204 64052 28244
rect 64012 27784 64052 27824
rect 63724 27364 63764 27404
rect 63916 27616 63956 27656
rect 64204 29128 64244 29168
rect 63244 26776 63284 26816
rect 62860 26524 62900 26564
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 64684 30640 64724 30680
rect 64588 29716 64628 29756
rect 67468 37948 67508 37988
rect 67660 37948 67700 37988
rect 67564 37360 67604 37400
rect 67276 36856 67316 36896
rect 67756 36856 67796 36896
rect 66124 36604 66164 36644
rect 65644 36016 65684 36056
rect 66604 36100 66644 36140
rect 66508 35848 66548 35888
rect 65644 35680 65684 35720
rect 67468 36688 67508 36728
rect 67276 36100 67316 36140
rect 67180 35848 67220 35888
rect 67372 35848 67412 35888
rect 66028 35512 66068 35552
rect 66700 35512 66740 35552
rect 67084 35512 67124 35552
rect 65644 35008 65684 35048
rect 65452 33748 65492 33788
rect 65548 33664 65588 33704
rect 65452 31900 65492 31940
rect 65836 34840 65876 34880
rect 65836 34672 65876 34712
rect 65740 34168 65780 34208
rect 65644 32824 65684 32864
rect 65644 32572 65684 32612
rect 66316 34336 66356 34376
rect 66700 34924 66740 34964
rect 66892 34672 66932 34712
rect 66124 34084 66164 34124
rect 65932 33832 65972 33872
rect 65836 33328 65876 33368
rect 66028 33328 66068 33368
rect 65932 32824 65972 32864
rect 66796 34168 66836 34208
rect 66604 33664 66644 33704
rect 66508 33496 66548 33536
rect 66220 32656 66260 32696
rect 65836 32152 65876 32192
rect 66316 32152 66356 32192
rect 65644 31564 65684 31604
rect 65356 31396 65396 31436
rect 65164 29716 65204 29756
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 64972 29044 65012 29084
rect 64684 28456 64724 28496
rect 64396 28288 64436 28328
rect 64588 28288 64628 28328
rect 64300 28204 64340 28244
rect 64972 28204 65012 28244
rect 64876 28120 64916 28160
rect 65740 31396 65780 31436
rect 66316 31396 66356 31436
rect 66220 31312 66260 31352
rect 66700 32824 66740 32864
rect 66700 32152 66740 32192
rect 67180 34840 67220 34880
rect 67756 36016 67796 36056
rect 67564 34924 67604 34964
rect 67276 34672 67316 34712
rect 67468 34672 67508 34712
rect 67372 34336 67412 34376
rect 67660 34840 67700 34880
rect 67948 38200 67988 38240
rect 68044 36604 68084 36644
rect 67948 35932 67988 35972
rect 67852 35764 67892 35804
rect 67852 34840 67892 34880
rect 66988 32824 67028 32864
rect 66892 31648 66932 31688
rect 66988 31312 67028 31352
rect 69292 38200 69332 38240
rect 70636 38200 70676 38240
rect 68908 38116 68948 38156
rect 68428 37360 68468 37400
rect 68236 37192 68276 37232
rect 68620 37192 68660 37232
rect 68524 36772 68564 36812
rect 68620 36688 68660 36728
rect 68812 36688 68852 36728
rect 68428 36016 68468 36056
rect 68236 35428 68276 35468
rect 68140 35344 68180 35384
rect 69100 37360 69140 37400
rect 71020 38116 71060 38156
rect 69388 37948 69428 37988
rect 69100 36688 69140 36728
rect 69100 35848 69140 35888
rect 68812 34840 68852 34880
rect 68812 34588 68852 34628
rect 69580 37192 69620 37232
rect 69580 36772 69620 36812
rect 69484 36016 69524 36056
rect 69676 35848 69716 35888
rect 69772 35764 69812 35804
rect 69964 35848 70004 35888
rect 69868 35680 69908 35720
rect 69292 35596 69332 35636
rect 69580 35596 69620 35636
rect 69196 33916 69236 33956
rect 67948 32152 67988 32192
rect 68236 30724 68276 30764
rect 65452 30136 65492 30176
rect 65452 29632 65492 29672
rect 66028 30640 66068 30680
rect 65740 29800 65780 29840
rect 65356 29044 65396 29084
rect 65548 29044 65588 29084
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 65164 27784 65204 27824
rect 65260 27700 65300 27740
rect 65356 27616 65396 27656
rect 64492 27532 64532 27572
rect 64396 27364 64436 27404
rect 65452 27532 65492 27572
rect 65260 27364 65300 27404
rect 64300 27112 64340 27152
rect 63820 26776 63860 26816
rect 63820 26104 63860 26144
rect 63916 25852 63956 25892
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 64780 26188 64820 26228
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 63532 25516 63572 25556
rect 64012 25516 64052 25556
rect 63436 25432 63476 25472
rect 62860 25264 62900 25304
rect 63148 25180 63188 25220
rect 63724 25432 63764 25472
rect 63628 25348 63668 25388
rect 63436 25012 63476 25052
rect 62668 24760 62708 24800
rect 62572 24424 62612 24464
rect 63052 24424 63092 24464
rect 62476 24340 62516 24380
rect 62956 24256 62996 24296
rect 62860 24172 62900 24212
rect 62092 24004 62132 24044
rect 62284 24004 62324 24044
rect 62476 23836 62516 23876
rect 62764 23836 62804 23876
rect 60076 23500 60116 23540
rect 63052 23920 63092 23960
rect 62956 23836 62996 23876
rect 63916 25096 63956 25136
rect 63820 24592 63860 24632
rect 64588 25012 64628 25052
rect 64108 24676 64148 24716
rect 64396 24508 64436 24548
rect 64972 25936 65012 25976
rect 66604 30304 66644 30344
rect 66220 29632 66260 29672
rect 65644 27784 65684 27824
rect 65836 28120 65876 28160
rect 65740 27700 65780 27740
rect 65356 26272 65396 26312
rect 65548 26272 65588 26312
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 64876 24676 64916 24716
rect 65260 24676 65300 24716
rect 64780 24592 64820 24632
rect 65452 26104 65492 26144
rect 65932 27784 65972 27824
rect 65740 27532 65780 27572
rect 65452 25936 65492 25976
rect 65740 26104 65780 26144
rect 65644 25852 65684 25892
rect 64972 24592 65012 24632
rect 65356 24592 65396 24632
rect 66412 26776 66452 26816
rect 65932 25096 65972 25136
rect 66412 25012 66452 25052
rect 66412 24676 66452 24716
rect 65932 24592 65972 24632
rect 65644 24508 65684 24548
rect 64684 24424 64724 24464
rect 65164 24424 65204 24464
rect 66124 24340 66164 24380
rect 65740 24088 65780 24128
rect 65260 24004 65300 24044
rect 65644 24004 65684 24044
rect 64876 23920 64916 23960
rect 65164 23920 65204 23960
rect 64492 23836 64532 23876
rect 64780 23836 64820 23876
rect 62860 23416 62900 23456
rect 63244 23584 63284 23624
rect 63244 23416 63284 23456
rect 63628 23584 63668 23624
rect 60455 22744 60495 22784
rect 66796 28624 66836 28664
rect 68428 29632 68468 29672
rect 67756 29212 67796 29252
rect 68428 29044 68468 29084
rect 68428 28540 68468 28580
rect 66988 28288 67028 28328
rect 67276 28288 67316 28328
rect 68140 28120 68180 28160
rect 68332 27784 68372 27824
rect 66892 27364 66932 27404
rect 67660 27280 67700 27320
rect 67564 26944 67604 26984
rect 67756 26776 67796 26816
rect 68428 27700 68468 27740
rect 69100 33076 69140 33116
rect 69004 32824 69044 32864
rect 69964 35344 70004 35384
rect 69676 34924 69716 34964
rect 69772 34840 69812 34880
rect 69580 34756 69620 34796
rect 68716 32656 68756 32696
rect 68908 32656 68948 32696
rect 69100 32656 69140 32696
rect 68812 32404 68852 32444
rect 68620 27784 68660 27824
rect 67660 26608 67700 26648
rect 67372 26356 67412 26396
rect 67276 26188 67316 26228
rect 67180 26104 67220 26144
rect 68428 26440 68468 26480
rect 67084 25180 67124 25220
rect 68236 26188 68276 26228
rect 67372 25096 67412 25136
rect 68332 25264 68372 25304
rect 67660 25012 67700 25052
rect 67564 24760 67604 24800
rect 67852 25012 67892 25052
rect 68332 25012 68372 25052
rect 67660 24592 67700 24632
rect 68140 24592 68180 24632
rect 67276 23752 67316 23792
rect 67564 23752 67604 23792
rect 68620 26776 68660 26816
rect 68620 26524 68660 26564
rect 68620 26188 68660 26228
rect 68620 25936 68660 25976
rect 68524 25264 68564 25304
rect 68524 23920 68564 23960
rect 67660 23668 67700 23708
rect 68044 23668 68084 23708
rect 69004 32152 69044 32192
rect 69100 31312 69140 31352
rect 69100 31144 69140 31184
rect 68908 28960 68948 29000
rect 68812 26440 68852 26480
rect 68812 26188 68852 26228
rect 69292 32068 69332 32108
rect 69484 32152 69524 32192
rect 69388 31984 69428 32024
rect 69964 33664 70004 33704
rect 69772 32656 69812 32696
rect 71116 37948 71156 37988
rect 70444 37360 70484 37400
rect 71404 37192 71444 37232
rect 70732 36856 70772 36896
rect 70444 36688 70484 36728
rect 70252 35932 70292 35972
rect 70348 35848 70388 35888
rect 70444 35344 70484 35384
rect 70348 35260 70388 35300
rect 70252 35092 70292 35132
rect 70444 35176 70484 35216
rect 70348 34588 70388 34628
rect 70060 31984 70100 32024
rect 69676 30052 69716 30092
rect 69292 29800 69332 29840
rect 69004 27784 69044 27824
rect 69196 28288 69236 28328
rect 69100 27532 69140 27572
rect 69100 27364 69140 27404
rect 69004 26440 69044 26480
rect 68908 23920 68948 23960
rect 68716 23752 68756 23792
rect 69100 26272 69140 26312
rect 69484 29800 69524 29840
rect 69772 29800 69812 29840
rect 69580 29716 69620 29756
rect 69772 29128 69812 29168
rect 70252 31900 70292 31940
rect 70636 35176 70676 35216
rect 70540 35092 70580 35132
rect 70636 34840 70676 34880
rect 71596 36772 71636 36812
rect 71596 36520 71636 36560
rect 70924 36436 70964 36476
rect 70828 36016 70868 36056
rect 70732 34420 70772 34460
rect 71404 35764 71444 35804
rect 70924 35428 70964 35468
rect 71308 35260 71348 35300
rect 70636 33916 70676 33956
rect 70540 32236 70580 32276
rect 71020 33916 71060 33956
rect 71212 34504 71252 34544
rect 71308 34420 71348 34460
rect 71116 33496 71156 33536
rect 74284 38200 74324 38240
rect 72076 36688 72116 36728
rect 73324 37528 73364 37568
rect 73132 37444 73172 37484
rect 72940 37108 72980 37148
rect 73228 37360 73268 37400
rect 73708 37444 73748 37484
rect 73516 37360 73556 37400
rect 73036 37024 73076 37064
rect 72940 36520 72980 36560
rect 72172 36436 72212 36476
rect 72172 36016 72212 36056
rect 71884 35848 71924 35888
rect 72076 35848 72116 35888
rect 71692 35512 71732 35552
rect 71788 35176 71828 35216
rect 71500 34756 71540 34796
rect 72652 35512 72692 35552
rect 71692 34504 71732 34544
rect 71500 34000 71540 34040
rect 71980 34336 72020 34376
rect 71788 34000 71828 34040
rect 70924 32824 70964 32864
rect 70732 32320 70772 32360
rect 70636 32152 70676 32192
rect 71116 32572 71156 32612
rect 71020 32236 71060 32276
rect 70732 32068 70772 32108
rect 70732 31480 70772 31520
rect 71212 31900 71252 31940
rect 71116 31480 71156 31520
rect 70540 30808 70580 30848
rect 70732 31060 70772 31100
rect 71020 31060 71060 31100
rect 70636 30724 70676 30764
rect 70540 30640 70580 30680
rect 70444 30388 70484 30428
rect 69964 29716 70004 29756
rect 69964 29464 70004 29504
rect 70348 29464 70388 29504
rect 70156 29212 70196 29252
rect 70828 30808 70868 30848
rect 71020 30640 71060 30680
rect 71020 30472 71060 30512
rect 70924 30388 70964 30428
rect 70636 29800 70676 29840
rect 70828 29464 70868 29504
rect 70540 29128 70580 29168
rect 70156 29044 70196 29084
rect 71116 29968 71156 30008
rect 71020 29800 71060 29840
rect 71788 33496 71828 33536
rect 71500 32824 71540 32864
rect 71788 32656 71828 32696
rect 71500 32320 71540 32360
rect 71692 32320 71732 32360
rect 71404 31732 71444 31772
rect 71404 31564 71444 31604
rect 71404 31312 71444 31352
rect 71692 31732 71732 31772
rect 71596 31480 71636 31520
rect 71980 34000 72020 34040
rect 72172 33664 72212 33704
rect 71980 33580 72020 33620
rect 71980 32656 72020 32696
rect 71980 32236 72020 32276
rect 71980 31984 72020 32024
rect 71884 31648 71924 31688
rect 71692 31060 71732 31100
rect 71596 30976 71636 31016
rect 71308 30808 71348 30848
rect 71308 30556 71348 30596
rect 71500 30808 71540 30848
rect 71500 29884 71540 29924
rect 71404 29464 71444 29504
rect 71788 30220 71828 30260
rect 72556 33664 72596 33704
rect 72844 34336 72884 34376
rect 72652 32992 72692 33032
rect 72460 32824 72500 32864
rect 73324 37192 73364 37232
rect 73036 36016 73076 36056
rect 73228 36016 73268 36056
rect 73132 35848 73172 35888
rect 73228 35512 73268 35552
rect 73996 37360 74036 37400
rect 73900 37192 73940 37232
rect 73036 32992 73076 33032
rect 72748 32236 72788 32276
rect 72940 32152 72980 32192
rect 72460 31984 72500 32024
rect 72076 31564 72116 31604
rect 73036 31900 73076 31940
rect 72172 30220 72212 30260
rect 71692 30052 71732 30092
rect 71884 29884 71924 29924
rect 72268 29968 72308 30008
rect 70636 29044 70676 29084
rect 71020 29044 71060 29084
rect 70348 28876 70388 28916
rect 70060 28792 70100 28832
rect 69868 28288 69908 28328
rect 70060 27952 70100 27992
rect 70060 27784 70100 27824
rect 69292 26776 69332 26816
rect 69580 27364 69620 27404
rect 69484 26356 69524 26396
rect 69388 26272 69428 26312
rect 69292 26188 69332 26228
rect 69388 26104 69428 26144
rect 69772 27616 69812 27656
rect 69772 27448 69812 27488
rect 69196 25852 69236 25892
rect 70252 28456 70292 28496
rect 70636 28540 70676 28580
rect 70828 28876 70868 28916
rect 71212 28792 71252 28832
rect 70540 27952 70580 27992
rect 70732 27952 70772 27992
rect 70252 27448 70292 27488
rect 70636 27784 70676 27824
rect 71116 28456 71156 28496
rect 71020 28288 71060 28328
rect 71212 27952 71252 27992
rect 70636 27448 70676 27488
rect 70540 26104 70580 26144
rect 71596 29044 71636 29084
rect 71500 28540 71540 28580
rect 71500 28120 71540 28160
rect 70444 26020 70484 26060
rect 70636 26020 70676 26060
rect 70540 25936 70580 25976
rect 70348 25852 70388 25892
rect 70348 25012 70388 25052
rect 71116 27280 71156 27320
rect 70924 27112 70964 27152
rect 71020 26272 71060 26312
rect 70732 25516 70772 25556
rect 70540 24928 70580 24968
rect 71020 24760 71060 24800
rect 71020 24592 71060 24632
rect 70156 23920 70196 23960
rect 70540 23920 70580 23960
rect 70828 23920 70868 23960
rect 70156 23752 70196 23792
rect 70444 23752 70484 23792
rect 71308 26188 71348 26228
rect 71692 27784 71732 27824
rect 71788 27616 71828 27656
rect 71596 27112 71636 27152
rect 71692 27028 71732 27068
rect 71884 27112 71924 27152
rect 71884 26608 71924 26648
rect 72268 26692 72308 26732
rect 71980 26440 72020 26480
rect 71788 26272 71828 26312
rect 71500 26188 71540 26228
rect 73036 26860 73076 26900
rect 71980 25852 72020 25892
rect 72652 25852 72692 25892
rect 71212 25432 71252 25472
rect 71404 25096 71444 25136
rect 71212 24928 71252 24968
rect 71308 24592 71348 24632
rect 71596 24760 71636 24800
rect 72844 25096 72884 25136
rect 73036 25096 73076 25136
rect 72460 25012 72500 25052
rect 72076 24676 72116 24716
rect 74572 37276 74612 37316
rect 74956 37276 74996 37316
rect 75052 37108 75092 37148
rect 74764 36688 74804 36728
rect 75244 37192 75284 37232
rect 75148 37024 75188 37064
rect 75052 36016 75092 36056
rect 74284 35932 74324 35972
rect 74476 35932 74516 35972
rect 73900 35848 73940 35888
rect 73708 35680 73748 35720
rect 74188 35176 74228 35216
rect 73420 32824 73460 32864
rect 73612 32824 73652 32864
rect 73900 32236 73940 32276
rect 73612 32152 73652 32192
rect 73228 30976 73268 31016
rect 73612 30808 73652 30848
rect 73708 29968 73748 30008
rect 73420 28708 73460 28748
rect 73228 25936 73268 25976
rect 73132 23920 73172 23960
rect 73324 23920 73364 23960
rect 73612 23920 73652 23960
rect 70924 23584 70964 23624
rect 71212 23584 71252 23624
rect 73804 28540 73844 28580
rect 73804 23920 73844 23960
rect 74092 29968 74132 30008
rect 76588 37360 76628 37400
rect 75532 37024 75572 37064
rect 74380 34924 74420 34964
rect 74284 27952 74324 27992
rect 75340 34336 75380 34376
rect 74476 33496 74516 33536
rect 74764 33412 74804 33452
rect 74860 32824 74900 32864
rect 74572 32236 74612 32276
rect 75148 32656 75188 32696
rect 74572 31144 74612 31184
rect 74476 26104 74516 26144
rect 74476 25936 74516 25976
rect 74380 25852 74420 25892
rect 74284 25516 74324 25556
rect 74476 25264 74516 25304
rect 74860 30976 74900 31016
rect 76108 37192 76148 37232
rect 76300 36772 76340 36812
rect 75724 36016 75764 36056
rect 75532 34336 75572 34376
rect 76876 37276 76916 37316
rect 76780 36772 76820 36812
rect 76684 36688 76724 36728
rect 76588 36520 76628 36560
rect 76780 36352 76820 36392
rect 75916 35848 75956 35888
rect 76204 35848 76244 35888
rect 75532 34168 75572 34208
rect 75820 34336 75860 34376
rect 75820 33748 75860 33788
rect 75436 32824 75476 32864
rect 76396 35848 76436 35888
rect 76012 35176 76052 35216
rect 76588 34672 76628 34712
rect 76396 34588 76436 34628
rect 76204 34504 76244 34544
rect 76588 34420 76628 34460
rect 76012 34168 76052 34208
rect 76684 34336 76724 34376
rect 76300 33832 76340 33872
rect 76204 33496 76244 33536
rect 76012 33412 76052 33452
rect 76012 32824 76052 32864
rect 75916 32656 75956 32696
rect 75820 32152 75860 32192
rect 75532 31228 75572 31268
rect 75340 30892 75380 30932
rect 75532 30892 75572 30932
rect 74764 30640 74804 30680
rect 74956 30640 74996 30680
rect 74860 30472 74900 30512
rect 75148 30640 75188 30680
rect 75052 30472 75092 30512
rect 74956 30388 74996 30428
rect 74956 30220 74996 30260
rect 75436 30808 75476 30848
rect 75436 30472 75476 30512
rect 75340 30220 75380 30260
rect 74860 29716 74900 29756
rect 74668 27028 74708 27068
rect 74860 26860 74900 26900
rect 74764 26776 74804 26816
rect 74860 26692 74900 26732
rect 74764 26356 74804 26396
rect 74668 26104 74708 26144
rect 75052 29884 75092 29924
rect 75532 30220 75572 30260
rect 75724 30220 75764 30260
rect 75532 29800 75572 29840
rect 75340 28708 75380 28748
rect 75436 28288 75476 28328
rect 75436 27952 75476 27992
rect 75052 27616 75092 27656
rect 76012 31732 76052 31772
rect 75916 31480 75956 31520
rect 76012 30640 76052 30680
rect 75916 30388 75956 30428
rect 76012 29800 76052 29840
rect 75916 29716 75956 29756
rect 76012 29464 76052 29504
rect 76300 30724 76340 30764
rect 76588 33664 76628 33704
rect 76684 33664 76724 33704
rect 76492 33412 76532 33452
rect 76684 33328 76724 33368
rect 76588 32152 76628 32192
rect 76684 31984 76724 32024
rect 76492 31060 76532 31100
rect 76588 30640 76628 30680
rect 76396 30472 76436 30512
rect 76204 30388 76244 30428
rect 76300 30304 76340 30344
rect 76204 29296 76244 29336
rect 75052 27364 75092 27404
rect 75244 27364 75284 27404
rect 74860 26188 74900 26228
rect 74956 26104 74996 26144
rect 74764 25936 74804 25976
rect 74476 24928 74516 24968
rect 74284 24592 74324 24632
rect 74572 24844 74612 24884
rect 74476 24508 74516 24548
rect 74092 24004 74132 24044
rect 74764 24592 74804 24632
rect 74860 24004 74900 24044
rect 75820 27028 75860 27068
rect 75628 26944 75668 26984
rect 75436 26860 75476 26900
rect 75628 26776 75668 26816
rect 75916 26776 75956 26816
rect 75820 26692 75860 26732
rect 75724 26608 75764 26648
rect 75148 25936 75188 25976
rect 75436 26104 75476 26144
rect 75820 26440 75860 26480
rect 75820 26104 75860 26144
rect 75916 25516 75956 25556
rect 76492 29464 76532 29504
rect 76396 28372 76436 28412
rect 77452 37360 77492 37400
rect 77356 37192 77396 37232
rect 77260 37108 77300 37148
rect 77068 36520 77108 36560
rect 77548 36772 77588 36812
rect 77260 36352 77300 36392
rect 77068 35848 77108 35888
rect 77068 35512 77108 35552
rect 76876 34672 76916 34712
rect 77068 34588 77108 34628
rect 76972 34504 77012 34544
rect 76972 34336 77012 34376
rect 76876 34252 76916 34292
rect 77452 35848 77492 35888
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 77836 37192 77876 37232
rect 78124 37276 78164 37316
rect 78412 37360 78452 37400
rect 78220 37108 78260 37148
rect 79468 37108 79508 37148
rect 78316 36688 78356 36728
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 77932 35680 77972 35720
rect 77644 34504 77684 34544
rect 78124 34336 78164 34376
rect 77260 33664 77300 33704
rect 77452 33664 77492 33704
rect 77356 33496 77396 33536
rect 76972 33412 77012 33452
rect 77164 33412 77204 33452
rect 77164 32992 77204 33032
rect 76972 32320 77012 32360
rect 76876 31648 76916 31688
rect 77164 31984 77204 32024
rect 76972 31480 77012 31520
rect 77452 32320 77492 32360
rect 77740 32992 77780 33032
rect 77740 32656 77780 32696
rect 78124 33496 78164 33536
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 79468 34336 79508 34376
rect 78412 33664 78452 33704
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 78124 32992 78164 33032
rect 78508 32992 78548 33032
rect 78220 32824 78260 32864
rect 78028 32656 78068 32696
rect 78028 31900 78068 31940
rect 77452 31312 77492 31352
rect 77452 30976 77492 31016
rect 77068 30892 77108 30932
rect 76972 30220 77012 30260
rect 77164 30640 77204 30680
rect 76684 28624 76724 28664
rect 77644 31060 77684 31100
rect 77644 30808 77684 30848
rect 77548 30472 77588 30512
rect 77164 29716 77204 29756
rect 77068 28624 77108 28664
rect 76588 28288 76628 28328
rect 76684 28036 76724 28076
rect 76876 28288 76916 28328
rect 76972 28204 77012 28244
rect 77356 28288 77396 28328
rect 77260 28204 77300 28244
rect 77164 28120 77204 28160
rect 77068 28036 77108 28076
rect 76300 26692 76340 26732
rect 76588 26776 76628 26816
rect 76204 26608 76244 26648
rect 76492 26608 76532 26648
rect 76300 25516 76340 25556
rect 76876 27616 76916 27656
rect 77068 27616 77108 27656
rect 76780 26104 76820 26144
rect 77356 26608 77396 26648
rect 77356 26104 77396 26144
rect 75724 24592 75764 24632
rect 75340 24508 75380 24548
rect 75916 24424 75956 24464
rect 75244 23836 75284 23876
rect 75532 23836 75572 23876
rect 75052 23752 75092 23792
rect 74860 23584 74900 23624
rect 75244 23584 75284 23624
rect 76492 25180 76532 25220
rect 76588 24592 76628 24632
rect 76396 24508 76436 24548
rect 76108 24424 76148 24464
rect 76108 23752 76148 23792
rect 76492 23752 76532 23792
rect 76876 25180 76916 25220
rect 77836 31312 77876 31352
rect 77836 30808 77876 30848
rect 77740 26104 77780 26144
rect 78412 31984 78452 32024
rect 79468 31900 79508 31940
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 79468 30808 79508 30848
rect 78028 30472 78068 30512
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 78124 28288 78164 28328
rect 79468 28288 79508 28328
rect 77932 25264 77972 25304
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 78508 26608 78548 26648
rect 79468 26608 79508 26648
rect 78316 25264 78356 25304
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 78988 24592 79028 24632
rect 79084 23752 79124 23792
rect 78796 23416 78836 23456
rect 79276 23416 79316 23456
rect 78604 22744 78644 22784
rect 78855 22744 78895 22784
rect 53068 17620 53108 17660
rect 53545 17284 53585 17324
rect 53655 17200 53695 17240
rect 53945 17200 53985 17240
rect 52876 17116 52916 17156
rect 54345 17116 54385 17156
rect 54455 17116 54495 17156
rect 52492 16948 52532 16988
rect 52396 16780 52436 16820
rect 54028 16780 54068 16820
rect 53068 16696 53108 16736
rect 52492 16612 52532 16652
rect 52012 15352 52052 15392
rect 52396 16192 52436 16232
rect 52780 16528 52820 16568
rect 52780 16276 52820 16316
rect 53740 16612 53780 16652
rect 53068 16218 53108 16232
rect 53068 16192 53108 16218
rect 53740 16360 53780 16400
rect 52684 15520 52724 15560
rect 52396 14932 52436 14972
rect 52684 14260 52724 14300
rect 52588 14176 52628 14216
rect 53164 14932 53204 14972
rect 53068 14176 53108 14216
rect 52684 14008 52724 14048
rect 54028 16192 54068 16232
rect 53644 15688 53684 15728
rect 54028 14764 54068 14804
rect 53644 14512 53684 14552
rect 53452 14092 53492 14132
rect 53356 13924 53396 13964
rect 52108 13840 52148 13880
rect 51916 13588 51956 13628
rect 52108 13252 52148 13292
rect 51916 12916 51956 12956
rect 50860 11824 50900 11864
rect 51724 11740 51764 11780
rect 51532 11656 51572 11696
rect 53260 13252 53300 13292
rect 53356 13168 53396 13208
rect 54988 17200 55028 17240
rect 55145 17200 55185 17240
rect 54700 16192 54740 16232
rect 55545 17200 55585 17240
rect 55945 17200 55985 17240
rect 55564 16444 55604 16484
rect 55468 16360 55508 16400
rect 55084 16276 55124 16316
rect 54316 15520 54356 15560
rect 54988 15520 55028 15560
rect 54700 14680 54740 14720
rect 54508 13672 54548 13712
rect 54316 13588 54356 13628
rect 53644 13336 53684 13376
rect 54316 13336 54356 13376
rect 53548 13168 53588 13208
rect 53452 13084 53492 13124
rect 54412 13168 54452 13208
rect 54988 14428 55028 14468
rect 55276 16192 55316 16232
rect 55180 16024 55220 16064
rect 55660 16192 55700 16232
rect 55756 16024 55796 16064
rect 55564 15856 55604 15896
rect 54700 13168 54740 13208
rect 55180 13252 55220 13292
rect 55084 13168 55124 13208
rect 56524 16108 56564 16148
rect 56044 15856 56084 15896
rect 56332 14680 56372 14720
rect 55948 14428 55988 14468
rect 55852 13756 55892 13796
rect 55756 13420 55796 13460
rect 55372 13168 55412 13208
rect 55276 13000 55316 13040
rect 56428 14092 56468 14132
rect 56236 13924 56276 13964
rect 56044 13168 56084 13208
rect 56524 13756 56564 13796
rect 56428 13588 56468 13628
rect 57945 17116 57985 17156
rect 57292 15940 57332 15980
rect 58345 17200 58385 17240
rect 58252 16192 58292 16232
rect 58540 16192 58580 16232
rect 57868 15856 57908 15896
rect 56908 14764 56948 14804
rect 57580 14680 57620 14720
rect 57676 14428 57716 14468
rect 57388 13924 57428 13964
rect 57100 13756 57140 13796
rect 56908 13672 56948 13712
rect 56812 13504 56852 13544
rect 56428 13168 56468 13208
rect 56332 13084 56372 13124
rect 53293 12244 53333 12284
rect 52588 11824 52628 11864
rect 52204 11656 52244 11696
rect 52396 11656 52436 11696
rect 50764 11572 50804 11612
rect 51244 11572 51284 11612
rect 51436 11572 51476 11612
rect 51916 11572 51956 11612
rect 50668 10984 50708 11024
rect 50956 11152 50996 11192
rect 50860 10984 50900 11024
rect 52300 11572 52340 11612
rect 52108 11152 52148 11192
rect 50284 9472 50324 9512
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 50476 7456 50516 7496
rect 51916 10900 51956 10940
rect 51436 9472 51476 9512
rect 52012 9640 52052 9680
rect 51724 9472 51764 9512
rect 51628 9388 51668 9428
rect 51148 8128 51188 8168
rect 49612 7120 49652 7160
rect 49996 7120 50036 7160
rect 50188 7120 50228 7160
rect 50860 7120 50900 7160
rect 51052 7120 51092 7160
rect 51724 7120 51764 7160
rect 48940 6280 48980 6320
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 48460 5608 48500 5648
rect 48268 4936 48308 4976
rect 48556 5020 48596 5060
rect 48844 4936 48884 4976
rect 49132 5440 49172 5480
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 50092 5608 50132 5648
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 49228 4852 49268 4892
rect 48556 4768 48596 4808
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 50764 4180 50804 4220
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 50188 3760 50228 3800
rect 51436 6448 51476 6488
rect 51244 6112 51284 6152
rect 51244 5608 51284 5648
rect 52300 10984 52340 11024
rect 52204 10060 52244 10100
rect 52108 9556 52148 9596
rect 52204 9472 52244 9512
rect 52492 10144 52532 10184
rect 53740 11740 53780 11780
rect 53644 11656 53684 11696
rect 52684 10984 52724 11024
rect 52396 9472 52436 9512
rect 52684 9640 52724 9680
rect 53164 10984 53204 11024
rect 53452 10984 53492 11024
rect 53068 10816 53108 10856
rect 53548 10900 53588 10940
rect 53164 10060 53204 10100
rect 53452 9724 53492 9764
rect 52876 9388 52916 9428
rect 52684 9052 52724 9092
rect 52300 8044 52340 8084
rect 52588 8044 52628 8084
rect 52396 6700 52436 6740
rect 52012 5524 52052 5564
rect 52492 6448 52532 6488
rect 53068 9472 53108 9512
rect 53356 9472 53396 9512
rect 52972 8548 53012 8588
rect 53164 9052 53204 9092
rect 53356 8548 53396 8588
rect 53548 8548 53588 8588
rect 53260 8044 53300 8084
rect 52972 7792 53012 7832
rect 52876 7456 52916 7496
rect 53067 7036 53107 7076
rect 52684 6448 52724 6488
rect 52588 5860 52628 5900
rect 54124 9724 54164 9764
rect 54316 9472 54356 9512
rect 54028 8968 54068 9008
rect 53740 8044 53780 8084
rect 53740 7792 53780 7832
rect 53644 7288 53684 7328
rect 54124 8044 54164 8084
rect 54796 12580 54836 12620
rect 55180 12244 55220 12284
rect 56620 13168 56660 13208
rect 56716 12916 56756 12956
rect 56620 12580 56660 12620
rect 57484 13084 57524 13124
rect 57772 14260 57812 14300
rect 58348 14428 58388 14468
rect 57964 14260 58004 14300
rect 57868 13420 57908 13460
rect 57868 13252 57908 13292
rect 57676 13000 57716 13040
rect 58924 14512 58964 14552
rect 58828 13672 58868 13712
rect 58252 13588 58292 13628
rect 58060 13000 58100 13040
rect 57388 12832 57428 12872
rect 57196 12664 57236 12704
rect 57484 11908 57524 11948
rect 56812 11824 56852 11864
rect 57292 11656 57332 11696
rect 57868 12832 57908 12872
rect 57676 12664 57716 12704
rect 57772 12412 57812 12452
rect 57676 11824 57716 11864
rect 57964 12160 58004 12200
rect 57964 11824 58004 11864
rect 56332 11236 56372 11276
rect 56332 10816 56372 10856
rect 56524 10396 56564 10436
rect 56716 9724 56756 9764
rect 54604 7876 54644 7916
rect 53452 7204 53492 7244
rect 52780 5776 52820 5816
rect 53356 7036 53396 7076
rect 52972 5860 53012 5900
rect 52396 5440 52436 5480
rect 51532 4348 51572 4388
rect 51820 4936 51860 4976
rect 51820 4684 51860 4724
rect 51724 4432 51764 4472
rect 51628 4264 51668 4304
rect 50860 3928 50900 3968
rect 51628 3760 51668 3800
rect 50956 3424 50996 3464
rect 52108 4096 52148 4136
rect 52108 3508 52148 3548
rect 52012 3424 52052 3464
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 52396 4684 52436 4724
rect 52684 4936 52724 4976
rect 52684 4348 52724 4388
rect 52588 4264 52628 4304
rect 52588 4096 52628 4136
rect 52780 4264 52820 4304
rect 53068 5608 53108 5648
rect 53164 5524 53204 5564
rect 53548 5608 53588 5648
rect 54220 7288 54260 7328
rect 54412 7288 54452 7328
rect 54892 7204 54932 7244
rect 54316 6700 54356 6740
rect 54220 6532 54260 6572
rect 53836 5692 53876 5732
rect 53740 5608 53780 5648
rect 53644 4852 53684 4892
rect 54604 6532 54644 6572
rect 54412 5776 54452 5816
rect 54796 5776 54836 5816
rect 54124 5692 54164 5732
rect 54700 5692 54740 5732
rect 54220 5608 54260 5648
rect 55948 8548 55988 8588
rect 57388 10228 57428 10268
rect 58156 12664 58196 12704
rect 58636 13420 58676 13460
rect 58444 13168 58484 13208
rect 58732 13168 58772 13208
rect 58540 13084 58580 13124
rect 58252 12160 58292 12200
rect 58060 10396 58100 10436
rect 57868 10312 57908 10352
rect 58348 11656 58388 11696
rect 58540 11656 58580 11696
rect 59020 12580 59060 12620
rect 60745 17116 60785 17156
rect 60940 17116 60980 17156
rect 59500 15856 59540 15896
rect 59500 14680 59540 14720
rect 59404 14344 59444 14384
rect 59308 13336 59348 13376
rect 59212 12496 59252 12536
rect 60844 16444 60884 16484
rect 59980 15352 60020 15392
rect 59692 12580 59732 12620
rect 59020 11992 59060 12032
rect 58924 11572 58964 11612
rect 58444 11152 58484 11192
rect 58348 10144 58388 10184
rect 58060 9640 58100 9680
rect 58060 8884 58100 8924
rect 57772 8800 57812 8840
rect 57964 8800 58004 8840
rect 57868 8464 57908 8504
rect 55564 7120 55604 7160
rect 55084 6448 55124 6488
rect 54892 5608 54932 5648
rect 54028 4936 54068 4976
rect 53836 4432 53876 4472
rect 53260 4096 53300 4136
rect 53644 4096 53684 4136
rect 55084 4096 55124 4136
rect 52972 3928 53012 3968
rect 52780 3844 52820 3884
rect 54796 3844 54836 3884
rect 53932 3592 53972 3632
rect 52780 3424 52820 3464
rect 55372 4180 55412 4220
rect 55180 3424 55220 3464
rect 8908 2668 8948 2708
rect 52300 2668 52340 2708
rect 4300 2584 4340 2624
rect 4780 2584 4820 2624
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 55468 3928 55508 3968
rect 55852 6448 55892 6488
rect 57004 6784 57044 6824
rect 57292 6448 57332 6488
rect 56908 6280 56948 6320
rect 56236 5608 56276 5648
rect 55660 4936 55700 4976
rect 55660 4768 55700 4808
rect 55948 4936 55988 4976
rect 56332 4936 56372 4976
rect 56140 4768 56180 4808
rect 57004 5692 57044 5732
rect 58252 9808 58292 9848
rect 58348 9640 58388 9680
rect 58348 9052 58388 9092
rect 58924 11152 58964 11192
rect 59500 11992 59540 12032
rect 59308 11572 59348 11612
rect 59308 11320 59348 11360
rect 58732 10228 58772 10268
rect 58924 10228 58964 10268
rect 59212 10312 59252 10352
rect 59404 11152 59444 11192
rect 59692 11992 59732 12032
rect 59788 10984 59828 11024
rect 59692 10228 59732 10268
rect 59308 9640 59348 9680
rect 58636 9472 58676 9512
rect 58732 8884 58772 8924
rect 58732 8716 58772 8756
rect 58444 8464 58484 8504
rect 58156 8380 58196 8420
rect 58060 8044 58100 8084
rect 58636 8632 58676 8672
rect 59020 8968 59060 9008
rect 59212 8716 59252 8756
rect 59116 8632 59156 8672
rect 59500 10060 59540 10100
rect 59596 9640 59636 9680
rect 59692 9472 59732 9512
rect 59500 8464 59540 8504
rect 58828 8380 58868 8420
rect 58540 8044 58580 8084
rect 58348 7708 58388 7748
rect 57964 6616 58004 6656
rect 58060 6532 58100 6572
rect 58156 6448 58196 6488
rect 58540 6532 58580 6572
rect 58828 7708 58868 7748
rect 58732 6616 58772 6656
rect 58060 6280 58100 6320
rect 58252 6280 58292 6320
rect 58060 6028 58100 6068
rect 57580 4936 57620 4976
rect 56716 4852 56756 4892
rect 56524 4768 56564 4808
rect 55852 4348 55892 4388
rect 55756 4180 55796 4220
rect 55660 4096 55700 4136
rect 55948 4012 55988 4052
rect 55852 3928 55892 3968
rect 55948 3592 55988 3632
rect 55948 3424 55988 3464
rect 54796 1912 54836 1952
rect 53548 1324 53588 1364
rect 55564 2080 55604 2120
rect 55756 2668 55796 2708
rect 55948 2584 55988 2624
rect 56236 4432 56276 4472
rect 56620 4012 56660 4052
rect 56332 3508 56372 3548
rect 57004 4432 57044 4472
rect 56812 4348 56852 4388
rect 56140 3172 56180 3212
rect 56716 3172 56756 3212
rect 55660 1912 55700 1952
rect 55564 1408 55604 1448
rect 55372 1324 55412 1364
rect 55948 2080 55988 2120
rect 56332 2416 56372 2456
rect 56716 2584 56756 2624
rect 56620 2500 56660 2540
rect 56524 2416 56564 2456
rect 56332 1492 56372 1532
rect 56236 1408 56276 1448
rect 55852 1072 55892 1112
rect 56236 1072 56276 1112
rect 57292 4348 57332 4388
rect 57100 4096 57140 4136
rect 57388 4264 57428 4304
rect 57964 4264 58004 4304
rect 58156 5608 58196 5648
rect 58540 4768 58580 4808
rect 58636 4264 58676 4304
rect 57196 3508 57236 3548
rect 57004 2500 57044 2540
rect 56812 2080 56852 2120
rect 57388 2668 57428 2708
rect 57292 2584 57332 2624
rect 56812 1492 56852 1532
rect 57196 1072 57236 1112
rect 58252 4096 58292 4136
rect 58156 2584 58196 2624
rect 57772 1912 57812 1952
rect 57484 1240 57524 1280
rect 58828 6448 58868 6488
rect 59308 6952 59348 6992
rect 59020 6532 59060 6572
rect 59596 7960 59636 8000
rect 59500 6700 59540 6740
rect 59308 6616 59348 6656
rect 59212 6448 59252 6488
rect 59500 6532 59540 6572
rect 59020 6028 59060 6068
rect 58924 5608 58964 5648
rect 58924 5440 58964 5480
rect 59404 5608 59444 5648
rect 59308 5440 59348 5480
rect 59404 5356 59444 5396
rect 59308 5188 59348 5228
rect 59212 4264 59252 4304
rect 58732 4180 58772 4220
rect 59116 4180 59156 4220
rect 59020 4096 59060 4136
rect 58828 3172 58868 3212
rect 58732 3088 58772 3128
rect 58924 2584 58964 2624
rect 59500 3676 59540 3716
rect 59308 3424 59348 3464
rect 59404 3172 59444 3212
rect 59404 2920 59444 2960
rect 59116 2836 59156 2876
rect 59212 2584 59252 2624
rect 58828 2416 58868 2456
rect 58924 2080 58964 2120
rect 58924 1660 58964 1700
rect 59308 1240 59348 1280
rect 59500 1240 59540 1280
rect 60748 16192 60788 16232
rect 60364 15436 60404 15476
rect 60172 15352 60212 15392
rect 60364 15184 60404 15224
rect 60172 14848 60212 14888
rect 60076 11068 60116 11108
rect 61228 16444 61268 16484
rect 61132 16192 61172 16232
rect 61708 16276 61748 16316
rect 60556 14764 60596 14804
rect 60556 14260 60596 14300
rect 60556 13000 60596 13040
rect 60940 15352 60980 15392
rect 60844 14680 60884 14720
rect 61420 14764 61460 14804
rect 61132 14596 61172 14636
rect 60940 13420 60980 13460
rect 60460 10480 60500 10520
rect 60460 10060 60500 10100
rect 60652 8632 60692 8672
rect 59692 5188 59732 5228
rect 59980 7120 60020 7160
rect 60076 7036 60116 7076
rect 60076 6700 60116 6740
rect 59980 6616 60020 6656
rect 59884 5356 59924 5396
rect 59788 4180 59828 4220
rect 59788 3676 59828 3716
rect 59692 2836 59732 2876
rect 60268 7120 60308 7160
rect 60172 6616 60212 6656
rect 60844 12664 60884 12704
rect 60940 11656 60980 11696
rect 61612 14008 61652 14048
rect 61516 13924 61556 13964
rect 61420 13252 61460 13292
rect 61516 13084 61556 13124
rect 61804 15520 61844 15560
rect 61900 14932 61940 14972
rect 61996 14512 62036 14552
rect 61996 14344 62036 14384
rect 61900 13420 61940 13460
rect 62188 14932 62228 14972
rect 62092 14176 62132 14216
rect 62188 14008 62228 14048
rect 61708 11992 61748 12032
rect 61036 11488 61076 11528
rect 61036 10984 61076 11024
rect 60844 9472 60884 9512
rect 60748 8128 60788 8168
rect 60652 7120 60692 7160
rect 60268 6280 60308 6320
rect 61420 6616 61460 6656
rect 61036 5608 61076 5648
rect 61516 5860 61556 5900
rect 62668 16192 62708 16232
rect 62572 15604 62612 15644
rect 62572 14764 62612 14804
rect 62476 14680 62516 14720
rect 62380 14512 62420 14552
rect 62764 14512 62804 14552
rect 63052 16192 63092 16232
rect 62956 15688 62996 15728
rect 62956 14848 62996 14888
rect 62380 14008 62420 14048
rect 62380 13336 62420 13376
rect 62476 13000 62516 13040
rect 62092 12664 62132 12704
rect 61996 12580 62036 12620
rect 61900 11320 61940 11360
rect 62284 12496 62324 12536
rect 62188 12412 62228 12452
rect 61996 10228 62036 10268
rect 61900 10144 61940 10184
rect 62188 10984 62228 11024
rect 62476 12076 62516 12116
rect 62188 9556 62228 9596
rect 62092 9472 62132 9512
rect 61900 8632 61940 8672
rect 62188 7708 62228 7748
rect 61900 7036 61940 7076
rect 62668 14176 62708 14216
rect 62572 11236 62612 11276
rect 62476 9724 62516 9764
rect 62956 13252 62996 13292
rect 62860 13084 62900 13124
rect 62764 12496 62804 12536
rect 62764 11656 62804 11696
rect 64588 17116 64628 17156
rect 64855 17116 64895 17156
rect 63724 16024 63764 16064
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 64684 16864 64724 16904
rect 65356 16948 65396 16988
rect 64972 16192 65012 16232
rect 65740 16360 65780 16400
rect 66604 17116 66644 17156
rect 66855 17116 66895 17156
rect 66124 15856 66164 15896
rect 64876 15772 64916 15812
rect 64108 15016 64148 15056
rect 63436 14764 63476 14804
rect 63724 14764 63764 14804
rect 63916 14764 63956 14804
rect 63244 13504 63284 13544
rect 63724 14512 63764 14552
rect 64300 14764 64340 14804
rect 63820 14428 63860 14468
rect 63916 14008 63956 14048
rect 63628 13924 63668 13964
rect 63820 13924 63860 13964
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 63628 12748 63668 12788
rect 63724 12496 63764 12536
rect 64876 14680 64916 14720
rect 65740 15520 65780 15560
rect 65260 14932 65300 14972
rect 65260 14764 65300 14804
rect 64492 14428 64532 14468
rect 65260 14428 65300 14468
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 64396 14008 64436 14048
rect 64780 13252 64820 13292
rect 64876 13168 64916 13208
rect 65452 14512 65492 14552
rect 65356 14344 65396 14384
rect 66220 15436 66260 15476
rect 64396 12748 64436 12788
rect 64012 12580 64052 12620
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 64588 12496 64628 12536
rect 63052 12076 63092 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 63340 11656 63380 11696
rect 63436 11572 63476 11612
rect 62956 11404 62996 11444
rect 62956 10984 62996 11024
rect 62860 9136 62900 9176
rect 63916 11656 63956 11696
rect 64204 11908 64244 11948
rect 64396 11656 64436 11696
rect 64780 11908 64820 11948
rect 65548 12496 65588 12536
rect 64012 11404 64052 11444
rect 63820 11320 63860 11360
rect 63820 10984 63860 11024
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 63436 10144 63476 10184
rect 63436 9472 63476 9512
rect 63628 10060 63668 10100
rect 63532 9304 63572 9344
rect 63724 9976 63764 10016
rect 63628 9220 63668 9260
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 63820 8884 63860 8924
rect 62860 8632 62900 8672
rect 63052 8632 63092 8672
rect 63916 8632 63956 8672
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 64684 10984 64724 11024
rect 64588 10900 64628 10940
rect 65068 10900 65108 10940
rect 64876 10732 64916 10772
rect 64588 10144 64628 10184
rect 64492 9976 64532 10016
rect 64972 9976 65012 10016
rect 65260 10732 65300 10772
rect 64108 9640 64148 9680
rect 64300 9304 64340 9344
rect 64588 8884 64628 8924
rect 64492 8800 64532 8840
rect 64396 8632 64436 8672
rect 63820 7960 63860 8000
rect 62284 6784 62324 6824
rect 61804 6112 61844 6152
rect 61612 5608 61652 5648
rect 60844 5356 60884 5396
rect 60172 5104 60212 5144
rect 60460 5104 60500 5144
rect 60172 4936 60212 4976
rect 59980 3424 60020 3464
rect 60364 2584 60404 2624
rect 60940 4936 60980 4976
rect 60844 4432 60884 4472
rect 60844 4180 60884 4220
rect 61612 4936 61652 4976
rect 62284 5524 62324 5564
rect 62380 5104 62420 5144
rect 62380 4600 62420 4640
rect 61516 4348 61556 4388
rect 62188 4348 62228 4388
rect 61228 4096 61268 4136
rect 63628 7708 63668 7748
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 63340 6280 63380 6320
rect 62572 5608 62612 5648
rect 62956 5608 62996 5648
rect 62764 4264 62804 4304
rect 62476 3844 62516 3884
rect 62092 3676 62132 3716
rect 60844 3004 60884 3044
rect 61804 3424 61844 3464
rect 59788 2416 59828 2456
rect 61516 2416 61556 2456
rect 60748 1240 60788 1280
rect 61708 1324 61748 1364
rect 62860 3592 62900 3632
rect 62572 1324 62612 1364
rect 62380 1240 62420 1280
rect 63148 5020 63188 5060
rect 64012 7036 64052 7076
rect 64012 6868 64052 6908
rect 64012 6532 64052 6572
rect 63628 6280 63668 6320
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 63724 5860 63764 5900
rect 63436 5608 63476 5648
rect 64204 5692 64244 5732
rect 64396 7960 64436 8000
rect 64588 7960 64628 8000
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 64780 9640 64820 9680
rect 64876 9556 64916 9596
rect 65452 10648 65492 10688
rect 65452 10144 65492 10184
rect 64780 9220 64820 9260
rect 64972 8800 65012 8840
rect 66700 15520 66740 15560
rect 66508 14260 66548 14300
rect 66892 15940 66932 15980
rect 66988 14428 67028 14468
rect 66796 11992 66836 12032
rect 66220 11824 66260 11864
rect 65644 9976 65684 10016
rect 66892 10060 66932 10100
rect 66508 9472 66548 9512
rect 66124 8800 66164 8840
rect 65068 8632 65108 8672
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 64972 8128 65012 8168
rect 65260 8044 65300 8084
rect 65068 7960 65108 8000
rect 65740 8044 65780 8084
rect 64684 7204 64724 7244
rect 64876 7036 64916 7076
rect 65068 7120 65108 7160
rect 64780 6952 64820 6992
rect 64972 6952 65012 6992
rect 65356 7036 65396 7076
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 64588 5776 64628 5816
rect 65068 5776 65108 5816
rect 64492 5692 64532 5732
rect 64396 5608 64436 5648
rect 64300 5188 64340 5228
rect 64012 4768 64052 4808
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 63436 4180 63476 4220
rect 63052 3088 63092 3128
rect 63052 1072 63092 1112
rect 64780 5608 64820 5648
rect 65164 5692 65204 5732
rect 64876 5440 64916 5480
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 66220 7960 66260 8000
rect 65836 7792 65876 7832
rect 65740 7204 65780 7244
rect 66124 7792 66164 7832
rect 66508 8632 66548 8672
rect 66124 7120 66164 7160
rect 65932 6952 65972 6992
rect 65548 5692 65588 5732
rect 65260 5188 65300 5228
rect 64684 5020 64724 5060
rect 64204 4768 64244 4808
rect 64012 3592 64052 3632
rect 63916 3424 63956 3464
rect 64108 3424 64148 3464
rect 64492 4600 64532 4640
rect 65260 4600 65300 4640
rect 64396 4264 64436 4304
rect 64300 3424 64340 3464
rect 64684 4516 64724 4556
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 63820 2584 63860 2624
rect 64588 3424 64628 3464
rect 64492 3088 64532 3128
rect 65836 5440 65876 5480
rect 66220 7036 66260 7076
rect 66028 6448 66068 6488
rect 66124 5692 66164 5732
rect 65932 4936 65972 4976
rect 65740 4768 65780 4808
rect 65836 4264 65876 4304
rect 65644 4180 65684 4220
rect 65260 4012 65300 4052
rect 66700 6952 66740 6992
rect 66412 5692 66452 5732
rect 66316 5608 66356 5648
rect 66604 5608 66644 5648
rect 66892 7036 66932 7076
rect 66892 6448 66932 6488
rect 66220 4516 66260 4556
rect 66124 4432 66164 4472
rect 65932 4012 65972 4052
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 65260 3424 65300 3464
rect 66604 4936 66644 4976
rect 66316 3508 66356 3548
rect 66508 3508 66548 3548
rect 64780 3340 64820 3380
rect 64684 3004 64724 3044
rect 64204 2920 64244 2960
rect 66892 4264 66932 4304
rect 66604 3424 66644 3464
rect 67660 16108 67700 16148
rect 67180 14764 67220 14804
rect 67276 14428 67316 14468
rect 67564 14428 67604 14468
rect 67468 14092 67508 14132
rect 67372 14008 67412 14048
rect 67276 13756 67316 13796
rect 67180 12748 67220 12788
rect 67660 13756 67700 13796
rect 67564 13252 67604 13292
rect 67948 15856 67988 15896
rect 67852 15772 67892 15812
rect 68236 16192 68276 16232
rect 67852 13672 67892 13712
rect 67372 11908 67412 11948
rect 67660 10648 67700 10688
rect 67276 10312 67316 10352
rect 67084 10228 67124 10268
rect 67276 8632 67316 8672
rect 66988 3676 67028 3716
rect 66124 2920 66164 2960
rect 64492 2668 64532 2708
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 64012 1324 64052 1364
rect 64108 1072 64148 1112
rect 61996 988 62036 1028
rect 67660 10228 67700 10268
rect 67852 10312 67892 10352
rect 67756 9136 67796 9176
rect 68140 14176 68180 14216
rect 68044 14092 68084 14132
rect 68524 16024 68564 16064
rect 68908 16192 68948 16232
rect 70156 16192 70196 16232
rect 71404 17116 71444 17156
rect 71655 17116 71695 17156
rect 69772 16108 69812 16148
rect 69388 16024 69428 16064
rect 70540 16024 70580 16064
rect 69292 15940 69332 15980
rect 68812 15520 68852 15560
rect 68716 15436 68756 15476
rect 68716 15268 68756 15308
rect 68620 14008 68660 14048
rect 68908 15268 68948 15308
rect 68908 14680 68948 14720
rect 68812 14092 68852 14132
rect 67948 7120 67988 7160
rect 67852 5860 67892 5900
rect 67660 4852 67700 4892
rect 67756 4684 67796 4724
rect 64780 2668 64820 2708
rect 64684 2584 64724 2624
rect 64876 2584 64916 2624
rect 65260 2584 65300 2624
rect 64684 2416 64724 2456
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 65260 2080 65300 2120
rect 64684 1240 64724 1280
rect 65740 1912 65780 1952
rect 65260 1324 65300 1364
rect 66028 1072 66068 1112
rect 66892 2500 66932 2540
rect 67468 2500 67508 2540
rect 67372 2416 67412 2456
rect 66892 2080 66932 2120
rect 67276 1912 67316 1952
rect 67564 1996 67604 2036
rect 67468 1912 67508 1952
rect 67948 2584 67988 2624
rect 68332 13756 68372 13796
rect 68140 13672 68180 13712
rect 68428 12832 68468 12872
rect 68620 13000 68660 13040
rect 68812 13168 68852 13208
rect 68812 13000 68852 13040
rect 68812 12832 68852 12872
rect 68716 12664 68756 12704
rect 69196 14344 69236 14384
rect 69100 14092 69140 14132
rect 69004 14008 69044 14048
rect 69196 13924 69236 13964
rect 69292 13252 69332 13292
rect 69100 13084 69140 13124
rect 69004 12664 69044 12704
rect 68908 11908 68948 11948
rect 68908 11488 68948 11528
rect 68428 10564 68468 10604
rect 68428 10396 68468 10436
rect 68332 10144 68372 10184
rect 69100 12328 69140 12368
rect 69292 12940 69332 12980
rect 70924 15856 70964 15896
rect 71116 15604 71156 15644
rect 70060 15520 70100 15560
rect 69868 15352 69908 15392
rect 70252 14176 70292 14216
rect 70060 14092 70100 14132
rect 69964 14008 70004 14048
rect 69676 13504 69716 13544
rect 70060 13504 70100 13544
rect 69484 13252 69524 13292
rect 69196 11488 69236 11528
rect 69100 10984 69140 11024
rect 69580 13168 69620 13208
rect 69676 12916 69716 12956
rect 69580 12244 69620 12284
rect 69772 12832 69812 12872
rect 69772 12244 69812 12284
rect 69676 11824 69716 11864
rect 70732 15436 70772 15476
rect 70828 15184 70868 15224
rect 70732 14848 70772 14888
rect 71020 15520 71060 15560
rect 71308 15184 71348 15224
rect 70828 14428 70868 14468
rect 70924 14260 70964 14300
rect 70444 13504 70484 13544
rect 70924 13672 70964 13712
rect 70444 13336 70484 13376
rect 70732 13336 70772 13376
rect 70540 13168 70580 13208
rect 70060 12832 70100 12872
rect 69964 12496 70004 12536
rect 70060 12328 70100 12368
rect 70636 12664 70676 12704
rect 70252 12328 70292 12368
rect 70540 12496 70580 12536
rect 70444 12412 70484 12452
rect 69004 10900 69044 10940
rect 69580 10900 69620 10940
rect 69772 11656 69812 11696
rect 69868 11488 69908 11528
rect 70636 11656 70676 11696
rect 70444 10984 70484 11024
rect 68812 10228 68852 10268
rect 68236 9976 68276 10016
rect 68524 10144 68564 10184
rect 71116 13168 71156 13208
rect 71212 12496 71252 12536
rect 69388 10480 69428 10520
rect 69580 10396 69620 10436
rect 69388 10312 69428 10352
rect 69100 10228 69140 10268
rect 68812 10060 68852 10100
rect 68919 10060 68959 10100
rect 68716 9976 68756 10016
rect 68140 8632 68180 8672
rect 68332 8044 68372 8084
rect 68428 7960 68468 8000
rect 68716 8800 68756 8840
rect 69484 10144 69524 10184
rect 69772 10312 69812 10352
rect 69676 10144 69716 10184
rect 70156 10564 70196 10604
rect 69868 9976 69908 10016
rect 69676 9892 69716 9932
rect 69580 9556 69620 9596
rect 69580 9220 69620 9260
rect 69484 8716 69524 8756
rect 69772 9388 69812 9428
rect 69772 9220 69812 9260
rect 69964 9472 70004 9512
rect 69964 9304 70004 9344
rect 69676 8632 69716 8672
rect 69868 8632 69908 8672
rect 70732 10312 70772 10352
rect 70348 10228 70388 10268
rect 70156 10060 70196 10100
rect 70444 10060 70484 10100
rect 70348 9556 70388 9596
rect 70252 9472 70292 9512
rect 70252 9220 70292 9260
rect 70156 8800 70196 8840
rect 69388 8044 69428 8084
rect 69772 8464 69812 8504
rect 69196 7036 69236 7076
rect 69100 6952 69140 6992
rect 69868 7708 69908 7748
rect 69580 7120 69620 7160
rect 68524 6280 68564 6320
rect 69388 6448 69428 6488
rect 69388 6280 69428 6320
rect 69292 5860 69332 5900
rect 69292 5692 69332 5732
rect 68716 4936 68756 4976
rect 68236 3424 68276 3464
rect 68332 3172 68372 3212
rect 68908 4684 68948 4724
rect 69100 4936 69140 4976
rect 69676 6448 69716 6488
rect 70636 9640 70676 9680
rect 70540 9304 70580 9344
rect 71020 10396 71060 10436
rect 70924 10144 70964 10184
rect 70828 9556 70868 9596
rect 70924 9472 70964 9512
rect 71116 9640 71156 9680
rect 71500 15604 71540 15644
rect 71596 14680 71636 14720
rect 71500 14008 71540 14048
rect 71692 12916 71732 12956
rect 72556 15772 72596 15812
rect 72172 15688 72212 15728
rect 73132 16192 73172 16232
rect 72748 15604 72788 15644
rect 72172 14512 72212 14552
rect 72268 13084 72308 13124
rect 71788 12748 71828 12788
rect 72844 12664 72884 12704
rect 71692 12496 71732 12536
rect 72556 11152 72596 11192
rect 71404 10648 71444 10688
rect 72940 10396 72980 10436
rect 71308 10144 71348 10184
rect 71788 10060 71828 10100
rect 72844 10060 72884 10100
rect 71788 9892 71828 9932
rect 71980 9640 72020 9680
rect 71308 9556 71348 9596
rect 71308 9304 71348 9344
rect 70636 8632 70676 8672
rect 70732 8548 70772 8588
rect 70348 7708 70388 7748
rect 70732 7708 70772 7748
rect 69964 7036 70004 7076
rect 69772 6280 69812 6320
rect 69772 5860 69812 5900
rect 70444 7120 70484 7160
rect 70060 6868 70100 6908
rect 70252 6868 70292 6908
rect 69004 4516 69044 4556
rect 68908 4432 68948 4472
rect 68812 4264 68852 4304
rect 69484 4180 69524 4220
rect 69292 4012 69332 4052
rect 69004 3592 69044 3632
rect 69388 3592 69428 3632
rect 70348 4936 70388 4976
rect 70252 4516 70292 4556
rect 69964 4180 70004 4220
rect 69868 3424 69908 3464
rect 68908 3088 68948 3128
rect 68716 3004 68756 3044
rect 70060 3424 70100 3464
rect 69964 3172 70004 3212
rect 69004 3004 69044 3044
rect 69868 3004 69908 3044
rect 68140 2416 68180 2456
rect 68236 2080 68276 2120
rect 68524 1996 68564 2036
rect 68044 1660 68084 1700
rect 67372 1072 67412 1112
rect 64204 988 64244 1028
rect 69196 2080 69236 2120
rect 69004 1828 69044 1868
rect 70060 1912 70100 1952
rect 70252 1912 70292 1952
rect 70924 8632 70964 8672
rect 70924 7120 70964 7160
rect 70828 5776 70868 5816
rect 70828 3508 70868 3548
rect 70924 1240 70964 1280
rect 69772 1072 69812 1112
rect 71116 8632 71156 8672
rect 71212 8548 71252 8588
rect 71884 9472 71924 9512
rect 71692 9388 71732 9428
rect 71404 8716 71444 8756
rect 71404 8128 71444 8168
rect 71404 7120 71444 7160
rect 71596 7960 71636 8000
rect 71980 9388 72020 9428
rect 71884 8632 71924 8672
rect 71308 7036 71348 7076
rect 71116 4936 71156 4976
rect 71404 5692 71444 5732
rect 71500 5608 71540 5648
rect 71884 7120 71924 7160
rect 71788 7036 71828 7076
rect 71788 5776 71828 5816
rect 71692 5692 71732 5732
rect 74284 15352 74324 15392
rect 73804 14680 73844 14720
rect 73708 14512 73748 14552
rect 73900 14512 73940 14552
rect 74380 14596 74420 14636
rect 74188 14344 74228 14384
rect 74380 14344 74420 14384
rect 73612 13588 73652 13628
rect 73516 12916 73556 12956
rect 73324 12664 73364 12704
rect 73996 10396 74036 10436
rect 73516 9136 73556 9176
rect 73612 8044 73652 8084
rect 72172 7120 72212 7160
rect 72268 5608 72308 5648
rect 71596 4936 71636 4976
rect 71500 4264 71540 4304
rect 71212 3508 71252 3548
rect 71404 3424 71444 3464
rect 71884 4936 71924 4976
rect 71692 4012 71732 4052
rect 71596 3424 71636 3464
rect 72076 5020 72116 5060
rect 72172 4936 72212 4976
rect 72076 3424 72116 3464
rect 72268 4348 72308 4388
rect 72460 4516 72500 4556
rect 72460 4348 72500 4388
rect 71980 3172 72020 3212
rect 71692 3088 71732 3128
rect 71788 3004 71828 3044
rect 71212 2584 71252 2624
rect 71212 2080 71252 2120
rect 73036 7876 73076 7916
rect 73612 5524 73652 5564
rect 72268 2836 72308 2876
rect 71980 2584 72020 2624
rect 72268 2500 72308 2540
rect 71116 1828 71156 1868
rect 71404 1324 71444 1364
rect 72652 2584 72692 2624
rect 72556 2164 72596 2204
rect 72652 1912 72692 1952
rect 72460 1324 72500 1364
rect 72076 1240 72116 1280
rect 71020 1072 71060 1112
rect 71212 1072 71252 1112
rect 71884 1072 71924 1112
rect 72460 1072 72500 1112
rect 72652 1072 72692 1112
rect 72940 2752 72980 2792
rect 73132 2668 73172 2708
rect 73132 2164 73172 2204
rect 73036 2080 73076 2120
rect 74956 16192 74996 16232
rect 75148 15520 75188 15560
rect 74668 15268 74708 15308
rect 74764 14764 74804 14804
rect 74668 14512 74708 14552
rect 74092 9472 74132 9512
rect 75532 14848 75572 14888
rect 75244 14680 75284 14720
rect 75052 14596 75092 14636
rect 74956 14512 74996 14552
rect 74956 14008 74996 14048
rect 74572 13756 74612 13796
rect 74668 13168 74708 13208
rect 74380 13084 74420 13124
rect 74284 13000 74324 13040
rect 75244 14008 75284 14048
rect 74860 13000 74900 13040
rect 74964 13000 75004 13040
rect 74476 12664 74516 12704
rect 74572 12328 74612 12368
rect 74764 12580 74804 12620
rect 75148 13168 75188 13208
rect 75244 13084 75284 13124
rect 75532 14428 75572 14468
rect 76972 16192 77012 16232
rect 76204 14848 76244 14888
rect 75724 14680 75764 14720
rect 76012 14344 76052 14384
rect 75820 13672 75860 13712
rect 75628 13588 75668 13628
rect 75436 13252 75476 13292
rect 75724 13252 75764 13292
rect 75052 12748 75092 12788
rect 74764 12328 74804 12368
rect 75052 11908 75092 11948
rect 74860 11320 74900 11360
rect 74668 10984 74708 11024
rect 75244 12748 75284 12788
rect 75820 13168 75860 13208
rect 76108 12664 76148 12704
rect 75532 12580 75572 12620
rect 75436 11656 75476 11696
rect 75340 11488 75380 11528
rect 75244 11320 75284 11360
rect 75244 11152 75284 11192
rect 74860 10900 74900 10940
rect 74764 10816 74804 10856
rect 74764 10480 74804 10520
rect 74764 10144 74804 10184
rect 74284 5776 74324 5816
rect 75148 10984 75188 11024
rect 75724 11908 75764 11948
rect 75629 11572 75669 11612
rect 76012 11488 76052 11528
rect 75916 11404 75956 11444
rect 75244 10900 75284 10940
rect 75340 10816 75380 10856
rect 75244 9472 75284 9512
rect 75820 10732 75860 10772
rect 76204 11656 76244 11696
rect 77164 14176 77204 14216
rect 76588 13336 76628 13376
rect 76396 12748 76436 12788
rect 77260 13336 77300 13376
rect 77164 13252 77204 13292
rect 76972 13084 77012 13124
rect 76684 12664 76724 12704
rect 76396 11404 76436 11444
rect 76684 11656 76724 11696
rect 77452 13336 77492 13376
rect 77740 16192 77780 16232
rect 77356 12916 77396 12956
rect 77164 11572 77204 11612
rect 76300 11236 76340 11276
rect 76588 11236 76628 11276
rect 75916 10396 75956 10436
rect 76300 10816 76340 10856
rect 75532 9976 75572 10016
rect 76012 9976 76052 10016
rect 75436 8968 75476 9008
rect 75724 9472 75764 9512
rect 75724 9220 75764 9260
rect 75436 7708 75476 7748
rect 75244 7120 75284 7160
rect 76012 9136 76052 9176
rect 75820 8968 75860 9008
rect 75916 8884 75956 8924
rect 75628 8548 75668 8588
rect 75724 7876 75764 7916
rect 75628 7708 75668 7748
rect 75532 7120 75572 7160
rect 75820 7624 75860 7664
rect 75820 7120 75860 7160
rect 76684 10732 76724 10772
rect 76588 10396 76628 10436
rect 76492 10228 76532 10268
rect 76203 9388 76243 9428
rect 76300 8884 76340 8924
rect 76492 9640 76532 9680
rect 76492 9220 76532 9260
rect 77260 11404 77300 11444
rect 77260 10900 77300 10940
rect 76972 10816 77012 10856
rect 76780 9472 76820 9512
rect 76684 9304 76724 9344
rect 76588 8548 76628 8588
rect 76300 8044 76340 8084
rect 76204 7960 76244 8000
rect 76396 7960 76436 8000
rect 76012 7708 76052 7748
rect 76108 7624 76148 7664
rect 76012 7204 76052 7244
rect 73804 3508 73844 3548
rect 74380 4432 74420 4472
rect 74860 4348 74900 4388
rect 74860 3424 74900 3464
rect 76012 6868 76052 6908
rect 76204 6868 76244 6908
rect 76012 5860 76052 5900
rect 75628 5608 75668 5648
rect 76492 7204 76532 7244
rect 76588 6868 76628 6908
rect 76588 5860 76628 5900
rect 76492 5776 76532 5816
rect 76204 5608 76244 5648
rect 76396 5608 76436 5648
rect 75148 4432 75188 4472
rect 75340 4012 75380 4052
rect 76300 5524 76340 5564
rect 76108 5104 76148 5144
rect 76492 5104 76532 5144
rect 76012 4264 76052 4304
rect 75436 3592 75476 3632
rect 75244 3508 75284 3548
rect 74668 3340 74708 3380
rect 73612 2668 73652 2708
rect 74380 2668 74420 2708
rect 73804 2584 73844 2624
rect 74188 2584 74228 2624
rect 74092 2500 74132 2540
rect 73324 1912 73364 1952
rect 73804 1912 73844 1952
rect 74188 2080 74228 2120
rect 73996 1828 74036 1868
rect 73228 1240 73268 1280
rect 74380 1996 74420 2036
rect 74092 1156 74132 1196
rect 73996 1072 74036 1112
rect 74572 1912 74612 1952
rect 75340 3088 75380 3128
rect 75148 2752 75188 2792
rect 75052 2584 75092 2624
rect 75916 4096 75956 4136
rect 75820 3172 75860 3212
rect 75724 3004 75764 3044
rect 75244 2500 75284 2540
rect 75244 1912 75284 1952
rect 75436 1912 75476 1952
rect 75628 1072 75668 1112
rect 76300 4096 76340 4136
rect 76492 4180 76532 4220
rect 76876 8800 76916 8840
rect 77068 9472 77108 9512
rect 78988 17116 79028 17156
rect 77740 10732 77780 10772
rect 77836 10228 77876 10268
rect 77836 10060 77876 10100
rect 77356 9640 77396 9680
rect 77452 9472 77492 9512
rect 77260 9388 77300 9428
rect 77644 9472 77684 9512
rect 77740 9220 77780 9260
rect 76972 8128 77012 8168
rect 77164 7960 77204 8000
rect 77068 7540 77108 7580
rect 77260 7372 77300 7412
rect 77740 8884 77780 8924
rect 77644 8800 77684 8840
rect 77452 8632 77492 8672
rect 77452 8128 77492 8168
rect 77548 7960 77588 8000
rect 77452 7540 77492 7580
rect 77452 7372 77492 7412
rect 77452 7120 77492 7160
rect 77836 8632 77876 8672
rect 77836 7204 77876 7244
rect 78124 12916 78164 12956
rect 78892 16192 78932 16232
rect 79372 17116 79412 17156
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 78604 14512 78644 14552
rect 79655 17116 79695 17156
rect 79180 14512 79220 14552
rect 78700 14176 78740 14216
rect 79372 14176 79412 14216
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 78316 12244 78356 12284
rect 79276 12244 79316 12284
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 78316 11572 78356 11612
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 78316 10144 78356 10184
rect 78028 10060 78068 10100
rect 79468 10060 79508 10100
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 79468 8884 79508 8924
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 77260 5608 77300 5648
rect 77740 5776 77780 5816
rect 76588 4096 76628 4136
rect 76492 3592 76532 3632
rect 76396 3424 76436 3464
rect 76588 3424 76628 3464
rect 76012 2836 76052 2876
rect 75916 1912 75956 1952
rect 77452 4768 77492 4808
rect 77260 4180 77300 4220
rect 77164 4012 77204 4052
rect 76972 3088 77012 3128
rect 76780 2836 76820 2876
rect 77836 4768 77876 4808
rect 77644 4264 77684 4304
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 79468 5776 79508 5816
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 79468 4180 79508 4220
rect 77644 3424 77684 3464
rect 77836 3088 77876 3128
rect 76876 2584 76916 2624
rect 77260 2836 77300 2876
rect 76204 2500 76244 2540
rect 76684 2500 76724 2540
rect 75820 1072 75860 1112
rect 76108 1072 76148 1112
rect 77164 2500 77204 2540
rect 77068 1996 77108 2036
rect 76876 1912 76916 1952
rect 78124 2836 78164 2876
rect 78028 2500 78068 2540
rect 77740 2332 77780 2372
rect 77740 2080 77780 2120
rect 78220 2752 78260 2792
rect 78604 3424 78644 3464
rect 78412 2332 78452 2372
rect 78316 1912 78356 1952
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 79180 2752 79220 2792
rect 77260 1828 77300 1868
rect 78220 1240 78260 1280
rect 78892 1912 78932 1952
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 79468 1240 79508 1280
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 67459 38200 67468 38240
rect 67508 38200 67948 38240
rect 67988 38200 67997 38240
rect 69283 38200 69292 38240
rect 69332 38200 70636 38240
rect 70676 38200 74284 38240
rect 74324 38200 74333 38240
rect 59299 38156 59357 38157
rect 58531 38116 58540 38156
rect 58580 38116 59308 38156
rect 59348 38116 67084 38156
rect 67124 38116 67133 38156
rect 68899 38116 68908 38156
rect 68948 38116 71020 38156
rect 71060 38116 71069 38156
rect 59299 38115 59357 38116
rect 56899 38032 56908 38072
rect 56948 38032 58252 38072
rect 58292 38032 58301 38072
rect 58915 37948 58924 37988
rect 58964 37948 59116 37988
rect 59156 37948 62572 37988
rect 62612 37948 62621 37988
rect 66307 37948 66316 37988
rect 66356 37948 67468 37988
rect 67508 37948 67517 37988
rect 67651 37948 67660 37988
rect 67700 37948 69388 37988
rect 69428 37948 71116 37988
rect 71156 37948 71165 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 73315 37528 73324 37568
rect 73364 37528 74132 37568
rect 0 37508 80 37528
rect 73123 37444 73132 37484
rect 73172 37444 73708 37484
rect 73748 37444 73757 37484
rect 55651 37360 55660 37400
rect 55700 37360 55948 37400
rect 55988 37360 55997 37400
rect 59491 37360 59500 37400
rect 59540 37360 59549 37400
rect 62371 37360 62380 37400
rect 62420 37360 64972 37400
rect 65012 37360 65644 37400
rect 65684 37360 65693 37400
rect 67555 37360 67564 37400
rect 67604 37360 68428 37400
rect 68468 37360 69100 37400
rect 69140 37360 70444 37400
rect 70484 37360 70493 37400
rect 73219 37360 73228 37400
rect 73268 37360 73516 37400
rect 73556 37360 73996 37400
rect 74036 37360 74045 37400
rect 58627 37276 58636 37316
rect 58676 37276 59404 37316
rect 59444 37276 59453 37316
rect 59500 37232 59540 37360
rect 73411 37316 73469 37317
rect 74092 37316 74132 37528
rect 74476 37360 76588 37400
rect 76628 37360 76637 37400
rect 77443 37360 77452 37400
rect 77492 37360 78412 37400
rect 78452 37360 78461 37400
rect 74476 37316 74516 37360
rect 59587 37276 59596 37316
rect 59636 37276 60268 37316
rect 60308 37276 60317 37316
rect 61123 37276 61132 37316
rect 61172 37276 62284 37316
rect 62324 37276 62333 37316
rect 73411 37276 73420 37316
rect 73460 37276 74516 37316
rect 74563 37276 74572 37316
rect 74612 37276 74956 37316
rect 74996 37276 76244 37316
rect 76867 37276 76876 37316
rect 76916 37276 78124 37316
rect 78164 37276 78173 37316
rect 73411 37275 73469 37276
rect 76204 37232 76244 37276
rect 56227 37192 56236 37232
rect 56276 37192 57580 37232
rect 57620 37192 57629 37232
rect 59299 37192 59308 37232
rect 59348 37192 59540 37232
rect 68227 37192 68236 37232
rect 68276 37192 68620 37232
rect 68660 37192 68669 37232
rect 69571 37192 69580 37232
rect 69620 37192 71404 37232
rect 71444 37192 71453 37232
rect 73315 37192 73324 37232
rect 73364 37192 73900 37232
rect 73940 37192 73949 37232
rect 75235 37192 75244 37232
rect 75284 37192 76108 37232
rect 76148 37192 76157 37232
rect 76204 37192 77356 37232
rect 77396 37192 77836 37232
rect 77876 37192 77885 37232
rect 72931 37108 72940 37148
rect 72980 37108 75052 37148
rect 75092 37108 75101 37148
rect 77251 37108 77260 37148
rect 77300 37108 78220 37148
rect 78260 37108 79468 37148
rect 79508 37108 79517 37148
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 67756 37024 73036 37064
rect 73076 37024 75148 37064
rect 75188 37024 75532 37064
rect 75572 37024 75581 37064
rect 58915 36940 58924 36980
rect 58964 36940 61804 36980
rect 61844 36940 61853 36980
rect 67756 36896 67796 37024
rect 73315 36896 73373 36897
rect 58819 36856 58828 36896
rect 58868 36856 58877 36896
rect 60355 36856 60364 36896
rect 60404 36856 61132 36896
rect 61172 36856 62380 36896
rect 62420 36856 62429 36896
rect 67267 36856 67276 36896
rect 67316 36856 67756 36896
rect 67796 36856 67805 36896
rect 70723 36856 70732 36896
rect 70772 36856 73324 36896
rect 73364 36856 73373 36896
rect 58828 36812 58868 36856
rect 73315 36855 73373 36856
rect 54691 36772 54700 36812
rect 54740 36772 55852 36812
rect 55892 36772 55901 36812
rect 57571 36772 57580 36812
rect 57620 36772 58444 36812
rect 58484 36772 58868 36812
rect 61708 36772 63340 36812
rect 63380 36772 63389 36812
rect 63907 36772 63916 36812
rect 63956 36772 63965 36812
rect 68515 36772 68524 36812
rect 68564 36772 69580 36812
rect 69620 36772 71596 36812
rect 71636 36772 71645 36812
rect 76291 36772 76300 36812
rect 76340 36772 76780 36812
rect 76820 36772 77548 36812
rect 77588 36772 77597 36812
rect 0 36728 80 36748
rect 33859 36728 33917 36729
rect 61708 36728 61748 36772
rect 63916 36728 63956 36772
rect 0 36688 33868 36728
rect 33908 36688 33917 36728
rect 55939 36688 55948 36728
rect 55988 36688 56428 36728
rect 56468 36688 57388 36728
rect 57428 36688 57437 36728
rect 58819 36688 58828 36728
rect 58868 36688 58877 36728
rect 60547 36688 60556 36728
rect 60596 36688 61708 36728
rect 61748 36688 61757 36728
rect 62371 36688 62380 36728
rect 62420 36688 63956 36728
rect 64003 36688 64012 36728
rect 64052 36688 65356 36728
rect 65396 36688 65405 36728
rect 67459 36688 67468 36728
rect 67508 36688 68620 36728
rect 68660 36688 68669 36728
rect 68803 36688 68812 36728
rect 68852 36688 69100 36728
rect 69140 36688 69149 36728
rect 70435 36688 70444 36728
rect 70484 36688 72076 36728
rect 72116 36688 74764 36728
rect 74804 36688 76684 36728
rect 76724 36688 78316 36728
rect 78356 36688 78365 36728
rect 0 36668 80 36688
rect 33859 36687 33917 36688
rect 58828 36644 58868 36688
rect 58828 36604 62956 36644
rect 62996 36604 63148 36644
rect 63188 36604 63197 36644
rect 63340 36604 64396 36644
rect 64436 36604 66124 36644
rect 66164 36604 68044 36644
rect 68084 36604 68093 36644
rect 56035 36520 56044 36560
rect 56084 36520 57292 36560
rect 57332 36520 57341 36560
rect 63340 36476 63380 36604
rect 71587 36520 71596 36560
rect 71636 36520 72940 36560
rect 72980 36520 72989 36560
rect 76579 36520 76588 36560
rect 76628 36520 77068 36560
rect 77108 36520 77117 36560
rect 56323 36436 56332 36476
rect 56372 36436 57100 36476
rect 57140 36436 57149 36476
rect 63235 36436 63244 36476
rect 63284 36436 63380 36476
rect 70915 36436 70924 36476
rect 70964 36436 72172 36476
rect 72212 36436 72221 36476
rect 76771 36352 76780 36392
rect 76820 36352 77260 36392
rect 77300 36352 77309 36392
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 59011 36184 59020 36224
rect 59060 36184 59500 36224
rect 59540 36184 59549 36224
rect 66595 36100 66604 36140
rect 66644 36100 67276 36140
rect 67316 36100 67325 36140
rect 49219 36016 49228 36056
rect 49268 36016 50572 36056
rect 50612 36016 50621 36056
rect 58627 36016 58636 36056
rect 58676 36016 59596 36056
rect 59636 36016 59645 36056
rect 64483 36016 64492 36056
rect 64532 36016 65644 36056
rect 65684 36016 67756 36056
rect 67796 36016 68428 36056
rect 68468 36016 68477 36056
rect 69475 36016 69484 36056
rect 69524 36016 70828 36056
rect 70868 36016 70877 36056
rect 72163 36016 72172 36056
rect 72212 36016 73036 36056
rect 73076 36016 73228 36056
rect 73268 36016 73277 36056
rect 75043 36016 75052 36056
rect 75092 36016 75724 36056
rect 75764 36016 75773 36056
rect 50371 35932 50380 35972
rect 50420 35932 50956 35972
rect 50996 35932 51005 35972
rect 53260 35932 57100 35972
rect 57140 35932 57149 35972
rect 59491 35932 59500 35972
rect 59540 35932 61900 35972
rect 61940 35932 61949 35972
rect 67939 35932 67948 35972
rect 67988 35932 70252 35972
rect 70292 35932 70301 35972
rect 71884 35932 74284 35972
rect 74324 35932 74333 35972
rect 74467 35932 74476 35972
rect 74516 35932 76436 35972
rect 0 35828 80 35908
rect 50956 35888 50996 35932
rect 53260 35888 53300 35932
rect 71884 35888 71924 35932
rect 76195 35888 76253 35889
rect 76396 35888 76436 35932
rect 50956 35848 53300 35888
rect 55651 35848 55660 35888
rect 55700 35848 56620 35888
rect 56660 35848 56669 35888
rect 58627 35848 58636 35888
rect 58676 35848 59116 35888
rect 59156 35848 59308 35888
rect 59348 35848 59357 35888
rect 64387 35848 64396 35888
rect 64436 35848 66508 35888
rect 66548 35848 66557 35888
rect 67171 35848 67180 35888
rect 67220 35848 67229 35888
rect 67363 35848 67372 35888
rect 67412 35848 69100 35888
rect 69140 35848 69676 35888
rect 69716 35848 69725 35888
rect 69955 35848 69964 35888
rect 70004 35848 70348 35888
rect 70388 35848 70397 35888
rect 71875 35848 71884 35888
rect 71924 35848 71933 35888
rect 72067 35848 72076 35888
rect 72116 35848 72125 35888
rect 73123 35848 73132 35888
rect 73172 35848 73900 35888
rect 73940 35848 75916 35888
rect 75956 35848 75965 35888
rect 76110 35848 76204 35888
rect 76244 35848 76253 35888
rect 76387 35848 76396 35888
rect 76436 35848 76445 35888
rect 77059 35848 77068 35888
rect 77108 35848 77452 35888
rect 77492 35848 77501 35888
rect 51043 35764 51052 35804
rect 51092 35764 51436 35804
rect 51476 35764 52300 35804
rect 52340 35764 52349 35804
rect 59203 35764 59212 35804
rect 59252 35764 59500 35804
rect 59540 35764 59549 35804
rect 67180 35720 67220 35848
rect 72076 35804 72116 35848
rect 76195 35847 76253 35848
rect 67843 35764 67852 35804
rect 67892 35764 69772 35804
rect 69812 35764 69821 35804
rect 69868 35764 71404 35804
rect 71444 35764 72116 35804
rect 69868 35720 69908 35764
rect 55843 35680 55852 35720
rect 55892 35680 58252 35720
rect 58292 35680 58924 35720
rect 58964 35680 58973 35720
rect 59587 35680 59596 35720
rect 59636 35680 61516 35720
rect 61556 35680 63380 35720
rect 65635 35680 65644 35720
rect 65684 35680 67220 35720
rect 69859 35680 69868 35720
rect 69908 35680 69917 35720
rect 73699 35680 73708 35720
rect 73748 35680 77932 35720
rect 77972 35680 77981 35720
rect 63340 35636 63380 35680
rect 73708 35636 73748 35680
rect 63340 35596 69292 35636
rect 69332 35596 69341 35636
rect 69571 35596 69580 35636
rect 69620 35596 73748 35636
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 55459 35512 55468 35552
rect 55508 35512 56140 35552
rect 56180 35512 56908 35552
rect 56948 35512 56957 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 66019 35512 66028 35552
rect 66068 35512 66700 35552
rect 66740 35512 67084 35552
rect 67124 35512 67133 35552
rect 71683 35512 71692 35552
rect 71732 35512 72652 35552
rect 72692 35512 72701 35552
rect 73219 35512 73228 35552
rect 73268 35512 77068 35552
rect 77108 35512 77117 35552
rect 68227 35428 68236 35468
rect 68276 35428 70924 35468
rect 70964 35428 70973 35468
rect 68131 35344 68140 35384
rect 68180 35344 68189 35384
rect 69955 35344 69964 35384
rect 70004 35344 70444 35384
rect 70484 35344 70493 35384
rect 51523 35260 51532 35300
rect 51572 35260 52780 35300
rect 52820 35260 54508 35300
rect 54548 35260 54557 35300
rect 62851 35216 62909 35217
rect 49699 35176 49708 35216
rect 49748 35176 53356 35216
rect 53396 35176 53405 35216
rect 56035 35176 56044 35216
rect 56084 35176 57196 35216
rect 57236 35176 57772 35216
rect 57812 35176 57821 35216
rect 62766 35176 62860 35216
rect 62900 35176 62909 35216
rect 68140 35216 68180 35344
rect 70339 35260 70348 35300
rect 70388 35260 71308 35300
rect 71348 35260 71357 35300
rect 68140 35176 70444 35216
rect 70484 35176 70493 35216
rect 70627 35176 70636 35216
rect 70676 35176 71788 35216
rect 71828 35176 71837 35216
rect 74179 35176 74188 35216
rect 74228 35176 76012 35216
rect 76052 35176 76061 35216
rect 62851 35175 62909 35176
rect 51811 35092 51820 35132
rect 51860 35092 53740 35132
rect 53780 35092 53789 35132
rect 54787 35092 54796 35132
rect 54836 35092 57484 35132
rect 57524 35092 57964 35132
rect 58004 35092 58828 35132
rect 58868 35092 58877 35132
rect 70243 35092 70252 35132
rect 70292 35092 70540 35132
rect 70580 35092 70589 35132
rect 0 34988 80 35068
rect 52099 35008 52108 35048
rect 52148 35008 55852 35048
rect 55892 35008 55901 35048
rect 61603 35008 61612 35048
rect 61652 35008 61900 35048
rect 61940 35008 65644 35048
rect 65684 35008 65693 35048
rect 61795 34924 61804 34964
rect 61844 34924 61996 34964
rect 62036 34924 62284 34964
rect 62324 34924 62764 34964
rect 62804 34924 62813 34964
rect 66691 34924 66700 34964
rect 66740 34924 67564 34964
rect 67604 34924 69676 34964
rect 69716 34924 74380 34964
rect 74420 34924 74429 34964
rect 54979 34840 54988 34880
rect 55028 34840 56140 34880
rect 56180 34840 57580 34880
rect 57620 34840 64532 34880
rect 65827 34840 65836 34880
rect 65876 34840 67180 34880
rect 67220 34840 67229 34880
rect 67651 34840 67660 34880
rect 67700 34840 67852 34880
rect 67892 34840 67901 34880
rect 68803 34840 68812 34880
rect 68852 34840 69716 34880
rect 69763 34840 69772 34880
rect 69812 34840 70636 34880
rect 70676 34840 70685 34880
rect 64492 34796 64532 34840
rect 69676 34796 69716 34840
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 64492 34756 69580 34796
rect 69620 34756 69629 34796
rect 69676 34756 71500 34796
rect 71540 34756 71549 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 61699 34672 61708 34712
rect 61748 34672 65836 34712
rect 65876 34672 65885 34712
rect 66883 34672 66892 34712
rect 66932 34672 67276 34712
rect 67316 34672 67325 34712
rect 67459 34672 67468 34712
rect 67508 34672 67517 34712
rect 76579 34672 76588 34712
rect 76628 34672 76876 34712
rect 76916 34672 76925 34712
rect 56323 34588 56332 34628
rect 56372 34588 56381 34628
rect 58723 34588 58732 34628
rect 58772 34588 59404 34628
rect 59444 34588 59453 34628
rect 63139 34588 63148 34628
rect 63188 34588 64012 34628
rect 64052 34588 64061 34628
rect 56332 34544 56372 34588
rect 67468 34544 67508 34672
rect 68803 34588 68812 34628
rect 68852 34588 70348 34628
rect 70388 34588 70397 34628
rect 76387 34588 76396 34628
rect 76436 34588 77068 34628
rect 77108 34588 77117 34628
rect 46147 34504 46156 34544
rect 46196 34504 49228 34544
rect 49268 34504 49277 34544
rect 51235 34504 51244 34544
rect 51284 34504 52204 34544
rect 52244 34504 52253 34544
rect 56236 34504 58060 34544
rect 58100 34504 58109 34544
rect 59779 34504 59788 34544
rect 59828 34504 61996 34544
rect 62036 34504 62045 34544
rect 67372 34504 67508 34544
rect 71203 34504 71212 34544
rect 71252 34504 71692 34544
rect 71732 34504 71741 34544
rect 76195 34504 76204 34544
rect 76244 34504 76972 34544
rect 77012 34504 77644 34544
rect 77684 34504 77693 34544
rect 48931 34336 48940 34376
rect 48980 34336 49516 34376
rect 49556 34336 50476 34376
rect 50516 34336 51436 34376
rect 51476 34336 51485 34376
rect 52195 34336 52204 34376
rect 52244 34336 56044 34376
rect 56084 34336 56093 34376
rect 52204 34292 52244 34336
rect 56236 34292 56276 34504
rect 67372 34376 67412 34504
rect 70723 34420 70732 34460
rect 70772 34420 71308 34460
rect 71348 34420 71357 34460
rect 73420 34420 76588 34460
rect 76628 34420 76637 34460
rect 73420 34376 73460 34420
rect 58051 34336 58060 34376
rect 58100 34336 58252 34376
rect 58292 34336 58301 34376
rect 61507 34336 61516 34376
rect 61556 34336 61996 34376
rect 62036 34336 62045 34376
rect 62179 34336 62188 34376
rect 62228 34336 62860 34376
rect 62900 34336 62909 34376
rect 66307 34336 66316 34376
rect 66356 34336 67372 34376
rect 67412 34336 67421 34376
rect 71971 34336 71980 34376
rect 72020 34336 72844 34376
rect 72884 34336 73460 34376
rect 75331 34336 75340 34376
rect 75380 34336 75532 34376
rect 75572 34336 75581 34376
rect 75811 34336 75820 34376
rect 75860 34336 76684 34376
rect 76724 34336 76972 34376
rect 77012 34336 77021 34376
rect 78115 34336 78124 34376
rect 78164 34336 79468 34376
rect 79508 34336 79517 34376
rect 78124 34292 78164 34336
rect 49219 34252 49228 34292
rect 49268 34252 50284 34292
rect 50324 34252 52244 34292
rect 56227 34252 56236 34292
rect 56276 34252 56285 34292
rect 62755 34252 62764 34292
rect 62804 34252 63148 34292
rect 63188 34252 63197 34292
rect 76867 34252 76876 34292
rect 76916 34252 78164 34292
rect 0 34148 80 34228
rect 47011 34168 47020 34208
rect 47060 34168 49036 34208
rect 49076 34168 49085 34208
rect 58627 34168 58636 34208
rect 58676 34168 59596 34208
rect 59636 34168 60364 34208
rect 60404 34168 60413 34208
rect 65731 34168 65740 34208
rect 65780 34168 66796 34208
rect 66836 34168 66845 34208
rect 75523 34168 75532 34208
rect 75572 34168 76012 34208
rect 76052 34168 76061 34208
rect 62755 34124 62813 34125
rect 59491 34084 59500 34124
rect 59540 34084 59980 34124
rect 60020 34084 60029 34124
rect 62179 34084 62188 34124
rect 62228 34084 62764 34124
rect 62804 34084 66124 34124
rect 66164 34084 66173 34124
rect 62755 34083 62813 34084
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 57763 34000 57772 34040
rect 57812 34000 58348 34040
rect 58388 34000 58397 34040
rect 61987 34000 61996 34040
rect 62036 34000 62380 34040
rect 62420 34000 62429 34040
rect 62476 34000 62900 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 71491 34000 71500 34040
rect 71540 34000 71788 34040
rect 71828 34000 71980 34040
rect 72020 34000 72029 34040
rect 58435 33916 58444 33956
rect 58484 33916 61612 33956
rect 61652 33916 61661 33956
rect 62476 33872 62516 34000
rect 62860 33956 62900 34000
rect 62860 33916 69196 33956
rect 69236 33916 69245 33956
rect 70627 33916 70636 33956
rect 70676 33916 71020 33956
rect 71060 33916 71069 33956
rect 76675 33872 76733 33873
rect 54019 33832 54028 33872
rect 54068 33832 54077 33872
rect 54403 33832 54412 33872
rect 54452 33832 62516 33872
rect 62659 33832 62668 33872
rect 62708 33832 62717 33872
rect 65923 33832 65932 33872
rect 65972 33832 65981 33872
rect 76291 33832 76300 33872
rect 76340 33832 76684 33872
rect 76724 33832 76733 33872
rect 54028 33788 54068 33832
rect 51619 33748 51628 33788
rect 51668 33748 53932 33788
rect 53972 33748 53981 33788
rect 54028 33748 54892 33788
rect 54932 33748 55316 33788
rect 58531 33748 58540 33788
rect 58580 33748 60268 33788
rect 60308 33748 61708 33788
rect 61748 33748 61757 33788
rect 55276 33704 55316 33748
rect 49027 33664 49036 33704
rect 49076 33664 49228 33704
rect 49268 33664 49277 33704
rect 54019 33664 54028 33704
rect 54068 33664 54700 33704
rect 54740 33664 54749 33704
rect 55267 33664 55276 33704
rect 55316 33664 55325 33704
rect 59683 33664 59692 33704
rect 59732 33664 60460 33704
rect 60500 33664 61900 33704
rect 61940 33664 62380 33704
rect 62420 33664 62429 33704
rect 62668 33620 62708 33832
rect 62851 33788 62909 33789
rect 62851 33748 62860 33788
rect 62900 33748 65452 33788
rect 65492 33748 65501 33788
rect 62851 33747 62909 33748
rect 63244 33704 63284 33748
rect 65932 33704 65972 33832
rect 76675 33831 76733 33832
rect 75811 33748 75820 33788
rect 75860 33748 77492 33788
rect 76963 33704 77021 33705
rect 77452 33704 77492 33748
rect 63235 33664 63244 33704
rect 63284 33664 63293 33704
rect 65539 33664 65548 33704
rect 65588 33664 66604 33704
rect 66644 33664 66653 33704
rect 69955 33664 69964 33704
rect 70004 33664 72172 33704
rect 72212 33664 72556 33704
rect 72596 33664 72605 33704
rect 76579 33664 76588 33704
rect 76628 33664 76684 33704
rect 76724 33664 76733 33704
rect 76963 33664 76972 33704
rect 77012 33664 77260 33704
rect 77300 33664 77309 33704
rect 77443 33664 77452 33704
rect 77492 33664 78412 33704
rect 78452 33664 78461 33704
rect 76963 33663 77021 33664
rect 71971 33620 72029 33621
rect 62668 33580 63148 33620
rect 63188 33580 63197 33620
rect 71886 33580 71980 33620
rect 72020 33580 72029 33620
rect 71971 33579 72029 33580
rect 52483 33496 52492 33536
rect 52532 33496 53452 33536
rect 53492 33496 54028 33536
rect 54068 33496 54077 33536
rect 59971 33496 59980 33536
rect 60020 33496 63052 33536
rect 63092 33496 66508 33536
rect 66548 33496 66557 33536
rect 71107 33496 71116 33536
rect 71156 33496 71788 33536
rect 71828 33496 74476 33536
rect 74516 33496 76204 33536
rect 76244 33496 76253 33536
rect 77347 33496 77356 33536
rect 77396 33496 78124 33536
rect 78164 33496 78173 33536
rect 48355 33412 48364 33452
rect 48404 33412 49228 33452
rect 49268 33412 49277 33452
rect 50467 33412 50476 33452
rect 50516 33412 51724 33452
rect 51764 33412 55180 33452
rect 55220 33412 55229 33452
rect 58339 33412 58348 33452
rect 58388 33412 58924 33452
rect 58964 33412 58973 33452
rect 74755 33412 74764 33452
rect 74804 33412 76012 33452
rect 76052 33412 76061 33452
rect 76483 33412 76492 33452
rect 76532 33412 76972 33452
rect 77012 33412 77164 33452
rect 77204 33412 77213 33452
rect 0 33308 80 33388
rect 76675 33368 76733 33369
rect 53731 33328 53740 33368
rect 53780 33328 54028 33368
rect 54068 33328 54316 33368
rect 54356 33328 54365 33368
rect 54499 33328 54508 33368
rect 54548 33328 61996 33368
rect 62036 33328 62045 33368
rect 65827 33328 65836 33368
rect 65876 33328 66028 33368
rect 66068 33328 66077 33368
rect 76590 33328 76684 33368
rect 76724 33328 76733 33368
rect 76675 33327 76733 33328
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 58915 33244 58924 33284
rect 58964 33244 59212 33284
rect 59252 33244 59261 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 46819 33160 46828 33200
rect 46868 33160 47020 33200
rect 47060 33160 47069 33200
rect 70627 33116 70685 33117
rect 43180 33076 58156 33116
rect 58196 33076 58205 33116
rect 58636 33076 59020 33116
rect 59060 33076 60940 33116
rect 60980 33076 60989 33116
rect 69091 33076 69100 33116
rect 69140 33076 70636 33116
rect 70676 33076 70685 33116
rect 43180 32948 43220 33076
rect 58636 33032 58676 33076
rect 70627 33075 70685 33076
rect 48739 32992 48748 33032
rect 48788 32992 50764 33032
rect 50804 32992 53644 33032
rect 53684 32992 53693 33032
rect 58627 32992 58636 33032
rect 58676 32992 58685 33032
rect 72643 32992 72652 33032
rect 72692 32992 73036 33032
rect 73076 32992 73085 33032
rect 77155 32992 77164 33032
rect 77204 32992 77740 33032
rect 77780 32992 77789 33032
rect 78115 32992 78124 33032
rect 78164 32992 78508 33032
rect 78548 32992 78557 33032
rect 42211 32908 42220 32948
rect 42260 32908 42700 32948
rect 42740 32908 43220 32948
rect 46051 32908 46060 32948
rect 46100 32908 46252 32948
rect 46292 32908 47788 32948
rect 47828 32908 47837 32948
rect 48643 32908 48652 32948
rect 48692 32908 49036 32948
rect 49076 32908 49085 32948
rect 63235 32908 63244 32948
rect 63284 32908 63293 32948
rect 47107 32824 47116 32864
rect 47156 32824 47884 32864
rect 47924 32824 47933 32864
rect 50563 32824 50572 32864
rect 50612 32824 53548 32864
rect 53588 32824 53597 32864
rect 54499 32824 54508 32864
rect 54548 32824 54796 32864
rect 54836 32824 54845 32864
rect 57571 32824 57580 32864
rect 57620 32824 58252 32864
rect 58292 32824 58301 32864
rect 61891 32824 61900 32864
rect 61940 32824 62476 32864
rect 62516 32824 63148 32864
rect 63188 32824 63197 32864
rect 42115 32656 42124 32696
rect 42164 32656 42892 32696
rect 42932 32656 50380 32696
rect 50420 32656 50429 32696
rect 50572 32612 50612 32824
rect 63244 32780 63284 32908
rect 65635 32824 65644 32864
rect 65684 32824 65932 32864
rect 65972 32824 65981 32864
rect 66691 32824 66700 32864
rect 66740 32824 66988 32864
rect 67028 32824 67037 32864
rect 68995 32824 69004 32864
rect 69044 32824 70924 32864
rect 70964 32824 71500 32864
rect 71540 32824 72460 32864
rect 72500 32824 72509 32864
rect 73411 32824 73420 32864
rect 73460 32824 73612 32864
rect 73652 32824 74860 32864
rect 74900 32824 75436 32864
rect 75476 32824 76012 32864
rect 76052 32824 78220 32864
rect 78260 32824 78269 32864
rect 50755 32740 50764 32780
rect 50804 32740 51244 32780
rect 51284 32740 52204 32780
rect 52244 32740 54412 32780
rect 54452 32740 54461 32780
rect 58147 32740 58156 32780
rect 58196 32740 58540 32780
rect 58580 32740 58589 32780
rect 61315 32740 61324 32780
rect 61364 32740 63916 32780
rect 63956 32740 63965 32780
rect 54595 32656 54604 32696
rect 54644 32656 57676 32696
rect 57716 32656 57725 32696
rect 62947 32656 62956 32696
rect 62996 32656 64108 32696
rect 64148 32656 64157 32696
rect 66211 32656 66220 32696
rect 66260 32656 68716 32696
rect 68756 32656 68908 32696
rect 68948 32656 68957 32696
rect 69091 32656 69100 32696
rect 69140 32656 69772 32696
rect 69812 32656 69821 32696
rect 71779 32656 71788 32696
rect 71828 32656 71980 32696
rect 72020 32656 72029 32696
rect 75139 32656 75148 32696
rect 75188 32656 75916 32696
rect 75956 32656 75965 32696
rect 77731 32656 77740 32696
rect 77780 32656 78028 32696
rect 78068 32656 78077 32696
rect 70915 32612 70973 32613
rect 71788 32612 71828 32656
rect 46435 32572 46444 32612
rect 46484 32572 47308 32612
rect 47348 32572 47357 32612
rect 48835 32572 48844 32612
rect 48884 32572 49324 32612
rect 49364 32572 50612 32612
rect 50659 32572 50668 32612
rect 50708 32572 51052 32612
rect 51092 32572 53548 32612
rect 53588 32572 53597 32612
rect 61987 32572 61996 32612
rect 62036 32572 62572 32612
rect 62612 32572 62621 32612
rect 63331 32572 63340 32612
rect 63380 32572 64588 32612
rect 64628 32572 65644 32612
rect 65684 32572 70924 32612
rect 70964 32572 70973 32612
rect 71107 32572 71116 32612
rect 71156 32572 71828 32612
rect 70915 32571 70973 32572
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 42403 32488 42412 32528
rect 42452 32488 44716 32528
rect 44756 32488 46924 32528
rect 46964 32488 46973 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 60931 32404 60940 32444
rect 60980 32404 68812 32444
rect 68852 32404 68861 32444
rect 49219 32360 49277 32361
rect 49134 32320 49228 32360
rect 49268 32320 49277 32360
rect 49411 32320 49420 32360
rect 49460 32320 50476 32360
rect 50516 32320 50956 32360
rect 50996 32320 51005 32360
rect 54412 32320 54700 32360
rect 54740 32320 54749 32360
rect 63235 32320 63244 32360
rect 63284 32320 64012 32360
rect 64052 32320 64061 32360
rect 70723 32320 70732 32360
rect 70772 32320 71500 32360
rect 71540 32320 71692 32360
rect 71732 32320 71741 32360
rect 76963 32320 76972 32360
rect 77012 32320 77452 32360
rect 77492 32320 77501 32360
rect 49219 32319 49277 32320
rect 44611 32152 44620 32192
rect 44660 32152 45004 32192
rect 45044 32152 47308 32192
rect 47348 32152 47980 32192
rect 48020 32152 48364 32192
rect 48404 32152 49132 32192
rect 49172 32152 49181 32192
rect 50083 32152 50092 32192
rect 50132 32152 51820 32192
rect 51860 32152 51869 32192
rect 53923 32152 53932 32192
rect 53972 32152 54220 32192
rect 54260 32152 54269 32192
rect 54412 32108 54452 32320
rect 54883 32236 54892 32276
rect 54932 32236 55372 32276
rect 55412 32236 56332 32276
rect 56372 32236 56381 32276
rect 59779 32236 59788 32276
rect 59828 32236 59868 32276
rect 62563 32236 62572 32276
rect 62612 32236 62956 32276
rect 62996 32236 63005 32276
rect 63427 32236 63436 32276
rect 63476 32236 64300 32276
rect 64340 32236 64349 32276
rect 70531 32236 70540 32276
rect 70580 32236 71020 32276
rect 71060 32236 71069 32276
rect 71971 32236 71980 32276
rect 72020 32236 72748 32276
rect 72788 32236 73900 32276
rect 73940 32236 74572 32276
rect 74612 32236 74621 32276
rect 55651 32192 55709 32193
rect 59788 32192 59828 32236
rect 54499 32152 54508 32192
rect 54548 32152 54988 32192
rect 55028 32152 55276 32192
rect 55316 32152 55325 32192
rect 55566 32152 55660 32192
rect 55700 32152 56812 32192
rect 56852 32152 56861 32192
rect 59107 32152 59116 32192
rect 59156 32152 59308 32192
rect 59348 32152 61612 32192
rect 61652 32152 61804 32192
rect 61844 32152 64492 32192
rect 64532 32152 64541 32192
rect 65251 32152 65260 32192
rect 65300 32152 65836 32192
rect 65876 32152 65885 32192
rect 66307 32152 66316 32192
rect 66356 32152 66700 32192
rect 66740 32152 66749 32192
rect 67939 32152 67948 32192
rect 67988 32152 69004 32192
rect 69044 32152 69484 32192
rect 69524 32152 70636 32192
rect 70676 32152 72940 32192
rect 72980 32152 73612 32192
rect 73652 32152 73661 32192
rect 75811 32152 75820 32192
rect 75860 32152 76588 32192
rect 76628 32152 76637 32192
rect 55651 32151 55709 32152
rect 70627 32108 70685 32109
rect 75820 32108 75860 32152
rect 48931 32068 48940 32108
rect 48980 32068 49996 32108
rect 50036 32068 50045 32108
rect 54403 32068 54412 32108
rect 54452 32068 54461 32108
rect 62755 32068 62764 32108
rect 62804 32068 63244 32108
rect 63284 32068 63293 32108
rect 69283 32068 69292 32108
rect 69332 32068 70636 32108
rect 70676 32068 70732 32108
rect 70772 32068 75860 32108
rect 70627 32067 70685 32068
rect 48739 31984 48748 32024
rect 48788 31984 49364 32024
rect 58243 31984 58252 32024
rect 58292 31984 59308 32024
rect 59348 31984 59357 32024
rect 69379 31984 69388 32024
rect 69428 31984 70060 32024
rect 70100 31984 70109 32024
rect 71971 31984 71980 32024
rect 72020 31984 72460 32024
rect 72500 31984 72509 32024
rect 73420 31984 76684 32024
rect 76724 31984 77164 32024
rect 77204 31984 78412 32024
rect 78452 31984 78461 32024
rect 49324 31940 49364 31984
rect 73420 31940 73460 31984
rect 46819 31900 46828 31940
rect 46868 31900 48460 31940
rect 48500 31900 48980 31940
rect 49324 31900 49612 31940
rect 49652 31900 49661 31940
rect 54403 31900 54412 31940
rect 54452 31900 54988 31940
rect 55028 31900 55037 31940
rect 59875 31900 59884 31940
rect 59924 31900 60748 31940
rect 60788 31900 60797 31940
rect 65443 31900 65452 31940
rect 65492 31900 70252 31940
rect 70292 31900 70301 31940
rect 71203 31900 71212 31940
rect 71252 31900 73036 31940
rect 73076 31900 73460 31940
rect 78019 31900 78028 31940
rect 78068 31900 79468 31940
rect 79508 31900 79517 31940
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 46339 31732 46348 31772
rect 46388 31732 46397 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 0 31628 80 31708
rect 46348 31688 46388 31732
rect 44803 31648 44812 31688
rect 44852 31648 46388 31688
rect 48940 31688 48980 31900
rect 49219 31816 49228 31856
rect 49268 31816 49516 31856
rect 49556 31816 49565 31856
rect 53539 31816 53548 31856
rect 53588 31816 62284 31856
rect 62324 31816 62333 31856
rect 63139 31816 63148 31856
rect 63188 31816 64108 31856
rect 64148 31816 64157 31856
rect 56035 31772 56093 31773
rect 71011 31772 71069 31773
rect 49987 31732 49996 31772
rect 50036 31732 50476 31772
rect 50516 31732 50860 31772
rect 50900 31732 50909 31772
rect 55939 31732 55948 31772
rect 55988 31732 56044 31772
rect 56084 31732 58348 31772
rect 58388 31732 58397 31772
rect 59299 31732 59308 31772
rect 59348 31732 59788 31772
rect 59828 31732 59837 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 71011 31732 71020 31772
rect 71060 31732 71404 31772
rect 71444 31732 71692 31772
rect 71732 31732 71741 31772
rect 76003 31732 76012 31772
rect 76052 31732 76061 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 56035 31731 56093 31732
rect 71011 31731 71069 31732
rect 71875 31688 71933 31689
rect 48940 31648 53300 31688
rect 63043 31648 63052 31688
rect 63092 31648 63132 31688
rect 66316 31648 66892 31688
rect 66932 31648 66941 31688
rect 71790 31648 71884 31688
rect 71924 31648 71933 31688
rect 76012 31688 76052 31732
rect 76012 31648 76876 31688
rect 76916 31648 77492 31688
rect 49219 31604 49277 31605
rect 46147 31564 46156 31604
rect 46196 31564 46732 31604
rect 46772 31564 46781 31604
rect 49027 31564 49036 31604
rect 49076 31564 49228 31604
rect 49268 31564 49277 31604
rect 53260 31604 53300 31648
rect 63052 31604 63092 31648
rect 53260 31564 57196 31604
rect 57236 31564 57245 31604
rect 59395 31564 59404 31604
rect 59444 31564 60844 31604
rect 60884 31564 65644 31604
rect 65684 31564 65693 31604
rect 49219 31563 49277 31564
rect 60067 31480 60076 31520
rect 60116 31480 61996 31520
rect 62036 31480 62045 31520
rect 66316 31436 66356 31648
rect 71875 31647 71933 31648
rect 71395 31604 71453 31605
rect 71971 31604 72029 31605
rect 76963 31604 77021 31605
rect 71310 31564 71404 31604
rect 71444 31564 71453 31604
rect 71952 31564 71980 31604
rect 72020 31564 72076 31604
rect 72116 31564 76972 31604
rect 77012 31564 77021 31604
rect 71395 31563 71453 31564
rect 71971 31563 72029 31564
rect 76963 31563 77021 31564
rect 70723 31480 70732 31520
rect 70772 31480 71116 31520
rect 71156 31480 71596 31520
rect 71636 31480 71645 31520
rect 75907 31480 75916 31520
rect 75956 31480 76972 31520
rect 77012 31480 77021 31520
rect 60643 31396 60652 31436
rect 60692 31396 65356 31436
rect 65396 31396 65405 31436
rect 65731 31396 65740 31436
rect 65780 31396 66316 31436
rect 66356 31396 66365 31436
rect 71971 31352 72029 31353
rect 77452 31352 77492 31648
rect 41443 31312 41452 31352
rect 41492 31312 45004 31352
rect 45044 31312 45053 31352
rect 46627 31312 46636 31352
rect 46676 31312 47212 31352
rect 47252 31312 49036 31352
rect 49076 31312 49085 31352
rect 49219 31312 49228 31352
rect 49268 31312 49708 31352
rect 49748 31312 50092 31352
rect 50132 31312 50141 31352
rect 50371 31312 50380 31352
rect 50420 31312 50860 31352
rect 50900 31312 50909 31352
rect 52387 31312 52396 31352
rect 52436 31312 54124 31352
rect 54164 31312 56620 31352
rect 56660 31312 57388 31352
rect 57428 31312 57580 31352
rect 57620 31312 59116 31352
rect 59156 31312 59165 31352
rect 59779 31312 59788 31352
rect 59828 31312 61900 31352
rect 61940 31312 63148 31352
rect 63188 31312 63197 31352
rect 66211 31312 66220 31352
rect 66260 31312 66988 31352
rect 67028 31312 69100 31352
rect 69140 31312 69149 31352
rect 71395 31312 71404 31352
rect 71444 31312 71980 31352
rect 72020 31312 72029 31352
rect 77443 31312 77452 31352
rect 77492 31312 77836 31352
rect 77876 31312 77885 31352
rect 71971 31311 72029 31312
rect 62755 31268 62813 31269
rect 75523 31268 75581 31269
rect 42883 31228 42892 31268
rect 42932 31228 43220 31268
rect 43459 31228 43468 31268
rect 43508 31228 50188 31268
rect 50228 31228 50237 31268
rect 60355 31228 60364 31268
rect 60404 31228 62572 31268
rect 62612 31228 62621 31268
rect 62755 31228 62764 31268
rect 62804 31228 63051 31268
rect 63091 31228 63100 31268
rect 75438 31228 75532 31268
rect 75572 31228 75581 31268
rect 43180 31184 43220 31228
rect 62755 31227 62813 31228
rect 75523 31227 75581 31228
rect 42307 31144 42316 31184
rect 42356 31144 42604 31184
rect 42644 31144 43084 31184
rect 43124 31144 43133 31184
rect 43180 31144 43852 31184
rect 43892 31144 43901 31184
rect 49507 31144 49516 31184
rect 49556 31144 49708 31184
rect 49748 31144 49757 31184
rect 49891 31144 49900 31184
rect 49940 31144 50476 31184
rect 50516 31144 50764 31184
rect 50804 31144 50813 31184
rect 55267 31144 55276 31184
rect 55316 31144 55564 31184
rect 55604 31144 55613 31184
rect 55747 31144 55756 31184
rect 55796 31144 56140 31184
rect 56180 31144 56189 31184
rect 59875 31144 59884 31184
rect 59924 31144 60556 31184
rect 60596 31144 60605 31184
rect 61027 31144 61036 31184
rect 61076 31144 63244 31184
rect 63284 31144 63293 31184
rect 69091 31144 69100 31184
rect 69140 31144 74572 31184
rect 74612 31144 74621 31184
rect 71395 31100 71453 31101
rect 41059 31060 41068 31100
rect 41108 31060 43468 31100
rect 43508 31060 43517 31100
rect 59683 31060 59692 31100
rect 59732 31060 60268 31100
rect 60308 31060 60317 31100
rect 70723 31060 70732 31100
rect 70772 31060 71020 31100
rect 71060 31060 71069 31100
rect 71395 31060 71404 31100
rect 71444 31060 71692 31100
rect 71732 31060 71741 31100
rect 76483 31060 76492 31100
rect 76532 31060 77644 31100
rect 77684 31060 77693 31100
rect 71395 31059 71453 31060
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 42499 30976 42508 31016
rect 42548 30976 44812 31016
rect 44852 30976 44861 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 55939 30976 55948 31016
rect 55988 30976 56140 31016
rect 56180 30976 56189 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 71587 30976 71596 31016
rect 71636 30976 73228 31016
rect 73268 30976 73277 31016
rect 74851 30976 74860 31016
rect 74900 30976 75380 31016
rect 75340 30932 75380 30976
rect 77164 30976 77452 31016
rect 77492 30976 77501 31016
rect 43171 30892 43180 30932
rect 43220 30892 45772 30932
rect 45812 30892 59020 30932
rect 59060 30892 59069 30932
rect 75331 30892 75340 30932
rect 75380 30892 75389 30932
rect 75523 30892 75532 30932
rect 75572 30892 77068 30932
rect 77108 30892 77117 30932
rect 0 30788 80 30868
rect 54787 30848 54845 30849
rect 40195 30808 40204 30848
rect 40244 30808 42796 30848
rect 42836 30808 42845 30848
rect 50563 30808 50572 30848
rect 50612 30808 51532 30848
rect 51572 30808 51581 30848
rect 54702 30808 54796 30848
rect 54836 30808 54845 30848
rect 57955 30808 57964 30848
rect 58004 30808 59596 30848
rect 59636 30808 60076 30848
rect 60116 30808 60125 30848
rect 70531 30808 70540 30848
rect 70580 30808 70828 30848
rect 70868 30808 70877 30848
rect 71299 30808 71308 30848
rect 71348 30808 71500 30848
rect 71540 30808 71549 30848
rect 73603 30808 73612 30848
rect 73652 30808 75436 30848
rect 75476 30808 75485 30848
rect 54787 30807 54845 30808
rect 40204 30724 41644 30764
rect 41684 30724 43372 30764
rect 43412 30724 43988 30764
rect 57667 30724 57676 30764
rect 57716 30724 62476 30764
rect 62516 30724 62525 30764
rect 68227 30724 68236 30764
rect 68276 30724 70636 30764
rect 70676 30724 70685 30764
rect 74956 30724 76300 30764
rect 76340 30724 76349 30764
rect 40204 30680 40244 30724
rect 43948 30680 43988 30724
rect 74956 30680 74996 30724
rect 77164 30680 77204 30976
rect 77635 30808 77644 30848
rect 77684 30808 77836 30848
rect 77876 30808 79468 30848
rect 79508 30808 79517 30848
rect 40195 30640 40204 30680
rect 40244 30640 40253 30680
rect 41731 30640 41740 30680
rect 41780 30640 42604 30680
rect 42644 30640 42653 30680
rect 43180 30640 43756 30680
rect 43796 30640 43805 30680
rect 43939 30640 43948 30680
rect 43988 30640 47212 30680
rect 47252 30640 47261 30680
rect 49315 30640 49324 30680
rect 49364 30640 49804 30680
rect 49844 30640 49853 30680
rect 50467 30640 50476 30680
rect 50516 30640 51244 30680
rect 51284 30640 51293 30680
rect 54787 30640 54796 30680
rect 54836 30640 55852 30680
rect 55892 30640 55901 30680
rect 58627 30640 58636 30680
rect 58676 30640 59980 30680
rect 60020 30640 60029 30680
rect 60172 30640 61036 30680
rect 61076 30640 61085 30680
rect 64675 30640 64684 30680
rect 64724 30640 66028 30680
rect 66068 30640 66077 30680
rect 70531 30640 70540 30680
rect 70580 30640 71020 30680
rect 71060 30640 74764 30680
rect 74804 30640 74813 30680
rect 74947 30640 74956 30680
rect 74996 30640 75005 30680
rect 75139 30640 75148 30680
rect 75188 30640 76012 30680
rect 76052 30640 76588 30680
rect 76628 30640 76637 30680
rect 77155 30640 77164 30680
rect 77204 30640 77213 30680
rect 40867 30596 40925 30597
rect 43180 30596 43220 30640
rect 60172 30596 60212 30640
rect 63235 30596 63293 30597
rect 40782 30556 40876 30596
rect 40916 30556 40925 30596
rect 41443 30556 41452 30596
rect 41492 30556 41501 30596
rect 42115 30556 42124 30596
rect 42164 30556 42316 30596
rect 42356 30556 42365 30596
rect 42412 30556 43220 30596
rect 59587 30556 59596 30596
rect 59636 30556 60212 30596
rect 60259 30556 60268 30596
rect 60308 30556 63244 30596
rect 63284 30556 63293 30596
rect 66028 30596 66068 30640
rect 77155 30596 77213 30597
rect 66028 30556 71308 30596
rect 71348 30556 77164 30596
rect 77204 30556 77213 30596
rect 40867 30555 40925 30556
rect 41452 30512 41492 30556
rect 42412 30512 42452 30556
rect 63235 30555 63293 30556
rect 77155 30555 77213 30556
rect 71875 30512 71933 30513
rect 41452 30472 41644 30512
rect 41684 30472 42452 30512
rect 42979 30472 42988 30512
rect 43028 30472 43756 30512
rect 43796 30472 43805 30512
rect 52867 30472 52876 30512
rect 52916 30472 54604 30512
rect 54644 30472 54653 30512
rect 71011 30472 71020 30512
rect 71060 30472 71884 30512
rect 71924 30472 71933 30512
rect 74851 30472 74860 30512
rect 74900 30472 75052 30512
rect 75092 30472 75436 30512
rect 75476 30472 76396 30512
rect 76436 30472 76445 30512
rect 77539 30472 77548 30512
rect 77588 30472 78028 30512
rect 78068 30472 78077 30512
rect 71875 30471 71933 30472
rect 62755 30428 62813 30429
rect 40771 30388 40780 30428
rect 40820 30388 42508 30428
rect 42548 30388 42557 30428
rect 50371 30388 50380 30428
rect 50420 30388 54028 30428
rect 54068 30388 55180 30428
rect 55220 30388 55229 30428
rect 60259 30388 60268 30428
rect 60308 30388 61132 30428
rect 61172 30388 61181 30428
rect 62755 30388 62764 30428
rect 62804 30388 62860 30428
rect 62900 30388 62909 30428
rect 70435 30388 70444 30428
rect 70484 30388 70924 30428
rect 70964 30388 74956 30428
rect 74996 30388 75005 30428
rect 75907 30388 75916 30428
rect 75956 30388 76204 30428
rect 76244 30388 76253 30428
rect 62755 30387 62813 30388
rect 51427 30344 51485 30345
rect 75523 30344 75581 30345
rect 42211 30304 42220 30344
rect 42260 30304 42796 30344
rect 42836 30304 42845 30344
rect 46339 30304 46348 30344
rect 46388 30304 47116 30344
rect 47156 30304 47165 30344
rect 50179 30304 50188 30344
rect 50228 30304 51436 30344
rect 51476 30304 51485 30344
rect 55459 30304 55468 30344
rect 55508 30304 56236 30344
rect 56276 30304 58540 30344
rect 58580 30304 66604 30344
rect 66644 30304 66653 30344
rect 75523 30304 75532 30344
rect 75572 30304 76300 30344
rect 76340 30304 76349 30344
rect 51427 30303 51485 30304
rect 75523 30303 75581 30304
rect 76963 30260 77021 30261
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 39715 30220 39724 30260
rect 39764 30220 40204 30260
rect 40244 30220 40253 30260
rect 44707 30220 44716 30260
rect 44756 30220 45004 30260
rect 45044 30220 45053 30260
rect 45955 30220 45964 30260
rect 46004 30220 46924 30260
rect 46964 30220 46973 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 50659 30220 50668 30260
rect 50708 30220 50956 30260
rect 50996 30220 51005 30260
rect 54691 30220 54700 30260
rect 54740 30220 54988 30260
rect 55028 30220 55037 30260
rect 60931 30220 60940 30260
rect 60980 30220 61420 30260
rect 61460 30220 61469 30260
rect 63043 30220 63052 30260
rect 63092 30220 63436 30260
rect 63476 30220 63485 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 71779 30220 71788 30260
rect 71828 30220 72172 30260
rect 72212 30220 72221 30260
rect 74947 30220 74956 30260
rect 74996 30220 75340 30260
rect 75380 30220 75389 30260
rect 75523 30220 75532 30260
rect 75572 30220 75724 30260
rect 75764 30220 75773 30260
rect 76878 30220 76972 30260
rect 77012 30220 77021 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 76963 30219 77021 30220
rect 55267 30176 55325 30177
rect 46051 30136 46060 30176
rect 46100 30136 46252 30176
rect 46292 30136 46301 30176
rect 51523 30136 51532 30176
rect 51572 30136 55084 30176
rect 55124 30136 55276 30176
rect 55316 30136 55325 30176
rect 63331 30136 63340 30176
rect 63380 30136 65452 30176
rect 65492 30136 65501 30176
rect 55267 30135 55325 30136
rect 55075 30092 55133 30093
rect 44611 30052 44620 30092
rect 44660 30052 45868 30092
rect 45908 30052 46348 30092
rect 46388 30052 46397 30092
rect 51427 30052 51436 30092
rect 51476 30052 55084 30092
rect 55124 30052 55133 30092
rect 59971 30052 59980 30092
rect 60020 30052 61228 30092
rect 61268 30052 62956 30092
rect 62996 30052 63005 30092
rect 69667 30052 69676 30092
rect 69716 30052 71692 30092
rect 71732 30052 71741 30092
rect 55075 30051 55133 30052
rect 0 29948 80 30028
rect 42115 29968 42124 30008
rect 42164 29968 43852 30008
rect 43892 29968 43901 30008
rect 51043 29968 51052 30008
rect 51092 29968 51340 30008
rect 51380 29968 51389 30008
rect 55555 29968 55564 30008
rect 55604 29968 56044 30008
rect 56084 29968 56093 30008
rect 60355 29968 60364 30008
rect 60404 29968 60748 30008
rect 60788 29968 60797 30008
rect 71107 29968 71116 30008
rect 71156 29968 72268 30008
rect 72308 29968 73708 30008
rect 73748 29968 74092 30008
rect 74132 29968 74141 30008
rect 55075 29924 55133 29925
rect 50371 29884 50380 29924
rect 50420 29884 51724 29924
rect 51764 29884 51773 29924
rect 53260 29884 54796 29924
rect 54836 29884 54845 29924
rect 55075 29884 55084 29924
rect 55124 29884 55852 29924
rect 55892 29884 55901 29924
rect 58819 29884 58828 29924
rect 58868 29884 59692 29924
rect 59732 29884 64012 29924
rect 64052 29884 64061 29924
rect 71491 29884 71500 29924
rect 71540 29884 71884 29924
rect 71924 29884 75052 29924
rect 75092 29884 75101 29924
rect 40003 29800 40012 29840
rect 40052 29800 40684 29840
rect 40724 29800 42412 29840
rect 42452 29800 42461 29840
rect 47587 29800 47596 29840
rect 47636 29800 48364 29840
rect 48404 29800 49036 29840
rect 49076 29800 52492 29840
rect 52532 29800 52541 29840
rect 41347 29716 41356 29756
rect 41396 29716 41836 29756
rect 41876 29716 43084 29756
rect 43124 29716 43220 29756
rect 46435 29716 46444 29756
rect 46484 29716 47212 29756
rect 47252 29716 47261 29756
rect 51043 29716 51052 29756
rect 51092 29716 51436 29756
rect 51476 29716 51485 29756
rect 41539 29632 41548 29672
rect 41588 29632 41740 29672
rect 41780 29632 41789 29672
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 43180 29252 43220 29716
rect 53260 29672 53300 29884
rect 55075 29883 55133 29884
rect 54691 29800 54700 29840
rect 54740 29800 55084 29840
rect 55124 29800 56236 29840
rect 56276 29800 56285 29840
rect 63148 29800 63628 29840
rect 63668 29800 63677 29840
rect 63811 29800 63820 29840
rect 63860 29800 65740 29840
rect 65780 29800 65789 29840
rect 69283 29800 69292 29840
rect 69332 29800 69484 29840
rect 69524 29800 69533 29840
rect 69763 29800 69772 29840
rect 69812 29800 70636 29840
rect 70676 29800 71020 29840
rect 71060 29800 71069 29840
rect 75523 29800 75532 29840
rect 75572 29800 76012 29840
rect 76052 29800 76061 29840
rect 63148 29756 63188 29800
rect 63139 29716 63148 29756
rect 63188 29716 63197 29756
rect 64579 29716 64588 29756
rect 64628 29716 65164 29756
rect 65204 29716 65213 29756
rect 69571 29716 69580 29756
rect 69620 29716 69964 29756
rect 70004 29716 70013 29756
rect 74851 29716 74860 29756
rect 74900 29716 75916 29756
rect 75956 29716 77164 29756
rect 77204 29716 77213 29756
rect 55651 29672 55709 29673
rect 56035 29672 56093 29673
rect 49123 29632 49132 29672
rect 49172 29632 49420 29672
rect 49460 29632 50572 29672
rect 50612 29632 53300 29672
rect 55566 29632 55660 29672
rect 55700 29632 55709 29672
rect 55950 29632 56044 29672
rect 56084 29632 56093 29672
rect 55651 29631 55709 29632
rect 56035 29631 56093 29632
rect 63235 29672 63293 29673
rect 63235 29632 63244 29672
rect 63284 29632 63340 29672
rect 63380 29632 63408 29672
rect 65443 29632 65452 29672
rect 65492 29632 66220 29672
rect 66260 29632 68428 29672
rect 68468 29632 68477 29672
rect 63235 29631 63293 29632
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 50275 29464 50284 29504
rect 50324 29464 50333 29504
rect 50947 29464 50956 29504
rect 50996 29464 51244 29504
rect 51284 29464 51293 29504
rect 59395 29464 59404 29504
rect 59444 29464 60172 29504
rect 60212 29464 60221 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 69955 29464 69964 29504
rect 70004 29464 70348 29504
rect 70388 29464 70397 29504
rect 70819 29464 70828 29504
rect 70868 29464 71404 29504
rect 71444 29464 73460 29504
rect 76003 29464 76012 29504
rect 76052 29464 76492 29504
rect 76532 29464 76541 29504
rect 50284 29336 50324 29464
rect 73420 29336 73460 29464
rect 43459 29296 43468 29336
rect 43508 29296 45004 29336
rect 45044 29296 45053 29336
rect 49507 29296 49516 29336
rect 49556 29296 49804 29336
rect 49844 29296 49853 29336
rect 50083 29296 50092 29336
rect 50132 29296 50324 29336
rect 59875 29296 59884 29336
rect 59924 29296 59964 29336
rect 73420 29296 76204 29336
rect 76244 29296 76253 29336
rect 59884 29252 59924 29296
rect 43180 29212 46156 29252
rect 46196 29212 51052 29252
rect 51092 29212 51101 29252
rect 51532 29212 53644 29252
rect 53684 29212 54028 29252
rect 54068 29212 54077 29252
rect 54124 29212 54316 29252
rect 54356 29212 54365 29252
rect 55939 29212 55948 29252
rect 55988 29212 56332 29252
rect 56372 29212 56381 29252
rect 59107 29212 59116 29252
rect 59156 29212 63380 29252
rect 67747 29212 67756 29252
rect 67796 29212 70156 29252
rect 70196 29212 70205 29252
rect 0 29108 80 29188
rect 40771 29128 40780 29168
rect 40820 29128 41452 29168
rect 41492 29128 41501 29168
rect 45091 29128 45100 29168
rect 45140 29128 46060 29168
rect 46100 29128 46109 29168
rect 49699 29128 49708 29168
rect 49748 29128 50860 29168
rect 50900 29128 50909 29168
rect 51532 29084 51572 29212
rect 54124 29168 54164 29212
rect 63340 29168 63380 29212
rect 51811 29128 51820 29168
rect 51860 29128 54164 29168
rect 54211 29128 54220 29168
rect 54260 29128 55180 29168
rect 55220 29128 55229 29168
rect 55363 29128 55372 29168
rect 55412 29128 55852 29168
rect 55892 29128 55901 29168
rect 60355 29128 60364 29168
rect 60404 29128 60844 29168
rect 60884 29128 60893 29168
rect 63340 29128 63532 29168
rect 63572 29128 63581 29168
rect 63907 29128 63916 29168
rect 63956 29128 64204 29168
rect 64244 29128 64253 29168
rect 69763 29128 69772 29168
rect 69812 29128 70540 29168
rect 70580 29128 70589 29168
rect 54220 29084 54260 29128
rect 50371 29044 50380 29084
rect 50420 29044 51340 29084
rect 51380 29044 51572 29084
rect 52483 29044 52492 29084
rect 52532 29044 54260 29084
rect 60547 29044 60556 29084
rect 60596 29044 61132 29084
rect 61172 29044 61181 29084
rect 63427 29044 63436 29084
rect 63476 29044 64012 29084
rect 64052 29044 64061 29084
rect 64963 29044 64972 29084
rect 65012 29044 65356 29084
rect 65396 29044 65548 29084
rect 65588 29044 65597 29084
rect 68419 29044 68428 29084
rect 68468 29044 69044 29084
rect 70147 29044 70156 29084
rect 70196 29044 70636 29084
rect 70676 29044 70685 29084
rect 71011 29044 71020 29084
rect 71060 29044 71596 29084
rect 71636 29044 71645 29084
rect 69004 29000 69044 29044
rect 71107 29000 71165 29001
rect 41059 28960 41068 29000
rect 41108 28960 41260 29000
rect 41300 28960 42028 29000
rect 42068 28960 42077 29000
rect 47779 28960 47788 29000
rect 47828 28960 49516 29000
rect 49556 28960 49565 29000
rect 50275 28960 50284 29000
rect 50324 28960 51724 29000
rect 51764 28960 53932 29000
rect 53972 28960 55084 29000
rect 55124 28960 55133 29000
rect 55564 28960 61076 29000
rect 62947 28960 62956 29000
rect 62996 28960 68908 29000
rect 68948 28960 68957 29000
rect 69004 28960 71116 29000
rect 71156 28960 71165 29000
rect 55564 28916 55604 28960
rect 41740 28876 42220 28916
rect 42260 28876 42269 28916
rect 47203 28876 47212 28916
rect 47252 28876 48748 28916
rect 48788 28876 55604 28916
rect 55651 28876 55660 28916
rect 55700 28876 55709 28916
rect 41740 28832 41780 28876
rect 41731 28792 41740 28832
rect 41780 28792 41789 28832
rect 49603 28792 49612 28832
rect 49652 28792 50572 28832
rect 50612 28792 50956 28832
rect 50996 28792 51005 28832
rect 54691 28792 54700 28832
rect 54740 28792 55564 28832
rect 55604 28792 55613 28832
rect 54787 28748 54845 28749
rect 55660 28748 55700 28876
rect 61036 28832 61076 28960
rect 71107 28959 71165 28960
rect 70339 28876 70348 28916
rect 70388 28876 70828 28916
rect 70868 28876 70877 28916
rect 61027 28792 61036 28832
rect 61076 28792 61085 28832
rect 70051 28792 70060 28832
rect 70100 28792 71212 28832
rect 71252 28792 71261 28832
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 40003 28708 40012 28748
rect 40052 28708 42316 28748
rect 42356 28708 42365 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 50467 28708 50476 28748
rect 50516 28708 54796 28748
rect 54836 28708 55948 28748
rect 55988 28708 55997 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 73411 28708 73420 28748
rect 73460 28708 75340 28748
rect 75380 28708 75389 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 50956 28664 50996 28708
rect 54787 28707 54845 28708
rect 51427 28664 51485 28665
rect 40387 28624 40396 28664
rect 40436 28624 41548 28664
rect 41588 28624 41597 28664
rect 50947 28624 50956 28664
rect 50996 28624 51036 28664
rect 51342 28624 51436 28664
rect 51476 28624 51485 28664
rect 56419 28624 56428 28664
rect 56468 28624 58732 28664
rect 58772 28624 66796 28664
rect 66836 28624 66845 28664
rect 76675 28624 76684 28664
rect 76724 28624 77068 28664
rect 77108 28624 77117 28664
rect 51427 28623 51485 28624
rect 39619 28540 39628 28580
rect 39668 28540 40436 28580
rect 41443 28540 41452 28580
rect 41492 28540 41932 28580
rect 41972 28540 41981 28580
rect 55267 28540 55276 28580
rect 55316 28540 55468 28580
rect 55508 28540 55517 28580
rect 59011 28540 59020 28580
rect 59060 28540 59404 28580
rect 59444 28540 68428 28580
rect 68468 28540 68477 28580
rect 70627 28540 70636 28580
rect 70676 28540 71500 28580
rect 71540 28540 73804 28580
rect 73844 28540 73853 28580
rect 40396 28496 40436 28540
rect 40387 28456 40396 28496
rect 40436 28456 40445 28496
rect 52963 28456 52972 28496
rect 53012 28456 54796 28496
rect 54836 28456 54845 28496
rect 60643 28456 60652 28496
rect 60692 28456 60701 28496
rect 63715 28456 63724 28496
rect 63764 28456 64684 28496
rect 64724 28456 64733 28496
rect 70243 28456 70252 28496
rect 70292 28456 71116 28496
rect 71156 28456 71165 28496
rect 55651 28412 55709 28413
rect 60652 28412 60692 28456
rect 40963 28372 40972 28412
rect 41012 28372 41260 28412
rect 41300 28372 41309 28412
rect 51715 28372 51724 28412
rect 51764 28372 55660 28412
rect 55700 28372 55709 28412
rect 55651 28371 55709 28372
rect 59884 28372 60692 28412
rect 76387 28372 76396 28412
rect 76436 28372 77396 28412
rect 0 28268 80 28348
rect 59884 28328 59924 28372
rect 64579 28328 64637 28329
rect 71011 28328 71069 28329
rect 77356 28328 77396 28372
rect 40387 28288 40396 28328
rect 40436 28288 41452 28328
rect 41492 28288 41501 28328
rect 45667 28288 45676 28328
rect 45716 28288 46348 28328
rect 46388 28288 46397 28328
rect 49987 28288 49996 28328
rect 50036 28288 51820 28328
rect 51860 28288 51869 28328
rect 52099 28288 52108 28328
rect 52148 28288 52588 28328
rect 52628 28288 52637 28328
rect 55651 28288 55660 28328
rect 55700 28288 56428 28328
rect 56468 28288 56477 28328
rect 59875 28288 59884 28328
rect 59924 28288 59933 28328
rect 60355 28288 60364 28328
rect 60404 28288 60652 28328
rect 60692 28288 60701 28328
rect 61699 28288 61708 28328
rect 61748 28288 63148 28328
rect 63188 28288 64396 28328
rect 64436 28288 64445 28328
rect 64579 28288 64588 28328
rect 64628 28288 64722 28328
rect 66979 28288 66988 28328
rect 67028 28288 67276 28328
rect 67316 28288 69196 28328
rect 69236 28288 69868 28328
rect 69908 28288 69917 28328
rect 70926 28288 71020 28328
rect 71060 28288 71069 28328
rect 75427 28288 75436 28328
rect 75476 28288 76588 28328
rect 76628 28288 76876 28328
rect 76916 28288 76925 28328
rect 77347 28288 77356 28328
rect 77396 28288 78124 28328
rect 78164 28288 79468 28328
rect 79508 28288 79517 28328
rect 64579 28287 64637 28288
rect 71011 28287 71069 28288
rect 38371 28204 38380 28244
rect 38420 28204 40972 28244
rect 41012 28204 41021 28244
rect 41539 28204 41548 28244
rect 41588 28204 42604 28244
rect 42644 28204 51052 28244
rect 51092 28204 51101 28244
rect 51148 28204 53300 28244
rect 64003 28204 64012 28244
rect 64052 28204 64300 28244
rect 64340 28204 64972 28244
rect 65012 28204 65021 28244
rect 76963 28204 76972 28244
rect 77012 28204 77260 28244
rect 77300 28204 77309 28244
rect 51148 28160 51188 28204
rect 53260 28160 53300 28204
rect 77155 28160 77213 28161
rect 48835 28120 48844 28160
rect 48884 28120 50092 28160
rect 50132 28120 50141 28160
rect 50563 28120 50572 28160
rect 50612 28120 51188 28160
rect 51235 28120 51244 28160
rect 51284 28120 52396 28160
rect 52436 28120 52445 28160
rect 53260 28120 55756 28160
rect 55796 28120 55805 28160
rect 57091 28120 57100 28160
rect 57140 28120 59308 28160
rect 59348 28120 59357 28160
rect 64867 28120 64876 28160
rect 64916 28120 65836 28160
rect 65876 28120 68140 28160
rect 68180 28120 71500 28160
rect 71540 28120 71549 28160
rect 77070 28120 77164 28160
rect 77204 28120 77213 28160
rect 77155 28119 77213 28120
rect 51235 28076 51293 28077
rect 50179 28036 50188 28076
rect 50228 28036 50380 28076
rect 50420 28036 50429 28076
rect 51235 28036 51244 28076
rect 51284 28036 58540 28076
rect 58580 28036 58589 28076
rect 76675 28036 76684 28076
rect 76724 28036 77068 28076
rect 77108 28036 77117 28076
rect 51235 28035 51293 28036
rect 50371 27992 50429 27993
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 50371 27952 50380 27992
rect 50420 27952 51860 27992
rect 52291 27952 52300 27992
rect 52340 27952 54508 27992
rect 54548 27952 63532 27992
rect 63572 27952 63581 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 70051 27952 70060 27992
rect 70100 27952 70540 27992
rect 70580 27952 70589 27992
rect 70723 27952 70732 27992
rect 70772 27952 71212 27992
rect 71252 27952 71261 27992
rect 73420 27952 74284 27992
rect 74324 27952 75436 27992
rect 75476 27952 75485 27992
rect 50371 27951 50429 27952
rect 51715 27908 51773 27909
rect 38659 27868 38668 27908
rect 38708 27868 48212 27908
rect 50371 27868 50380 27908
rect 50420 27868 50668 27908
rect 50708 27868 51244 27908
rect 51284 27868 51293 27908
rect 51630 27868 51724 27908
rect 51764 27868 51773 27908
rect 51820 27908 51860 27952
rect 73420 27908 73460 27952
rect 51820 27868 60940 27908
rect 60980 27868 60989 27908
rect 70060 27868 73460 27908
rect 48172 27824 48212 27868
rect 51715 27867 51773 27868
rect 70060 27824 70100 27868
rect 41347 27784 41356 27824
rect 41396 27784 44140 27824
rect 44180 27784 44189 27824
rect 44995 27784 45004 27824
rect 45044 27784 45964 27824
rect 46004 27784 46444 27824
rect 46484 27784 46493 27824
rect 47203 27784 47212 27824
rect 47252 27784 47692 27824
rect 47732 27784 47741 27824
rect 48172 27784 58444 27824
rect 58484 27784 58493 27824
rect 59203 27784 59212 27824
rect 59252 27784 59692 27824
rect 59732 27784 59741 27824
rect 59875 27784 59884 27824
rect 59924 27784 59933 27824
rect 61891 27784 61900 27824
rect 61940 27784 64012 27824
rect 64052 27784 64061 27824
rect 65155 27784 65164 27824
rect 65204 27784 65644 27824
rect 65684 27784 65932 27824
rect 65972 27784 65981 27824
rect 68323 27784 68332 27824
rect 68372 27784 68620 27824
rect 68660 27784 69004 27824
rect 69044 27784 70060 27824
rect 70100 27784 70109 27824
rect 70627 27784 70636 27824
rect 70676 27784 71692 27824
rect 71732 27784 71741 27824
rect 37699 27700 37708 27740
rect 37748 27700 40396 27740
rect 40436 27700 40445 27740
rect 40963 27656 41021 27657
rect 39811 27616 39820 27656
rect 39860 27616 40300 27656
rect 40340 27616 40349 27656
rect 40878 27616 40972 27656
rect 41012 27616 43276 27656
rect 43316 27616 43325 27656
rect 40963 27615 41021 27616
rect 0 27428 80 27508
rect 40867 27488 40925 27489
rect 43468 27488 43508 27784
rect 43555 27700 43564 27740
rect 43604 27700 45580 27740
rect 45620 27700 45629 27740
rect 46531 27700 46540 27740
rect 46580 27700 47788 27740
rect 47828 27700 47837 27740
rect 51715 27700 51724 27740
rect 51764 27700 52108 27740
rect 52148 27700 52157 27740
rect 55171 27700 55180 27740
rect 55220 27700 56812 27740
rect 56852 27700 56861 27740
rect 59884 27656 59924 27784
rect 65251 27700 65260 27740
rect 65300 27700 65740 27740
rect 65780 27700 65789 27740
rect 68419 27700 68428 27740
rect 68468 27700 73460 27740
rect 47395 27616 47404 27656
rect 47444 27616 47692 27656
rect 47732 27616 47741 27656
rect 51907 27616 51916 27656
rect 51956 27616 52204 27656
rect 52244 27616 52253 27656
rect 55939 27616 55948 27656
rect 55988 27616 56332 27656
rect 56372 27616 56381 27656
rect 59299 27616 59308 27656
rect 59348 27616 59924 27656
rect 60835 27616 60844 27656
rect 60884 27616 61132 27656
rect 61172 27616 61181 27656
rect 63907 27616 63916 27656
rect 63956 27616 65356 27656
rect 65396 27616 65405 27656
rect 69763 27616 69772 27656
rect 69812 27616 71788 27656
rect 71828 27616 71837 27656
rect 73420 27572 73460 27700
rect 75043 27616 75052 27656
rect 75092 27616 76876 27656
rect 76916 27616 77068 27656
rect 77108 27616 77117 27656
rect 76195 27572 76253 27573
rect 46339 27532 46348 27572
rect 46388 27532 47308 27572
rect 47348 27532 47357 27572
rect 47779 27532 47788 27572
rect 47828 27532 49420 27572
rect 49460 27532 49469 27572
rect 52387 27532 52396 27572
rect 52436 27532 55372 27572
rect 55412 27532 55421 27572
rect 59779 27532 59788 27572
rect 59828 27532 60268 27572
rect 60308 27532 63436 27572
rect 63476 27532 64492 27572
rect 64532 27532 64541 27572
rect 65443 27532 65452 27572
rect 65492 27532 65740 27572
rect 65780 27532 65789 27572
rect 69091 27532 69100 27572
rect 69140 27532 69149 27572
rect 73420 27532 76204 27572
rect 76244 27532 76253 27572
rect 40867 27448 40876 27488
rect 40916 27448 43220 27488
rect 43468 27448 52052 27488
rect 40867 27447 40925 27448
rect 41251 27404 41309 27405
rect 43180 27404 43220 27448
rect 50371 27404 50429 27405
rect 40483 27364 40492 27404
rect 40532 27364 41068 27404
rect 41108 27364 41260 27404
rect 41300 27364 41309 27404
rect 41539 27364 41548 27404
rect 41588 27364 43084 27404
rect 43124 27364 43133 27404
rect 43180 27364 50380 27404
rect 50420 27364 50429 27404
rect 41251 27363 41309 27364
rect 50371 27363 50429 27364
rect 51715 27404 51773 27405
rect 51715 27364 51724 27404
rect 51764 27364 51820 27404
rect 51860 27364 51869 27404
rect 51715 27363 51773 27364
rect 52012 27320 52052 27448
rect 52396 27404 52436 27532
rect 52771 27488 52829 27489
rect 69100 27488 69140 27532
rect 76195 27531 76253 27532
rect 52771 27448 52780 27488
rect 52820 27448 60460 27488
rect 60500 27448 61324 27488
rect 61364 27448 61373 27488
rect 69100 27448 69772 27488
rect 69812 27448 69821 27488
rect 70243 27448 70252 27488
rect 70292 27448 70636 27488
rect 70676 27448 70685 27488
rect 52771 27447 52829 27448
rect 52099 27364 52108 27404
rect 52148 27364 52436 27404
rect 59491 27364 59500 27404
rect 59540 27364 59980 27404
rect 60020 27364 60029 27404
rect 63340 27364 63724 27404
rect 63764 27364 63773 27404
rect 64387 27364 64396 27404
rect 64436 27364 65260 27404
rect 65300 27364 66892 27404
rect 66932 27364 66941 27404
rect 69091 27364 69100 27404
rect 69140 27364 69580 27404
rect 69620 27364 69629 27404
rect 75043 27364 75052 27404
rect 75092 27364 75244 27404
rect 75284 27364 75293 27404
rect 63340 27320 63380 27364
rect 52012 27280 57964 27320
rect 58004 27280 58013 27320
rect 60931 27280 60940 27320
rect 60980 27280 61228 27320
rect 61268 27280 63380 27320
rect 63724 27320 63764 27364
rect 71107 27320 71165 27321
rect 63724 27280 67660 27320
rect 67700 27280 67709 27320
rect 71022 27280 71116 27320
rect 71156 27280 71165 27320
rect 71107 27279 71165 27280
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 39619 27196 39628 27236
rect 39668 27196 41260 27236
rect 41300 27196 41309 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 49603 27196 49612 27236
rect 49652 27196 50092 27236
rect 50132 27196 53356 27236
rect 53396 27196 53405 27236
rect 59779 27196 59788 27236
rect 59828 27196 60748 27236
rect 60788 27196 62860 27236
rect 62900 27196 62909 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 40483 27112 40492 27152
rect 40532 27112 43372 27152
rect 43412 27112 60364 27152
rect 60404 27112 60413 27152
rect 61996 27112 64300 27152
rect 64340 27112 64349 27152
rect 70915 27112 70924 27152
rect 70964 27112 71596 27152
rect 71636 27112 71884 27152
rect 71924 27112 71933 27152
rect 61996 27068 62036 27112
rect 40867 27028 40876 27068
rect 40916 27028 41740 27068
rect 41780 27028 41789 27068
rect 44899 27028 44908 27068
rect 44948 27028 45100 27068
rect 45140 27028 45149 27068
rect 54211 27028 54220 27068
rect 54260 27028 55660 27068
rect 55700 27028 55709 27068
rect 58147 27028 58156 27068
rect 58196 27028 58444 27068
rect 58484 27028 59884 27068
rect 59924 27028 61996 27068
rect 62036 27028 62045 27068
rect 62275 27028 62284 27068
rect 62324 27028 71692 27068
rect 71732 27028 71741 27068
rect 74659 27028 74668 27068
rect 74708 27028 75820 27068
rect 75860 27028 75869 27068
rect 50275 26984 50333 26985
rect 32995 26944 33004 26984
rect 33044 26944 34252 26984
rect 34292 26944 34301 26984
rect 41443 26944 41452 26984
rect 41492 26944 44756 26984
rect 45283 26944 45292 26984
rect 45332 26944 45676 26984
rect 45716 26944 45725 26984
rect 46051 26944 46060 26984
rect 46100 26944 46636 26984
rect 46676 26944 46685 26984
rect 50190 26944 50284 26984
rect 50324 26944 50333 26984
rect 51235 26944 51244 26984
rect 51284 26944 51628 26984
rect 51668 26944 51677 26984
rect 57667 26944 57676 26984
rect 57716 26944 58252 26984
rect 58292 26944 67564 26984
rect 67604 26944 67613 26984
rect 75619 26944 75628 26984
rect 75668 26944 75708 26984
rect 44716 26900 44756 26944
rect 50275 26943 50333 26944
rect 51523 26900 51581 26901
rect 75628 26900 75668 26944
rect 35011 26860 35020 26900
rect 35060 26860 35596 26900
rect 35636 26860 35645 26900
rect 38851 26860 38860 26900
rect 38900 26860 39052 26900
rect 39092 26860 41644 26900
rect 41684 26860 43220 26900
rect 44707 26860 44716 26900
rect 44756 26860 47596 26900
rect 47636 26860 47645 26900
rect 51523 26860 51532 26900
rect 51572 26860 53260 26900
rect 53300 26860 53309 26900
rect 59107 26860 59116 26900
rect 59156 26860 59980 26900
rect 60020 26860 60029 26900
rect 60835 26860 60844 26900
rect 60884 26860 62284 26900
rect 62324 26860 62333 26900
rect 73027 26860 73036 26900
rect 73076 26860 74860 26900
rect 74900 26860 74909 26900
rect 75427 26860 75436 26900
rect 75476 26860 75956 26900
rect 35203 26776 35212 26816
rect 35252 26776 35692 26816
rect 35732 26776 35741 26816
rect 40099 26776 40108 26816
rect 40148 26776 40780 26816
rect 40820 26776 40829 26816
rect 43180 26732 43220 26860
rect 51523 26859 51581 26860
rect 75916 26816 75956 26860
rect 43267 26776 43276 26816
rect 43316 26776 46444 26816
rect 46484 26776 46636 26816
rect 46676 26776 47212 26816
rect 47252 26776 47261 26816
rect 48259 26776 48268 26816
rect 48308 26776 49612 26816
rect 49652 26776 49661 26816
rect 50275 26776 50284 26816
rect 50324 26776 51476 26816
rect 51523 26776 51532 26816
rect 51572 26776 52300 26816
rect 52340 26776 52349 26816
rect 52396 26776 57484 26816
rect 57524 26776 57533 26816
rect 58819 26776 58828 26816
rect 58868 26776 63244 26816
rect 63284 26776 63820 26816
rect 63860 26776 63869 26816
rect 66403 26776 66412 26816
rect 66452 26776 67756 26816
rect 67796 26776 67805 26816
rect 68611 26776 68620 26816
rect 68660 26776 69292 26816
rect 69332 26776 69341 26816
rect 74755 26776 74764 26816
rect 74804 26776 75628 26816
rect 75668 26776 75677 26816
rect 75907 26776 75916 26816
rect 75956 26776 76588 26816
rect 76628 26776 76637 26816
rect 39715 26692 39724 26732
rect 39764 26692 39916 26732
rect 39956 26692 40204 26732
rect 40244 26692 40253 26732
rect 40387 26692 40396 26732
rect 40436 26692 41740 26732
rect 41780 26692 41789 26732
rect 43180 26692 49516 26732
rect 49556 26692 49565 26732
rect 50179 26692 50188 26732
rect 50228 26692 50572 26732
rect 50612 26692 50621 26732
rect 0 26588 80 26668
rect 40396 26648 40436 26692
rect 51436 26648 51476 26776
rect 39619 26608 39628 26648
rect 39668 26608 40436 26648
rect 44995 26608 45004 26648
rect 45044 26608 45676 26648
rect 45716 26608 47980 26648
rect 48020 26608 48029 26648
rect 48739 26608 48748 26648
rect 48788 26608 50764 26648
rect 50804 26608 50813 26648
rect 51436 26608 52300 26648
rect 52340 26608 52349 26648
rect 38947 26564 39005 26565
rect 52396 26564 52436 26776
rect 53251 26692 53260 26732
rect 53300 26692 60556 26732
rect 60596 26692 72268 26732
rect 72308 26692 72317 26732
rect 74851 26692 74860 26732
rect 74900 26692 75820 26732
rect 75860 26692 76300 26732
rect 76340 26692 76349 26732
rect 55459 26608 55468 26648
rect 55508 26608 56044 26648
rect 56084 26608 56093 26648
rect 59107 26608 59116 26648
rect 59156 26608 59500 26648
rect 59540 26608 59692 26648
rect 59732 26608 59741 26648
rect 67651 26608 67660 26648
rect 67700 26608 68660 26648
rect 71875 26608 71884 26648
rect 71924 26608 75724 26648
rect 75764 26608 76204 26648
rect 76244 26608 76253 26648
rect 76483 26608 76492 26648
rect 76532 26608 77356 26648
rect 77396 26608 78508 26648
rect 78548 26608 79468 26648
rect 79508 26608 79517 26648
rect 68620 26564 68660 26608
rect 38947 26524 38956 26564
rect 38996 26524 52436 26564
rect 52492 26524 61324 26564
rect 61364 26524 61373 26564
rect 62851 26524 62860 26564
rect 62900 26524 68468 26564
rect 68611 26524 68620 26564
rect 68660 26524 68669 26564
rect 38947 26523 39005 26524
rect 52492 26480 52532 26524
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 50179 26440 50188 26480
rect 50228 26440 52532 26480
rect 52963 26480 53021 26481
rect 68428 26480 68468 26524
rect 52963 26440 52972 26480
rect 53012 26440 58924 26480
rect 58964 26440 58973 26480
rect 59683 26440 59692 26480
rect 59732 26440 60076 26480
rect 60116 26440 60125 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 68419 26440 68428 26480
rect 68468 26440 68477 26480
rect 68803 26440 68812 26480
rect 68852 26440 69004 26480
rect 69044 26440 69053 26480
rect 71971 26440 71980 26480
rect 72020 26440 75820 26480
rect 75860 26440 75869 26480
rect 52963 26439 53021 26440
rect 34924 26356 37036 26396
rect 37076 26356 37085 26396
rect 40675 26356 40684 26396
rect 40724 26356 41452 26396
rect 41492 26356 44044 26396
rect 44084 26356 59308 26396
rect 59348 26356 59357 26396
rect 67363 26356 67372 26396
rect 67412 26356 69484 26396
rect 69524 26356 74764 26396
rect 74804 26356 74813 26396
rect 34924 26312 34964 26356
rect 34915 26272 34924 26312
rect 34964 26272 34973 26312
rect 35779 26272 35788 26312
rect 35828 26272 35837 26312
rect 49411 26272 49420 26312
rect 49460 26272 50188 26312
rect 50228 26272 50237 26312
rect 50659 26272 50668 26312
rect 50708 26272 52108 26312
rect 52148 26272 52157 26312
rect 52291 26272 52300 26312
rect 52340 26272 52588 26312
rect 52628 26272 57004 26312
rect 57044 26272 59020 26312
rect 59060 26272 59069 26312
rect 60259 26272 60268 26312
rect 60308 26272 60460 26312
rect 60500 26272 61228 26312
rect 61268 26272 61277 26312
rect 65347 26272 65356 26312
rect 65396 26272 65548 26312
rect 65588 26272 68276 26312
rect 69091 26272 69100 26312
rect 69140 26272 69388 26312
rect 69428 26272 69437 26312
rect 71011 26272 71020 26312
rect 71060 26272 71788 26312
rect 71828 26272 71837 26312
rect 35788 26144 35828 26272
rect 68236 26228 68276 26272
rect 39235 26188 39244 26228
rect 39284 26188 39820 26228
rect 39860 26188 40300 26228
rect 40340 26188 40349 26228
rect 43171 26188 43180 26228
rect 43220 26188 60652 26228
rect 60692 26188 60701 26228
rect 61603 26188 61612 26228
rect 61652 26188 64780 26228
rect 64820 26188 64829 26228
rect 67267 26188 67276 26228
rect 67316 26188 67325 26228
rect 68227 26188 68236 26228
rect 68276 26188 68285 26228
rect 68611 26188 68620 26228
rect 68660 26188 68812 26228
rect 68852 26188 68861 26228
rect 69283 26188 69292 26228
rect 69332 26188 71308 26228
rect 71348 26188 71500 26228
rect 71540 26188 71549 26228
rect 73420 26188 74860 26228
rect 74900 26188 74909 26228
rect 41251 26144 41309 26145
rect 67276 26144 67316 26188
rect 73420 26144 73460 26188
rect 34435 26104 34444 26144
rect 34484 26104 35308 26144
rect 35348 26104 35357 26144
rect 35788 26104 36268 26144
rect 36308 26104 36317 26144
rect 36451 26104 36460 26144
rect 36500 26104 38380 26144
rect 38420 26104 38429 26144
rect 41166 26104 41260 26144
rect 41300 26104 41309 26144
rect 43651 26104 43660 26144
rect 43700 26104 45100 26144
rect 45140 26104 45149 26144
rect 49603 26104 49612 26144
rect 49652 26104 49996 26144
rect 50036 26104 50045 26144
rect 51427 26104 51436 26144
rect 51476 26104 51724 26144
rect 51764 26104 55468 26144
rect 55508 26104 55517 26144
rect 55747 26104 55756 26144
rect 55796 26104 57292 26144
rect 57332 26104 57341 26144
rect 58531 26104 58540 26144
rect 58580 26104 59500 26144
rect 59540 26104 59884 26144
rect 59924 26104 59933 26144
rect 60067 26104 60076 26144
rect 60116 26104 60460 26144
rect 60500 26104 60509 26144
rect 63811 26104 63820 26144
rect 63860 26104 65452 26144
rect 65492 26104 65501 26144
rect 65731 26104 65740 26144
rect 65780 26104 67180 26144
rect 67220 26104 67229 26144
rect 67276 26104 69388 26144
rect 69428 26104 70540 26144
rect 70580 26104 73460 26144
rect 74467 26104 74476 26144
rect 74516 26104 74668 26144
rect 74708 26104 74717 26144
rect 74947 26104 74956 26144
rect 74996 26104 75436 26144
rect 75476 26104 75485 26144
rect 75811 26104 75820 26144
rect 75860 26104 76780 26144
rect 76820 26104 76829 26144
rect 77347 26104 77356 26144
rect 77396 26104 77740 26144
rect 77780 26104 77789 26144
rect 41251 26103 41309 26104
rect 38947 26060 39005 26061
rect 52867 26060 52925 26061
rect 61027 26060 61085 26061
rect 7180 26020 38092 26060
rect 38132 26020 38141 26060
rect 38862 26020 38956 26060
rect 38996 26020 39005 26060
rect 47107 26020 47116 26060
rect 47156 26020 48076 26060
rect 48116 26020 48125 26060
rect 52483 26020 52492 26060
rect 52532 26020 52541 26060
rect 52867 26020 52876 26060
rect 52916 26020 57676 26060
rect 57716 26020 57725 26060
rect 60942 26020 61036 26060
rect 61076 26020 61085 26060
rect 61219 26020 61228 26060
rect 61268 26020 70444 26060
rect 70484 26020 70493 26060
rect 70540 26020 70636 26060
rect 70676 26020 70685 26060
rect 7180 25976 7220 26020
rect 38947 26019 39005 26020
rect 835 25936 844 25976
rect 884 25936 7220 25976
rect 32227 25936 32236 25976
rect 32276 25936 33196 25976
rect 33236 25936 34444 25976
rect 34484 25936 34493 25976
rect 35203 25936 35212 25976
rect 35252 25936 36460 25976
rect 36500 25936 36509 25976
rect 44899 25936 44908 25976
rect 44948 25936 45772 25976
rect 45812 25936 47020 25976
rect 47060 25936 48268 25976
rect 48308 25936 48317 25976
rect 48547 25936 48556 25976
rect 48596 25936 49132 25976
rect 49172 25936 49181 25976
rect 44908 25892 44948 25936
rect 52492 25892 52532 26020
rect 52867 26019 52925 26020
rect 61027 26019 61085 26020
rect 70540 25976 70580 26020
rect 54883 25936 54892 25976
rect 54932 25936 56236 25976
rect 56276 25936 56285 25976
rect 57379 25936 57388 25976
rect 57428 25936 58348 25976
rect 58388 25936 58397 25976
rect 59395 25936 59404 25976
rect 59444 25936 61132 25976
rect 61172 25936 61181 25976
rect 64963 25936 64972 25976
rect 65012 25936 65452 25976
rect 65492 25936 65501 25976
rect 68611 25936 68620 25976
rect 68660 25936 70540 25976
rect 70580 25936 70589 25976
rect 73219 25936 73228 25976
rect 73268 25936 74476 25976
rect 74516 25936 74525 25976
rect 74755 25936 74764 25976
rect 74804 25936 75148 25976
rect 75188 25936 75197 25976
rect 33379 25852 33388 25892
rect 33428 25852 33868 25892
rect 33908 25852 33917 25892
rect 35107 25852 35116 25892
rect 35156 25852 35980 25892
rect 36020 25852 36029 25892
rect 36163 25852 36172 25892
rect 36212 25852 37228 25892
rect 37268 25852 38476 25892
rect 38516 25852 38860 25892
rect 38900 25852 38909 25892
rect 43651 25852 43660 25892
rect 43700 25852 44948 25892
rect 45571 25852 45580 25892
rect 45620 25852 46060 25892
rect 46100 25852 46109 25892
rect 51811 25852 51820 25892
rect 51860 25852 54700 25892
rect 54740 25852 54749 25892
rect 60739 25852 60748 25892
rect 60788 25852 63916 25892
rect 63956 25852 65644 25892
rect 65684 25852 65693 25892
rect 69187 25852 69196 25892
rect 69236 25852 70348 25892
rect 70388 25852 71980 25892
rect 72020 25852 72652 25892
rect 72692 25852 74380 25892
rect 74420 25852 74429 25892
rect 0 25808 80 25828
rect 0 25768 652 25808
rect 692 25768 701 25808
rect 58915 25768 58924 25808
rect 58964 25768 60844 25808
rect 60884 25768 60893 25808
rect 0 25748 80 25768
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 39523 25684 39532 25724
rect 39572 25684 40780 25724
rect 40820 25684 40829 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 39139 25600 39148 25640
rect 39188 25600 43220 25640
rect 46627 25600 46636 25640
rect 46676 25600 46924 25640
rect 46964 25600 46973 25640
rect 47971 25600 47980 25640
rect 48020 25600 58732 25640
rect 58772 25600 58781 25640
rect 40963 25556 41021 25557
rect 39523 25516 39532 25556
rect 39572 25516 40012 25556
rect 40052 25516 40061 25556
rect 40387 25516 40396 25556
rect 40436 25516 40972 25556
rect 41012 25516 41021 25556
rect 43180 25556 43220 25600
rect 43180 25516 49324 25556
rect 49364 25516 49612 25556
rect 49652 25516 49661 25556
rect 63523 25516 63532 25556
rect 63572 25516 64012 25556
rect 64052 25516 64061 25556
rect 70723 25516 70732 25556
rect 70772 25516 73460 25556
rect 74275 25516 74284 25556
rect 74324 25516 75916 25556
rect 75956 25516 76300 25556
rect 76340 25516 76349 25556
rect 40963 25515 41021 25516
rect 35875 25432 35884 25472
rect 35924 25432 35933 25472
rect 38083 25432 38092 25472
rect 38132 25432 43220 25472
rect 45187 25432 45196 25472
rect 45236 25432 45484 25472
rect 45524 25432 45533 25472
rect 46051 25432 46060 25472
rect 46100 25432 46444 25472
rect 46484 25432 46493 25472
rect 63427 25432 63436 25472
rect 63476 25432 63724 25472
rect 63764 25432 63773 25472
rect 71203 25432 71212 25472
rect 71252 25432 71261 25472
rect 31747 25348 31756 25388
rect 31796 25348 34580 25388
rect 34540 25304 34580 25348
rect 35884 25304 35924 25432
rect 43180 25388 43220 25432
rect 39427 25348 39436 25388
rect 39476 25348 40108 25388
rect 40148 25348 40157 25388
rect 43180 25348 44852 25388
rect 44899 25348 44908 25388
rect 44948 25348 46732 25388
rect 46772 25348 46781 25388
rect 54691 25348 54700 25388
rect 54740 25348 63628 25388
rect 63668 25348 63677 25388
rect 44812 25304 44852 25348
rect 55267 25304 55325 25305
rect 30979 25264 30988 25304
rect 31028 25264 32812 25304
rect 32852 25264 33868 25304
rect 33908 25264 33917 25304
rect 34531 25264 34540 25304
rect 34580 25264 34589 25304
rect 35587 25264 35596 25304
rect 35636 25264 35924 25304
rect 37219 25264 37228 25304
rect 37268 25264 39340 25304
rect 39380 25264 39389 25304
rect 39619 25264 39628 25304
rect 39668 25264 39820 25304
rect 39860 25264 39869 25304
rect 42115 25264 42124 25304
rect 42164 25264 42988 25304
rect 43028 25264 43660 25304
rect 43700 25264 43709 25304
rect 44812 25264 45524 25304
rect 45571 25264 45580 25304
rect 45620 25264 46540 25304
rect 46580 25264 46589 25304
rect 49987 25264 49996 25304
rect 50036 25264 50668 25304
rect 50708 25264 50717 25304
rect 52099 25264 52108 25304
rect 52148 25264 55276 25304
rect 55316 25264 55325 25304
rect 55459 25264 55468 25304
rect 55508 25264 56236 25304
rect 56276 25264 56285 25304
rect 58627 25264 58636 25304
rect 58676 25264 61516 25304
rect 61556 25264 62860 25304
rect 62900 25264 62909 25304
rect 68323 25264 68332 25304
rect 68372 25264 68524 25304
rect 68564 25264 68573 25304
rect 45484 25220 45524 25264
rect 55267 25263 55325 25264
rect 64579 25220 64637 25221
rect 32995 25180 33004 25220
rect 33044 25180 33140 25220
rect 33475 25180 33484 25220
rect 33524 25180 34636 25220
rect 34676 25180 36076 25220
rect 36116 25180 36125 25220
rect 38467 25180 38476 25220
rect 38516 25180 39724 25220
rect 39764 25180 39773 25220
rect 40003 25180 40012 25220
rect 40052 25180 40204 25220
rect 40244 25180 44044 25220
rect 44084 25180 45388 25220
rect 45428 25180 45437 25220
rect 45484 25180 52588 25220
rect 52628 25180 52637 25220
rect 59203 25180 59212 25220
rect 59252 25180 59500 25220
rect 59540 25180 59549 25220
rect 59683 25180 59692 25220
rect 59732 25180 63148 25220
rect 63188 25180 64588 25220
rect 64628 25180 67084 25220
rect 67124 25180 67133 25220
rect 33100 25136 33140 25180
rect 64579 25179 64637 25180
rect 71212 25136 71252 25432
rect 73420 25220 73460 25516
rect 74467 25264 74476 25304
rect 74516 25264 77932 25304
rect 77972 25264 78316 25304
rect 78356 25264 78365 25304
rect 73420 25180 76492 25220
rect 76532 25180 76876 25220
rect 76916 25180 76925 25220
rect 835 25096 844 25136
rect 884 25096 3916 25136
rect 3956 25096 3965 25136
rect 31651 25096 31660 25136
rect 31700 25096 32140 25136
rect 32180 25096 32189 25136
rect 33100 25096 33292 25136
rect 33332 25096 33341 25136
rect 38371 25096 38380 25136
rect 38420 25096 54700 25136
rect 54740 25096 54749 25136
rect 55459 25096 55468 25136
rect 55508 25096 55756 25136
rect 55796 25096 55805 25136
rect 57091 25096 57100 25136
rect 57140 25096 58060 25136
rect 58100 25096 58109 25136
rect 58435 25096 58444 25136
rect 58484 25096 60364 25136
rect 60404 25096 60413 25136
rect 60643 25096 60652 25136
rect 60692 25096 60940 25136
rect 60980 25096 60989 25136
rect 63340 25096 63916 25136
rect 63956 25096 65932 25136
rect 65972 25096 65981 25136
rect 67363 25096 67372 25136
rect 67412 25096 68372 25136
rect 71212 25096 71404 25136
rect 71444 25096 72844 25136
rect 72884 25096 73036 25136
rect 73076 25096 73085 25136
rect 63340 25052 63380 25096
rect 68332 25052 68372 25096
rect 33091 25012 33100 25052
rect 33140 25012 35692 25052
rect 35732 25012 35741 25052
rect 39139 25012 39148 25052
rect 39188 25012 39916 25052
rect 39956 25012 44140 25052
rect 44180 25012 45484 25052
rect 45524 25012 45533 25052
rect 46435 25012 46444 25052
rect 46484 25012 48172 25052
rect 48212 25012 49420 25052
rect 49460 25012 60404 25052
rect 60451 25012 60460 25052
rect 60500 25012 63380 25052
rect 63427 25012 63436 25052
rect 63476 25012 64588 25052
rect 64628 25012 66412 25052
rect 66452 25012 66461 25052
rect 67651 25012 67660 25052
rect 67700 25012 67852 25052
rect 67892 25012 67901 25052
rect 68323 25012 68332 25052
rect 68372 25012 70348 25052
rect 70388 25012 72460 25052
rect 72500 25012 72509 25052
rect 0 24968 80 24988
rect 51427 24968 51485 24969
rect 59299 24968 59357 24969
rect 60364 24968 60404 25012
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 35587 24928 35596 24968
rect 35636 24928 40492 24968
rect 40532 24928 40541 24968
rect 40588 24928 40876 24968
rect 40916 24928 40925 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 50371 24928 50380 24968
rect 50420 24928 50572 24968
rect 50612 24928 50621 24968
rect 51427 24928 51436 24968
rect 51476 24928 59308 24968
rect 59348 24928 59357 24968
rect 59875 24928 59884 24968
rect 59924 24928 60268 24968
rect 60308 24928 60317 24968
rect 60364 24928 61708 24968
rect 61748 24928 61757 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 70531 24928 70540 24968
rect 70580 24928 71212 24968
rect 71252 24928 74476 24968
rect 74516 24928 74525 24968
rect 0 24908 80 24928
rect 30787 24884 30845 24885
rect 40588 24884 40628 24928
rect 51427 24927 51485 24928
rect 59299 24927 59357 24928
rect 30787 24844 30796 24884
rect 30836 24844 31852 24884
rect 31892 24844 33484 24884
rect 33524 24844 33533 24884
rect 35011 24844 35020 24884
rect 35060 24844 36556 24884
rect 36596 24844 36605 24884
rect 40579 24844 40588 24884
rect 40628 24844 40637 24884
rect 41155 24844 41164 24884
rect 41204 24844 43220 24884
rect 46819 24844 46828 24884
rect 46868 24844 47020 24884
rect 47060 24844 47069 24884
rect 50659 24844 50668 24884
rect 50708 24844 51148 24884
rect 51188 24844 51724 24884
rect 51764 24844 51773 24884
rect 51907 24844 51916 24884
rect 51956 24844 74572 24884
rect 74612 24844 74621 24884
rect 30787 24843 30845 24844
rect 43180 24800 43220 24844
rect 29731 24760 29740 24800
rect 29780 24760 32236 24800
rect 32276 24760 32285 24800
rect 35875 24760 35884 24800
rect 35924 24760 36268 24800
rect 36308 24760 37996 24800
rect 38036 24760 38045 24800
rect 43180 24760 43276 24800
rect 43316 24760 59308 24800
rect 59348 24760 59357 24800
rect 59587 24760 59596 24800
rect 59636 24760 60364 24800
rect 60404 24760 62668 24800
rect 62708 24760 67564 24800
rect 67604 24760 67613 24800
rect 71011 24760 71020 24800
rect 71060 24760 71596 24800
rect 71636 24760 71645 24800
rect 7459 24676 7468 24716
rect 7508 24676 55180 24716
rect 55220 24676 55229 24716
rect 58051 24676 58060 24716
rect 58100 24676 59500 24716
rect 59540 24676 59788 24716
rect 59828 24676 59837 24716
rect 60163 24676 60172 24716
rect 60212 24676 60748 24716
rect 60788 24676 60797 24716
rect 64099 24676 64108 24716
rect 64148 24676 64876 24716
rect 64916 24676 65260 24716
rect 65300 24676 65309 24716
rect 66403 24676 66412 24716
rect 66452 24676 72076 24716
rect 72116 24676 72125 24716
rect 50275 24632 50333 24633
rect 32419 24592 32428 24632
rect 32468 24592 33196 24632
rect 33236 24592 33245 24632
rect 34156 24592 36172 24632
rect 36212 24592 36940 24632
rect 36980 24592 36989 24632
rect 39907 24592 39916 24632
rect 39956 24592 41164 24632
rect 41204 24592 41213 24632
rect 42307 24592 42316 24632
rect 42356 24592 44428 24632
rect 44468 24592 44477 24632
rect 49699 24592 49708 24632
rect 49748 24592 50284 24632
rect 50324 24592 50380 24632
rect 50420 24592 50429 24632
rect 51331 24592 51340 24632
rect 51380 24592 52108 24632
rect 52148 24592 52157 24632
rect 52867 24592 52876 24632
rect 52916 24592 53548 24632
rect 53588 24592 56140 24632
rect 56180 24592 58636 24632
rect 58676 24592 58685 24632
rect 59011 24592 59020 24632
rect 59060 24592 59692 24632
rect 59732 24592 59884 24632
rect 59924 24592 59933 24632
rect 60451 24592 60460 24632
rect 60500 24592 61132 24632
rect 61172 24592 61181 24632
rect 63811 24592 63820 24632
rect 63860 24592 64780 24632
rect 64820 24592 64829 24632
rect 64963 24592 64972 24632
rect 65012 24592 65356 24632
rect 65396 24592 65405 24632
rect 65923 24592 65932 24632
rect 65972 24592 67660 24632
rect 67700 24592 67709 24632
rect 68131 24592 68140 24632
rect 68180 24592 68189 24632
rect 71011 24592 71020 24632
rect 71060 24592 71308 24632
rect 71348 24592 71357 24632
rect 74275 24592 74284 24632
rect 74324 24592 74764 24632
rect 74804 24592 74813 24632
rect 75715 24592 75724 24632
rect 75764 24592 76588 24632
rect 76628 24592 78988 24632
rect 79028 24592 79037 24632
rect 34156 24548 34196 24592
rect 50275 24591 50333 24592
rect 50371 24548 50429 24549
rect 68140 24548 68180 24592
rect 33859 24508 33868 24548
rect 33908 24508 34196 24548
rect 40195 24508 40204 24548
rect 40244 24508 40684 24548
rect 40724 24508 40733 24548
rect 40867 24508 40876 24548
rect 40916 24508 41068 24548
rect 41108 24508 41117 24548
rect 49603 24508 49612 24548
rect 49652 24508 49996 24548
rect 50036 24508 50045 24548
rect 50371 24508 50380 24548
rect 50420 24508 50860 24548
rect 50900 24508 51436 24548
rect 51476 24508 51820 24548
rect 51860 24508 56332 24548
rect 56372 24508 56381 24548
rect 64387 24508 64396 24548
rect 64436 24508 65644 24548
rect 65684 24508 68180 24548
rect 74467 24508 74476 24548
rect 74516 24508 75340 24548
rect 75380 24508 76396 24548
rect 76436 24508 76445 24548
rect 34156 24464 34196 24508
rect 50371 24507 50429 24508
rect 34147 24424 34156 24464
rect 34196 24424 34205 24464
rect 37027 24424 37036 24464
rect 37076 24424 39628 24464
rect 39668 24424 40012 24464
rect 40052 24424 40061 24464
rect 44899 24424 44908 24464
rect 44948 24424 45868 24464
rect 45908 24424 45917 24464
rect 50467 24424 50476 24464
rect 50516 24424 51532 24464
rect 51572 24424 51581 24464
rect 57187 24424 57196 24464
rect 57236 24424 62284 24464
rect 62324 24424 62333 24464
rect 62563 24424 62572 24464
rect 62612 24424 63052 24464
rect 63092 24424 63101 24464
rect 64675 24424 64684 24464
rect 64724 24424 65164 24464
rect 65204 24424 65213 24464
rect 75907 24424 75916 24464
rect 75956 24424 76108 24464
rect 76148 24424 76157 24464
rect 40099 24340 40108 24380
rect 40148 24340 41644 24380
rect 41684 24340 41693 24380
rect 43180 24340 57676 24380
rect 57716 24340 57725 24380
rect 59971 24340 59980 24380
rect 60020 24340 60364 24380
rect 60404 24340 60413 24380
rect 62467 24340 62476 24380
rect 62516 24340 66124 24380
rect 66164 24340 66173 24380
rect 43180 24296 43220 24340
rect 32707 24256 32716 24296
rect 32756 24256 35212 24296
rect 35252 24256 43220 24296
rect 44227 24256 44236 24296
rect 44276 24256 44716 24296
rect 44756 24256 45196 24296
rect 45236 24256 45388 24296
rect 45428 24256 45437 24296
rect 54019 24256 54028 24296
rect 54068 24256 62956 24296
rect 62996 24256 63005 24296
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 51811 24172 51820 24212
rect 51860 24172 62860 24212
rect 62900 24172 62909 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 35683 24088 35692 24128
rect 35732 24088 37516 24128
rect 37556 24088 39244 24128
rect 39284 24088 39293 24128
rect 48748 24088 62132 24128
rect 62179 24088 62188 24128
rect 62228 24088 65740 24128
rect 65780 24088 65789 24128
rect 0 24068 80 24088
rect 48748 24044 48788 24088
rect 52579 24044 52637 24045
rect 62092 24044 62132 24088
rect 43180 24004 46636 24044
rect 46676 24004 46685 24044
rect 48739 24004 48748 24044
rect 48788 24004 48797 24044
rect 50083 24004 50092 24044
rect 50132 24004 50764 24044
rect 50804 24004 50813 24044
rect 52579 24004 52588 24044
rect 52628 24004 52684 24044
rect 52724 24004 52733 24044
rect 55555 24004 55564 24044
rect 55604 24004 55756 24044
rect 55796 24004 55805 24044
rect 62083 24004 62092 24044
rect 62132 24004 62141 24044
rect 62275 24004 62284 24044
rect 62324 24004 65260 24044
rect 65300 24004 65644 24044
rect 65684 24004 65693 24044
rect 74083 24004 74092 24044
rect 74132 24004 74860 24044
rect 74900 24004 74909 24044
rect 40963 23960 41021 23961
rect 43180 23960 43220 24004
rect 52579 24003 52637 24004
rect 50563 23960 50621 23961
rect 29539 23920 29548 23960
rect 29588 23920 30892 23960
rect 30932 23920 35116 23960
rect 35156 23920 35165 23960
rect 36163 23920 36172 23960
rect 36212 23920 38860 23960
rect 38900 23920 38909 23960
rect 40867 23920 40876 23960
rect 40916 23920 40972 23960
rect 41012 23920 41021 23960
rect 41443 23920 41452 23960
rect 41492 23920 43220 23960
rect 44995 23920 45004 23960
rect 45044 23920 45196 23960
rect 45236 23920 46156 23960
rect 46196 23920 46205 23960
rect 50478 23920 50572 23960
rect 50612 23920 50621 23960
rect 50851 23920 50860 23960
rect 50900 23920 51244 23960
rect 51284 23920 51293 23960
rect 55843 23920 55852 23960
rect 55892 23920 57292 23960
rect 57332 23920 62900 23960
rect 63043 23920 63052 23960
rect 63092 23920 64876 23960
rect 64916 23920 65164 23960
rect 65204 23920 65213 23960
rect 68515 23920 68524 23960
rect 68564 23920 68908 23960
rect 68948 23920 68957 23960
rect 70147 23920 70156 23960
rect 70196 23920 70540 23960
rect 70580 23920 70828 23960
rect 70868 23920 70877 23960
rect 73123 23920 73132 23960
rect 73172 23920 73181 23960
rect 73315 23920 73324 23960
rect 73364 23920 73612 23960
rect 73652 23920 73804 23960
rect 73844 23920 73853 23960
rect 40963 23919 41021 23920
rect 50563 23919 50621 23920
rect 40483 23876 40541 23877
rect 835 23836 844 23876
rect 884 23836 1996 23876
rect 2036 23836 2045 23876
rect 32131 23836 32140 23876
rect 32180 23836 32716 23876
rect 32756 23836 32765 23876
rect 40398 23836 40492 23876
rect 40532 23836 40541 23876
rect 40675 23836 40684 23876
rect 40724 23836 41260 23876
rect 41300 23836 42220 23876
rect 42260 23836 50188 23876
rect 50228 23836 50237 23876
rect 50371 23836 50380 23876
rect 50420 23836 50956 23876
rect 50996 23836 51005 23876
rect 51532 23836 62476 23876
rect 62516 23836 62764 23876
rect 62804 23836 62813 23876
rect 40483 23835 40541 23836
rect 51139 23792 51197 23793
rect 51532 23792 51572 23836
rect 62860 23792 62900 23920
rect 73132 23876 73172 23920
rect 62947 23836 62956 23876
rect 62996 23836 64492 23876
rect 64532 23836 64780 23876
rect 64820 23836 64829 23876
rect 73132 23836 75244 23876
rect 75284 23836 75532 23876
rect 75572 23836 75581 23876
rect 79075 23792 79133 23793
rect 31651 23752 31660 23792
rect 31700 23752 32236 23792
rect 32276 23752 32285 23792
rect 36067 23752 36076 23792
rect 36116 23752 36652 23792
rect 36692 23752 37324 23792
rect 37364 23752 37373 23792
rect 38083 23752 38092 23792
rect 38132 23752 38764 23792
rect 38804 23752 40780 23792
rect 40820 23752 40829 23792
rect 44611 23752 44620 23792
rect 44660 23752 45964 23792
rect 46004 23752 46013 23792
rect 47587 23752 47596 23792
rect 47636 23752 48268 23792
rect 48308 23752 49324 23792
rect 49364 23752 49373 23792
rect 51054 23752 51148 23792
rect 51188 23752 51197 23792
rect 51523 23752 51532 23792
rect 51572 23752 51581 23792
rect 52099 23752 52108 23792
rect 52148 23752 52588 23792
rect 52628 23752 52637 23792
rect 54691 23752 54700 23792
rect 54740 23752 58060 23792
rect 58100 23752 58348 23792
rect 58388 23752 58397 23792
rect 62860 23752 67276 23792
rect 67316 23752 67564 23792
rect 67604 23752 67613 23792
rect 68707 23752 68716 23792
rect 68756 23752 70156 23792
rect 70196 23752 70444 23792
rect 70484 23752 70493 23792
rect 75043 23752 75052 23792
rect 75092 23752 76108 23792
rect 76148 23752 76492 23792
rect 76532 23752 76541 23792
rect 78990 23752 79084 23792
rect 79124 23752 79133 23792
rect 51139 23751 51197 23752
rect 79075 23751 79133 23752
rect 58435 23708 58493 23709
rect 31075 23668 31084 23708
rect 31124 23668 31468 23708
rect 31508 23668 33004 23708
rect 33044 23668 33053 23708
rect 41731 23668 41740 23708
rect 41780 23668 45004 23708
rect 45044 23668 45053 23708
rect 48067 23668 48076 23708
rect 48116 23668 50764 23708
rect 50804 23668 50813 23708
rect 58350 23668 58444 23708
rect 58484 23668 58493 23708
rect 67651 23668 67660 23708
rect 67700 23668 68044 23708
rect 68084 23668 68093 23708
rect 58435 23667 58493 23668
rect 56323 23624 56381 23625
rect 835 23584 844 23624
rect 884 23584 1420 23624
rect 1460 23584 1469 23624
rect 1795 23584 1804 23624
rect 1844 23584 2188 23624
rect 2228 23584 27380 23624
rect 36259 23584 36268 23624
rect 36308 23584 38956 23624
rect 38996 23584 39005 23624
rect 43939 23584 43948 23624
rect 43988 23584 44428 23624
rect 44468 23584 44477 23624
rect 50083 23584 50092 23624
rect 50132 23584 50141 23624
rect 51427 23584 51436 23624
rect 51476 23584 54124 23624
rect 54164 23584 56332 23624
rect 56372 23584 56381 23624
rect 27340 23540 27380 23584
rect 50092 23540 50132 23584
rect 56323 23583 56381 23584
rect 56515 23624 56573 23625
rect 70915 23624 70973 23625
rect 56515 23584 56524 23624
rect 56564 23584 63244 23624
rect 63284 23584 63628 23624
rect 63668 23584 63677 23624
rect 70830 23584 70924 23624
rect 70964 23584 71212 23624
rect 71252 23584 71261 23624
rect 74851 23584 74860 23624
rect 74900 23584 75244 23624
rect 75284 23584 75293 23624
rect 56515 23583 56573 23584
rect 70915 23583 70973 23584
rect 60547 23540 60605 23541
rect 27340 23500 43372 23540
rect 43412 23500 44524 23540
rect 44564 23500 44573 23540
rect 50092 23500 50228 23540
rect 40963 23456 41021 23457
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 31171 23416 31180 23456
rect 31220 23416 31372 23456
rect 31412 23416 31421 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 40099 23416 40108 23456
rect 40148 23416 40972 23456
rect 41012 23416 41021 23456
rect 44995 23416 45004 23456
rect 45044 23416 46060 23456
rect 46100 23416 46109 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 40963 23415 41021 23416
rect 50188 23372 50228 23500
rect 56524 23500 57292 23540
rect 57332 23500 57580 23540
rect 57620 23500 57629 23540
rect 57955 23500 57964 23540
rect 58004 23500 60076 23540
rect 60116 23500 60556 23540
rect 60596 23500 60605 23540
rect 56524 23456 56564 23500
rect 60547 23499 60605 23500
rect 56803 23456 56861 23457
rect 51811 23416 51820 23456
rect 51860 23416 56564 23456
rect 56611 23416 56620 23456
rect 56660 23416 56812 23456
rect 56852 23416 56861 23456
rect 57667 23416 57676 23456
rect 57716 23416 58060 23456
rect 58100 23416 58109 23456
rect 62851 23416 62860 23456
rect 62900 23416 63244 23456
rect 63284 23416 63293 23456
rect 78787 23416 78796 23456
rect 78836 23416 79276 23456
rect 79316 23416 79325 23456
rect 56803 23415 56861 23416
rect 56035 23372 56093 23373
rect 36259 23332 36268 23372
rect 36308 23332 37036 23372
rect 37076 23332 37085 23372
rect 46147 23332 46156 23372
rect 46196 23332 46636 23372
rect 46676 23332 46685 23372
rect 49996 23332 50228 23372
rect 50659 23332 50668 23372
rect 50708 23332 50717 23372
rect 50851 23332 50860 23372
rect 50900 23332 55892 23372
rect 55950 23332 56044 23372
rect 56084 23332 56093 23372
rect 0 23288 80 23308
rect 49996 23288 50036 23332
rect 50668 23288 50708 23332
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 32611 23248 32620 23288
rect 32660 23248 32908 23288
rect 32948 23248 32957 23288
rect 36835 23248 36844 23288
rect 36884 23248 37900 23288
rect 37940 23248 37949 23288
rect 40867 23248 40876 23288
rect 40916 23248 41356 23288
rect 41396 23248 41405 23288
rect 44899 23248 44908 23288
rect 44948 23248 44957 23288
rect 49027 23248 49036 23288
rect 49076 23248 49996 23288
rect 50036 23248 50045 23288
rect 50091 23248 50100 23288
rect 50140 23248 50708 23288
rect 52771 23248 52780 23288
rect 52820 23248 54316 23288
rect 54356 23248 54365 23288
rect 0 23228 80 23248
rect 44908 23204 44948 23248
rect 51139 23204 51197 23205
rect 55267 23204 55325 23205
rect 1507 23164 1516 23204
rect 1556 23164 2132 23204
rect 28963 23164 28972 23204
rect 29012 23164 29548 23204
rect 29588 23164 29597 23204
rect 32131 23164 32140 23204
rect 32180 23164 35788 23204
rect 35828 23164 37324 23204
rect 37364 23164 37652 23204
rect 41635 23164 41644 23204
rect 41684 23164 44620 23204
rect 44660 23164 46636 23204
rect 46676 23164 46685 23204
rect 50380 23164 50476 23204
rect 50516 23164 50764 23204
rect 50804 23164 50813 23204
rect 51139 23164 51148 23204
rect 51188 23164 51340 23204
rect 51380 23164 51389 23204
rect 52003 23164 52012 23204
rect 52052 23164 53644 23204
rect 53684 23164 53693 23204
rect 54787 23164 54796 23204
rect 54836 23164 55276 23204
rect 55316 23164 55325 23204
rect 55852 23204 55892 23332
rect 56035 23331 56093 23332
rect 56419 23288 56477 23289
rect 56334 23248 56428 23288
rect 56468 23248 56477 23288
rect 56419 23247 56477 23248
rect 55852 23164 56908 23204
rect 56948 23164 57196 23204
rect 57236 23164 57245 23204
rect 2092 23120 2132 23164
rect 1411 23080 1420 23120
rect 1460 23080 1900 23120
rect 1940 23080 1949 23120
rect 2083 23080 2092 23120
rect 2132 23080 4108 23120
rect 4148 23080 4780 23120
rect 4820 23080 4829 23120
rect 28387 23080 28396 23120
rect 28436 23080 31028 23120
rect 31171 23080 31180 23120
rect 31220 23080 31852 23120
rect 31892 23080 31901 23120
rect 32227 23080 32236 23120
rect 32276 23080 32716 23120
rect 32756 23080 32765 23120
rect 30988 22952 31028 23080
rect 37612 23060 37652 23164
rect 38467 23080 38476 23120
rect 38516 23080 39148 23120
rect 39188 23080 39197 23120
rect 45283 23080 45292 23120
rect 45332 23080 45484 23120
rect 45524 23080 48748 23120
rect 48788 23080 48797 23120
rect 48931 23080 48940 23120
rect 48980 23080 49900 23120
rect 49940 23080 50284 23120
rect 50324 23080 50333 23120
rect 31747 22996 31756 23036
rect 31796 22996 32140 23036
rect 32180 22996 32189 23036
rect 37603 23020 37612 23060
rect 37652 23020 37661 23060
rect 50380 23036 50420 23164
rect 51139 23163 51197 23164
rect 55267 23163 55325 23164
rect 52483 23120 52541 23121
rect 50659 23080 50668 23120
rect 50708 23080 51436 23120
rect 51476 23080 51485 23120
rect 52398 23080 52492 23120
rect 52532 23080 52541 23120
rect 52675 23080 52684 23120
rect 52724 23080 54604 23120
rect 54644 23080 54653 23120
rect 52483 23079 52541 23080
rect 45091 22996 45100 23036
rect 45140 22996 45580 23036
rect 45620 22996 45629 23036
rect 49795 22996 49804 23036
rect 49844 22996 50420 23036
rect 50563 23036 50621 23037
rect 50563 22996 50572 23036
rect 50612 22996 51244 23036
rect 51284 22996 51293 23036
rect 52195 22996 52204 23036
rect 52244 22996 54055 23036
rect 54095 22996 54104 23036
rect 50563 22995 50621 22996
rect 50764 22952 50804 22996
rect 53251 22952 53309 22953
rect 30979 22912 30988 22952
rect 31028 22912 31037 22952
rect 37123 22912 37132 22952
rect 37172 22912 37996 22952
rect 38036 22912 38045 22952
rect 41539 22912 41548 22952
rect 41588 22912 42028 22952
rect 42068 22912 42077 22952
rect 50755 22912 50764 22952
rect 50804 22912 50844 22952
rect 52291 22912 52300 22952
rect 52340 22912 52972 22952
rect 53012 22912 53021 22952
rect 53251 22912 53260 22952
rect 53300 22912 54455 22952
rect 54495 22912 54504 22952
rect 53251 22911 53309 22912
rect 58819 22868 58877 22869
rect 1699 22828 1708 22868
rect 1748 22828 2764 22868
rect 2804 22828 2813 22868
rect 52675 22828 52684 22868
rect 52724 22828 53545 22868
rect 53585 22828 53594 22868
rect 58819 22828 58828 22868
rect 58895 22828 58963 22868
rect 58819 22827 58877 22828
rect 54883 22784 54941 22785
rect 60547 22784 60605 22785
rect 52387 22744 52396 22784
rect 52436 22744 53945 22784
rect 53985 22744 53994 22784
rect 54846 22744 54855 22784
rect 54932 22744 54990 22784
rect 60432 22744 60455 22784
rect 60495 22744 60556 22784
rect 60596 22744 60605 22784
rect 78595 22744 78604 22784
rect 78644 22744 78855 22784
rect 78895 22744 78904 22784
rect 54883 22743 54941 22744
rect 60547 22743 60605 22744
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 36451 22576 36460 22616
rect 36500 22576 36748 22616
rect 36788 22576 37228 22616
rect 37268 22576 37277 22616
rect 43180 22576 51820 22616
rect 51860 22576 51869 22616
rect 30787 22532 30845 22533
rect 43180 22532 43220 22576
rect 28291 22492 28300 22532
rect 28340 22492 30796 22532
rect 30836 22492 30845 22532
rect 35203 22492 35212 22532
rect 35252 22492 43220 22532
rect 43555 22492 43564 22532
rect 43604 22492 47980 22532
rect 48020 22492 48029 22532
rect 50371 22492 50380 22532
rect 50420 22492 51148 22532
rect 51188 22492 51197 22532
rect 30787 22491 30845 22492
rect 0 22448 80 22468
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 27619 22408 27628 22448
rect 27668 22408 27916 22448
rect 27956 22408 30700 22448
rect 30740 22408 31564 22448
rect 31604 22408 32908 22448
rect 32948 22408 32957 22448
rect 0 22388 80 22408
rect 27715 22364 27773 22365
rect 27630 22324 27724 22364
rect 27764 22324 27773 22364
rect 28195 22324 28204 22364
rect 28244 22324 31180 22364
rect 31220 22324 31660 22364
rect 31700 22324 31709 22364
rect 27715 22323 27773 22324
rect 28483 22280 28541 22281
rect 28398 22240 28492 22280
rect 28532 22240 28541 22280
rect 29827 22240 29836 22280
rect 29876 22240 30604 22280
rect 30644 22240 31564 22280
rect 31604 22240 31613 22280
rect 31747 22240 31756 22280
rect 31796 22240 32332 22280
rect 32372 22240 32381 22280
rect 39235 22240 39244 22280
rect 39284 22240 40780 22280
rect 40820 22240 40829 22280
rect 42403 22240 42412 22280
rect 42452 22240 43660 22280
rect 43700 22240 43709 22280
rect 45475 22240 45484 22280
rect 45524 22240 46252 22280
rect 46292 22240 46301 22280
rect 46723 22240 46732 22280
rect 46772 22240 48556 22280
rect 48596 22240 50092 22280
rect 50132 22240 50141 22280
rect 52108 22240 52684 22280
rect 52724 22240 52733 22280
rect 28483 22239 28541 22240
rect 51907 22196 51965 22197
rect 52108 22196 52148 22240
rect 52579 22196 52637 22197
rect 32227 22156 32236 22196
rect 32276 22156 32812 22196
rect 32852 22156 32861 22196
rect 35683 22156 35692 22196
rect 35732 22156 36268 22196
rect 36308 22156 36317 22196
rect 38083 22156 38092 22196
rect 38132 22156 51916 22196
rect 51956 22156 51965 22196
rect 52099 22156 52108 22196
rect 52148 22156 52157 22196
rect 52494 22156 52588 22196
rect 52628 22156 52876 22196
rect 52916 22156 52925 22196
rect 51907 22155 51965 22156
rect 52579 22155 52637 22156
rect 38947 22112 39005 22113
rect 28675 22072 28684 22112
rect 28724 22072 29644 22112
rect 29684 22072 29693 22112
rect 30019 22072 30028 22112
rect 30068 22072 38956 22112
rect 38996 22072 40204 22112
rect 40244 22072 40253 22112
rect 38947 22071 39005 22072
rect 6979 21988 6988 22028
rect 7028 21988 52300 22028
rect 52340 21988 52349 22028
rect 27715 21944 27773 21945
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 27715 21904 27724 21944
rect 27764 21904 30028 21944
rect 30068 21904 30077 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 36163 21904 36172 21944
rect 36212 21904 36221 21944
rect 41347 21904 41356 21944
rect 41396 21904 43564 21944
rect 43604 21904 43613 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 27715 21903 27773 21904
rect 32899 21820 32908 21860
rect 32948 21820 32957 21860
rect 32908 21776 32948 21820
rect 36172 21776 36212 21904
rect 50371 21820 50380 21860
rect 50420 21820 50572 21860
rect 50612 21820 50621 21860
rect 29059 21736 29068 21776
rect 29108 21736 29117 21776
rect 32908 21736 36212 21776
rect 36547 21736 36556 21776
rect 36596 21736 36605 21776
rect 43180 21736 45292 21776
rect 45332 21736 45341 21776
rect 45667 21736 45676 21776
rect 45716 21736 45725 21776
rect 23203 21652 23212 21692
rect 23252 21652 28204 21692
rect 28244 21652 28253 21692
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 27811 21568 27820 21608
rect 27860 21568 28588 21608
rect 28628 21568 28637 21608
rect 28867 21568 28876 21608
rect 28916 21568 28925 21608
rect 0 21548 80 21568
rect 28876 21524 28916 21568
rect 1891 21484 1900 21524
rect 1940 21484 3052 21524
rect 3092 21484 3101 21524
rect 4003 21484 4012 21524
rect 4052 21484 4396 21524
rect 4436 21484 4445 21524
rect 26947 21484 26956 21524
rect 26996 21484 28916 21524
rect 29068 21440 29108 21736
rect 31459 21652 31468 21692
rect 31508 21652 32332 21692
rect 32372 21652 35212 21692
rect 35252 21652 35261 21692
rect 29443 21568 29452 21608
rect 29492 21568 32140 21608
rect 32180 21568 32620 21608
rect 32660 21568 35788 21608
rect 35828 21568 36076 21608
rect 36116 21568 36125 21608
rect 36172 21524 36212 21736
rect 36556 21692 36596 21736
rect 43180 21692 43220 21736
rect 36556 21652 36748 21692
rect 36788 21652 38092 21692
rect 38132 21652 38141 21692
rect 40675 21652 40684 21692
rect 40724 21652 41260 21692
rect 41300 21652 41309 21692
rect 42403 21652 42412 21692
rect 42452 21652 43220 21692
rect 44035 21608 44093 21609
rect 36259 21568 36268 21608
rect 36308 21568 36460 21608
rect 36500 21568 36509 21608
rect 39139 21568 39148 21608
rect 39188 21568 42508 21608
rect 42548 21568 42557 21608
rect 43950 21568 44044 21608
rect 44084 21568 44093 21608
rect 44803 21568 44812 21608
rect 44852 21568 45292 21608
rect 45332 21568 45341 21608
rect 44035 21567 44093 21568
rect 45676 21524 45716 21736
rect 99920 21692 100000 21726
rect 50371 21652 50380 21692
rect 50420 21652 51052 21692
rect 51092 21652 51101 21692
rect 99888 21652 100000 21692
rect 52291 21608 52349 21609
rect 53059 21608 53117 21609
rect 49027 21568 49036 21608
rect 49076 21568 49612 21608
rect 49652 21568 50956 21608
rect 50996 21568 51005 21608
rect 52206 21568 52300 21608
rect 52340 21568 52349 21608
rect 52579 21568 52588 21608
rect 52628 21568 53068 21608
rect 53108 21568 53117 21608
rect 99920 21586 100000 21652
rect 52291 21567 52349 21568
rect 53059 21567 53117 21568
rect 36163 21484 36172 21524
rect 36212 21484 36221 21524
rect 45379 21484 45388 21524
rect 45428 21484 45716 21524
rect 45859 21484 45868 21524
rect 45908 21484 49420 21524
rect 49460 21484 49469 21524
rect 50659 21484 50668 21524
rect 50708 21484 50860 21524
rect 50900 21484 50909 21524
rect 3235 21400 3244 21440
rect 3284 21400 3628 21440
rect 3668 21400 27148 21440
rect 27188 21400 27197 21440
rect 28483 21400 28492 21440
rect 28532 21400 31756 21440
rect 31796 21400 43220 21440
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 28003 21148 28012 21188
rect 28052 21148 28300 21188
rect 28340 21148 28349 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 43180 21104 43220 21400
rect 46540 21356 46580 21484
rect 50371 21440 50429 21441
rect 49507 21400 49516 21440
rect 49556 21400 50380 21440
rect 50420 21400 50429 21440
rect 50371 21399 50429 21400
rect 46531 21316 46540 21356
rect 46580 21316 46589 21356
rect 47683 21316 47692 21356
rect 47732 21316 48844 21356
rect 48884 21316 48893 21356
rect 45379 21232 45388 21272
rect 45428 21232 48364 21272
rect 48404 21232 51532 21272
rect 51572 21232 51581 21272
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 3619 21064 3628 21104
rect 3668 21064 3820 21104
rect 3860 21064 3869 21104
rect 38371 21064 38380 21104
rect 38420 21064 41588 21104
rect 43180 21064 50764 21104
rect 50804 21064 50813 21104
rect 41548 21020 41588 21064
rect 30307 20980 30316 21020
rect 30356 20980 40492 21020
rect 40532 20980 40541 21020
rect 41539 20980 41548 21020
rect 41588 20980 41597 21020
rect 50275 20980 50284 21020
rect 50324 20980 51916 21020
rect 51956 20980 52684 21020
rect 52724 20980 52733 21020
rect 26179 20896 26188 20936
rect 26228 20896 27532 20936
rect 27572 20896 27581 20936
rect 27724 20896 38380 20936
rect 38420 20896 38429 20936
rect 39043 20896 39052 20936
rect 39092 20896 42412 20936
rect 42452 20896 43948 20936
rect 43988 20896 45004 20936
rect 45044 20896 45053 20936
rect 27724 20852 27764 20896
rect 931 20812 940 20852
rect 980 20812 5068 20852
rect 5108 20812 5117 20852
rect 25891 20812 25900 20852
rect 25940 20812 26380 20852
rect 26420 20812 26429 20852
rect 27139 20812 27148 20852
rect 27188 20812 27764 20852
rect 28963 20812 28972 20852
rect 29012 20812 43084 20852
rect 43124 20812 43660 20852
rect 43700 20812 43709 20852
rect 0 20768 80 20788
rect 26380 20768 26420 20812
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 835 20728 844 20768
rect 884 20728 3532 20768
rect 3572 20728 3581 20768
rect 26380 20728 27340 20768
rect 27380 20728 27389 20768
rect 27619 20728 27628 20768
rect 27668 20728 27916 20768
rect 27956 20728 27965 20768
rect 28483 20728 28492 20768
rect 28532 20728 28876 20768
rect 28916 20728 28925 20768
rect 38467 20728 38476 20768
rect 38516 20728 38956 20768
rect 38996 20728 39005 20768
rect 39139 20728 39148 20768
rect 39188 20728 39436 20768
rect 39476 20728 39485 20768
rect 42499 20728 42508 20768
rect 42548 20728 44140 20768
rect 44180 20728 44908 20768
rect 44948 20728 44957 20768
rect 45475 20728 45484 20768
rect 45524 20728 46060 20768
rect 46100 20728 46109 20768
rect 0 20708 80 20728
rect 40867 20684 40925 20685
rect 4387 20644 4396 20684
rect 4436 20644 40876 20684
rect 40916 20644 40925 20684
rect 40867 20643 40925 20644
rect 3715 20560 3724 20600
rect 3764 20560 22828 20600
rect 22868 20560 22877 20600
rect 26659 20560 26668 20600
rect 26708 20560 26956 20600
rect 26996 20560 27005 20600
rect 27331 20560 27340 20600
rect 27380 20560 31372 20600
rect 31412 20560 39436 20600
rect 39476 20560 39485 20600
rect 42883 20560 42892 20600
rect 42932 20560 43084 20600
rect 43124 20560 43133 20600
rect 43180 20560 43276 20600
rect 43316 20560 43325 20600
rect 44995 20560 45004 20600
rect 45044 20560 52300 20600
rect 52340 20560 52349 20600
rect 43180 20516 43220 20560
rect 3619 20476 3628 20516
rect 3668 20476 5356 20516
rect 5396 20476 5405 20516
rect 30787 20476 30796 20516
rect 30836 20476 32716 20516
rect 32756 20476 36076 20516
rect 36116 20476 36125 20516
rect 42787 20476 42796 20516
rect 42836 20476 43220 20516
rect 51619 20476 51628 20516
rect 51668 20476 52588 20516
rect 52628 20476 52637 20516
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 32515 20224 32524 20264
rect 32564 20224 32573 20264
rect 37603 20224 37612 20264
rect 37652 20224 38284 20264
rect 38324 20224 38333 20264
rect 32524 20180 32564 20224
rect 25507 20140 25516 20180
rect 25556 20140 26764 20180
rect 26804 20140 27820 20180
rect 27860 20140 27869 20180
rect 32524 20140 33004 20180
rect 33044 20140 33053 20180
rect 39331 20140 39340 20180
rect 39380 20140 40972 20180
rect 41012 20140 41021 20180
rect 43075 20140 43084 20180
rect 43124 20140 43276 20180
rect 43316 20140 43325 20180
rect 44899 20140 44908 20180
rect 44948 20140 47212 20180
rect 47252 20140 47596 20180
rect 47636 20140 48940 20180
rect 48980 20140 50860 20180
rect 50900 20140 51532 20180
rect 51572 20140 51581 20180
rect 33859 20096 33917 20097
rect 2659 20056 2668 20096
rect 2708 20056 11116 20096
rect 11156 20056 11165 20096
rect 11683 20056 11692 20096
rect 11732 20056 17300 20096
rect 26563 20056 26572 20096
rect 26612 20056 29548 20096
rect 29588 20056 29597 20096
rect 33859 20056 33868 20096
rect 33908 20056 39148 20096
rect 39188 20056 39197 20096
rect 44227 20056 44236 20096
rect 44276 20056 45676 20096
rect 45716 20056 45725 20096
rect 17260 20012 17300 20056
rect 33859 20055 33917 20056
rect 99920 20012 100000 20089
rect 1987 19972 1996 20012
rect 2036 19972 10828 20012
rect 10868 19972 10877 20012
rect 17260 19972 26420 20012
rect 42595 19972 42604 20012
rect 42644 19972 43084 20012
rect 43124 19972 43852 20012
rect 43892 19972 43901 20012
rect 44323 19972 44332 20012
rect 44372 19972 45292 20012
rect 45332 19972 45341 20012
rect 99888 19972 100000 20012
rect 0 19928 80 19948
rect 26380 19928 26420 19972
rect 99920 19949 100000 19972
rect 41731 19928 41789 19929
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 26371 19888 26380 19928
rect 26420 19888 26429 19928
rect 26563 19888 26572 19928
rect 26612 19888 26956 19928
rect 26996 19888 27005 19928
rect 32899 19888 32908 19928
rect 32948 19888 34444 19928
rect 34484 19888 34828 19928
rect 34868 19888 34877 19928
rect 36259 19888 36268 19928
rect 36308 19888 37708 19928
rect 37748 19888 37757 19928
rect 38083 19888 38092 19928
rect 38132 19888 38141 19928
rect 38275 19888 38284 19928
rect 38324 19888 38668 19928
rect 38708 19888 38717 19928
rect 40771 19888 40780 19928
rect 40820 19888 41740 19928
rect 41780 19888 41789 19928
rect 44035 19888 44044 19928
rect 44084 19888 44716 19928
rect 44756 19888 44765 19928
rect 0 19868 80 19888
rect 38092 19844 38132 19888
rect 41731 19887 41789 19888
rect 4867 19804 4876 19844
rect 4916 19804 21772 19844
rect 21812 19804 21821 19844
rect 23491 19804 23500 19844
rect 23540 19804 23692 19844
rect 23732 19804 28972 19844
rect 29012 19804 29021 19844
rect 29539 19804 29548 19844
rect 29588 19804 35020 19844
rect 35060 19804 37516 19844
rect 37556 19804 38132 19844
rect 38467 19804 38476 19844
rect 38516 19804 39052 19844
rect 39092 19804 39101 19844
rect 42691 19804 42700 19844
rect 42740 19804 42988 19844
rect 43028 19804 43037 19844
rect 5059 19720 5068 19760
rect 5108 19720 43276 19760
rect 43316 19720 43325 19760
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 34915 19636 34924 19676
rect 34964 19636 37900 19676
rect 37940 19636 39532 19676
rect 39572 19636 39581 19676
rect 40387 19636 40396 19676
rect 40436 19636 42508 19676
rect 42548 19636 42557 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 48931 19636 48940 19676
rect 48980 19636 49612 19676
rect 49652 19636 49661 19676
rect 34924 19592 34964 19636
rect 9571 19552 9580 19592
rect 9620 19552 10924 19592
rect 10964 19552 10973 19592
rect 32995 19552 33004 19592
rect 33044 19552 34964 19592
rect 40771 19552 40780 19592
rect 40820 19552 41644 19592
rect 41684 19552 41693 19592
rect 44515 19552 44524 19592
rect 44564 19552 51532 19592
rect 51572 19552 51581 19592
rect 51811 19508 51869 19509
rect 14659 19468 14668 19508
rect 14708 19468 51820 19508
rect 51860 19468 51869 19508
rect 51811 19467 51869 19468
rect 39331 19424 39389 19425
rect 29059 19384 29068 19424
rect 29108 19384 29260 19424
rect 29300 19384 29309 19424
rect 32035 19384 32044 19424
rect 32084 19384 32093 19424
rect 32899 19384 32908 19424
rect 32948 19384 33292 19424
rect 33332 19384 33341 19424
rect 39331 19384 39340 19424
rect 39380 19384 39436 19424
rect 39476 19384 39485 19424
rect 41251 19384 41260 19424
rect 41300 19384 41932 19424
rect 41972 19384 41981 19424
rect 43180 19384 47500 19424
rect 47540 19384 49652 19424
rect 21763 19300 21772 19340
rect 21812 19300 27724 19340
rect 27764 19300 27773 19340
rect 30211 19300 30220 19340
rect 30260 19300 31660 19340
rect 31700 19300 31852 19340
rect 31892 19300 31901 19340
rect 10051 19216 10060 19256
rect 10100 19216 13516 19256
rect 13556 19216 31084 19256
rect 31124 19216 31133 19256
rect 11875 19132 11884 19172
rect 11924 19132 12268 19172
rect 12308 19132 12317 19172
rect 22339 19132 22348 19172
rect 22388 19132 25900 19172
rect 25940 19132 29012 19172
rect 29059 19132 29068 19172
rect 29108 19132 29932 19172
rect 29972 19132 29981 19172
rect 0 19088 80 19108
rect 22540 19088 22580 19132
rect 28972 19088 29012 19132
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 22531 19048 22540 19088
rect 22580 19048 22620 19088
rect 25411 19048 25420 19088
rect 25460 19048 26476 19088
rect 26516 19048 26525 19088
rect 28972 19048 30124 19088
rect 30164 19048 31948 19088
rect 31988 19048 31997 19088
rect 0 19028 80 19048
rect 32044 19004 32084 19384
rect 39331 19383 39389 19384
rect 43180 19340 43220 19384
rect 40387 19300 40396 19340
rect 40436 19300 43220 19340
rect 45283 19300 45292 19340
rect 45332 19300 49268 19340
rect 38947 19216 38956 19256
rect 38996 19216 39436 19256
rect 39476 19216 39485 19256
rect 40972 19088 41012 19300
rect 42307 19216 42316 19256
rect 42356 19216 42796 19256
rect 42836 19216 42845 19256
rect 49027 19216 49036 19256
rect 49076 19216 49085 19256
rect 41443 19132 41452 19172
rect 41492 19132 42124 19172
rect 42164 19132 42173 19172
rect 40963 19048 40972 19088
rect 41012 19048 41021 19088
rect 43660 19048 44620 19088
rect 44660 19048 44669 19088
rect 21955 18964 21964 19004
rect 22004 18964 22252 19004
rect 22292 18964 25804 19004
rect 25844 18964 29452 19004
rect 29492 18964 30028 19004
rect 30068 18964 30077 19004
rect 31843 18964 31852 19004
rect 31892 18964 32084 19004
rect 43660 18920 43700 19048
rect 49036 18920 49076 19216
rect 49228 18920 49268 19300
rect 49612 18920 49652 19384
rect 51715 19088 51773 19089
rect 51715 19048 51724 19088
rect 51764 19048 52012 19088
rect 52052 19048 52061 19088
rect 51715 19047 51773 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 24451 18880 24460 18920
rect 24500 18880 30316 18920
rect 30356 18880 30365 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 43075 18880 43084 18920
rect 43124 18880 43700 18920
rect 43843 18880 43852 18920
rect 43892 18880 44332 18920
rect 44372 18880 44381 18920
rect 49027 18880 49036 18920
rect 49076 18880 49085 18920
rect 49219 18880 49228 18920
rect 49268 18880 49277 18920
rect 49603 18880 49612 18920
rect 49652 18880 49661 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 50563 18836 50621 18837
rect 25987 18796 25996 18836
rect 26036 18796 27244 18836
rect 27284 18796 28588 18836
rect 28628 18796 28637 18836
rect 36268 18796 50572 18836
rect 50612 18796 50621 18836
rect 36268 18752 36308 18796
rect 50563 18795 50621 18796
rect 51715 18752 51773 18753
rect 8899 18712 8908 18752
rect 8948 18712 11020 18752
rect 11060 18712 11069 18752
rect 22435 18712 22444 18752
rect 22484 18712 23020 18752
rect 23060 18712 25036 18752
rect 25076 18712 25085 18752
rect 25699 18712 25708 18752
rect 25748 18712 26188 18752
rect 26228 18712 26237 18752
rect 28963 18712 28972 18752
rect 29012 18712 29740 18752
rect 29780 18712 29789 18752
rect 32227 18712 32236 18752
rect 32276 18712 32620 18752
rect 32660 18712 33868 18752
rect 33908 18712 33917 18752
rect 35308 18712 36308 18752
rect 39427 18712 39436 18752
rect 39476 18712 41164 18752
rect 41204 18712 41213 18752
rect 42019 18712 42028 18752
rect 42068 18712 43660 18752
rect 43700 18712 44140 18752
rect 44180 18712 44189 18752
rect 48643 18712 48652 18752
rect 48692 18712 49036 18752
rect 49076 18712 51724 18752
rect 51764 18712 51773 18752
rect 35308 18668 35348 18712
rect 51715 18711 51773 18712
rect 7180 18628 12076 18668
rect 12116 18628 24844 18668
rect 24884 18628 24893 18668
rect 26284 18628 26860 18668
rect 26900 18628 30700 18668
rect 30740 18628 33004 18668
rect 33044 18628 33053 18668
rect 33187 18628 33196 18668
rect 33236 18628 35308 18668
rect 35348 18628 35357 18668
rect 35779 18628 35788 18668
rect 35828 18628 36172 18668
rect 36212 18628 36221 18668
rect 38371 18628 38380 18668
rect 38420 18628 40204 18668
rect 40244 18628 40253 18668
rect 42595 18628 42604 18668
rect 42644 18628 43180 18668
rect 43220 18628 44428 18668
rect 44468 18628 44477 18668
rect 44611 18628 44620 18668
rect 44660 18628 45196 18668
rect 45236 18628 46060 18668
rect 46100 18628 46109 18668
rect 46828 18628 49132 18668
rect 49172 18628 49324 18668
rect 49364 18628 49373 18668
rect 7180 18584 7220 18628
rect 26284 18584 26324 18628
rect 46828 18584 46868 18628
rect 4867 18544 4876 18584
rect 4916 18544 5356 18584
rect 5396 18544 7220 18584
rect 22147 18544 22156 18584
rect 22196 18544 23404 18584
rect 23444 18544 26324 18584
rect 26371 18544 26380 18584
rect 26420 18544 26764 18584
rect 26804 18544 27820 18584
rect 27860 18544 27869 18584
rect 31171 18544 31180 18584
rect 31220 18544 31660 18584
rect 31700 18544 34252 18584
rect 34292 18544 34301 18584
rect 35683 18544 35692 18584
rect 35732 18544 38612 18584
rect 38659 18544 38668 18584
rect 38708 18544 40012 18584
rect 40052 18544 41068 18584
rect 41108 18544 41117 18584
rect 42115 18544 42124 18584
rect 42164 18544 42796 18584
rect 42836 18544 42845 18584
rect 43939 18544 43948 18584
rect 43988 18544 45484 18584
rect 45524 18544 45533 18584
rect 46819 18544 46828 18584
rect 46868 18544 46877 18584
rect 47683 18544 47692 18584
rect 47732 18544 48844 18584
rect 48884 18544 48893 18584
rect 22339 18500 22397 18501
rect 23683 18500 23741 18501
rect 38572 18500 38612 18544
rect 52387 18500 52445 18501
rect 1699 18460 1708 18500
rect 1748 18460 10924 18500
rect 10964 18460 12268 18500
rect 12308 18460 14668 18500
rect 14708 18460 14717 18500
rect 22254 18460 22348 18500
rect 22388 18460 22397 18500
rect 22339 18459 22397 18460
rect 23020 18460 23692 18500
rect 23732 18460 23741 18500
rect 24835 18460 24844 18500
rect 24884 18460 26092 18500
rect 26132 18460 26141 18500
rect 28963 18460 28972 18500
rect 29012 18460 32140 18500
rect 32180 18460 32189 18500
rect 32323 18460 32332 18500
rect 32372 18460 34156 18500
rect 34196 18460 35500 18500
rect 35540 18460 36460 18500
rect 36500 18460 37420 18500
rect 37460 18460 37469 18500
rect 38563 18460 38572 18500
rect 38612 18460 40396 18500
rect 40436 18460 40445 18500
rect 42883 18460 42892 18500
rect 42932 18460 43084 18500
rect 43124 18460 43133 18500
rect 47491 18460 47500 18500
rect 47540 18460 47788 18500
rect 47828 18460 47837 18500
rect 49795 18460 49804 18500
rect 49844 18460 50572 18500
rect 50612 18460 50621 18500
rect 51523 18460 51532 18500
rect 51572 18460 52396 18500
rect 52436 18460 52445 18500
rect 23020 18416 23060 18460
rect 23683 18459 23741 18460
rect 28972 18416 29012 18460
rect 52387 18459 52445 18460
rect 4099 18376 4108 18416
rect 4148 18376 23060 18416
rect 25507 18376 25516 18416
rect 25556 18376 29012 18416
rect 32419 18376 32428 18416
rect 32468 18376 35692 18416
rect 35732 18376 35741 18416
rect 41539 18376 41548 18416
rect 41588 18376 42028 18416
rect 42068 18376 42508 18416
rect 42548 18376 42557 18416
rect 46243 18376 46252 18416
rect 46292 18376 47020 18416
rect 47060 18376 47069 18416
rect 21955 18292 21964 18332
rect 22004 18292 22924 18332
rect 22964 18292 22973 18332
rect 23971 18292 23980 18332
rect 24020 18292 24748 18332
rect 24788 18292 27436 18332
rect 27476 18292 28396 18332
rect 28436 18292 30508 18332
rect 30548 18292 31564 18332
rect 31604 18292 31613 18332
rect 42211 18292 42220 18332
rect 42260 18292 42412 18332
rect 42452 18292 42461 18332
rect 42883 18292 42892 18332
rect 42932 18292 46828 18332
rect 46868 18292 46877 18332
rect 50467 18292 50476 18332
rect 50516 18292 51340 18332
rect 51380 18292 51389 18332
rect 0 18248 80 18268
rect 50371 18248 50429 18249
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 24259 18208 24268 18248
rect 24308 18208 27916 18248
rect 27956 18208 29644 18248
rect 29684 18208 32812 18248
rect 32852 18208 32861 18248
rect 36355 18208 36364 18248
rect 36404 18208 36652 18248
rect 36692 18208 38572 18248
rect 38612 18208 50380 18248
rect 50420 18208 50429 18248
rect 0 18188 80 18208
rect 50371 18207 50429 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 23875 18124 23884 18164
rect 23924 18124 24076 18164
rect 24116 18124 31852 18164
rect 31892 18124 31901 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 41635 18124 41644 18164
rect 41684 18124 42124 18164
rect 42164 18124 42892 18164
rect 42932 18124 42941 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 24547 18040 24556 18080
rect 24596 18040 29356 18080
rect 29396 18040 29405 18080
rect 43075 18040 43084 18080
rect 43124 18040 43220 18080
rect 46819 18040 46828 18080
rect 46868 18040 49516 18080
rect 49556 18040 49565 18080
rect 29356 17912 29396 18040
rect 43180 17996 43220 18040
rect 52003 17996 52061 17997
rect 32707 17956 32716 17996
rect 32756 17956 33388 17996
rect 33428 17956 33437 17996
rect 36460 17956 37036 17996
rect 37076 17956 38284 17996
rect 38324 17956 38333 17996
rect 41731 17956 41740 17996
rect 41780 17956 41789 17996
rect 43180 17956 51244 17996
rect 51284 17956 52012 17996
rect 52052 17956 52061 17996
rect 36460 17912 36500 17956
rect 41740 17912 41780 17956
rect 52003 17955 52061 17956
rect 29356 17872 33140 17912
rect 36451 17872 36460 17912
rect 36500 17872 36509 17912
rect 41740 17872 46484 17912
rect 33100 17828 33140 17872
rect 46444 17828 46484 17872
rect 22732 17788 24268 17828
rect 24308 17788 24317 17828
rect 31372 17788 32428 17828
rect 32468 17788 32477 17828
rect 33100 17788 34348 17828
rect 34388 17788 34397 17828
rect 36835 17788 36844 17828
rect 36884 17788 38956 17828
rect 38996 17788 39005 17828
rect 42595 17788 42604 17828
rect 42644 17788 43948 17828
rect 43988 17788 43997 17828
rect 46435 17788 46444 17828
rect 46484 17788 48940 17828
rect 48980 17788 48989 17828
rect 49507 17788 49516 17828
rect 49556 17788 49804 17828
rect 49844 17788 49853 17828
rect 22732 17744 22772 17788
rect 31372 17744 31412 17788
rect 22723 17704 22732 17744
rect 22772 17704 22781 17744
rect 22915 17704 22924 17744
rect 22964 17704 23692 17744
rect 23732 17704 23741 17744
rect 29827 17704 29836 17744
rect 29876 17704 31372 17744
rect 31412 17704 31421 17744
rect 31555 17704 31564 17744
rect 31604 17704 32332 17744
rect 32372 17704 32381 17744
rect 33187 17704 33196 17744
rect 33236 17704 33484 17744
rect 33524 17704 33533 17744
rect 39811 17704 39820 17744
rect 39860 17704 41932 17744
rect 41972 17704 41981 17744
rect 42787 17704 42796 17744
rect 42836 17704 44044 17744
rect 44084 17704 44093 17744
rect 45955 17704 45964 17744
rect 46004 17704 46252 17744
rect 46292 17704 46540 17744
rect 46580 17704 48748 17744
rect 48788 17704 48797 17744
rect 49603 17704 49612 17744
rect 49652 17704 49661 17744
rect 50083 17704 50092 17744
rect 50132 17704 50380 17744
rect 50420 17704 51916 17744
rect 51956 17704 51965 17744
rect 29836 17660 29876 17704
rect 49612 17660 49652 17704
rect 52195 17660 52253 17661
rect 23203 17620 23212 17660
rect 23252 17620 26668 17660
rect 26708 17620 29876 17660
rect 29923 17620 29932 17660
rect 29972 17620 30316 17660
rect 30356 17620 30365 17660
rect 32131 17620 32140 17660
rect 32180 17620 34388 17660
rect 42691 17620 42700 17660
rect 42740 17620 43084 17660
rect 43124 17620 43133 17660
rect 45571 17620 45580 17660
rect 45620 17620 45660 17660
rect 49612 17620 51148 17660
rect 51188 17620 51197 17660
rect 52195 17620 52204 17660
rect 52244 17620 53068 17660
rect 53108 17620 53117 17660
rect 25795 17576 25853 17577
rect 29539 17576 29597 17577
rect 34348 17576 34388 17620
rect 45580 17576 45620 17620
rect 52195 17619 52253 17620
rect 23107 17536 23116 17576
rect 23156 17536 23596 17576
rect 23636 17536 25804 17576
rect 25844 17536 25853 17576
rect 27427 17536 27436 17576
rect 27476 17536 29548 17576
rect 29588 17536 29597 17576
rect 34339 17536 34348 17576
rect 34388 17536 34397 17576
rect 44899 17536 44908 17576
rect 44948 17536 50476 17576
rect 50516 17536 50525 17576
rect 25795 17535 25853 17536
rect 29539 17535 29597 17536
rect 49603 17492 49661 17493
rect 53059 17492 53117 17493
rect 23779 17452 23788 17492
rect 23828 17452 25324 17492
rect 25364 17452 27244 17492
rect 27284 17452 28780 17492
rect 28820 17452 30220 17492
rect 30260 17452 31756 17492
rect 31796 17452 36844 17492
rect 36884 17452 36893 17492
rect 45571 17452 45580 17492
rect 45620 17452 47500 17492
rect 47540 17452 47549 17492
rect 49603 17452 49612 17492
rect 49652 17452 52300 17492
rect 52340 17452 53068 17492
rect 53108 17452 53117 17492
rect 49603 17451 49661 17452
rect 53059 17451 53117 17452
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 21955 17368 21964 17408
rect 22004 17368 31276 17408
rect 31316 17368 31325 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 45475 17368 45484 17408
rect 45524 17368 47596 17408
rect 47636 17368 47645 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 50668 17368 52492 17408
rect 52532 17368 52684 17408
rect 52724 17368 52733 17408
rect 0 17348 80 17368
rect 32707 17324 32765 17325
rect 41155 17324 41213 17325
rect 50668 17324 50708 17368
rect 30403 17284 30412 17324
rect 30452 17284 30604 17324
rect 30644 17284 32716 17324
rect 32756 17284 32765 17324
rect 32899 17284 32908 17324
rect 32948 17284 33964 17324
rect 34004 17284 35116 17324
rect 35156 17284 35596 17324
rect 35636 17284 38284 17324
rect 38324 17284 38333 17324
rect 41070 17284 41164 17324
rect 41204 17284 41213 17324
rect 49411 17284 49420 17324
rect 49460 17284 50668 17324
rect 50708 17284 50717 17324
rect 52579 17284 52588 17324
rect 52628 17284 53545 17324
rect 53585 17284 53594 17324
rect 32707 17283 32765 17284
rect 41155 17283 41213 17284
rect 51619 17240 51677 17241
rect 53923 17240 53981 17241
rect 55075 17240 55133 17241
rect 55459 17240 55517 17241
rect 55651 17240 55709 17241
rect 58243 17240 58301 17241
rect 42211 17200 42220 17240
rect 42260 17200 42300 17240
rect 42979 17200 42988 17240
rect 43028 17200 44332 17240
rect 44372 17200 47500 17240
rect 47540 17200 47549 17240
rect 49603 17200 49612 17240
rect 49652 17200 49661 17240
rect 50371 17200 50380 17240
rect 50420 17200 51436 17240
rect 51476 17200 51485 17240
rect 51619 17200 51628 17240
rect 51668 17200 51762 17240
rect 52771 17200 52780 17240
rect 52820 17200 53655 17240
rect 53695 17200 53704 17240
rect 53923 17200 53932 17240
rect 53985 17200 54067 17240
rect 54960 17200 54988 17240
rect 55028 17200 55084 17240
rect 55124 17200 55145 17240
rect 55185 17200 55219 17240
rect 55459 17200 55468 17240
rect 55508 17200 55545 17240
rect 55585 17200 55603 17240
rect 55651 17200 55660 17240
rect 55700 17200 55945 17240
rect 55985 17200 55994 17240
rect 58243 17200 58252 17240
rect 58292 17200 58345 17240
rect 58385 17200 58394 17240
rect 42220 17156 42260 17200
rect 49612 17156 49652 17200
rect 51619 17199 51677 17200
rect 53923 17199 53981 17200
rect 55075 17199 55133 17200
rect 55459 17199 55517 17200
rect 55651 17199 55709 17200
rect 58243 17199 58301 17200
rect 51907 17156 51965 17157
rect 52579 17156 52637 17157
rect 53059 17156 53117 17157
rect 57859 17156 57917 17157
rect 2371 17116 2380 17156
rect 2420 17116 3340 17156
rect 3380 17116 23500 17156
rect 23540 17116 23549 17156
rect 30115 17116 30124 17156
rect 30164 17116 30508 17156
rect 30548 17116 30557 17156
rect 34051 17116 34060 17156
rect 34100 17116 38092 17156
rect 38132 17116 38141 17156
rect 41923 17116 41932 17156
rect 41972 17116 42604 17156
rect 42644 17116 42653 17156
rect 45763 17116 45772 17156
rect 45812 17116 46156 17156
rect 46196 17116 46205 17156
rect 49219 17116 49228 17156
rect 49268 17116 51724 17156
rect 51764 17116 51773 17156
rect 51907 17116 51916 17156
rect 51956 17116 52300 17156
rect 52340 17116 52349 17156
rect 52494 17116 52588 17156
rect 52628 17116 52876 17156
rect 52916 17116 52925 17156
rect 53059 17116 53068 17156
rect 53108 17116 54345 17156
rect 54385 17116 54394 17156
rect 54446 17116 54455 17156
rect 54495 17116 54548 17156
rect 51907 17115 51965 17116
rect 52579 17115 52637 17116
rect 53059 17115 53117 17116
rect 54508 17072 54548 17116
rect 57859 17116 57868 17156
rect 57908 17116 57945 17156
rect 57985 17116 58003 17156
rect 60736 17116 60745 17156
rect 60785 17116 60940 17156
rect 60980 17116 60989 17156
rect 64579 17116 64588 17156
rect 64628 17116 64855 17156
rect 64895 17116 64904 17156
rect 66595 17116 66604 17156
rect 66644 17116 66855 17156
rect 66895 17116 66904 17156
rect 71395 17116 71404 17156
rect 71444 17116 71655 17156
rect 71695 17116 71704 17156
rect 78979 17116 78988 17156
rect 79028 17116 79372 17156
rect 79412 17116 79655 17156
rect 79695 17116 79704 17156
rect 57859 17115 57917 17116
rect 4195 17032 4204 17072
rect 4244 17032 4588 17072
rect 4628 17032 5164 17072
rect 5204 17032 5213 17072
rect 33571 17032 33580 17072
rect 33620 17032 34100 17072
rect 41059 17032 41068 17072
rect 41108 17032 41836 17072
rect 41876 17032 41885 17072
rect 42883 17032 42892 17072
rect 42932 17032 43948 17072
rect 43988 17032 43997 17072
rect 44707 17032 44716 17072
rect 44756 17032 45388 17072
rect 45428 17032 47020 17072
rect 47060 17032 48364 17072
rect 48404 17032 48413 17072
rect 49987 17032 49996 17072
rect 50036 17032 50764 17072
rect 50804 17032 50813 17072
rect 51043 17032 51052 17072
rect 51092 17032 51628 17072
rect 51668 17032 51677 17072
rect 52387 17032 52396 17072
rect 52436 17032 54548 17072
rect 23395 16948 23404 16988
rect 23444 16948 24556 16988
rect 24596 16948 24605 16988
rect 22339 16904 22397 16905
rect 2179 16864 2188 16904
rect 2228 16864 2956 16904
rect 2996 16864 22348 16904
rect 22388 16864 22397 16904
rect 22339 16863 22397 16864
rect 34060 16820 34100 17032
rect 41443 16948 41452 16988
rect 41492 16948 43124 16988
rect 45091 16948 45100 16988
rect 45140 16948 45180 16988
rect 45667 16948 45676 16988
rect 45716 16948 48652 16988
rect 48692 16948 50804 16988
rect 52483 16948 52492 16988
rect 52532 16948 65356 16988
rect 65396 16948 65405 16988
rect 39715 16904 39773 16905
rect 43084 16904 43124 16948
rect 45100 16904 45140 16948
rect 50764 16904 50804 16948
rect 37123 16864 37132 16904
rect 37172 16864 39724 16904
rect 39764 16864 39773 16904
rect 43075 16864 43084 16904
rect 43124 16864 43133 16904
rect 43747 16864 43756 16904
rect 43796 16864 44140 16904
rect 44180 16864 47308 16904
rect 47348 16864 47357 16904
rect 49891 16864 49900 16904
rect 49940 16864 50188 16904
rect 50228 16864 50668 16904
rect 50708 16864 50717 16904
rect 50764 16864 64684 16904
rect 64724 16864 64733 16904
rect 39715 16863 39773 16864
rect 36643 16820 36701 16821
rect 34060 16780 36652 16820
rect 36692 16780 36701 16820
rect 46051 16780 46060 16820
rect 46100 16780 47116 16820
rect 47156 16780 47165 16820
rect 50467 16780 50476 16820
rect 50516 16780 51244 16820
rect 51284 16780 51293 16820
rect 52387 16780 52396 16820
rect 52436 16780 54028 16820
rect 54068 16780 54077 16820
rect 34060 16736 34100 16780
rect 36643 16779 36701 16780
rect 50476 16736 50516 16780
rect 34051 16696 34060 16736
rect 34100 16696 34109 16736
rect 43363 16696 43372 16736
rect 43412 16696 44524 16736
rect 44564 16696 50516 16736
rect 51907 16696 51916 16736
rect 51956 16696 53068 16736
rect 53108 16696 53117 16736
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 4003 16612 4012 16652
rect 4052 16612 5068 16652
rect 5108 16612 11788 16652
rect 11828 16612 11837 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 43075 16612 43084 16652
rect 43124 16612 43220 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 52483 16612 52492 16652
rect 52532 16612 53740 16652
rect 53780 16612 53789 16652
rect 0 16568 80 16588
rect 43180 16568 43220 16612
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 2563 16528 2572 16568
rect 2612 16528 10636 16568
rect 10676 16528 10685 16568
rect 43180 16528 47884 16568
rect 47924 16528 49612 16568
rect 49652 16528 51628 16568
rect 51668 16528 51677 16568
rect 52771 16528 52780 16568
rect 52820 16528 53300 16568
rect 0 16508 80 16528
rect 3340 16484 3380 16528
rect 51628 16484 51668 16528
rect 53260 16484 53300 16528
rect 3331 16444 3340 16484
rect 3380 16444 3420 16484
rect 4387 16444 4396 16484
rect 4436 16444 6988 16484
rect 7028 16444 7037 16484
rect 33859 16444 33868 16484
rect 33908 16444 34252 16484
rect 34292 16444 34732 16484
rect 34772 16444 34781 16484
rect 37315 16444 37324 16484
rect 37364 16444 37996 16484
rect 38036 16444 38045 16484
rect 39235 16444 39244 16484
rect 39284 16444 42412 16484
rect 42452 16444 44140 16484
rect 44180 16444 44189 16484
rect 51628 16444 52916 16484
rect 53260 16444 55564 16484
rect 55604 16444 55613 16484
rect 60835 16444 60844 16484
rect 60884 16444 61228 16484
rect 61268 16444 61277 16484
rect 52675 16400 52733 16401
rect 37507 16360 37516 16400
rect 37556 16360 38476 16400
rect 38516 16360 38525 16400
rect 42787 16360 42796 16400
rect 42836 16360 43084 16400
rect 43124 16360 43133 16400
rect 45091 16360 45100 16400
rect 45140 16360 46292 16400
rect 50563 16360 50572 16400
rect 50612 16360 51724 16400
rect 51764 16360 52684 16400
rect 52724 16360 52733 16400
rect 46252 16316 46292 16360
rect 52675 16359 52733 16360
rect 52876 16316 52916 16444
rect 53731 16360 53740 16400
rect 53780 16360 55468 16400
rect 55508 16360 65740 16400
rect 65780 16360 65789 16400
rect 61699 16316 61757 16317
rect 3811 16276 3820 16316
rect 3860 16276 4204 16316
rect 4244 16276 24460 16316
rect 24500 16276 24509 16316
rect 32995 16276 33004 16316
rect 33044 16276 33772 16316
rect 33812 16276 36844 16316
rect 36884 16276 40108 16316
rect 40148 16276 40157 16316
rect 42499 16276 42508 16316
rect 42548 16276 43173 16316
rect 43213 16276 45292 16316
rect 45332 16276 45341 16316
rect 46243 16276 46252 16316
rect 46292 16276 47404 16316
rect 47444 16276 48268 16316
rect 48308 16276 48317 16316
rect 48643 16276 48652 16316
rect 48692 16276 49420 16316
rect 49460 16276 49469 16316
rect 51427 16276 51436 16316
rect 51476 16276 52780 16316
rect 52820 16276 52829 16316
rect 52876 16276 55084 16316
rect 55124 16276 55133 16316
rect 61614 16276 61708 16316
rect 61748 16276 61757 16316
rect 61699 16275 61757 16276
rect 54691 16232 54749 16233
rect 55459 16232 55517 16233
rect 37027 16192 37036 16232
rect 37076 16192 37708 16232
rect 37748 16192 37757 16232
rect 46051 16192 46060 16232
rect 46100 16192 47212 16232
rect 47252 16192 47261 16232
rect 47491 16192 47500 16232
rect 47540 16192 49900 16232
rect 49940 16192 51244 16232
rect 51284 16192 51532 16232
rect 51572 16192 51581 16232
rect 51811 16192 51820 16232
rect 51860 16192 52396 16232
rect 52436 16192 52445 16232
rect 53059 16192 53068 16232
rect 53108 16192 54028 16232
rect 54068 16192 54077 16232
rect 54606 16192 54700 16232
rect 54740 16192 54749 16232
rect 55267 16192 55276 16232
rect 55316 16192 55468 16232
rect 55508 16192 55517 16232
rect 54691 16191 54749 16192
rect 55459 16191 55517 16192
rect 55651 16232 55709 16233
rect 58243 16232 58301 16233
rect 58531 16232 58589 16233
rect 64963 16232 65021 16233
rect 70147 16232 70205 16233
rect 78883 16232 78941 16233
rect 55651 16192 55660 16232
rect 55700 16192 55794 16232
rect 58158 16192 58252 16232
rect 58292 16192 58301 16232
rect 58446 16192 58540 16232
rect 58580 16192 58589 16232
rect 60739 16192 60748 16232
rect 60788 16192 61132 16232
rect 61172 16192 61181 16232
rect 62659 16192 62668 16232
rect 62708 16192 63052 16232
rect 63092 16192 63101 16232
rect 64878 16192 64972 16232
rect 65012 16192 65021 16232
rect 68227 16192 68236 16232
rect 68276 16192 68908 16232
rect 68948 16192 68957 16232
rect 70062 16192 70156 16232
rect 70196 16192 70205 16232
rect 73123 16192 73132 16232
rect 73172 16192 74956 16232
rect 74996 16192 75005 16232
rect 76963 16192 76972 16232
rect 77012 16192 77740 16232
rect 77780 16192 77789 16232
rect 78798 16192 78892 16232
rect 78932 16192 78941 16232
rect 55651 16191 55709 16192
rect 58243 16191 58301 16192
rect 58531 16191 58589 16192
rect 64963 16191 65021 16192
rect 70147 16191 70205 16192
rect 78883 16191 78941 16192
rect 45283 16108 45292 16148
rect 45332 16108 56524 16148
rect 56564 16108 56573 16148
rect 67651 16108 67660 16148
rect 67700 16108 69772 16148
rect 69812 16108 69821 16148
rect 53251 16064 53309 16065
rect 67651 16064 67709 16065
rect 3619 16024 3628 16064
rect 3668 16024 3916 16064
rect 3956 16024 11692 16064
rect 11732 16024 11741 16064
rect 39811 16024 39820 16064
rect 39860 16024 42604 16064
rect 42644 16024 43220 16064
rect 45475 16024 45484 16064
rect 45524 16024 45772 16064
rect 45812 16024 45821 16064
rect 53251 16024 53260 16064
rect 53300 16024 55180 16064
rect 55220 16024 55229 16064
rect 55747 16024 55756 16064
rect 55796 16024 63724 16064
rect 63764 16024 63773 16064
rect 67651 16024 67660 16064
rect 67700 16024 68524 16064
rect 68564 16024 68573 16064
rect 69379 16024 69388 16064
rect 69428 16024 70540 16064
rect 70580 16024 70589 16064
rect 43180 15980 43220 16024
rect 53251 16023 53309 16024
rect 67651 16023 67709 16024
rect 40195 15940 40204 15980
rect 40244 15940 40492 15980
rect 40532 15940 40541 15980
rect 41827 15940 41836 15980
rect 41876 15940 42028 15980
rect 42068 15940 42077 15980
rect 43180 15940 57292 15980
rect 57332 15940 57341 15980
rect 66883 15940 66892 15980
rect 66932 15940 69292 15980
rect 69332 15940 69341 15980
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 31075 15856 31084 15896
rect 31124 15856 33964 15896
rect 34004 15856 34013 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 39907 15856 39916 15896
rect 39956 15856 40300 15896
rect 40340 15856 40349 15896
rect 43363 15856 43372 15896
rect 43412 15856 46060 15896
rect 46100 15856 46109 15896
rect 47299 15856 47308 15896
rect 47348 15856 47500 15896
rect 47540 15856 48268 15896
rect 48308 15856 48317 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 51331 15856 51340 15896
rect 51380 15856 51820 15896
rect 51860 15856 51869 15896
rect 55555 15856 55564 15896
rect 55604 15856 56044 15896
rect 56084 15856 57868 15896
rect 57908 15856 57917 15896
rect 59491 15856 59500 15896
rect 59540 15856 66124 15896
rect 66164 15856 66173 15896
rect 67939 15856 67948 15896
rect 67988 15856 70924 15896
rect 70964 15856 70973 15896
rect 4003 15772 4012 15812
rect 4052 15772 4204 15812
rect 4244 15772 4253 15812
rect 33475 15772 33484 15812
rect 33524 15772 35596 15812
rect 35636 15772 36364 15812
rect 36404 15772 36413 15812
rect 64867 15772 64876 15812
rect 64916 15772 67852 15812
rect 67892 15772 72556 15812
rect 72596 15772 72605 15812
rect 0 15728 80 15748
rect 41731 15728 41789 15729
rect 52195 15728 52253 15729
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 2947 15688 2956 15728
rect 2996 15688 3820 15728
rect 3860 15688 4396 15728
rect 4436 15688 4445 15728
rect 33187 15688 33196 15728
rect 33236 15688 33245 15728
rect 34819 15688 34828 15728
rect 34868 15688 35212 15728
rect 35252 15688 36268 15728
rect 36308 15688 37228 15728
rect 37268 15688 37277 15728
rect 40579 15688 40588 15728
rect 40628 15688 40637 15728
rect 41731 15688 41740 15728
rect 41780 15688 52204 15728
rect 52244 15688 53644 15728
rect 53684 15688 53693 15728
rect 62947 15688 62956 15728
rect 62996 15688 63005 15728
rect 63340 15688 72172 15728
rect 72212 15688 72221 15728
rect 0 15668 80 15688
rect 33196 15644 33236 15688
rect 2851 15604 2860 15644
rect 2900 15604 3532 15644
rect 3572 15604 3581 15644
rect 31843 15604 31852 15644
rect 31892 15604 32140 15644
rect 32180 15604 32189 15644
rect 33196 15604 35116 15644
rect 35156 15604 35165 15644
rect 36931 15604 36940 15644
rect 36980 15604 37804 15644
rect 37844 15604 38380 15644
rect 38420 15604 38429 15644
rect 40588 15560 40628 15688
rect 41731 15687 41789 15688
rect 52195 15687 52253 15688
rect 62956 15644 62996 15688
rect 63340 15644 63380 15688
rect 62563 15604 62572 15644
rect 62612 15604 63380 15644
rect 71107 15604 71116 15644
rect 71156 15604 71500 15644
rect 71540 15604 72748 15644
rect 72788 15604 72797 15644
rect 1795 15520 1804 15560
rect 1844 15520 3148 15560
rect 3188 15520 3197 15560
rect 4579 15520 4588 15560
rect 4628 15520 4780 15560
rect 4820 15520 5068 15560
rect 5108 15520 5117 15560
rect 29443 15520 29452 15560
rect 29492 15520 32428 15560
rect 32468 15520 33620 15560
rect 34339 15520 34348 15560
rect 34388 15520 34924 15560
rect 34964 15520 34973 15560
rect 35971 15520 35980 15560
rect 36020 15520 37516 15560
rect 37556 15520 38572 15560
rect 38612 15520 38621 15560
rect 39139 15520 39148 15560
rect 39188 15520 40204 15560
rect 40244 15520 40492 15560
rect 40532 15520 40541 15560
rect 40588 15520 40876 15560
rect 40916 15520 40925 15560
rect 42019 15520 42028 15560
rect 42068 15520 42508 15560
rect 42548 15520 42988 15560
rect 43028 15520 43180 15560
rect 43220 15520 43229 15560
rect 47875 15520 47884 15560
rect 47924 15520 48172 15560
rect 48212 15520 48221 15560
rect 50563 15520 50572 15560
rect 50612 15520 51052 15560
rect 51092 15520 51101 15560
rect 52675 15520 52684 15560
rect 52724 15520 54316 15560
rect 54356 15520 54988 15560
rect 55028 15520 55037 15560
rect 61795 15520 61804 15560
rect 61844 15520 65740 15560
rect 65780 15520 66700 15560
rect 66740 15520 68812 15560
rect 68852 15520 68861 15560
rect 70051 15520 70060 15560
rect 70100 15520 71020 15560
rect 71060 15520 71069 15560
rect 73420 15520 75148 15560
rect 75188 15520 75197 15560
rect 33580 15476 33620 15520
rect 42028 15476 42068 15520
rect 52963 15476 53021 15477
rect 73420 15476 73460 15520
rect 33571 15436 33580 15476
rect 33620 15436 35404 15476
rect 35444 15436 36460 15476
rect 36500 15436 36509 15476
rect 40003 15436 40012 15476
rect 40052 15436 42068 15476
rect 46435 15436 46444 15476
rect 46484 15436 50380 15476
rect 50420 15436 50429 15476
rect 52963 15436 52972 15476
rect 53012 15436 60364 15476
rect 60404 15436 60413 15476
rect 66211 15436 66220 15476
rect 66260 15436 68716 15476
rect 68756 15436 70004 15476
rect 70723 15436 70732 15476
rect 70772 15436 73460 15476
rect 52963 15435 53021 15436
rect 69964 15392 70004 15436
rect 30211 15352 30220 15392
rect 30260 15352 31564 15392
rect 31604 15352 31613 15392
rect 34147 15352 34156 15392
rect 34196 15352 34924 15392
rect 34964 15352 34973 15392
rect 36547 15352 36556 15392
rect 36596 15352 36844 15392
rect 36884 15352 36893 15392
rect 51235 15352 51244 15392
rect 51284 15352 52012 15392
rect 52052 15352 52061 15392
rect 59971 15352 59980 15392
rect 60020 15352 60172 15392
rect 60212 15352 60940 15392
rect 60980 15352 69868 15392
rect 69908 15352 69917 15392
rect 69964 15352 74284 15392
rect 74324 15352 74333 15392
rect 69868 15308 69908 15352
rect 7363 15268 7372 15308
rect 7412 15268 45004 15308
rect 45044 15268 45053 15308
rect 68707 15268 68716 15308
rect 68756 15268 68908 15308
rect 68948 15268 68957 15308
rect 69868 15268 74668 15308
rect 74708 15268 74717 15308
rect 51619 15224 51677 15225
rect 8611 15184 8620 15224
rect 8660 15184 51628 15224
rect 51668 15184 51677 15224
rect 51619 15183 51677 15184
rect 52771 15224 52829 15225
rect 52771 15184 52780 15224
rect 52820 15184 60364 15224
rect 60404 15184 60413 15224
rect 70819 15184 70828 15224
rect 70868 15184 71308 15224
rect 71348 15184 71357 15224
rect 52771 15183 52829 15184
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 35683 15100 35692 15140
rect 35732 15100 36844 15140
rect 36884 15100 36893 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 47299 15016 47308 15056
rect 47348 15016 48076 15056
rect 48116 15016 50380 15056
rect 50420 15016 64108 15056
rect 64148 15016 64157 15056
rect 835 14932 844 14972
rect 884 14932 1516 14972
rect 1556 14932 1565 14972
rect 31747 14932 31756 14972
rect 31796 14932 32716 14972
rect 32756 14932 32908 14972
rect 32948 14932 32957 14972
rect 52387 14932 52396 14972
rect 52436 14932 53164 14972
rect 53204 14932 53213 14972
rect 61891 14932 61900 14972
rect 61940 14932 62188 14972
rect 62228 14932 65260 14972
rect 65300 14932 65309 14972
rect 0 14888 80 14908
rect 63331 14888 63389 14889
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 1987 14848 1996 14888
rect 2036 14848 2572 14888
rect 2612 14848 2621 14888
rect 33091 14848 33100 14888
rect 33140 14848 34348 14888
rect 34388 14848 35212 14888
rect 35252 14848 35261 14888
rect 60163 14848 60172 14888
rect 60212 14848 62708 14888
rect 62947 14848 62956 14888
rect 62996 14848 63340 14888
rect 63380 14848 70732 14888
rect 70772 14848 70781 14888
rect 75523 14848 75532 14888
rect 75572 14848 76204 14888
rect 76244 14848 76253 14888
rect 0 14828 80 14848
rect 60556 14804 60596 14848
rect 62668 14804 62708 14848
rect 63331 14847 63389 14848
rect 67171 14804 67229 14805
rect 2179 14764 2188 14804
rect 2228 14764 4876 14804
rect 4916 14764 4925 14804
rect 32035 14764 32044 14804
rect 32084 14764 33388 14804
rect 33428 14764 35116 14804
rect 35156 14764 35165 14804
rect 54019 14764 54028 14804
rect 54068 14764 56908 14804
rect 56948 14764 56957 14804
rect 60547 14764 60556 14804
rect 60596 14764 60605 14804
rect 61411 14764 61420 14804
rect 61460 14764 62572 14804
rect 62612 14764 62621 14804
rect 62668 14764 63436 14804
rect 63476 14764 63724 14804
rect 63764 14764 63773 14804
rect 63907 14764 63916 14804
rect 63956 14764 64300 14804
rect 64340 14764 65260 14804
rect 65300 14764 65309 14804
rect 67086 14764 67180 14804
rect 67220 14764 74764 14804
rect 74804 14764 74813 14804
rect 67171 14763 67229 14764
rect 54691 14720 54749 14721
rect 1315 14680 1324 14720
rect 1364 14680 2380 14720
rect 2420 14680 3340 14720
rect 3380 14680 3389 14720
rect 31459 14680 31468 14720
rect 31508 14680 34348 14720
rect 34388 14680 35308 14720
rect 35348 14680 35980 14720
rect 36020 14680 36029 14720
rect 36739 14680 36748 14720
rect 36788 14680 37228 14720
rect 37268 14680 37277 14720
rect 38083 14680 38092 14720
rect 38132 14680 39436 14720
rect 39476 14680 39485 14720
rect 40003 14680 40012 14720
rect 40052 14680 40061 14720
rect 42211 14680 42220 14720
rect 42260 14680 42700 14720
rect 42740 14680 42749 14720
rect 42979 14680 42988 14720
rect 43028 14680 43276 14720
rect 43316 14680 43325 14720
rect 46147 14680 46156 14720
rect 46196 14680 46540 14720
rect 46580 14680 48076 14720
rect 48116 14680 48125 14720
rect 54606 14680 54700 14720
rect 54740 14680 54749 14720
rect 56323 14680 56332 14720
rect 56372 14680 57580 14720
rect 57620 14680 59500 14720
rect 59540 14680 59549 14720
rect 60835 14680 60844 14720
rect 60884 14680 62476 14720
rect 62516 14680 62525 14720
rect 63340 14680 64876 14720
rect 64916 14680 64925 14720
rect 68899 14680 68908 14720
rect 68948 14680 71596 14720
rect 71636 14680 71645 14720
rect 73795 14680 73804 14720
rect 73844 14680 75244 14720
rect 75284 14680 75724 14720
rect 75764 14680 75773 14720
rect 40012 14636 40052 14680
rect 54691 14679 54749 14680
rect 63340 14636 63380 14680
rect 1699 14596 1708 14636
rect 1748 14596 3244 14636
rect 3284 14596 4012 14636
rect 4052 14596 4061 14636
rect 39331 14596 39340 14636
rect 39380 14596 40052 14636
rect 61123 14596 61132 14636
rect 61172 14596 63380 14636
rect 74371 14596 74380 14636
rect 74420 14596 75052 14636
rect 75092 14596 75101 14636
rect 32611 14552 32669 14553
rect 32227 14512 32236 14552
rect 32276 14512 32620 14552
rect 32660 14512 32669 14552
rect 39715 14512 39724 14552
rect 39764 14512 39773 14552
rect 53635 14512 53644 14552
rect 53684 14512 58924 14552
rect 58964 14512 58973 14552
rect 61987 14512 61996 14552
rect 62036 14512 62380 14552
rect 62420 14512 62429 14552
rect 62755 14512 62764 14552
rect 62804 14512 62813 14552
rect 63715 14512 63724 14552
rect 63764 14512 65452 14552
rect 65492 14512 70868 14552
rect 72163 14512 72172 14552
rect 72212 14512 73708 14552
rect 73748 14512 73757 14552
rect 73891 14512 73900 14552
rect 73940 14512 74668 14552
rect 74708 14512 74717 14552
rect 74947 14512 74956 14552
rect 74996 14512 76052 14552
rect 78595 14512 78604 14552
rect 78644 14512 79180 14552
rect 79220 14512 79229 14552
rect 32611 14511 32669 14512
rect 2947 14428 2956 14468
rect 2996 14428 3244 14468
rect 3284 14428 3293 14468
rect 31747 14428 31756 14468
rect 31796 14428 32428 14468
rect 32468 14428 32477 14468
rect 37315 14428 37324 14468
rect 37364 14428 38572 14468
rect 38612 14428 38621 14468
rect 39724 14384 39764 14512
rect 62764 14468 62804 14512
rect 68323 14468 68381 14469
rect 70828 14468 70868 14512
rect 76012 14468 76052 14512
rect 78604 14468 78644 14512
rect 54979 14428 54988 14468
rect 55028 14428 55948 14468
rect 55988 14428 57676 14468
rect 57716 14428 58348 14468
rect 58388 14428 58397 14468
rect 61996 14428 63820 14468
rect 63860 14428 63869 14468
rect 64483 14428 64492 14468
rect 64532 14428 65260 14468
rect 65300 14428 66988 14468
rect 67028 14428 67276 14468
rect 67316 14428 67325 14468
rect 67555 14428 67564 14468
rect 67604 14428 68332 14468
rect 68372 14428 68381 14468
rect 70819 14428 70828 14468
rect 70868 14428 75532 14468
rect 75572 14428 75581 14468
rect 76012 14428 78644 14468
rect 52003 14384 52061 14385
rect 58348 14384 58388 14428
rect 61996 14384 62036 14428
rect 68323 14427 68381 14428
rect 76012 14384 76052 14428
rect 2179 14344 2188 14384
rect 2228 14344 2476 14384
rect 2516 14344 2525 14384
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 37411 14344 37420 14384
rect 37460 14344 39148 14384
rect 39188 14344 39764 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 52003 14344 52012 14384
rect 52052 14344 53300 14384
rect 58348 14344 59404 14384
rect 59444 14344 59453 14384
rect 61987 14344 61996 14384
rect 62036 14344 62045 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 65347 14344 65356 14384
rect 65396 14344 69140 14384
rect 69187 14344 69196 14384
rect 69236 14344 74188 14384
rect 74228 14344 74237 14384
rect 74371 14344 74380 14384
rect 74420 14344 74429 14384
rect 76003 14344 76012 14384
rect 76052 14344 76061 14384
rect 52003 14343 52061 14344
rect 53260 14300 53300 14344
rect 69100 14300 69140 14344
rect 39331 14260 39340 14300
rect 39380 14260 41356 14300
rect 41396 14260 41405 14300
rect 46915 14260 46924 14300
rect 46964 14260 51724 14300
rect 51764 14260 51773 14300
rect 52675 14260 52684 14300
rect 52724 14260 53204 14300
rect 53260 14260 57772 14300
rect 57812 14260 57821 14300
rect 57955 14260 57964 14300
rect 58004 14260 60556 14300
rect 60596 14260 66508 14300
rect 66548 14260 66557 14300
rect 69100 14260 70924 14300
rect 70964 14260 70973 14300
rect 53164 14216 53204 14260
rect 1507 14176 1516 14216
rect 1556 14176 3532 14216
rect 3572 14176 4204 14216
rect 4244 14176 7276 14216
rect 7316 14176 8620 14216
rect 8660 14176 8669 14216
rect 31843 14176 31852 14216
rect 31892 14176 33772 14216
rect 33812 14176 33821 14216
rect 39811 14176 39820 14216
rect 39860 14176 41164 14216
rect 41204 14176 42700 14216
rect 42740 14176 43220 14216
rect 45955 14176 45964 14216
rect 46004 14176 47020 14216
rect 47060 14176 47404 14216
rect 47444 14176 47453 14216
rect 51235 14176 51244 14216
rect 51284 14176 52588 14216
rect 52628 14176 53068 14216
rect 53108 14176 53117 14216
rect 53164 14176 56468 14216
rect 62083 14176 62092 14216
rect 62132 14176 62668 14216
rect 62708 14176 62717 14216
rect 68131 14176 68140 14216
rect 68180 14176 70252 14216
rect 70292 14176 70301 14216
rect 43180 14132 43220 14176
rect 56428 14132 56468 14176
rect 31267 14092 31276 14132
rect 31316 14092 32236 14132
rect 32276 14092 37132 14132
rect 37172 14092 39628 14132
rect 39668 14092 39677 14132
rect 42595 14092 42604 14132
rect 42644 14092 42892 14132
rect 42932 14092 42941 14132
rect 43171 14092 43180 14132
rect 43220 14092 43229 14132
rect 50563 14092 50572 14132
rect 50612 14092 53452 14132
rect 53492 14092 53501 14132
rect 56419 14092 56428 14132
rect 56468 14092 56477 14132
rect 67459 14092 67468 14132
rect 67508 14092 68044 14132
rect 68084 14092 68093 14132
rect 68803 14092 68812 14132
rect 68852 14092 69100 14132
rect 69140 14092 70060 14132
rect 70100 14092 70109 14132
rect 0 14048 80 14068
rect 38572 14048 38612 14092
rect 52387 14048 52445 14049
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 1699 14008 1708 14048
rect 1748 14008 2092 14048
rect 2132 14008 2668 14048
rect 2708 14008 3628 14048
rect 3668 14008 3820 14048
rect 3860 14008 3869 14048
rect 30211 14008 30220 14048
rect 30260 14008 31564 14048
rect 31604 14008 37324 14048
rect 37364 14008 37373 14048
rect 38563 14008 38572 14048
rect 38612 14008 38652 14048
rect 38755 14008 38764 14048
rect 38804 14008 39148 14048
rect 39188 14008 39197 14048
rect 40387 14008 40396 14048
rect 40436 14008 41548 14048
rect 41588 14008 43660 14048
rect 43700 14008 43709 14048
rect 44611 14008 44620 14048
rect 44660 14008 46156 14048
rect 46196 14008 46205 14048
rect 46339 14008 46348 14048
rect 46388 14008 47788 14048
rect 47828 14008 47837 14048
rect 52387 14008 52396 14048
rect 52436 14008 52684 14048
rect 52724 14008 52733 14048
rect 61603 14008 61612 14048
rect 61652 14008 62188 14048
rect 62228 14008 62237 14048
rect 62371 14008 62380 14048
rect 62420 14008 63916 14048
rect 63956 14008 64396 14048
rect 64436 14008 67372 14048
rect 67412 14008 67421 14048
rect 68611 14008 68620 14048
rect 68660 14008 69004 14048
rect 69044 14008 69053 14048
rect 69955 14008 69964 14048
rect 70004 14008 71500 14048
rect 71540 14008 71549 14048
rect 0 13988 80 14008
rect 52387 14007 52445 14008
rect 69187 13964 69245 13965
rect 1987 13924 1996 13964
rect 2036 13924 2284 13964
rect 2324 13924 2572 13964
rect 2612 13924 2621 13964
rect 31939 13924 31948 13964
rect 31988 13924 32620 13964
rect 32660 13924 32669 13964
rect 39235 13924 39244 13964
rect 39284 13924 41260 13964
rect 41300 13924 41309 13964
rect 53347 13924 53356 13964
rect 53396 13924 56236 13964
rect 56276 13924 57388 13964
rect 57428 13924 57437 13964
rect 61507 13924 61516 13964
rect 61556 13924 63628 13964
rect 63668 13924 63820 13964
rect 63860 13924 63869 13964
rect 69102 13924 69196 13964
rect 69236 13924 69245 13964
rect 69187 13923 69245 13924
rect 74380 13880 74420 14344
rect 77155 14176 77164 14216
rect 77204 14176 78700 14216
rect 78740 14176 79372 14216
rect 79412 14176 79421 14216
rect 74947 14008 74956 14048
rect 74996 14008 75244 14048
rect 75284 14008 75293 14048
rect 40099 13840 40108 13880
rect 40148 13840 41932 13880
rect 41972 13840 41981 13880
rect 43459 13840 43468 13880
rect 43508 13840 43852 13880
rect 43892 13840 43901 13880
rect 52099 13840 52108 13880
rect 52148 13840 74612 13880
rect 68323 13796 68381 13797
rect 74572 13796 74612 13840
rect 45187 13756 45196 13796
rect 45236 13756 55852 13796
rect 55892 13756 55901 13796
rect 56044 13756 56524 13796
rect 56564 13756 57100 13796
rect 57140 13756 57149 13796
rect 67267 13756 67276 13796
rect 67316 13756 67660 13796
rect 67700 13756 67709 13796
rect 68238 13756 68332 13796
rect 68372 13756 68381 13796
rect 74563 13756 74572 13796
rect 74612 13756 74621 13796
rect 56044 13712 56084 13756
rect 68323 13755 68381 13756
rect 50755 13672 50764 13712
rect 50804 13672 51436 13712
rect 51476 13672 51485 13712
rect 54499 13672 54508 13712
rect 54548 13672 56084 13712
rect 56899 13672 56908 13712
rect 56948 13672 58828 13712
rect 58868 13672 58877 13712
rect 67843 13672 67852 13712
rect 67892 13672 68140 13712
rect 68180 13672 68189 13712
rect 70915 13672 70924 13712
rect 70964 13672 75820 13712
rect 75860 13672 75869 13712
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 42403 13588 42412 13628
rect 42452 13588 42700 13628
rect 42740 13588 42749 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 50467 13588 50476 13628
rect 50516 13588 50956 13628
rect 50996 13588 51005 13628
rect 51907 13588 51916 13628
rect 51956 13588 54316 13628
rect 54356 13588 54365 13628
rect 56419 13588 56428 13628
rect 56468 13588 58252 13628
rect 58292 13588 58301 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 73603 13588 73612 13628
rect 73652 13588 75628 13628
rect 75668 13588 75677 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 70435 13544 70493 13545
rect 32803 13504 32812 13544
rect 32852 13504 33100 13544
rect 33140 13504 33149 13544
rect 43267 13504 43276 13544
rect 43316 13504 45484 13544
rect 45524 13504 56812 13544
rect 56852 13504 56861 13544
rect 59212 13504 63244 13544
rect 63284 13504 63293 13544
rect 69667 13504 69676 13544
rect 69716 13504 70060 13544
rect 70100 13504 70444 13544
rect 70484 13504 70493 13544
rect 43180 13420 46004 13460
rect 47587 13420 47596 13460
rect 47636 13420 48844 13460
rect 48884 13420 48893 13460
rect 51619 13420 51628 13460
rect 51668 13420 55756 13460
rect 55796 13420 55805 13460
rect 57859 13420 57868 13460
rect 57908 13420 58636 13460
rect 58676 13420 58685 13460
rect 43180 13376 43220 13420
rect 45964 13376 46004 13420
rect 59212 13376 59252 13504
rect 70435 13503 70493 13504
rect 60931 13420 60940 13460
rect 60980 13420 61900 13460
rect 61940 13420 61949 13460
rect 36739 13336 36748 13376
rect 36788 13336 39340 13376
rect 39380 13336 43220 13376
rect 45859 13336 45868 13376
rect 45908 13336 45917 13376
rect 45964 13336 53644 13376
rect 53684 13336 53693 13376
rect 54307 13336 54316 13376
rect 54356 13336 59252 13376
rect 59299 13336 59308 13376
rect 59348 13336 62380 13376
rect 62420 13336 62429 13376
rect 70435 13336 70444 13376
rect 70484 13336 70732 13376
rect 70772 13336 76588 13376
rect 76628 13336 76637 13376
rect 77251 13336 77260 13376
rect 77300 13336 77452 13376
rect 77492 13336 77501 13376
rect 45868 13292 45908 13336
rect 1219 13252 1228 13292
rect 1268 13252 3532 13292
rect 3572 13252 3581 13292
rect 32611 13252 32620 13292
rect 32660 13252 34924 13292
rect 34964 13252 35500 13292
rect 35540 13252 35549 13292
rect 43651 13252 43660 13292
rect 43700 13252 44332 13292
rect 44372 13252 44716 13292
rect 44756 13252 45580 13292
rect 45620 13252 46540 13292
rect 46580 13252 47404 13292
rect 47444 13252 49228 13292
rect 49268 13252 49277 13292
rect 50851 13252 50860 13292
rect 50900 13252 52108 13292
rect 52148 13252 53260 13292
rect 53300 13252 53309 13292
rect 55171 13252 55180 13292
rect 55220 13252 56468 13292
rect 57859 13252 57868 13292
rect 57908 13252 61420 13292
rect 61460 13252 62956 13292
rect 62996 13252 64780 13292
rect 64820 13252 64829 13292
rect 67555 13252 67564 13292
rect 67604 13252 69292 13292
rect 69332 13252 69341 13292
rect 69475 13252 69484 13292
rect 69524 13252 75436 13292
rect 75476 13252 75485 13292
rect 75715 13252 75724 13292
rect 75764 13252 77164 13292
rect 77204 13252 77213 13292
rect 0 13208 80 13228
rect 49228 13208 49268 13252
rect 56428 13208 56468 13252
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 2755 13168 2764 13208
rect 2804 13168 2956 13208
rect 2996 13168 4396 13208
rect 4436 13168 5164 13208
rect 5204 13168 5213 13208
rect 31651 13168 31660 13208
rect 31700 13168 32812 13208
rect 32852 13168 32861 13208
rect 35011 13168 35020 13208
rect 35060 13168 38668 13208
rect 38708 13168 38717 13208
rect 41635 13168 41644 13208
rect 41684 13168 42796 13208
rect 42836 13168 42845 13208
rect 45667 13168 45676 13208
rect 45716 13168 46156 13208
rect 46196 13168 46205 13208
rect 48067 13168 48076 13208
rect 48116 13168 48125 13208
rect 49228 13168 49708 13208
rect 49748 13168 50476 13208
rect 50516 13168 53356 13208
rect 53396 13168 53405 13208
rect 53539 13168 53548 13208
rect 53588 13168 54412 13208
rect 54452 13168 54461 13208
rect 54691 13168 54700 13208
rect 54740 13168 55084 13208
rect 55124 13168 55133 13208
rect 55363 13168 55372 13208
rect 55412 13168 56044 13208
rect 56084 13168 56093 13208
rect 56419 13168 56428 13208
rect 56468 13168 56477 13208
rect 56611 13168 56620 13208
rect 56660 13168 58444 13208
rect 58484 13168 58732 13208
rect 58772 13168 58781 13208
rect 62860 13168 64876 13208
rect 64916 13168 64925 13208
rect 68803 13168 68812 13208
rect 68852 13168 69580 13208
rect 69620 13168 69629 13208
rect 70531 13168 70540 13208
rect 70580 13168 71116 13208
rect 71156 13168 74612 13208
rect 74659 13168 74668 13208
rect 74708 13168 75148 13208
rect 75188 13168 75820 13208
rect 75860 13168 75869 13208
rect 0 13148 80 13168
rect 48076 13124 48116 13168
rect 62860 13124 62900 13168
rect 70540 13124 70580 13168
rect 74572 13124 74612 13168
rect 35203 13084 35212 13124
rect 35252 13084 35980 13124
rect 36020 13084 38476 13124
rect 38516 13084 38525 13124
rect 40291 13084 40300 13124
rect 40340 13084 41548 13124
rect 41588 13084 41597 13124
rect 46435 13084 46444 13124
rect 46484 13084 47980 13124
rect 48020 13084 48029 13124
rect 48076 13084 49324 13124
rect 49364 13084 49373 13124
rect 53443 13084 53452 13124
rect 53492 13084 56332 13124
rect 56372 13084 57484 13124
rect 57524 13084 57533 13124
rect 58531 13084 58540 13124
rect 58580 13084 61516 13124
rect 61556 13084 62860 13124
rect 62900 13084 62909 13124
rect 69091 13084 69100 13124
rect 69140 13084 70580 13124
rect 72259 13084 72268 13124
rect 72308 13084 74380 13124
rect 74420 13084 74429 13124
rect 74572 13084 75244 13124
rect 75284 13084 76972 13124
rect 77012 13084 77021 13124
rect 74956 13040 74996 13084
rect 4204 13000 4492 13040
rect 4532 13000 4541 13040
rect 45763 13000 45772 13040
rect 45812 13000 48076 13040
rect 48116 13000 48125 13040
rect 55267 13000 55276 13040
rect 55316 13000 56756 13040
rect 57667 13000 57676 13040
rect 57716 13000 58060 13040
rect 58100 13000 60556 13040
rect 60596 13000 62476 13040
rect 62516 13000 62525 13040
rect 68611 13000 68620 13040
rect 68660 13000 68812 13040
rect 68852 13000 68861 13040
rect 74275 13000 74284 13040
rect 74324 13000 74860 13040
rect 74900 13000 74909 13040
rect 74955 13000 74964 13040
rect 75004 13000 75013 13040
rect 4204 12872 4244 13000
rect 56716 12980 56756 13000
rect 56716 12956 56796 12980
rect 42307 12916 42316 12956
rect 42356 12916 43276 12956
rect 43316 12916 43564 12956
rect 43604 12916 43613 12956
rect 45379 12916 45388 12956
rect 45428 12916 45868 12956
rect 45908 12916 45917 12956
rect 51235 12916 51244 12956
rect 51284 12916 51916 12956
rect 51956 12916 51965 12956
rect 56707 12916 56716 12956
rect 56756 12940 56796 12956
rect 69283 12940 69292 12980
rect 69332 12956 69341 12980
rect 69332 12940 69676 12956
rect 56756 12916 56765 12940
rect 69292 12916 69676 12940
rect 69716 12916 70196 12956
rect 71683 12916 71692 12956
rect 71732 12916 73516 12956
rect 73556 12916 77356 12956
rect 77396 12916 78124 12956
rect 78164 12916 78173 12956
rect 70156 12872 70196 12916
rect 2467 12832 2476 12872
rect 2516 12832 4108 12872
rect 4148 12832 4244 12872
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 57379 12832 57388 12872
rect 57428 12832 57868 12872
rect 57908 12832 57917 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 68419 12832 68428 12872
rect 68468 12832 68812 12872
rect 68852 12832 68861 12872
rect 69763 12832 69772 12872
rect 69812 12832 70060 12872
rect 70100 12832 70109 12872
rect 70156 12832 73460 12872
rect 2659 12748 2668 12788
rect 2708 12748 4972 12788
rect 5012 12748 5021 12788
rect 47491 12748 47500 12788
rect 47540 12748 47788 12788
rect 47828 12748 47837 12788
rect 63619 12748 63628 12788
rect 63668 12748 64396 12788
rect 64436 12748 67180 12788
rect 67220 12748 71788 12788
rect 71828 12748 71837 12788
rect 36547 12704 36605 12705
rect 1411 12664 1420 12704
rect 1460 12664 2380 12704
rect 2420 12664 2429 12704
rect 36462 12664 36556 12704
rect 36596 12664 36605 12704
rect 47683 12664 47692 12704
rect 47732 12664 48172 12704
rect 48212 12664 48221 12704
rect 49507 12664 49516 12704
rect 49556 12664 49708 12704
rect 49748 12664 49757 12704
rect 57187 12664 57196 12704
rect 57236 12664 57676 12704
rect 57716 12664 58156 12704
rect 58196 12664 58205 12704
rect 60835 12664 60844 12704
rect 60884 12664 62092 12704
rect 62132 12664 62141 12704
rect 68707 12664 68716 12704
rect 68756 12664 69004 12704
rect 69044 12664 69053 12704
rect 70627 12664 70636 12704
rect 70676 12664 72844 12704
rect 72884 12664 73324 12704
rect 73364 12664 73373 12704
rect 36547 12663 36605 12664
rect 73420 12620 73460 12832
rect 76387 12788 76445 12789
rect 75043 12748 75052 12788
rect 75092 12748 75244 12788
rect 75284 12748 75293 12788
rect 76302 12748 76396 12788
rect 76436 12748 76445 12788
rect 76387 12747 76445 12748
rect 74467 12664 74476 12704
rect 74516 12664 76108 12704
rect 76148 12664 76684 12704
rect 76724 12664 76733 12704
rect 48259 12580 48268 12620
rect 48308 12580 51628 12620
rect 51668 12580 51677 12620
rect 54787 12580 54796 12620
rect 54836 12580 56620 12620
rect 56660 12580 56669 12620
rect 59011 12580 59020 12620
rect 59060 12580 59692 12620
rect 59732 12580 59741 12620
rect 61987 12580 61996 12620
rect 62036 12580 64012 12620
rect 64052 12580 64061 12620
rect 73420 12580 74764 12620
rect 74804 12580 75532 12620
rect 75572 12580 75581 12620
rect 41731 12536 41789 12537
rect 49516 12536 49556 12580
rect 4771 12496 4780 12536
rect 4820 12496 5452 12536
rect 5492 12496 29932 12536
rect 29972 12496 29981 12536
rect 31363 12496 31372 12536
rect 31412 12496 40684 12536
rect 40724 12496 41740 12536
rect 41780 12496 41789 12536
rect 41923 12496 41932 12536
rect 41972 12496 42508 12536
rect 42548 12496 42557 12536
rect 48643 12496 48652 12536
rect 48692 12496 49036 12536
rect 49076 12496 49085 12536
rect 49507 12496 49516 12536
rect 49556 12496 49565 12536
rect 53260 12496 59212 12536
rect 59252 12496 59261 12536
rect 62275 12496 62284 12536
rect 62324 12496 62764 12536
rect 62804 12496 63724 12536
rect 63764 12496 63773 12536
rect 64579 12496 64588 12536
rect 64628 12496 65548 12536
rect 65588 12496 65597 12536
rect 69955 12496 69964 12536
rect 70004 12496 70540 12536
rect 70580 12496 70589 12536
rect 71203 12496 71212 12536
rect 71252 12496 71692 12536
rect 71732 12496 71741 12536
rect 41731 12495 41789 12496
rect 2947 12452 3005 12453
rect 1315 12412 1324 12452
rect 1364 12412 2956 12452
rect 2996 12412 3005 12452
rect 42019 12412 42028 12452
rect 42068 12412 42988 12452
rect 43028 12412 43037 12452
rect 49123 12412 49132 12452
rect 49172 12412 49420 12452
rect 49460 12412 49469 12452
rect 2947 12411 3005 12412
rect 0 12368 80 12388
rect 53260 12368 53300 12496
rect 57763 12452 57821 12453
rect 64588 12452 64628 12496
rect 57678 12412 57772 12452
rect 57812 12412 57821 12452
rect 62179 12412 62188 12452
rect 62228 12412 64628 12452
rect 70435 12412 70444 12452
rect 70484 12412 70493 12452
rect 57763 12411 57821 12412
rect 70444 12368 70484 12412
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 2563 12328 2572 12368
rect 2612 12328 2764 12368
rect 2804 12328 2813 12368
rect 5347 12328 5356 12368
rect 5396 12328 5836 12368
rect 5876 12328 5885 12368
rect 35587 12328 35596 12368
rect 35636 12328 36268 12368
rect 36308 12328 36748 12368
rect 36788 12328 36797 12368
rect 39523 12328 39532 12368
rect 39572 12328 41548 12368
rect 41588 12328 53300 12368
rect 69091 12328 69100 12368
rect 69140 12328 70060 12368
rect 70100 12328 70109 12368
rect 70243 12328 70252 12368
rect 70292 12328 70484 12368
rect 74563 12328 74572 12368
rect 74612 12328 74764 12368
rect 74804 12328 74813 12368
rect 0 12308 80 12328
rect 547 12244 556 12284
rect 596 12244 1516 12284
rect 1556 12244 1565 12284
rect 53284 12244 53293 12284
rect 53333 12244 55180 12284
rect 55220 12244 55229 12284
rect 69571 12244 69580 12284
rect 69620 12244 69772 12284
rect 69812 12244 69821 12284
rect 78307 12244 78316 12284
rect 78356 12244 79276 12284
rect 79316 12244 79325 12284
rect 57955 12160 57964 12200
rect 58004 12160 58252 12200
rect 58292 12160 58301 12200
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 62467 12076 62476 12116
rect 62516 12076 63052 12116
rect 63092 12076 63101 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 38851 11992 38860 12032
rect 38900 11992 39148 12032
rect 39188 11992 39197 12032
rect 42595 11992 42604 12032
rect 42644 11992 44812 12032
rect 44852 11992 59020 12032
rect 59060 11992 59069 12032
rect 59491 11992 59500 12032
rect 59540 11992 59692 12032
rect 59732 11992 61708 12032
rect 61748 11992 66796 12032
rect 66836 11992 66845 12032
rect 52867 11948 52925 11949
rect 33859 11908 33868 11948
rect 33908 11908 34828 11948
rect 34868 11908 34877 11948
rect 36163 11908 36172 11948
rect 36212 11908 38092 11948
rect 38132 11908 38141 11948
rect 45283 11908 45292 11948
rect 45332 11908 48268 11948
rect 48308 11908 48317 11948
rect 52867 11908 52876 11948
rect 52916 11908 57484 11948
rect 57524 11908 64148 11948
rect 64195 11908 64204 11948
rect 64244 11908 64780 11948
rect 64820 11908 64829 11948
rect 67363 11908 67372 11948
rect 67412 11908 68908 11948
rect 68948 11908 68957 11948
rect 75043 11908 75052 11948
rect 75092 11908 75724 11948
rect 75764 11908 75773 11948
rect 52867 11907 52925 11908
rect 64108 11864 64148 11908
rect 35011 11824 35020 11864
rect 35060 11824 36268 11864
rect 36308 11824 36652 11864
rect 36692 11824 36701 11864
rect 48547 11824 48556 11864
rect 48596 11824 49228 11864
rect 49268 11824 49277 11864
rect 50851 11824 50860 11864
rect 50900 11824 52588 11864
rect 52628 11824 52637 11864
rect 56803 11824 56812 11864
rect 56852 11824 57676 11864
rect 57716 11824 57964 11864
rect 58004 11824 58013 11864
rect 64108 11824 66220 11864
rect 66260 11824 66269 11864
rect 69667 11824 69676 11864
rect 69716 11824 69725 11864
rect 3619 11780 3677 11781
rect 1123 11740 1132 11780
rect 1172 11740 3628 11780
rect 3668 11740 3677 11780
rect 51715 11740 51724 11780
rect 51764 11740 53740 11780
rect 53780 11740 53789 11780
rect 3619 11739 3677 11740
rect 5635 11656 5644 11696
rect 5684 11656 6220 11696
rect 6260 11656 6269 11696
rect 34819 11656 34828 11696
rect 34868 11656 35308 11696
rect 35348 11656 35357 11696
rect 36835 11656 36844 11696
rect 36884 11656 37996 11696
rect 38036 11656 38860 11696
rect 38900 11656 38909 11696
rect 41539 11656 41548 11696
rect 41588 11656 41597 11696
rect 41827 11656 41836 11696
rect 41876 11656 42604 11696
rect 42644 11656 42653 11696
rect 45859 11656 45868 11696
rect 45908 11656 47884 11696
rect 47924 11656 47933 11696
rect 48451 11656 48460 11696
rect 48500 11656 49036 11696
rect 49076 11656 49085 11696
rect 49219 11656 49228 11696
rect 49268 11656 50092 11696
rect 50132 11656 50284 11696
rect 50324 11656 50333 11696
rect 51523 11656 51532 11696
rect 51572 11656 52204 11696
rect 52244 11656 52253 11696
rect 52387 11656 52396 11696
rect 52436 11656 53644 11696
rect 53684 11656 53693 11696
rect 57283 11656 57292 11696
rect 57332 11656 58348 11696
rect 58388 11656 58540 11696
rect 58580 11656 58589 11696
rect 60931 11656 60940 11696
rect 60980 11656 62764 11696
rect 62804 11656 62813 11696
rect 63331 11656 63340 11696
rect 63380 11656 63389 11696
rect 63436 11656 63916 11696
rect 63956 11656 64396 11696
rect 64436 11656 64445 11696
rect 41548 11612 41588 11656
rect 43075 11612 43133 11613
rect 35491 11572 35500 11612
rect 35540 11572 37612 11612
rect 37652 11572 37661 11612
rect 38083 11572 38092 11612
rect 38132 11572 39436 11612
rect 39476 11572 39485 11612
rect 41548 11572 43084 11612
rect 43124 11572 43276 11612
rect 43316 11572 43325 11612
rect 48355 11572 48364 11612
rect 48404 11572 49516 11612
rect 49556 11572 50764 11612
rect 50804 11572 51244 11612
rect 51284 11572 51293 11612
rect 51427 11572 51436 11612
rect 51476 11572 51916 11612
rect 51956 11572 52300 11612
rect 52340 11572 52349 11612
rect 58915 11572 58924 11612
rect 58964 11572 59308 11612
rect 59348 11572 59357 11612
rect 43075 11571 43133 11572
rect 0 11528 80 11548
rect 63340 11528 63380 11656
rect 63436 11612 63476 11656
rect 69676 11612 69716 11824
rect 69763 11656 69772 11696
rect 69812 11656 70636 11696
rect 70676 11656 70685 11696
rect 75427 11656 75436 11696
rect 75476 11656 76204 11696
rect 76244 11656 76684 11696
rect 76724 11656 76733 11696
rect 63427 11572 63436 11612
rect 63476 11572 63485 11612
rect 68908 11572 69716 11612
rect 75620 11572 75629 11612
rect 75669 11572 77164 11612
rect 77204 11572 78316 11612
rect 78356 11572 78365 11612
rect 68908 11528 68948 11572
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 2947 11488 2956 11528
rect 2996 11488 3532 11528
rect 3572 11488 3724 11528
rect 3764 11488 3773 11528
rect 4003 11488 4012 11528
rect 4052 11488 4684 11528
rect 4724 11488 4733 11528
rect 35395 11488 35404 11528
rect 35444 11488 37516 11528
rect 37556 11488 37565 11528
rect 61027 11488 61036 11528
rect 61076 11488 63380 11528
rect 68899 11488 68908 11528
rect 68948 11488 68957 11528
rect 69187 11488 69196 11528
rect 69236 11488 69868 11528
rect 69908 11488 69917 11528
rect 75331 11488 75340 11528
rect 75380 11488 76012 11528
rect 76052 11488 76061 11528
rect 0 11468 80 11488
rect 70435 11444 70493 11445
rect 62947 11404 62956 11444
rect 62996 11404 64012 11444
rect 64052 11404 64061 11444
rect 70435 11404 70444 11444
rect 70484 11404 75916 11444
rect 75956 11404 76396 11444
rect 76436 11404 77260 11444
rect 77300 11404 77309 11444
rect 70435 11403 70493 11404
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 38851 11320 38860 11360
rect 38900 11320 39532 11360
rect 39572 11320 39581 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 59299 11320 59308 11360
rect 59348 11320 61900 11360
rect 61940 11320 63820 11360
rect 63860 11320 63869 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 74851 11320 74860 11360
rect 74900 11320 75244 11360
rect 75284 11320 75293 11360
rect 56323 11236 56332 11276
rect 56372 11236 62572 11276
rect 62612 11236 62621 11276
rect 76291 11236 76300 11276
rect 76340 11236 76588 11276
rect 76628 11236 76637 11276
rect 1891 11152 1900 11192
rect 1940 11152 2188 11192
rect 2228 11152 2237 11192
rect 3427 11152 3436 11192
rect 3476 11152 5108 11192
rect 42595 11152 42604 11192
rect 42644 11152 46828 11192
rect 46868 11152 46877 11192
rect 50179 11152 50188 11192
rect 50228 11152 50956 11192
rect 50996 11152 52108 11192
rect 52148 11152 52157 11192
rect 58435 11152 58444 11192
rect 58484 11152 58924 11192
rect 58964 11152 59404 11192
rect 59444 11152 59453 11192
rect 72547 11152 72556 11192
rect 72596 11152 75244 11192
rect 75284 11152 75293 11192
rect 1795 11068 1804 11108
rect 1844 11068 3532 11108
rect 3572 11068 3581 11108
rect 5068 11024 5108 11152
rect 36547 11108 36605 11109
rect 36462 11068 36556 11108
rect 36596 11068 39340 11108
rect 39380 11068 39389 11108
rect 43939 11068 43948 11108
rect 43988 11068 46732 11108
rect 46772 11068 60076 11108
rect 60116 11068 60125 11108
rect 36547 11067 36605 11068
rect 1315 10984 1324 11024
rect 1364 10984 2324 11024
rect 2467 10984 2476 11024
rect 2516 10984 4012 11024
rect 4052 10984 4061 11024
rect 5059 10984 5068 11024
rect 5108 10984 7372 11024
rect 7412 10984 7421 11024
rect 35971 10984 35980 11024
rect 36020 10984 36748 11024
rect 36788 10984 36797 11024
rect 37027 10984 37036 11024
rect 37076 10984 37085 11024
rect 37699 10984 37708 11024
rect 37748 10984 38956 11024
rect 38996 10984 39005 11024
rect 48931 10984 48940 11024
rect 48980 10984 50188 11024
rect 50228 10984 50237 11024
rect 50659 10984 50668 11024
rect 50708 10984 50860 11024
rect 50900 10984 52300 11024
rect 52340 10984 52349 11024
rect 52675 10984 52684 11024
rect 52724 10984 52733 11024
rect 53155 10984 53164 11024
rect 53204 10984 53452 11024
rect 53492 10984 53501 11024
rect 59779 10984 59788 11024
rect 59828 10984 61036 11024
rect 61076 10984 61085 11024
rect 62179 10984 62188 11024
rect 62228 10984 62956 11024
rect 62996 10984 63005 11024
rect 63811 10984 63820 11024
rect 63860 10984 64684 11024
rect 64724 10984 64733 11024
rect 69091 10984 69100 11024
rect 69140 10984 70444 11024
rect 70484 10984 70493 11024
rect 74659 10984 74668 11024
rect 74708 10984 75148 11024
rect 75188 10984 75197 11024
rect 2284 10856 2324 10984
rect 37036 10940 37076 10984
rect 52003 10940 52061 10941
rect 37036 10900 39148 10940
rect 39188 10900 39532 10940
rect 39572 10900 39581 10940
rect 42307 10900 42316 10940
rect 42356 10900 44140 10940
rect 44180 10900 46252 10940
rect 46292 10900 46924 10940
rect 46964 10900 46973 10940
rect 51907 10900 51916 10940
rect 51956 10900 52012 10940
rect 52052 10900 52061 10940
rect 52684 10940 52724 10984
rect 52684 10900 53548 10940
rect 53588 10900 53597 10940
rect 64579 10900 64588 10940
rect 64628 10900 65068 10940
rect 65108 10900 65117 10940
rect 68995 10900 69004 10940
rect 69044 10900 69580 10940
rect 69620 10900 74860 10940
rect 74900 10900 75244 10940
rect 75284 10900 75293 10940
rect 77251 10900 77260 10940
rect 77300 10900 77309 10940
rect 2275 10816 2284 10856
rect 2324 10816 2333 10856
rect 1027 10732 1036 10772
rect 1076 10732 1085 10772
rect 0 10688 80 10708
rect 1036 10688 1076 10732
rect 0 10648 1076 10688
rect 0 10628 80 10648
rect 44332 10604 44372 10900
rect 52003 10899 52061 10900
rect 76387 10856 76445 10857
rect 77260 10856 77300 10900
rect 53059 10816 53068 10856
rect 53108 10816 56332 10856
rect 56372 10816 56381 10856
rect 74755 10816 74764 10856
rect 74804 10816 75340 10856
rect 75380 10816 75389 10856
rect 76291 10816 76300 10856
rect 76340 10816 76396 10856
rect 76436 10816 76445 10856
rect 76963 10816 76972 10856
rect 77012 10816 77300 10856
rect 76387 10815 76445 10816
rect 64867 10732 64876 10772
rect 64916 10732 65260 10772
rect 65300 10732 65309 10772
rect 75811 10732 75820 10772
rect 75860 10732 76684 10772
rect 76724 10732 77740 10772
rect 77780 10732 77789 10772
rect 46819 10648 46828 10688
rect 46868 10648 49420 10688
rect 49460 10648 49469 10688
rect 65443 10648 65452 10688
rect 65492 10648 67660 10688
rect 67700 10648 71404 10688
rect 71444 10648 71453 10688
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 44323 10564 44332 10604
rect 44372 10564 44381 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 68419 10564 68428 10604
rect 68468 10564 70156 10604
rect 70196 10564 73460 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 73420 10520 73460 10564
rect 42019 10480 42028 10520
rect 42068 10480 43220 10520
rect 47107 10480 47116 10520
rect 47156 10480 49228 10520
rect 49268 10480 60460 10520
rect 60500 10480 60509 10520
rect 69379 10480 69388 10520
rect 69428 10480 69437 10520
rect 73420 10480 74764 10520
rect 74804 10480 74813 10520
rect 43180 10436 43220 10480
rect 69388 10436 69428 10480
rect 1699 10396 1708 10436
rect 1748 10396 2476 10436
rect 2516 10396 2525 10436
rect 43180 10396 49516 10436
rect 49556 10396 49565 10436
rect 56515 10396 56524 10436
rect 56564 10396 58060 10436
rect 58100 10396 58109 10436
rect 68419 10396 68428 10436
rect 68468 10396 69428 10436
rect 69571 10396 69580 10436
rect 69620 10396 71020 10436
rect 71060 10396 72940 10436
rect 72980 10396 73996 10436
rect 74036 10396 74045 10436
rect 75907 10396 75916 10436
rect 75956 10396 76588 10436
rect 76628 10396 76637 10436
rect 2851 10312 2860 10352
rect 2900 10312 3052 10352
rect 3092 10312 3101 10352
rect 57859 10312 57868 10352
rect 57908 10312 59212 10352
rect 59252 10312 59261 10352
rect 67267 10312 67276 10352
rect 67316 10312 67852 10352
rect 67892 10312 67901 10352
rect 68332 10312 69332 10352
rect 69379 10312 69388 10352
rect 69428 10312 69772 10352
rect 69812 10312 70732 10352
rect 70772 10312 70781 10352
rect 58915 10268 58973 10269
rect 67651 10268 67709 10269
rect 3235 10228 3244 10268
rect 3284 10228 4876 10268
rect 4916 10228 4925 10268
rect 41635 10228 41644 10268
rect 41684 10228 41932 10268
rect 41972 10228 41981 10268
rect 42211 10228 42220 10268
rect 42260 10228 43220 10268
rect 43843 10228 43852 10268
rect 43892 10228 44140 10268
rect 44180 10228 44189 10268
rect 57379 10228 57388 10268
rect 57428 10228 58732 10268
rect 58772 10228 58781 10268
rect 58830 10228 58924 10268
rect 58964 10228 58973 10268
rect 59683 10228 59692 10268
rect 59732 10228 61996 10268
rect 62036 10228 67084 10268
rect 67124 10228 67133 10268
rect 67566 10228 67660 10268
rect 67700 10228 67709 10268
rect 43180 10184 43220 10228
rect 58732 10184 58772 10228
rect 58915 10227 58973 10228
rect 67651 10227 67709 10228
rect 68332 10184 68372 10312
rect 69292 10268 69332 10312
rect 69763 10268 69821 10269
rect 68803 10228 68812 10268
rect 68852 10228 69100 10268
rect 69140 10228 69149 10268
rect 69292 10228 69772 10268
rect 69812 10228 70348 10268
rect 70388 10228 70397 10268
rect 76483 10228 76492 10268
rect 76532 10228 77836 10268
rect 77876 10228 77885 10268
rect 69763 10227 69821 10228
rect 36451 10144 36460 10184
rect 36500 10144 37228 10184
rect 37268 10144 37277 10184
rect 41827 10144 41836 10184
rect 41876 10144 42316 10184
rect 42356 10144 42365 10184
rect 43180 10144 44812 10184
rect 44852 10144 46348 10184
rect 46388 10144 48940 10184
rect 48980 10144 48989 10184
rect 49795 10144 49804 10184
rect 49844 10144 52492 10184
rect 52532 10144 52541 10184
rect 58252 10144 58348 10184
rect 58388 10144 58397 10184
rect 58732 10144 61900 10184
rect 61940 10144 63436 10184
rect 63476 10144 63485 10184
rect 64579 10144 64588 10184
rect 64628 10144 65452 10184
rect 65492 10144 65501 10184
rect 68323 10144 68332 10184
rect 68372 10144 68381 10184
rect 68515 10144 68524 10184
rect 68564 10144 69484 10184
rect 69524 10144 69676 10184
rect 69716 10144 69725 10184
rect 70915 10144 70924 10184
rect 70964 10144 71308 10184
rect 71348 10144 71357 10184
rect 73420 10144 74764 10184
rect 74804 10144 78316 10184
rect 78356 10144 78365 10184
rect 39331 10100 39389 10101
rect 835 10060 844 10100
rect 884 10060 1516 10100
rect 1556 10060 1565 10100
rect 39246 10060 39340 10100
rect 39380 10060 39389 10100
rect 40963 10060 40972 10100
rect 41012 10060 41740 10100
rect 41780 10060 41789 10100
rect 52195 10060 52204 10100
rect 52244 10060 53164 10100
rect 53204 10060 53213 10100
rect 39331 10059 39389 10060
rect 50851 10016 50909 10017
rect 5059 9976 5068 10016
rect 5108 9976 7180 10016
rect 7220 9976 50860 10016
rect 50900 9976 50909 10016
rect 50851 9975 50909 9976
rect 0 9848 80 9868
rect 43171 9848 43229 9849
rect 58252 9848 58292 10144
rect 70435 10100 70493 10101
rect 73420 10100 73460 10144
rect 59491 10060 59500 10100
rect 59540 10060 60460 10100
rect 60500 10060 63628 10100
rect 63668 10060 63677 10100
rect 66883 10060 66892 10100
rect 66932 10060 68812 10100
rect 68852 10060 68861 10100
rect 68910 10060 68919 10100
rect 68959 10060 70156 10100
rect 70196 10060 70205 10100
rect 70350 10060 70444 10100
rect 70484 10060 70493 10100
rect 71779 10060 71788 10100
rect 71828 10060 72844 10100
rect 72884 10060 73460 10100
rect 77827 10060 77836 10100
rect 77876 10060 78028 10100
rect 78068 10060 79468 10100
rect 79508 10060 79517 10100
rect 69868 10016 69908 10060
rect 70435 10059 70493 10060
rect 63715 9976 63724 10016
rect 63764 9976 64492 10016
rect 64532 9976 64541 10016
rect 64963 9976 64972 10016
rect 65012 9976 65644 10016
rect 65684 9976 65693 10016
rect 68227 9976 68236 10016
rect 68276 9976 68716 10016
rect 68756 9976 68765 10016
rect 69859 9976 69868 10016
rect 69908 9976 69948 10016
rect 75523 9976 75532 10016
rect 75572 9976 76012 10016
rect 76052 9976 76061 10016
rect 69667 9892 69676 9932
rect 69716 9892 71788 9932
rect 71828 9892 71837 9932
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 2861 9808 2870 9848
rect 2910 9808 3436 9848
rect 3476 9808 3485 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 43171 9808 43180 9848
rect 43220 9808 44236 9848
rect 44276 9808 44285 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 58243 9808 58252 9848
rect 58292 9808 58301 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 0 9788 80 9808
rect 43171 9807 43229 9808
rect 40108 9724 42988 9764
rect 43028 9724 43037 9764
rect 53443 9724 53452 9764
rect 53492 9724 54124 9764
rect 54164 9724 56716 9764
rect 56756 9724 62476 9764
rect 62516 9724 62525 9764
rect 40108 9512 40148 9724
rect 40675 9640 40684 9680
rect 40724 9640 42700 9680
rect 42740 9640 42749 9680
rect 43075 9640 43084 9680
rect 43124 9640 43660 9680
rect 43700 9640 43852 9680
rect 43892 9640 43901 9680
rect 51436 9640 52012 9680
rect 52052 9640 52684 9680
rect 52724 9640 52733 9680
rect 58051 9640 58060 9680
rect 58100 9640 58348 9680
rect 58388 9640 58397 9680
rect 59299 9640 59308 9680
rect 59348 9640 59596 9680
rect 59636 9640 59645 9680
rect 64099 9640 64108 9680
rect 64148 9640 64780 9680
rect 64820 9640 64829 9680
rect 70627 9640 70636 9680
rect 70676 9640 71060 9680
rect 71107 9640 71116 9680
rect 71156 9640 71980 9680
rect 72020 9640 76492 9680
rect 76532 9640 76541 9680
rect 77347 9640 77356 9680
rect 77396 9640 77405 9680
rect 40867 9556 40876 9596
rect 40916 9556 41260 9596
rect 41300 9556 42988 9596
rect 43028 9556 43037 9596
rect 51436 9512 51476 9640
rect 71020 9596 71060 9640
rect 52099 9556 52108 9596
rect 52148 9556 52436 9596
rect 62179 9556 62188 9596
rect 62228 9556 64876 9596
rect 64916 9556 64925 9596
rect 69571 9556 69580 9596
rect 69620 9556 70348 9596
rect 70388 9556 70828 9596
rect 70868 9556 70877 9596
rect 71020 9556 71308 9596
rect 71348 9556 71357 9596
rect 52396 9512 52436 9556
rect 3715 9472 3724 9512
rect 3764 9472 4588 9512
rect 4628 9472 4637 9512
rect 40099 9472 40108 9512
rect 40148 9472 40157 9512
rect 40771 9472 40780 9512
rect 40820 9472 41356 9512
rect 41396 9472 42892 9512
rect 42932 9472 45484 9512
rect 45524 9472 45533 9512
rect 46723 9472 46732 9512
rect 46772 9472 47116 9512
rect 47156 9472 47165 9512
rect 50275 9472 50284 9512
rect 50324 9472 51436 9512
rect 51476 9472 51485 9512
rect 51715 9472 51724 9512
rect 51764 9472 52204 9512
rect 52244 9472 52253 9512
rect 52387 9472 52396 9512
rect 52436 9472 53068 9512
rect 53108 9472 53117 9512
rect 53260 9472 53356 9512
rect 53396 9472 54316 9512
rect 54356 9472 54365 9512
rect 58627 9472 58636 9512
rect 58676 9472 59692 9512
rect 59732 9472 59741 9512
rect 60835 9472 60844 9512
rect 60884 9472 62092 9512
rect 62132 9472 63436 9512
rect 63476 9472 66508 9512
rect 66548 9472 66557 9512
rect 69955 9472 69964 9512
rect 70004 9472 70013 9512
rect 70243 9472 70252 9512
rect 70292 9472 70924 9512
rect 70964 9472 70973 9512
rect 71875 9472 71884 9512
rect 71924 9472 74092 9512
rect 74132 9472 74141 9512
rect 75235 9472 75244 9512
rect 75284 9472 75724 9512
rect 75764 9472 75773 9512
rect 76771 9472 76780 9512
rect 76820 9472 77068 9512
rect 77108 9472 77117 9512
rect 53260 9428 53300 9472
rect 69964 9428 70004 9472
rect 835 9388 844 9428
rect 884 9388 4148 9428
rect 44227 9388 44236 9428
rect 44276 9388 47020 9428
rect 47060 9388 47980 9428
rect 48020 9388 48029 9428
rect 51619 9388 51628 9428
rect 51668 9388 52876 9428
rect 52916 9388 53300 9428
rect 69763 9388 69772 9428
rect 69812 9388 69908 9428
rect 69964 9388 71348 9428
rect 71683 9388 71692 9428
rect 71732 9388 71980 9428
rect 72020 9388 72029 9428
rect 76194 9388 76203 9428
rect 76243 9388 77260 9428
rect 77300 9388 77309 9428
rect 4108 9344 4148 9388
rect 2755 9304 2764 9344
rect 2804 9304 3532 9344
rect 3572 9304 3581 9344
rect 4099 9304 4108 9344
rect 4148 9304 4157 9344
rect 41539 9304 41548 9344
rect 41588 9304 41932 9344
rect 41972 9304 41981 9344
rect 42979 9304 42988 9344
rect 43028 9304 45580 9344
rect 45620 9304 45629 9344
rect 63523 9304 63532 9344
rect 63572 9304 64300 9344
rect 64340 9304 64349 9344
rect 69868 9260 69908 9388
rect 71308 9344 71348 9388
rect 69955 9304 69964 9344
rect 70004 9304 70540 9344
rect 70580 9304 70589 9344
rect 71299 9304 71308 9344
rect 71348 9304 71357 9344
rect 75724 9304 76684 9344
rect 76724 9304 76733 9344
rect 75724 9260 75764 9304
rect 77356 9260 77396 9640
rect 77443 9472 77452 9512
rect 77492 9472 77644 9512
rect 77684 9472 77693 9512
rect 42307 9220 42316 9260
rect 42356 9220 44044 9260
rect 44084 9220 44524 9260
rect 44564 9220 44573 9260
rect 46339 9220 46348 9260
rect 46388 9220 46732 9260
rect 46772 9220 46781 9260
rect 63619 9220 63628 9260
rect 63668 9220 64780 9260
rect 64820 9220 64829 9260
rect 69571 9220 69580 9260
rect 69620 9220 69772 9260
rect 69812 9220 69821 9260
rect 69868 9220 70252 9260
rect 70292 9220 70301 9260
rect 75715 9220 75724 9260
rect 75764 9220 75773 9260
rect 76483 9220 76492 9260
rect 76532 9220 77740 9260
rect 77780 9220 77789 9260
rect 835 9136 844 9176
rect 884 9136 1612 9176
rect 1652 9136 1661 9176
rect 62851 9136 62860 9176
rect 62900 9136 67756 9176
rect 67796 9136 67805 9176
rect 73507 9136 73516 9176
rect 73556 9136 76012 9176
rect 76052 9136 76061 9176
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 52675 9052 52684 9092
rect 52724 9052 53164 9092
rect 53204 9052 58348 9092
rect 58388 9052 58397 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 0 9008 80 9028
rect 2563 9008 2621 9009
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 2478 8968 2572 9008
rect 2612 8968 2621 9008
rect 54019 8968 54028 9008
rect 54068 8968 59020 9008
rect 59060 8968 59069 9008
rect 75427 8968 75436 9008
rect 75476 8968 75820 9008
rect 75860 8968 75869 9008
rect 0 8948 80 8968
rect 2563 8967 2621 8968
rect 2755 8884 2764 8924
rect 2804 8884 3340 8924
rect 3380 8884 3389 8924
rect 58051 8884 58060 8924
rect 58100 8884 58732 8924
rect 58772 8884 58781 8924
rect 63811 8884 63820 8924
rect 63860 8884 64588 8924
rect 64628 8884 64637 8924
rect 75907 8884 75916 8924
rect 75956 8884 76300 8924
rect 76340 8884 76349 8924
rect 77731 8884 77740 8924
rect 77780 8884 79468 8924
rect 79508 8884 79517 8924
rect 2947 8840 3005 8841
rect 2928 8800 2956 8840
rect 2996 8800 3052 8840
rect 3092 8800 5068 8840
rect 5108 8800 5117 8840
rect 57763 8800 57772 8840
rect 57812 8800 57821 8840
rect 57955 8800 57964 8840
rect 58004 8800 58772 8840
rect 64483 8800 64492 8840
rect 64532 8800 64972 8840
rect 65012 8800 66124 8840
rect 66164 8800 66173 8840
rect 68707 8800 68716 8840
rect 68756 8800 70156 8840
rect 70196 8800 70205 8840
rect 76867 8800 76876 8840
rect 76916 8800 77644 8840
rect 77684 8800 77693 8840
rect 2947 8799 3005 8800
rect 1699 8716 1708 8756
rect 1748 8716 2956 8756
rect 2996 8716 3148 8756
rect 3188 8716 3197 8756
rect 41539 8716 41548 8756
rect 41588 8716 42508 8756
rect 42548 8716 42557 8756
rect 44131 8716 44140 8756
rect 44180 8716 46924 8756
rect 46964 8716 48460 8756
rect 48500 8716 48509 8756
rect 2371 8632 2380 8672
rect 2420 8632 3724 8672
rect 3764 8632 3773 8672
rect 42787 8632 42796 8672
rect 42836 8632 45388 8672
rect 45428 8632 46636 8672
rect 46676 8632 48076 8672
rect 48116 8632 48125 8672
rect 57772 8588 57812 8800
rect 58732 8756 58772 8800
rect 58723 8716 58732 8756
rect 58772 8716 59212 8756
rect 59252 8716 59261 8756
rect 69475 8716 69484 8756
rect 69524 8716 71404 8756
rect 71444 8716 71453 8756
rect 58627 8632 58636 8672
rect 58676 8632 59116 8672
rect 59156 8632 59540 8672
rect 60643 8632 60652 8672
rect 60692 8632 61900 8672
rect 61940 8632 62860 8672
rect 62900 8632 62909 8672
rect 63043 8632 63052 8672
rect 63092 8632 63916 8672
rect 63956 8632 63965 8672
rect 64387 8632 64396 8672
rect 64436 8632 65068 8672
rect 65108 8632 65117 8672
rect 66499 8632 66508 8672
rect 66548 8632 67276 8672
rect 67316 8632 68140 8672
rect 68180 8632 69676 8672
rect 69716 8632 69725 8672
rect 69859 8632 69868 8672
rect 69908 8632 70636 8672
rect 70676 8632 70924 8672
rect 70964 8632 70973 8672
rect 71107 8632 71116 8672
rect 71156 8632 71884 8672
rect 71924 8632 71933 8672
rect 77443 8632 77452 8672
rect 77492 8632 77836 8672
rect 77876 8632 77885 8672
rect 1027 8548 1036 8588
rect 1076 8548 2284 8588
rect 2324 8548 2333 8588
rect 44803 8548 44812 8588
rect 44852 8548 46828 8588
rect 46868 8548 46877 8588
rect 48547 8548 48556 8588
rect 48596 8548 49036 8588
rect 49076 8548 49085 8588
rect 52963 8548 52972 8588
rect 53012 8548 53356 8588
rect 53396 8548 53548 8588
rect 53588 8548 53597 8588
rect 55939 8548 55948 8588
rect 55988 8548 57812 8588
rect 51331 8504 51389 8505
rect 59500 8504 59540 8632
rect 70723 8548 70732 8588
rect 70772 8548 71212 8588
rect 71252 8548 71261 8588
rect 75619 8548 75628 8588
rect 75668 8548 76588 8588
rect 76628 8548 76637 8588
rect 69763 8504 69821 8505
rect 2659 8464 2668 8504
rect 2708 8464 2804 8504
rect 4099 8464 4108 8504
rect 4148 8464 7468 8504
rect 7508 8464 51340 8504
rect 51380 8464 51389 8504
rect 57859 8464 57868 8504
rect 57908 8464 58444 8504
rect 58484 8464 58493 8504
rect 59491 8464 59500 8504
rect 59540 8464 59549 8504
rect 69678 8464 69772 8504
rect 69812 8464 69821 8504
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 0 8108 80 8128
rect 2764 8084 2804 8464
rect 51331 8463 51389 8464
rect 69763 8463 69821 8464
rect 58147 8380 58156 8420
rect 58196 8380 58828 8420
rect 58868 8380 58877 8420
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 46828 8212 49036 8252
rect 49076 8212 49085 8252
rect 46828 8168 46868 8212
rect 44131 8128 44140 8168
rect 44180 8128 44908 8168
rect 44948 8128 44957 8168
rect 46243 8128 46252 8168
rect 46292 8128 46828 8168
rect 46868 8128 46877 8168
rect 47011 8128 47020 8168
rect 47060 8128 47500 8168
rect 47540 8128 47692 8168
rect 47732 8128 47741 8168
rect 48259 8128 48268 8168
rect 48308 8128 48844 8168
rect 48884 8128 51148 8168
rect 51188 8128 60748 8168
rect 60788 8128 60797 8168
rect 64963 8128 64972 8168
rect 65012 8128 66260 8168
rect 71395 8128 71404 8168
rect 71444 8128 71636 8168
rect 76963 8128 76972 8168
rect 77012 8128 77452 8168
rect 77492 8128 77501 8168
rect 47020 8084 47060 8128
rect 2755 8044 2764 8084
rect 2804 8044 2813 8084
rect 42403 8044 42412 8084
rect 42452 8044 44428 8084
rect 44468 8044 47060 8084
rect 52291 8044 52300 8084
rect 52340 8044 52588 8084
rect 52628 8044 53260 8084
rect 53300 8044 53309 8084
rect 53731 8044 53740 8084
rect 53780 8044 54124 8084
rect 54164 8044 54173 8084
rect 58051 8044 58060 8084
rect 58100 8044 58540 8084
rect 58580 8044 58589 8084
rect 63820 8044 65260 8084
rect 65300 8044 65740 8084
rect 65780 8044 65789 8084
rect 2563 8000 2621 8001
rect 4771 8000 4829 8001
rect 48931 8000 48989 8001
rect 63820 8000 63860 8044
rect 66220 8000 66260 8128
rect 68323 8044 68332 8084
rect 68372 8044 69388 8084
rect 69428 8044 69437 8084
rect 71596 8000 71636 8128
rect 73603 8044 73612 8084
rect 73652 8044 76300 8084
rect 76340 8044 76349 8084
rect 2478 7960 2572 8000
rect 2612 7960 2621 8000
rect 2869 7960 2878 8000
rect 2918 7960 3724 8000
rect 3764 7960 3773 8000
rect 4291 7960 4300 8000
rect 4340 7960 4780 8000
rect 4820 7960 4829 8000
rect 45667 7960 45676 8000
rect 45716 7960 46540 8000
rect 46580 7960 46732 8000
rect 46772 7960 46781 8000
rect 47299 7960 47308 8000
rect 47348 7960 48556 8000
rect 48596 7960 48605 8000
rect 48846 7960 48940 8000
rect 48980 7960 48989 8000
rect 49411 7960 49420 8000
rect 49460 7960 59596 8000
rect 59636 7960 59645 8000
rect 63811 7960 63820 8000
rect 63860 7960 63869 8000
rect 64387 7960 64396 8000
rect 64436 7960 64588 8000
rect 64628 7960 65068 8000
rect 65108 7960 65117 8000
rect 66211 7960 66220 8000
rect 66260 7960 68428 8000
rect 68468 7960 68477 8000
rect 71587 7960 71596 8000
rect 71636 7960 71645 8000
rect 75724 7960 76204 8000
rect 76244 7960 76253 8000
rect 76387 7960 76396 8000
rect 76436 7960 77164 8000
rect 77204 7960 77548 8000
rect 77588 7960 77597 8000
rect 2563 7959 2621 7960
rect 4771 7959 4829 7960
rect 48931 7959 48989 7960
rect 75724 7916 75764 7960
rect 54595 7876 54604 7916
rect 54644 7876 73036 7916
rect 73076 7876 73085 7916
rect 75715 7876 75724 7916
rect 75764 7876 75773 7916
rect 52963 7792 52972 7832
rect 53012 7792 53740 7832
rect 53780 7792 53789 7832
rect 65827 7792 65836 7832
rect 65876 7792 66124 7832
rect 66164 7792 66173 7832
rect 3619 7748 3677 7749
rect 931 7708 940 7748
rect 980 7708 1516 7748
rect 1556 7708 1565 7748
rect 3534 7708 3628 7748
rect 3668 7708 4972 7748
rect 5012 7708 7180 7748
rect 7220 7708 7229 7748
rect 45379 7708 45388 7748
rect 45428 7708 47500 7748
rect 47540 7708 47549 7748
rect 48259 7708 48268 7748
rect 48308 7708 48460 7748
rect 48500 7708 48509 7748
rect 48739 7708 48748 7748
rect 48788 7708 49076 7748
rect 58339 7708 58348 7748
rect 58388 7708 58828 7748
rect 58868 7708 58877 7748
rect 62179 7708 62188 7748
rect 62228 7708 63628 7748
rect 63668 7708 63677 7748
rect 69859 7708 69868 7748
rect 69908 7708 70348 7748
rect 70388 7708 70732 7748
rect 70772 7708 70781 7748
rect 75427 7708 75436 7748
rect 75476 7708 75628 7748
rect 75668 7708 76012 7748
rect 76052 7708 76061 7748
rect 3619 7707 3677 7708
rect 1027 7624 1036 7664
rect 1076 7624 1996 7664
rect 2036 7624 2878 7664
rect 2918 7624 2927 7664
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 49036 7412 49076 7708
rect 75811 7624 75820 7664
rect 75860 7624 76108 7664
rect 76148 7624 76157 7664
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 77059 7540 77068 7580
rect 77108 7540 77452 7580
rect 77492 7540 77501 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 50467 7456 50476 7496
rect 50516 7456 52876 7496
rect 52916 7456 52925 7496
rect 47491 7372 47500 7412
rect 47540 7372 47788 7412
rect 47828 7372 47980 7412
rect 48020 7372 48364 7412
rect 48404 7372 48413 7412
rect 49027 7372 49036 7412
rect 49076 7372 49085 7412
rect 77251 7372 77260 7412
rect 77300 7372 77452 7412
rect 77492 7372 77501 7412
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 53635 7288 53644 7328
rect 53684 7288 54220 7328
rect 54260 7288 54269 7328
rect 54403 7288 54412 7328
rect 54452 7288 54492 7328
rect 0 7268 80 7288
rect 48931 7244 48989 7245
rect 54412 7244 54452 7288
rect 547 7204 556 7244
rect 596 7204 844 7244
rect 884 7204 893 7244
rect 48739 7204 48748 7244
rect 48788 7204 48940 7244
rect 48980 7204 48989 7244
rect 53443 7204 53452 7244
rect 53492 7204 54892 7244
rect 54932 7204 54941 7244
rect 64675 7204 64684 7244
rect 64724 7204 65740 7244
rect 65780 7204 65789 7244
rect 76003 7204 76012 7244
rect 76052 7204 76492 7244
rect 76532 7204 76541 7244
rect 77452 7204 77836 7244
rect 77876 7204 77885 7244
rect 48931 7203 48989 7204
rect 77452 7160 77492 7204
rect 46627 7120 46636 7160
rect 46676 7120 47116 7160
rect 47156 7120 48364 7160
rect 48404 7120 49612 7160
rect 49652 7120 49996 7160
rect 50036 7120 50188 7160
rect 50228 7120 50860 7160
rect 50900 7120 51052 7160
rect 51092 7120 51724 7160
rect 51764 7120 55564 7160
rect 55604 7120 55613 7160
rect 59971 7120 59980 7160
rect 60020 7120 60212 7160
rect 60259 7120 60268 7160
rect 60308 7120 60652 7160
rect 60692 7120 60701 7160
rect 65059 7120 65068 7160
rect 65108 7120 66124 7160
rect 66164 7120 66173 7160
rect 67939 7120 67948 7160
rect 67988 7120 69580 7160
rect 69620 7120 70444 7160
rect 70484 7120 70493 7160
rect 70915 7120 70924 7160
rect 70964 7120 71404 7160
rect 71444 7120 71453 7160
rect 71875 7120 71884 7160
rect 71924 7120 72172 7160
rect 72212 7120 72221 7160
rect 75235 7120 75244 7160
rect 75284 7120 75532 7160
rect 75572 7120 75820 7160
rect 75860 7120 75869 7160
rect 77443 7120 77452 7160
rect 77492 7120 77501 7160
rect 60172 7076 60212 7120
rect 2371 7036 2380 7076
rect 2420 7036 4108 7076
rect 4148 7036 4492 7076
rect 4532 7036 4541 7076
rect 53058 7036 53067 7076
rect 53107 7036 53356 7076
rect 53396 7036 53405 7076
rect 59308 7036 60076 7076
rect 60116 7036 60125 7076
rect 60172 7036 61900 7076
rect 61940 7036 61949 7076
rect 64003 7036 64012 7076
rect 64052 7036 64876 7076
rect 64916 7036 64925 7076
rect 65347 7036 65356 7076
rect 65396 7036 66220 7076
rect 66260 7036 66269 7076
rect 66883 7036 66892 7076
rect 66932 7036 69196 7076
rect 69236 7036 69245 7076
rect 69955 7036 69964 7076
rect 70004 7036 71308 7076
rect 71348 7036 71788 7076
rect 71828 7036 71837 7076
rect 59308 6992 59348 7036
rect 59299 6952 59308 6992
rect 59348 6952 59357 6992
rect 64771 6952 64780 6992
rect 64820 6952 64829 6992
rect 64963 6952 64972 6992
rect 65012 6952 65932 6992
rect 65972 6952 66700 6992
rect 66740 6952 66749 6992
rect 69091 6952 69100 6992
rect 69140 6952 69908 6992
rect 64780 6908 64820 6952
rect 64003 6868 64012 6908
rect 64052 6868 64820 6908
rect 69868 6908 69908 6952
rect 69868 6868 70060 6908
rect 70100 6868 70252 6908
rect 70292 6868 70301 6908
rect 76003 6868 76012 6908
rect 76052 6868 76204 6908
rect 76244 6868 76588 6908
rect 76628 6868 76637 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 56995 6784 57004 6824
rect 57044 6784 62284 6824
rect 62324 6784 62333 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 2851 6700 2860 6740
rect 2900 6700 4876 6740
rect 4916 6700 4925 6740
rect 52387 6700 52396 6740
rect 52436 6700 54316 6740
rect 54356 6700 54365 6740
rect 59491 6700 59500 6740
rect 59540 6700 60076 6740
rect 60116 6700 60125 6740
rect 57955 6616 57964 6656
rect 58004 6616 58732 6656
rect 58772 6616 58781 6656
rect 59299 6616 59308 6656
rect 59348 6616 59980 6656
rect 60020 6616 60172 6656
rect 60212 6616 61420 6656
rect 61460 6616 61469 6656
rect 3523 6532 3532 6572
rect 3572 6532 4492 6572
rect 4532 6532 4541 6572
rect 46819 6532 46828 6572
rect 46868 6532 47924 6572
rect 54211 6532 54220 6572
rect 54260 6532 54604 6572
rect 54644 6532 54653 6572
rect 58051 6532 58060 6572
rect 58100 6532 58540 6572
rect 58580 6532 58589 6572
rect 59011 6532 59020 6572
rect 59060 6532 59500 6572
rect 59540 6532 64012 6572
rect 64052 6532 64061 6572
rect 0 6488 80 6508
rect 47884 6488 47924 6532
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 2659 6448 2668 6488
rect 2708 6448 2804 6488
rect 3043 6448 3052 6488
rect 3092 6448 4204 6488
rect 4244 6448 5068 6488
rect 5108 6448 7372 6488
rect 7412 6448 7421 6488
rect 45571 6448 45580 6488
rect 45620 6448 47404 6488
rect 47444 6448 47453 6488
rect 47875 6448 47884 6488
rect 47924 6448 47933 6488
rect 51427 6448 51436 6488
rect 51476 6448 52492 6488
rect 52532 6448 52541 6488
rect 52675 6448 52684 6488
rect 52724 6448 55084 6488
rect 55124 6448 55852 6488
rect 55892 6448 57292 6488
rect 57332 6448 58156 6488
rect 58196 6448 58205 6488
rect 58819 6448 58828 6488
rect 58868 6448 59212 6488
rect 59252 6448 59261 6488
rect 66019 6448 66028 6488
rect 66068 6448 66892 6488
rect 66932 6448 66941 6488
rect 69379 6448 69388 6488
rect 69428 6448 69676 6488
rect 69716 6448 69725 6488
rect 0 6428 80 6448
rect 1315 6280 1324 6320
rect 1364 6280 2188 6320
rect 2228 6280 2237 6320
rect 2467 6280 2476 6320
rect 2516 6280 2668 6320
rect 2708 6280 2717 6320
rect 2764 6236 2804 6448
rect 45475 6364 45484 6404
rect 45524 6364 47308 6404
rect 47348 6364 47357 6404
rect 47884 6320 47924 6448
rect 47884 6280 48940 6320
rect 48980 6280 48989 6320
rect 56899 6280 56908 6320
rect 56948 6280 58060 6320
rect 58100 6280 58109 6320
rect 58243 6280 58252 6320
rect 58292 6280 60268 6320
rect 60308 6280 60317 6320
rect 63331 6280 63340 6320
rect 63380 6280 63628 6320
rect 63668 6280 63677 6320
rect 68515 6280 68524 6320
rect 68564 6280 69388 6320
rect 69428 6280 69772 6320
rect 69812 6280 69821 6320
rect 2668 6196 2804 6236
rect 2668 6068 2708 6196
rect 51235 6112 51244 6152
rect 51284 6112 61804 6152
rect 61844 6112 61853 6152
rect 2659 6028 2668 6068
rect 2708 6028 2717 6068
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 58051 6028 58060 6068
rect 58100 6028 59020 6068
rect 59060 6028 59069 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 52579 5860 52588 5900
rect 52628 5860 52972 5900
rect 53012 5860 53021 5900
rect 61507 5860 61516 5900
rect 61556 5860 63724 5900
rect 63764 5860 67852 5900
rect 67892 5860 67901 5900
rect 69283 5860 69292 5900
rect 69332 5860 69772 5900
rect 69812 5860 69821 5900
rect 76003 5860 76012 5900
rect 76052 5860 76588 5900
rect 76628 5860 76637 5900
rect 4099 5776 4108 5816
rect 4148 5776 4157 5816
rect 47395 5776 47404 5816
rect 47444 5776 47596 5816
rect 47636 5776 47645 5816
rect 52771 5776 52780 5816
rect 52820 5776 52829 5816
rect 54403 5776 54412 5816
rect 54452 5776 54796 5816
rect 54836 5776 54845 5816
rect 64579 5776 64588 5816
rect 64628 5776 65068 5816
rect 65108 5776 65117 5816
rect 70819 5776 70828 5816
rect 70868 5776 71788 5816
rect 71828 5776 71837 5816
rect 74275 5776 74284 5816
rect 74324 5776 74333 5816
rect 76483 5776 76492 5816
rect 76532 5776 77740 5816
rect 77780 5776 79468 5816
rect 79508 5776 79517 5816
rect 4108 5732 4148 5776
rect 1795 5692 1804 5732
rect 1844 5692 2956 5732
rect 2996 5692 3628 5732
rect 3668 5692 4148 5732
rect 52780 5732 52820 5776
rect 52780 5692 53836 5732
rect 53876 5692 53885 5732
rect 54115 5692 54124 5732
rect 54164 5692 54700 5732
rect 54740 5692 57004 5732
rect 57044 5692 57053 5732
rect 64195 5692 64204 5732
rect 64244 5692 64492 5732
rect 64532 5692 65164 5732
rect 65204 5692 65213 5732
rect 65539 5692 65548 5732
rect 65588 5692 66124 5732
rect 66164 5692 66412 5732
rect 66452 5692 66461 5732
rect 69283 5692 69292 5732
rect 69332 5692 71404 5732
rect 71444 5692 71692 5732
rect 71732 5692 71741 5732
rect 0 5648 80 5668
rect 74284 5648 74324 5776
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 2467 5608 2476 5648
rect 2516 5608 4108 5648
rect 4148 5608 6220 5648
rect 6260 5608 6269 5648
rect 47299 5608 47308 5648
rect 47348 5608 47357 5648
rect 48451 5608 48460 5648
rect 48500 5608 50092 5648
rect 50132 5608 51244 5648
rect 51284 5608 51293 5648
rect 53059 5608 53068 5648
rect 53108 5608 53548 5648
rect 53588 5608 53740 5648
rect 53780 5608 54220 5648
rect 54260 5608 54269 5648
rect 54883 5608 54892 5648
rect 54932 5608 56236 5648
rect 56276 5608 58156 5648
rect 58196 5608 58924 5648
rect 58964 5608 58973 5648
rect 59395 5608 59404 5648
rect 59444 5608 61036 5648
rect 61076 5608 61085 5648
rect 61603 5608 61612 5648
rect 61652 5608 62572 5648
rect 62612 5608 62956 5648
rect 62996 5608 63436 5648
rect 63476 5608 64396 5648
rect 64436 5608 64445 5648
rect 64771 5608 64780 5648
rect 64820 5608 66316 5648
rect 66356 5608 66604 5648
rect 66644 5608 66653 5648
rect 71491 5608 71500 5648
rect 71540 5608 72268 5648
rect 72308 5608 74324 5648
rect 75619 5608 75628 5648
rect 75668 5608 76204 5648
rect 76244 5608 76253 5648
rect 76387 5608 76396 5648
rect 76436 5608 77260 5648
rect 77300 5608 77309 5648
rect 0 5588 80 5608
rect 47308 5480 47348 5608
rect 61036 5564 61076 5608
rect 49132 5524 52012 5564
rect 52052 5524 53164 5564
rect 53204 5524 53213 5564
rect 61036 5524 62284 5564
rect 62324 5524 62333 5564
rect 73603 5524 73612 5564
rect 73652 5524 76300 5564
rect 76340 5524 76349 5564
rect 49132 5480 49172 5524
rect 52396 5480 52436 5524
rect 7363 5440 7372 5480
rect 7412 5440 43220 5480
rect 47308 5440 47500 5480
rect 47540 5440 47549 5480
rect 49123 5440 49132 5480
rect 49172 5440 49181 5480
rect 52387 5440 52396 5480
rect 52436 5440 52476 5480
rect 58915 5440 58924 5480
rect 58964 5440 59308 5480
rect 59348 5440 59357 5480
rect 64867 5440 64876 5480
rect 64916 5440 65836 5480
rect 65876 5440 65885 5480
rect 43180 5396 43220 5440
rect 51043 5396 51101 5397
rect 43180 5356 51052 5396
rect 51092 5356 51101 5396
rect 59395 5356 59404 5396
rect 59444 5356 59884 5396
rect 59924 5356 60844 5396
rect 60884 5356 60893 5396
rect 51043 5355 51101 5356
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 59299 5188 59308 5228
rect 59348 5188 59692 5228
rect 59732 5188 59741 5228
rect 64291 5188 64300 5228
rect 64340 5188 65260 5228
rect 65300 5188 65309 5228
rect 1219 5104 1228 5144
rect 1268 5104 2284 5144
rect 2324 5104 2333 5144
rect 2467 5104 2476 5144
rect 2516 5104 2525 5144
rect 60163 5104 60172 5144
rect 60212 5104 60460 5144
rect 60500 5104 62380 5144
rect 62420 5104 62429 5144
rect 76099 5104 76108 5144
rect 76148 5104 76492 5144
rect 76532 5104 76541 5144
rect 2476 5060 2516 5104
rect 2284 5020 2516 5060
rect 45859 5020 45868 5060
rect 45908 5020 47308 5060
rect 47348 5020 47357 5060
rect 48547 5020 48556 5060
rect 48596 5020 48636 5060
rect 51820 5020 53300 5060
rect 63139 5020 63148 5060
rect 63188 5020 64684 5060
rect 64724 5020 64733 5060
rect 70348 5020 72076 5060
rect 72116 5020 72125 5060
rect 1795 4852 1804 4892
rect 1844 4852 2188 4892
rect 2228 4852 2237 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 2284 4724 2324 5020
rect 48556 4976 48596 5020
rect 51820 4976 51860 5020
rect 53260 4976 53300 5020
rect 70348 4976 70388 5020
rect 48259 4936 48268 4976
rect 48308 4936 48844 4976
rect 48884 4936 48893 4976
rect 51811 4936 51820 4976
rect 51860 4936 51869 4976
rect 52675 4936 52684 4976
rect 52724 4936 52733 4976
rect 53260 4936 54028 4976
rect 54068 4936 55660 4976
rect 55700 4936 55709 4976
rect 55939 4936 55948 4976
rect 55988 4936 56332 4976
rect 56372 4936 56381 4976
rect 57571 4936 57580 4976
rect 57620 4936 60172 4976
rect 60212 4936 60940 4976
rect 60980 4936 61612 4976
rect 61652 4936 61661 4976
rect 65923 4936 65932 4976
rect 65972 4936 66604 4976
rect 66644 4936 66653 4976
rect 68707 4936 68716 4976
rect 68756 4936 69100 4976
rect 69140 4936 70348 4976
rect 70388 4936 70397 4976
rect 71107 4936 71116 4976
rect 71156 4936 71596 4976
rect 71636 4936 71645 4976
rect 71875 4936 71884 4976
rect 71924 4936 72172 4976
rect 72212 4936 72221 4976
rect 52684 4892 52724 4936
rect 49219 4852 49228 4892
rect 49268 4852 49277 4892
rect 52684 4852 53644 4892
rect 53684 4852 56716 4892
rect 56756 4852 56765 4892
rect 63340 4852 67660 4892
rect 67700 4852 67709 4892
rect 49228 4808 49268 4852
rect 63340 4808 63380 4852
rect 2371 4768 2380 4808
rect 2420 4768 3820 4808
rect 3860 4768 4780 4808
rect 4820 4768 4829 4808
rect 47395 4768 47404 4808
rect 47444 4768 48556 4808
rect 48596 4768 49268 4808
rect 55651 4768 55660 4808
rect 55700 4768 56140 4808
rect 56180 4768 56189 4808
rect 56515 4768 56524 4808
rect 56564 4768 58540 4808
rect 58580 4768 63380 4808
rect 64003 4768 64012 4808
rect 64052 4768 64204 4808
rect 64244 4768 65740 4808
rect 65780 4768 65789 4808
rect 77443 4768 77452 4808
rect 77492 4768 77836 4808
rect 77876 4768 77885 4808
rect 2284 4684 2476 4724
rect 2516 4684 2525 4724
rect 51811 4684 51820 4724
rect 51860 4684 52396 4724
rect 52436 4684 52445 4724
rect 67747 4684 67756 4724
rect 67796 4684 68908 4724
rect 68948 4684 68957 4724
rect 1891 4600 1900 4640
rect 1940 4600 2284 4640
rect 2324 4600 2333 4640
rect 62371 4600 62380 4640
rect 62420 4600 64436 4640
rect 64483 4600 64492 4640
rect 64532 4600 65260 4640
rect 65300 4600 65309 4640
rect 64396 4556 64436 4600
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 64396 4516 64684 4556
rect 64724 4516 66220 4556
rect 66260 4516 66269 4556
rect 68908 4516 69004 4556
rect 69044 4516 70252 4556
rect 70292 4516 72460 4556
rect 72500 4516 72509 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 68908 4472 68948 4516
rect 51715 4432 51724 4472
rect 51764 4432 53836 4472
rect 53876 4432 56236 4472
rect 56276 4432 57004 4472
rect 57044 4432 57053 4472
rect 60835 4432 60844 4472
rect 60884 4432 66124 4472
rect 66164 4432 66173 4472
rect 68899 4432 68908 4472
rect 68948 4432 68957 4472
rect 72268 4432 74380 4472
rect 74420 4432 75148 4472
rect 75188 4432 75197 4472
rect 72268 4388 72308 4432
rect 51523 4348 51532 4388
rect 51572 4348 52684 4388
rect 52724 4348 52733 4388
rect 55843 4348 55852 4388
rect 55892 4348 56812 4388
rect 56852 4348 57292 4388
rect 57332 4348 57341 4388
rect 61507 4348 61516 4388
rect 61556 4348 62188 4388
rect 62228 4348 62237 4388
rect 72259 4348 72268 4388
rect 72308 4348 72317 4388
rect 72451 4348 72460 4388
rect 72500 4348 74860 4388
rect 74900 4348 74909 4388
rect 70147 4304 70205 4305
rect 72268 4304 72308 4348
rect 51619 4264 51628 4304
rect 51668 4264 52588 4304
rect 52628 4264 52637 4304
rect 52771 4264 52780 4304
rect 52820 4264 52829 4304
rect 57379 4264 57388 4304
rect 57428 4264 57964 4304
rect 58004 4264 58013 4304
rect 58627 4264 58636 4304
rect 58676 4264 59212 4304
rect 59252 4264 62764 4304
rect 62804 4264 64396 4304
rect 64436 4264 64445 4304
rect 65827 4264 65836 4304
rect 65876 4264 66892 4304
rect 66932 4264 68812 4304
rect 68852 4264 70156 4304
rect 70196 4264 70205 4304
rect 71491 4264 71500 4304
rect 71540 4264 72308 4304
rect 76003 4264 76012 4304
rect 76052 4264 77644 4304
rect 77684 4264 77693 4304
rect 52780 4220 52820 4264
rect 70147 4263 70205 4264
rect 50755 4180 50764 4220
rect 50804 4180 55372 4220
rect 55412 4180 55756 4220
rect 55796 4180 55805 4220
rect 58723 4180 58732 4220
rect 58772 4180 59116 4220
rect 59156 4180 59165 4220
rect 59779 4180 59788 4220
rect 59828 4180 60844 4220
rect 60884 4180 63436 4220
rect 63476 4180 65644 4220
rect 65684 4180 65693 4220
rect 69475 4180 69484 4220
rect 69524 4180 69964 4220
rect 70004 4180 70013 4220
rect 76483 4180 76492 4220
rect 76532 4180 77260 4220
rect 77300 4180 79468 4220
rect 79508 4180 79517 4220
rect 4771 4136 4829 4137
rect 2083 4096 2092 4136
rect 2132 4096 2878 4136
rect 2918 4096 3916 4136
rect 3956 4096 3965 4136
rect 4579 4096 4588 4136
rect 4628 4096 4780 4136
rect 4820 4096 4829 4136
rect 52099 4096 52108 4136
rect 52148 4096 52588 4136
rect 52628 4096 53260 4136
rect 53300 4096 53309 4136
rect 53635 4096 53644 4136
rect 53684 4096 55084 4136
rect 55124 4096 55133 4136
rect 55651 4096 55660 4136
rect 55700 4096 57100 4136
rect 57140 4096 57149 4136
rect 58243 4096 58252 4136
rect 58292 4096 59020 4136
rect 59060 4096 61228 4136
rect 61268 4096 61277 4136
rect 75907 4096 75916 4136
rect 75956 4096 76300 4136
rect 76340 4096 76588 4136
rect 76628 4096 76637 4136
rect 4771 4095 4829 4096
rect 3811 4012 3820 4052
rect 3860 4012 5260 4052
rect 5300 4012 5309 4052
rect 55939 4012 55948 4052
rect 55988 4012 56620 4052
rect 56660 4012 56669 4052
rect 65251 4012 65260 4052
rect 65300 4012 65932 4052
rect 65972 4012 65981 4052
rect 69283 4012 69292 4052
rect 69332 4012 71692 4052
rect 71732 4012 71741 4052
rect 75331 4012 75340 4052
rect 75380 4012 77164 4052
rect 77204 4012 77213 4052
rect 0 3968 80 3988
rect 0 3928 1036 3968
rect 1076 3928 1085 3968
rect 50851 3928 50860 3968
rect 50900 3928 52972 3968
rect 53012 3928 55468 3968
rect 55508 3928 55852 3968
rect 55892 3928 55901 3968
rect 0 3908 80 3928
rect 52771 3844 52780 3884
rect 52820 3844 54796 3884
rect 54836 3844 62476 3884
rect 62516 3844 62525 3884
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 50179 3760 50188 3800
rect 50228 3760 51628 3800
rect 51668 3760 51677 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 59491 3676 59500 3716
rect 59540 3676 59788 3716
rect 59828 3676 62092 3716
rect 62132 3676 66988 3716
rect 67028 3676 67037 3716
rect 4003 3592 4012 3632
rect 4052 3592 4396 3632
rect 4436 3592 4445 3632
rect 53923 3592 53932 3632
rect 53972 3592 55948 3632
rect 55988 3592 55997 3632
rect 62851 3592 62860 3632
rect 62900 3592 64012 3632
rect 64052 3592 64061 3632
rect 68995 3592 69004 3632
rect 69044 3592 69388 3632
rect 69428 3592 69437 3632
rect 75427 3592 75436 3632
rect 75476 3592 76492 3632
rect 76532 3592 76541 3632
rect 50956 3508 52108 3548
rect 52148 3508 52157 3548
rect 56323 3508 56332 3548
rect 56372 3508 57196 3548
rect 57236 3508 57245 3548
rect 63916 3508 66316 3548
rect 66356 3508 66508 3548
rect 66548 3508 66557 3548
rect 70819 3508 70828 3548
rect 70868 3508 71212 3548
rect 71252 3508 71261 3548
rect 73795 3508 73804 3548
rect 73844 3508 75244 3548
rect 75284 3508 75293 3548
rect 50956 3464 50996 3508
rect 63916 3464 63956 3508
rect 2947 3424 2956 3464
rect 2996 3424 5068 3464
rect 5108 3424 5117 3464
rect 5251 3424 5260 3464
rect 5300 3424 7468 3464
rect 7508 3424 7517 3464
rect 50947 3424 50956 3464
rect 50996 3424 51005 3464
rect 52003 3424 52012 3464
rect 52052 3424 52780 3464
rect 52820 3424 52829 3464
rect 55171 3424 55180 3464
rect 55220 3424 55948 3464
rect 55988 3424 55997 3464
rect 59299 3424 59308 3464
rect 59348 3424 59980 3464
rect 60020 3424 61804 3464
rect 61844 3424 61853 3464
rect 63907 3424 63916 3464
rect 63956 3424 63965 3464
rect 64099 3424 64108 3464
rect 64148 3424 64300 3464
rect 64340 3424 64349 3464
rect 64579 3424 64588 3464
rect 64628 3424 65260 3464
rect 65300 3424 65309 3464
rect 66595 3424 66604 3464
rect 66644 3424 66653 3464
rect 68227 3424 68236 3464
rect 68276 3424 69868 3464
rect 69908 3424 69917 3464
rect 70051 3424 70060 3464
rect 70100 3424 71404 3464
rect 71444 3424 71596 3464
rect 71636 3424 72076 3464
rect 72116 3424 72125 3464
rect 74851 3424 74860 3464
rect 74900 3424 76396 3464
rect 76436 3424 76445 3464
rect 76579 3424 76588 3464
rect 76628 3424 77644 3464
rect 77684 3424 78604 3464
rect 78644 3424 78653 3464
rect 66604 3380 66644 3424
rect 76588 3380 76628 3424
rect 1219 3340 1228 3380
rect 1268 3340 2092 3380
rect 2132 3340 2141 3380
rect 64771 3340 64780 3380
rect 64820 3340 66644 3380
rect 74659 3340 74668 3380
rect 74708 3340 76628 3380
rect 4771 3296 4829 3297
rect 4579 3256 4588 3296
rect 4628 3256 4780 3296
rect 4820 3256 4829 3296
rect 4771 3255 4829 3256
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 56131 3172 56140 3212
rect 56180 3172 56716 3212
rect 56756 3172 56765 3212
rect 58819 3172 58828 3212
rect 58868 3172 59404 3212
rect 59444 3172 59453 3212
rect 68323 3172 68332 3212
rect 68372 3172 69964 3212
rect 70004 3172 71980 3212
rect 72020 3172 75820 3212
rect 75860 3172 75869 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 58723 3088 58732 3128
rect 58772 3088 63052 3128
rect 63092 3088 64492 3128
rect 64532 3088 64541 3128
rect 68899 3088 68908 3128
rect 68948 3088 71692 3128
rect 71732 3088 75340 3128
rect 75380 3088 76972 3128
rect 77012 3088 77836 3128
rect 77876 3088 77885 3128
rect 0 3068 80 3088
rect 64675 3044 64733 3045
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 59404 3004 60844 3044
rect 60884 3004 60893 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 64590 3004 64684 3044
rect 64724 3004 64733 3044
rect 68707 3004 68716 3044
rect 68756 3004 69004 3044
rect 69044 3004 69053 3044
rect 69859 3004 69868 3044
rect 69908 3004 71788 3044
rect 71828 3004 75724 3044
rect 75764 3004 75773 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 59404 2960 59444 3004
rect 64675 3003 64733 3004
rect 59395 2920 59404 2960
rect 59444 2920 59453 2960
rect 64195 2920 64204 2960
rect 64244 2920 66124 2960
rect 66164 2920 66173 2960
rect 59107 2836 59116 2876
rect 59156 2836 59692 2876
rect 59732 2836 59741 2876
rect 72259 2836 72268 2876
rect 72308 2836 76012 2876
rect 76052 2836 76780 2876
rect 76820 2836 76829 2876
rect 77251 2836 77260 2876
rect 77300 2836 78124 2876
rect 78164 2836 78173 2876
rect 835 2752 844 2792
rect 884 2752 1516 2792
rect 1556 2752 1565 2792
rect 72931 2752 72940 2792
rect 72980 2752 75148 2792
rect 75188 2752 75197 2792
rect 78211 2752 78220 2792
rect 78260 2752 79180 2792
rect 79220 2752 79229 2792
rect 1699 2668 1708 2708
rect 1748 2668 3148 2708
rect 3188 2668 8908 2708
rect 8948 2668 8957 2708
rect 52291 2668 52300 2708
rect 52340 2668 55756 2708
rect 55796 2668 57388 2708
rect 57428 2668 57437 2708
rect 64483 2668 64492 2708
rect 64532 2668 64780 2708
rect 64820 2668 64829 2708
rect 73123 2668 73132 2708
rect 73172 2668 73612 2708
rect 73652 2668 74380 2708
rect 74420 2668 74429 2708
rect 2563 2584 2572 2624
rect 2612 2584 4300 2624
rect 4340 2584 4780 2624
rect 4820 2584 4829 2624
rect 55939 2584 55948 2624
rect 55988 2584 56716 2624
rect 56756 2584 57292 2624
rect 57332 2584 58156 2624
rect 58196 2584 58205 2624
rect 58915 2584 58924 2624
rect 58964 2584 59212 2624
rect 59252 2584 60364 2624
rect 60404 2584 60413 2624
rect 63811 2584 63820 2624
rect 63860 2584 64684 2624
rect 64724 2584 64733 2624
rect 64867 2584 64876 2624
rect 64916 2584 65260 2624
rect 65300 2584 65309 2624
rect 67939 2584 67948 2624
rect 67988 2584 71212 2624
rect 71252 2584 71261 2624
rect 71971 2584 71980 2624
rect 72020 2584 72652 2624
rect 72692 2584 73804 2624
rect 73844 2584 73853 2624
rect 74179 2584 74188 2624
rect 74228 2584 75052 2624
rect 75092 2584 76876 2624
rect 76916 2584 76925 2624
rect 71212 2540 71252 2584
rect 1411 2500 1420 2540
rect 1460 2500 2476 2540
rect 2516 2500 2525 2540
rect 56611 2500 56620 2540
rect 56660 2500 57004 2540
rect 57044 2500 57053 2540
rect 66883 2500 66892 2540
rect 66932 2500 67468 2540
rect 67508 2500 67517 2540
rect 71212 2500 72268 2540
rect 72308 2500 72317 2540
rect 74083 2500 74092 2540
rect 74132 2500 75244 2540
rect 75284 2500 75293 2540
rect 76195 2500 76204 2540
rect 76244 2500 76684 2540
rect 76724 2500 77164 2540
rect 77204 2500 78028 2540
rect 78068 2500 78077 2540
rect 64675 2456 64733 2457
rect 56323 2416 56332 2456
rect 56372 2416 56524 2456
rect 56564 2416 56573 2456
rect 58819 2416 58828 2456
rect 58868 2416 59788 2456
rect 59828 2416 61516 2456
rect 61556 2416 61565 2456
rect 64590 2416 64684 2456
rect 64724 2416 64733 2456
rect 67363 2416 67372 2456
rect 67412 2416 68140 2456
rect 68180 2416 68189 2456
rect 64675 2415 64733 2416
rect 77731 2332 77740 2372
rect 77780 2332 78412 2372
rect 78452 2332 78461 2372
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 0 2228 80 2248
rect 72547 2164 72556 2204
rect 72596 2164 73132 2204
rect 73172 2164 73181 2204
rect 55555 2080 55564 2120
rect 55604 2080 55948 2120
rect 55988 2080 55997 2120
rect 56803 2080 56812 2120
rect 56852 2080 58924 2120
rect 58964 2080 58973 2120
rect 65251 2080 65260 2120
rect 65300 2080 66892 2120
rect 66932 2080 66941 2120
rect 68227 2080 68236 2120
rect 68276 2080 69196 2120
rect 69236 2080 71212 2120
rect 71252 2080 73036 2120
rect 73076 2080 73085 2120
rect 74179 2080 74188 2120
rect 74228 2080 74420 2120
rect 74380 2036 74420 2080
rect 75244 2080 77740 2120
rect 77780 2080 77789 2120
rect 67555 1996 67564 2036
rect 67604 1996 68524 2036
rect 68564 1996 68573 2036
rect 74371 1996 74380 2036
rect 74420 1996 74429 2036
rect 75244 1952 75284 2080
rect 77059 1996 77068 2036
rect 77108 1996 78932 2036
rect 78892 1952 78932 1996
rect 54787 1912 54796 1952
rect 54836 1912 55660 1952
rect 55700 1912 57772 1952
rect 57812 1912 57821 1952
rect 65731 1912 65740 1952
rect 65780 1912 67276 1952
rect 67316 1912 67468 1952
rect 67508 1912 70060 1952
rect 70100 1912 70252 1952
rect 70292 1912 72652 1952
rect 72692 1912 73324 1952
rect 73364 1912 73373 1952
rect 73795 1912 73804 1952
rect 73844 1912 74572 1952
rect 74612 1912 74621 1952
rect 75235 1912 75244 1952
rect 75284 1912 75293 1952
rect 75427 1912 75436 1952
rect 75476 1912 75916 1952
rect 75956 1912 75965 1952
rect 76867 1912 76876 1952
rect 76916 1912 78316 1952
rect 78356 1912 78365 1952
rect 78883 1912 78892 1952
rect 78932 1912 78941 1952
rect 68995 1828 69004 1868
rect 69044 1828 71116 1868
rect 71156 1828 73996 1868
rect 74036 1828 77260 1868
rect 77300 1828 77309 1868
rect 58915 1660 58924 1700
rect 58964 1660 68044 1700
rect 68084 1660 68093 1700
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 56323 1492 56332 1532
rect 56372 1492 56812 1532
rect 56852 1492 56861 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 55555 1408 55564 1448
rect 55604 1408 56236 1448
rect 56276 1408 56285 1448
rect 53539 1324 53548 1364
rect 53588 1324 55372 1364
rect 55412 1324 55421 1364
rect 61699 1324 61708 1364
rect 61748 1324 62572 1364
rect 62612 1324 62621 1364
rect 64003 1324 64012 1364
rect 64052 1324 65260 1364
rect 65300 1324 65309 1364
rect 71395 1324 71404 1364
rect 71444 1324 72460 1364
rect 72500 1324 72509 1364
rect 57475 1240 57484 1280
rect 57524 1240 59308 1280
rect 59348 1240 59357 1280
rect 59491 1240 59500 1280
rect 59540 1240 60748 1280
rect 60788 1240 60797 1280
rect 62371 1240 62380 1280
rect 62420 1240 64684 1280
rect 64724 1240 64733 1280
rect 70915 1240 70924 1280
rect 70964 1240 72076 1280
rect 72116 1240 73228 1280
rect 73268 1240 73277 1280
rect 78211 1240 78220 1280
rect 78260 1240 79468 1280
rect 79508 1240 79517 1280
rect 73420 1156 74092 1196
rect 74132 1156 74141 1196
rect 73420 1112 73460 1156
rect 55843 1072 55852 1112
rect 55892 1072 56236 1112
rect 56276 1072 57196 1112
rect 57236 1072 57245 1112
rect 63043 1072 63052 1112
rect 63092 1072 64108 1112
rect 64148 1072 64157 1112
rect 66019 1072 66028 1112
rect 66068 1072 67372 1112
rect 67412 1072 67421 1112
rect 69763 1072 69772 1112
rect 69812 1072 71020 1112
rect 71060 1072 71212 1112
rect 71252 1072 71261 1112
rect 71875 1072 71884 1112
rect 71924 1072 72460 1112
rect 72500 1072 72509 1112
rect 72643 1072 72652 1112
rect 72692 1072 73460 1112
rect 73987 1072 73996 1112
rect 74036 1072 75628 1112
rect 75668 1072 75677 1112
rect 75811 1072 75820 1112
rect 75860 1072 76108 1112
rect 76148 1072 76157 1112
rect 61987 988 61996 1028
rect 62036 988 64204 1028
rect 64244 988 64253 1028
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 59308 38116 59348 38156
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 73420 37276 73460 37316
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 73324 36856 73364 36896
rect 33868 36688 33908 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 76204 35848 76244 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 62860 35176 62900 35216
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 62764 34084 62804 34124
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 76684 33832 76724 33872
rect 62860 33748 62900 33788
rect 76972 33664 77012 33704
rect 71980 33580 72020 33620
rect 76684 33328 76724 33368
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 70636 33076 70676 33116
rect 70924 32572 70964 32612
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 49228 32320 49268 32360
rect 55660 32152 55700 32192
rect 70636 32068 70676 32108
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 56044 31732 56084 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 71020 31732 71060 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 71884 31648 71924 31688
rect 49228 31564 49268 31604
rect 71404 31564 71444 31604
rect 71980 31564 72020 31604
rect 76972 31564 77012 31604
rect 71980 31312 72020 31352
rect 62764 31228 62804 31268
rect 75532 31228 75572 31268
rect 71404 31060 71444 31100
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 54796 30808 54836 30848
rect 40876 30556 40916 30596
rect 63244 30556 63284 30596
rect 77164 30556 77204 30596
rect 71884 30472 71924 30512
rect 62764 30388 62804 30428
rect 51436 30304 51476 30344
rect 75532 30304 75572 30344
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 76972 30220 77012 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 55276 30136 55316 30176
rect 55084 30052 55124 30092
rect 55084 29884 55124 29924
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 55660 29632 55700 29672
rect 56044 29632 56084 29672
rect 63244 29632 63284 29672
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 71116 28960 71156 29000
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 54796 28708 54836 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 51436 28624 51476 28664
rect 55660 28372 55700 28412
rect 64588 28288 64628 28328
rect 71020 28288 71060 28328
rect 77164 28120 77204 28160
rect 51244 28036 51284 28076
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 50380 27952 50420 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 51724 27868 51764 27908
rect 40972 27616 41012 27656
rect 76204 27532 76244 27572
rect 40876 27448 40916 27488
rect 41260 27364 41300 27404
rect 50380 27364 50420 27404
rect 51724 27364 51764 27404
rect 52780 27448 52820 27488
rect 71116 27280 71156 27320
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 50284 26944 50324 26984
rect 51532 26860 51572 26900
rect 38956 26524 38996 26564
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 52972 26440 53012 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 41260 26104 41300 26144
rect 38956 26020 38996 26060
rect 52876 26020 52916 26060
rect 61036 26020 61076 26060
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 40972 25516 41012 25556
rect 55276 25264 55316 25304
rect 64588 25180 64628 25220
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 51436 24928 51476 24968
rect 59308 24928 59348 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 30796 24844 30836 24884
rect 50284 24592 50324 24632
rect 50380 24508 50420 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 52588 24004 52628 24044
rect 40972 23920 41012 23960
rect 50572 23920 50612 23960
rect 40492 23836 40532 23876
rect 51148 23752 51188 23792
rect 79084 23752 79124 23792
rect 58444 23668 58484 23708
rect 56332 23584 56372 23624
rect 56524 23584 56564 23624
rect 70924 23584 70964 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 40972 23416 41012 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 60556 23500 60596 23540
rect 56812 23416 56852 23456
rect 56044 23332 56084 23372
rect 51148 23164 51188 23204
rect 55276 23164 55316 23204
rect 56428 23248 56468 23288
rect 52492 23080 52532 23120
rect 50572 22996 50612 23036
rect 53260 22912 53300 22952
rect 58828 22828 58855 22868
rect 58855 22828 58868 22868
rect 54892 22744 54895 22784
rect 54895 22744 54932 22784
rect 60556 22744 60596 22784
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 30796 22492 30836 22532
rect 27724 22324 27764 22364
rect 28492 22240 28532 22280
rect 51916 22156 51956 22196
rect 52588 22156 52628 22196
rect 38956 22072 38996 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 27724 21904 27764 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 44044 21568 44084 21608
rect 52300 21568 52340 21608
rect 53068 21568 53108 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 50380 21400 50420 21440
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 40876 20644 40916 20684
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 33868 20056 33908 20096
rect 41740 19888 41780 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 51820 19468 51860 19508
rect 39340 19384 39380 19424
rect 51724 19048 51764 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 50572 18796 50612 18836
rect 51724 18712 51764 18752
rect 22348 18460 22388 18500
rect 23692 18460 23732 18500
rect 52396 18460 52436 18500
rect 50380 18208 50420 18248
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 52012 17956 52052 17996
rect 52204 17620 52244 17660
rect 25804 17536 25844 17576
rect 29548 17536 29588 17576
rect 49612 17452 49652 17492
rect 53068 17452 53108 17492
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 32716 17284 32756 17324
rect 41164 17284 41204 17324
rect 51628 17200 51668 17240
rect 53932 17200 53945 17240
rect 53945 17200 53972 17240
rect 55084 17200 55124 17240
rect 55468 17200 55508 17240
rect 55660 17200 55700 17240
rect 58252 17200 58292 17240
rect 51916 17116 51956 17156
rect 52588 17116 52628 17156
rect 53068 17116 53108 17156
rect 57868 17116 57908 17156
rect 22348 16864 22388 16904
rect 39724 16864 39764 16904
rect 36652 16780 36692 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 52684 16360 52724 16400
rect 61708 16276 61748 16316
rect 54700 16192 54740 16232
rect 55468 16192 55508 16232
rect 55660 16192 55700 16232
rect 58252 16192 58292 16232
rect 58540 16192 58580 16232
rect 64972 16192 65012 16232
rect 70156 16192 70196 16232
rect 78892 16192 78932 16232
rect 53260 16024 53300 16064
rect 67660 16024 67700 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 41740 15688 41780 15728
rect 52204 15688 52244 15728
rect 52972 15436 53012 15476
rect 51628 15184 51668 15224
rect 52780 15184 52820 15224
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 63340 14848 63380 14888
rect 67180 14764 67220 14804
rect 54700 14680 54740 14720
rect 32620 14512 32660 14552
rect 68332 14428 68372 14468
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 52012 14344 52052 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 52396 14008 52436 14048
rect 69196 13924 69236 13964
rect 68332 13756 68372 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 70444 13504 70484 13544
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 36556 12664 36596 12704
rect 76396 12748 76436 12788
rect 41740 12496 41780 12536
rect 2956 12412 2996 12452
rect 57772 12412 57812 12452
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 52876 11908 52916 11948
rect 3628 11740 3668 11780
rect 43084 11572 43124 11612
rect 70444 11404 70484 11444
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 36556 11068 36596 11108
rect 52012 10900 52052 10940
rect 76396 10816 76436 10856
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 58924 10228 58964 10268
rect 67660 10228 67700 10268
rect 69772 10228 69812 10268
rect 39340 10060 39380 10100
rect 50860 9976 50900 10016
rect 70444 10060 70484 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 43180 9808 43220 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 2572 8968 2612 9008
rect 2956 8800 2996 8840
rect 51340 8464 51380 8504
rect 69772 8464 69812 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 2572 7960 2612 8000
rect 4780 7960 4820 8000
rect 48940 7960 48980 8000
rect 3628 7708 3668 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 48940 7204 48980 7244
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 51052 5356 51092 5396
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 70156 4264 70196 4304
rect 4780 4096 4820 4136
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 4780 3256 4820 3296
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 64684 3004 64724 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 64684 2416 64724 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 59308 38156 59348 38165
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 33868 36728 33908 36737
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 30796 24884 30836 24893
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 30796 22532 30836 24844
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 30796 22483 30836 22492
rect 27724 22364 27764 22373
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 27724 21944 27764 22324
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 27724 18593 27764 21904
rect 28492 22280 28532 22289
rect 22347 18584 22389 18593
rect 22347 18544 22348 18584
rect 22388 18544 22389 18584
rect 22347 18535 22389 18544
rect 27723 18584 27765 18593
rect 27723 18544 27724 18584
rect 27764 18544 27765 18584
rect 27723 18535 27765 18544
rect 22348 18500 22388 18535
rect 28492 18509 28532 22240
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 33868 20096 33908 36688
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 49228 32360 49268 32369
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 49228 31604 49268 32320
rect 49228 31555 49268 31564
rect 55660 32192 55700 32201
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 54796 30848 54836 30857
rect 40876 30596 40916 30605
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 40876 27488 40916 30556
rect 51436 30344 51476 30353
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 51436 28664 51476 30304
rect 54796 28748 54836 30808
rect 55276 30176 55316 30185
rect 55084 30092 55124 30101
rect 55084 29924 55124 30052
rect 55084 29875 55124 29884
rect 54796 28699 54836 28708
rect 51436 28615 51476 28624
rect 51244 28076 51284 28085
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 50380 27992 50420 28001
rect 38956 26564 38996 26573
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 38956 26060 38996 26524
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 38956 22112 38996 26020
rect 40491 23876 40533 23885
rect 40491 23836 40492 23876
rect 40532 23836 40533 23876
rect 40491 23827 40533 23836
rect 40492 23742 40532 23827
rect 38956 22063 38996 22072
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 40876 20684 40916 27448
rect 40972 27656 41012 27665
rect 40972 25556 41012 27616
rect 41260 27404 41300 27413
rect 41260 26144 41300 27364
rect 50380 27404 50420 27952
rect 50420 27364 50516 27404
rect 50380 27355 50420 27364
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 50284 26984 50324 26993
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 41260 26095 41300 26104
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 40972 23960 41012 25516
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 50284 24632 50324 26944
rect 50284 24583 50324 24592
rect 50380 24548 50420 24557
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 40972 23456 41012 23920
rect 44043 23876 44085 23885
rect 44043 23836 44044 23876
rect 44084 23836 44085 23876
rect 44043 23827 44085 23836
rect 40972 23407 41012 23416
rect 44044 21608 44084 23827
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 44044 21559 44084 21568
rect 50380 21440 50420 24508
rect 50380 21391 50420 21400
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 40876 20635 40916 20644
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 33868 20047 33908 20056
rect 41740 19928 41780 19937
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 39340 19424 39380 19433
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 22348 16904 22388 18460
rect 23691 18500 23733 18509
rect 23691 18460 23692 18500
rect 23732 18460 23733 18500
rect 23691 18451 23733 18460
rect 28491 18500 28533 18509
rect 28491 18460 28492 18500
rect 28532 18460 28533 18500
rect 28491 18451 28533 18460
rect 23692 18366 23732 18451
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 29547 17660 29589 17669
rect 29547 17620 29548 17660
rect 29588 17620 29589 17660
rect 29547 17611 29589 17620
rect 25803 17576 25845 17585
rect 25803 17536 25804 17576
rect 25844 17536 25845 17576
rect 25803 17527 25845 17536
rect 29548 17576 29588 17611
rect 25804 17442 25844 17527
rect 29548 17525 29588 17536
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 32716 17324 32756 17333
rect 32716 16997 32756 17284
rect 32715 16988 32757 16997
rect 32715 16948 32716 16988
rect 32756 16948 32757 16988
rect 32715 16939 32757 16948
rect 22348 16855 22388 16864
rect 36651 16820 36693 16829
rect 36651 16780 36652 16820
rect 36692 16780 36693 16820
rect 36651 16771 36693 16780
rect 36652 16686 36692 16771
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 32619 14552 32661 14561
rect 32619 14512 32620 14552
rect 32660 14512 32661 14552
rect 32619 14503 32661 14512
rect 32620 14418 32660 14503
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 36556 12704 36596 12713
rect 2956 12452 2996 12461
rect 2572 9008 2612 9017
rect 2572 8000 2612 8968
rect 2956 8840 2996 12412
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 3628 11780 3668 11789
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 2956 8791 2996 8800
rect 2572 7951 2612 7960
rect 3628 7748 3668 11740
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 36556 11108 36596 12664
rect 36556 11059 36596 11068
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 39340 10100 39380 19384
rect 41164 17324 41204 17333
rect 41164 17165 41204 17284
rect 41163 17156 41205 17165
rect 41163 17116 41164 17156
rect 41204 17116 41205 17156
rect 41163 17107 41205 17116
rect 39723 16904 39765 16913
rect 39723 16864 39724 16904
rect 39764 16864 39765 16904
rect 39723 16855 39765 16864
rect 39724 16770 39764 16855
rect 41740 15728 41780 19888
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 50380 18248 50420 18257
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 49611 17660 49653 17669
rect 49611 17620 49612 17660
rect 49652 17620 49653 17660
rect 49611 17611 49653 17620
rect 49612 17492 49652 17611
rect 49612 17443 49652 17452
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 48939 17156 48981 17165
rect 48939 17116 48940 17156
rect 48980 17116 48981 17156
rect 48939 17107 48981 17116
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 48940 16577 48980 17107
rect 50380 16997 50420 18208
rect 49035 16988 49077 16997
rect 49035 16948 49036 16988
rect 49076 16948 49077 16988
rect 49035 16939 49077 16948
rect 50379 16988 50421 16997
rect 50379 16948 50380 16988
rect 50420 16948 50421 16988
rect 50379 16939 50421 16948
rect 49036 16661 49076 16939
rect 49035 16652 49077 16661
rect 49035 16612 49036 16652
rect 49076 16612 49077 16652
rect 49035 16603 49077 16612
rect 48939 16568 48981 16577
rect 48939 16528 48940 16568
rect 48980 16528 48981 16568
rect 48939 16519 48981 16528
rect 50476 16325 50516 27364
rect 50572 23960 50612 23969
rect 50572 23036 50612 23920
rect 51148 23792 51188 23801
rect 51051 23372 51093 23381
rect 51051 23332 51052 23372
rect 51092 23332 51093 23372
rect 51051 23323 51093 23332
rect 50859 23204 50901 23213
rect 50859 23164 50860 23204
rect 50900 23164 50901 23204
rect 50859 23155 50901 23164
rect 50572 22987 50612 22996
rect 50572 18836 50612 18845
rect 50572 17165 50612 18796
rect 50571 17156 50613 17165
rect 50571 17116 50572 17156
rect 50612 17116 50613 17156
rect 50571 17107 50613 17116
rect 50475 16316 50517 16325
rect 50475 16276 50476 16316
rect 50516 16276 50517 16316
rect 50475 16267 50517 16276
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 41740 12536 41780 15688
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 41740 12487 41780 12496
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 39340 10051 39380 10060
rect 43084 11612 43124 11621
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 43084 9848 43124 11572
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 50860 10016 50900 23155
rect 50860 9967 50900 9976
rect 43180 9848 43220 9857
rect 43084 9808 43180 9848
rect 34592 9799 34960 9808
rect 43180 9780 43220 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 3628 7699 3668 7708
rect 4780 8000 4820 8009
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4780 4136 4820 7960
rect 48940 8000 48980 8009
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 48940 7244 48980 7960
rect 48940 7195 48980 7204
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 51052 5396 51092 23323
rect 51148 23204 51188 23752
rect 51148 23155 51188 23164
rect 51244 14813 51284 28036
rect 51724 27908 51764 27917
rect 51724 27404 51764 27868
rect 51724 27355 51764 27364
rect 52780 27488 52820 27497
rect 51532 26900 51572 26909
rect 51436 24968 51476 24977
rect 51339 23288 51381 23297
rect 51339 23248 51340 23288
rect 51380 23248 51381 23288
rect 51339 23239 51381 23248
rect 51243 14804 51285 14813
rect 51243 14764 51244 14804
rect 51284 14764 51285 14804
rect 51243 14755 51285 14764
rect 51340 8504 51380 23239
rect 51436 13049 51476 24928
rect 51532 14897 51572 26860
rect 52588 24044 52628 24053
rect 52588 23801 52628 24004
rect 52587 23792 52629 23801
rect 52587 23752 52588 23792
rect 52628 23752 52629 23792
rect 52587 23743 52629 23752
rect 51819 23456 51861 23465
rect 51819 23416 51820 23456
rect 51860 23416 51861 23456
rect 51819 23407 51861 23416
rect 51820 19508 51860 23407
rect 52299 23120 52341 23129
rect 52299 23080 52300 23120
rect 52340 23080 52341 23120
rect 52299 23071 52341 23080
rect 52492 23120 52532 23129
rect 51915 22868 51957 22877
rect 51915 22828 51916 22868
rect 51956 22828 51957 22868
rect 51915 22819 51957 22828
rect 51916 22196 51956 22819
rect 51916 22147 51956 22156
rect 52300 21608 52340 23071
rect 52300 21559 52340 21568
rect 51820 19459 51860 19468
rect 51724 19088 51764 19097
rect 51724 18752 51764 19048
rect 51628 17240 51668 17249
rect 51628 15224 51668 17200
rect 51724 16241 51764 18712
rect 52396 18500 52436 18509
rect 52012 17996 52052 18005
rect 51915 17576 51957 17585
rect 51915 17536 51916 17576
rect 51956 17536 51957 17576
rect 51915 17527 51957 17536
rect 51916 17249 51956 17527
rect 51915 17240 51957 17249
rect 51915 17200 51916 17240
rect 51956 17200 51957 17240
rect 51915 17191 51957 17200
rect 51916 17156 51956 17191
rect 51916 17106 51956 17116
rect 51723 16232 51765 16241
rect 51723 16192 51724 16232
rect 51764 16192 51765 16232
rect 51723 16183 51765 16192
rect 51628 15175 51668 15184
rect 51531 14888 51573 14897
rect 51531 14848 51532 14888
rect 51572 14848 51573 14888
rect 51531 14839 51573 14848
rect 52012 14384 52052 17956
rect 52204 17660 52244 17669
rect 52204 15728 52244 17620
rect 52204 15679 52244 15688
rect 51435 13040 51477 13049
rect 51435 13000 51436 13040
rect 51476 13000 51477 13040
rect 51435 12991 51477 13000
rect 52012 10940 52052 14344
rect 52396 14048 52436 18460
rect 52492 14729 52532 23080
rect 52588 22196 52628 23743
rect 52588 22147 52628 22156
rect 52588 17156 52628 17167
rect 52588 17081 52628 17116
rect 52587 17072 52629 17081
rect 52587 17032 52588 17072
rect 52628 17032 52629 17072
rect 52587 17023 52629 17032
rect 52684 16400 52724 16409
rect 52684 16073 52724 16360
rect 52683 16064 52725 16073
rect 52683 16024 52684 16064
rect 52724 16024 52725 16064
rect 52683 16015 52725 16024
rect 52780 15224 52820 27448
rect 52972 26480 53012 26489
rect 52780 15175 52820 15184
rect 52876 26060 52916 26069
rect 52491 14720 52533 14729
rect 52491 14680 52492 14720
rect 52532 14680 52533 14720
rect 52491 14671 52533 14680
rect 52396 13999 52436 14008
rect 52876 11948 52916 26020
rect 52972 15476 53012 26440
rect 55276 25304 55316 30136
rect 55660 29672 55700 32152
rect 55660 28412 55700 29632
rect 56044 31772 56084 31781
rect 56044 29672 56084 31732
rect 56044 29623 56084 29632
rect 55660 28363 55700 28372
rect 55276 25255 55316 25264
rect 59308 24968 59348 38116
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 73420 37316 73460 37325
rect 73324 37276 73420 37316
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 73324 36896 73364 37276
rect 73420 37267 73460 37276
rect 73324 36847 73364 36856
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 76204 35888 76244 35897
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 62860 35216 62900 35225
rect 62764 34124 62804 34133
rect 62764 31268 62804 34084
rect 62860 33788 62900 35176
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 62860 33739 62900 33748
rect 71980 33620 72020 33629
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 70636 33116 70676 33125
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 70636 32108 70676 33076
rect 70636 32059 70676 32068
rect 70924 32612 70964 32621
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 62764 30428 62804 31228
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 62764 30379 62804 30388
rect 63244 30596 63284 30605
rect 63244 29672 63284 30556
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 63244 29623 63284 29632
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 64588 28328 64628 28337
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 59308 24919 59348 24928
rect 61036 26060 61076 26069
rect 61036 23885 61076 26020
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 64588 25220 64628 28288
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 64588 25171 64628 25180
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 61035 23876 61077 23885
rect 61035 23836 61036 23876
rect 61076 23836 61077 23876
rect 61035 23827 61077 23836
rect 58444 23708 58484 23717
rect 56332 23624 56372 23633
rect 56524 23624 56564 23633
rect 56372 23584 56524 23624
rect 56332 23575 56372 23584
rect 56524 23575 56564 23584
rect 56811 23456 56853 23465
rect 56811 23416 56812 23456
rect 56852 23416 56853 23456
rect 56811 23407 56853 23416
rect 56043 23372 56085 23381
rect 56043 23332 56044 23372
rect 56084 23332 56085 23372
rect 56043 23323 56085 23332
rect 56044 23238 56084 23323
rect 56812 23322 56852 23407
rect 56427 23288 56469 23297
rect 56427 23248 56428 23288
rect 56468 23248 56469 23288
rect 56427 23239 56469 23248
rect 55275 23204 55317 23213
rect 55275 23164 55276 23204
rect 55316 23164 55317 23204
rect 55275 23155 55317 23164
rect 54795 23120 54837 23129
rect 54795 23080 54796 23120
rect 54836 23080 54837 23120
rect 54795 23071 54837 23080
rect 53260 22952 53300 22961
rect 53068 22912 53260 22952
rect 53068 21608 53108 22912
rect 53260 22903 53300 22912
rect 54796 22784 54836 23071
rect 55276 23070 55316 23155
rect 56428 23154 56468 23239
rect 58444 22877 58484 23668
rect 70924 23624 70964 32572
rect 71020 31772 71060 31781
rect 71020 28328 71060 31732
rect 71884 31688 71924 31697
rect 71404 31604 71444 31613
rect 71404 31100 71444 31564
rect 71404 31051 71444 31060
rect 71884 30512 71924 31648
rect 71980 31604 72020 33580
rect 71980 31352 72020 31564
rect 71980 31303 72020 31312
rect 71884 30463 71924 30472
rect 75532 31268 75572 31277
rect 75532 30344 75572 31228
rect 75532 30295 75572 30304
rect 71020 28279 71060 28288
rect 71116 29000 71156 29009
rect 71116 27320 71156 28960
rect 76204 27572 76244 35848
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 76684 33872 76724 33881
rect 76684 33368 76724 33832
rect 76684 33319 76724 33328
rect 76972 33704 77012 33713
rect 76972 31604 77012 33664
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 76972 30260 77012 31564
rect 76972 30211 77012 30220
rect 77164 30596 77204 30605
rect 77164 28160 77204 30556
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 77164 28111 77204 28120
rect 76204 27523 76244 27532
rect 71116 27271 71156 27280
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 79083 23792 79125 23801
rect 79083 23752 79084 23792
rect 79124 23752 79125 23792
rect 79083 23743 79125 23752
rect 79084 23658 79124 23743
rect 70924 23575 70964 23584
rect 60556 23540 60596 23549
rect 58828 22877 58868 22962
rect 58443 22868 58485 22877
rect 58443 22828 58444 22868
rect 58484 22828 58485 22868
rect 58443 22819 58485 22828
rect 58827 22868 58869 22877
rect 58827 22828 58828 22868
rect 58868 22828 58869 22868
rect 58827 22819 58869 22828
rect 54892 22784 54932 22793
rect 54796 22744 54892 22784
rect 54892 22735 54932 22744
rect 60556 22784 60596 23500
rect 60556 22735 60596 22744
rect 53068 21559 53108 21568
rect 53068 17492 53108 17501
rect 53068 17156 53108 17452
rect 53931 17240 53973 17249
rect 53931 17200 53932 17240
rect 53972 17200 53973 17240
rect 53931 17191 53973 17200
rect 55084 17240 55124 17251
rect 53068 17107 53108 17116
rect 53932 17106 53972 17191
rect 55084 17165 55124 17200
rect 55468 17240 55508 17249
rect 55083 17156 55125 17165
rect 55083 17116 55084 17156
rect 55124 17116 55125 17156
rect 55083 17107 55125 17116
rect 55468 16997 55508 17200
rect 55660 17240 55700 17249
rect 55467 16988 55509 16997
rect 55467 16948 55468 16988
rect 55508 16948 55509 16988
rect 55467 16939 55509 16948
rect 54699 16652 54741 16661
rect 54699 16612 54700 16652
rect 54740 16612 54741 16652
rect 54699 16603 54741 16612
rect 54700 16232 54740 16603
rect 54700 16183 54740 16192
rect 55468 16232 55508 16939
rect 55660 16577 55700 17200
rect 58252 17240 58292 17249
rect 57868 17156 57908 17165
rect 57868 16913 57908 17116
rect 57867 16904 57909 16913
rect 57867 16864 57868 16904
rect 57908 16864 57909 16904
rect 57867 16855 57909 16864
rect 58252 16745 58292 17200
rect 78891 17072 78933 17081
rect 78891 17032 78892 17072
rect 78932 17032 78933 17072
rect 78891 17023 78933 17032
rect 58251 16736 58293 16745
rect 58251 16696 58252 16736
rect 58292 16696 58293 16736
rect 58251 16687 58293 16696
rect 55659 16568 55701 16577
rect 55659 16528 55660 16568
rect 55700 16528 55701 16568
rect 55659 16519 55701 16528
rect 55468 16183 55508 16192
rect 55660 16232 55700 16519
rect 55660 16183 55700 16192
rect 58252 16232 58292 16687
rect 61707 16316 61749 16325
rect 61707 16276 61708 16316
rect 61748 16276 61749 16316
rect 61707 16267 61749 16276
rect 58252 16183 58292 16192
rect 58540 16232 58580 16241
rect 53259 16064 53301 16073
rect 53259 16024 53260 16064
rect 53300 16024 53301 16064
rect 53259 16015 53301 16024
rect 53260 15930 53300 16015
rect 52972 15427 53012 15436
rect 54699 14720 54741 14729
rect 54699 14680 54700 14720
rect 54740 14680 54741 14720
rect 54699 14671 54741 14680
rect 54700 14586 54740 14671
rect 58540 14561 58580 16192
rect 61708 16182 61748 16267
rect 64971 16232 65013 16241
rect 64971 16192 64972 16232
rect 65012 16192 65013 16232
rect 64971 16183 65013 16192
rect 70156 16232 70196 16241
rect 64972 16098 65012 16183
rect 67660 16064 67700 16073
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 63339 14888 63381 14897
rect 63339 14848 63340 14888
rect 63380 14848 63381 14888
rect 63339 14839 63381 14848
rect 58923 14804 58965 14813
rect 58923 14764 58924 14804
rect 58964 14764 58965 14804
rect 58923 14755 58965 14764
rect 58539 14552 58581 14561
rect 58539 14512 58540 14552
rect 58580 14512 58581 14552
rect 58539 14503 58581 14512
rect 57771 13964 57813 13973
rect 57771 13924 57772 13964
rect 57812 13924 57813 13964
rect 57771 13915 57813 13924
rect 57772 13049 57812 13915
rect 57771 13040 57813 13049
rect 57771 13000 57772 13040
rect 57812 13000 57813 13040
rect 57771 12991 57813 13000
rect 57772 12452 57812 12991
rect 57772 12403 57812 12412
rect 52876 11899 52916 11908
rect 52012 10891 52052 10900
rect 58924 10268 58964 14755
rect 63340 14754 63380 14839
rect 67179 14804 67221 14813
rect 67179 14764 67180 14804
rect 67220 14764 67221 14804
rect 67179 14755 67221 14764
rect 67180 14670 67220 14755
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 58924 10219 58964 10228
rect 67660 10268 67700 16024
rect 68332 14468 68372 14477
rect 68332 13796 68372 14428
rect 69195 13964 69237 13973
rect 69195 13924 69196 13964
rect 69236 13924 69237 13964
rect 69195 13915 69237 13924
rect 69196 13830 69236 13915
rect 68332 13747 68372 13756
rect 67660 10219 67700 10228
rect 69772 10268 69812 10277
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 51340 8455 51380 8464
rect 69772 8504 69812 10228
rect 69772 8455 69812 8464
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 51052 5347 51092 5356
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 70156 4304 70196 16192
rect 78892 16232 78932 17023
rect 78892 16183 78932 16192
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 70444 13544 70484 13553
rect 70444 11444 70484 13504
rect 70444 10100 70484 11404
rect 76396 12788 76436 12797
rect 76396 10856 76436 12748
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 76396 10807 76436 10816
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 70444 10051 70484 10060
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 70156 4255 70196 4264
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4780 3296 4820 4096
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 4780 3247 4820 3256
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 64684 3044 64724 3053
rect 64684 2456 64724 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 64684 2407 64724 2416
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 22348 18544 22388 18584
rect 27724 18544 27764 18584
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 40492 23836 40532 23876
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 44044 23836 44084 23876
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 23692 18460 23732 18500
rect 28492 18460 28532 18500
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 29548 17620 29588 17660
rect 25804 17536 25844 17576
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 32716 16948 32756 16988
rect 36652 16780 36692 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 32620 14512 32660 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 41164 17116 41204 17156
rect 39724 16864 39764 16904
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 49612 17620 49652 17660
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 48940 17116 48980 17156
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 49036 16948 49076 16988
rect 50380 16948 50420 16988
rect 49036 16612 49076 16652
rect 48940 16528 48980 16568
rect 51052 23332 51092 23372
rect 50860 23164 50900 23204
rect 50572 17116 50612 17156
rect 50476 16276 50516 16316
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 51340 23248 51380 23288
rect 51244 14764 51284 14804
rect 52588 23752 52628 23792
rect 51820 23416 51860 23456
rect 52300 23080 52340 23120
rect 51916 22828 51956 22868
rect 51916 17536 51956 17576
rect 51916 17200 51956 17240
rect 51724 16192 51764 16232
rect 51532 14848 51572 14888
rect 51436 13000 51476 13040
rect 52588 17032 52628 17072
rect 52684 16024 52724 16064
rect 52492 14680 52532 14720
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 61036 23836 61076 23876
rect 56812 23416 56852 23456
rect 56044 23332 56084 23372
rect 56428 23248 56468 23288
rect 55276 23164 55316 23204
rect 54796 23080 54836 23120
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 79084 23752 79124 23792
rect 58444 22828 58484 22868
rect 58828 22828 58868 22868
rect 53932 17200 53972 17240
rect 55084 17116 55124 17156
rect 55468 16948 55508 16988
rect 54700 16612 54740 16652
rect 57868 16864 57908 16904
rect 78892 17032 78932 17072
rect 58252 16696 58292 16736
rect 55660 16528 55700 16568
rect 61708 16276 61748 16316
rect 53260 16024 53300 16064
rect 54700 14680 54740 14720
rect 64972 16192 65012 16232
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 63340 14848 63380 14888
rect 58924 14764 58964 14804
rect 58540 14512 58580 14552
rect 57772 13924 57812 13964
rect 57772 13000 57812 13040
rect 67180 14764 67220 14804
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 69196 13924 69236 13964
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 19463 38576 19510 38618
rect 19634 38576 19678 38618
rect 19802 38576 19849 38618
rect 19463 38536 19472 38576
rect 19634 38536 19636 38576
rect 19676 38536 19678 38576
rect 19840 38536 19849 38576
rect 19463 38494 19510 38536
rect 19634 38494 19678 38536
rect 19802 38494 19849 38536
rect 34583 38576 34630 38618
rect 34754 38576 34798 38618
rect 34922 38576 34969 38618
rect 34583 38536 34592 38576
rect 34754 38536 34756 38576
rect 34796 38536 34798 38576
rect 34960 38536 34969 38576
rect 34583 38494 34630 38536
rect 34754 38494 34798 38536
rect 34922 38494 34969 38536
rect 49703 38576 49750 38618
rect 49874 38576 49918 38618
rect 50042 38576 50089 38618
rect 49703 38536 49712 38576
rect 49874 38536 49876 38576
rect 49916 38536 49918 38576
rect 50080 38536 50089 38576
rect 49703 38494 49750 38536
rect 49874 38494 49918 38536
rect 50042 38494 50089 38536
rect 64823 38576 64870 38618
rect 64994 38576 65038 38618
rect 65162 38576 65209 38618
rect 64823 38536 64832 38576
rect 64994 38536 64996 38576
rect 65036 38536 65038 38576
rect 65200 38536 65209 38576
rect 64823 38494 64870 38536
rect 64994 38494 65038 38536
rect 65162 38494 65209 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 18223 37820 18270 37862
rect 18394 37820 18438 37862
rect 18562 37820 18609 37862
rect 18223 37780 18232 37820
rect 18394 37780 18396 37820
rect 18436 37780 18438 37820
rect 18600 37780 18609 37820
rect 18223 37738 18270 37780
rect 18394 37738 18438 37780
rect 18562 37738 18609 37780
rect 33343 37820 33390 37862
rect 33514 37820 33558 37862
rect 33682 37820 33729 37862
rect 33343 37780 33352 37820
rect 33514 37780 33516 37820
rect 33556 37780 33558 37820
rect 33720 37780 33729 37820
rect 33343 37738 33390 37780
rect 33514 37738 33558 37780
rect 33682 37738 33729 37780
rect 48463 37820 48510 37862
rect 48634 37820 48678 37862
rect 48802 37820 48849 37862
rect 48463 37780 48472 37820
rect 48634 37780 48636 37820
rect 48676 37780 48678 37820
rect 48840 37780 48849 37820
rect 48463 37738 48510 37780
rect 48634 37738 48678 37780
rect 48802 37738 48849 37780
rect 63583 37820 63630 37862
rect 63754 37820 63798 37862
rect 63922 37820 63969 37862
rect 63583 37780 63592 37820
rect 63754 37780 63756 37820
rect 63796 37780 63798 37820
rect 63960 37780 63969 37820
rect 63583 37738 63630 37780
rect 63754 37738 63798 37780
rect 63922 37738 63969 37780
rect 78703 37820 78750 37862
rect 78874 37820 78918 37862
rect 79042 37820 79089 37862
rect 78703 37780 78712 37820
rect 78874 37780 78876 37820
rect 78916 37780 78918 37820
rect 79080 37780 79089 37820
rect 78703 37738 78750 37780
rect 78874 37738 78918 37780
rect 79042 37738 79089 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 19463 37064 19510 37106
rect 19634 37064 19678 37106
rect 19802 37064 19849 37106
rect 19463 37024 19472 37064
rect 19634 37024 19636 37064
rect 19676 37024 19678 37064
rect 19840 37024 19849 37064
rect 19463 36982 19510 37024
rect 19634 36982 19678 37024
rect 19802 36982 19849 37024
rect 34583 37064 34630 37106
rect 34754 37064 34798 37106
rect 34922 37064 34969 37106
rect 34583 37024 34592 37064
rect 34754 37024 34756 37064
rect 34796 37024 34798 37064
rect 34960 37024 34969 37064
rect 34583 36982 34630 37024
rect 34754 36982 34798 37024
rect 34922 36982 34969 37024
rect 49703 37064 49750 37106
rect 49874 37064 49918 37106
rect 50042 37064 50089 37106
rect 49703 37024 49712 37064
rect 49874 37024 49876 37064
rect 49916 37024 49918 37064
rect 50080 37024 50089 37064
rect 49703 36982 49750 37024
rect 49874 36982 49918 37024
rect 50042 36982 50089 37024
rect 64823 37064 64870 37106
rect 64994 37064 65038 37106
rect 65162 37064 65209 37106
rect 64823 37024 64832 37064
rect 64994 37024 64996 37064
rect 65036 37024 65038 37064
rect 65200 37024 65209 37064
rect 64823 36982 64870 37024
rect 64994 36982 65038 37024
rect 65162 36982 65209 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 18223 36308 18270 36350
rect 18394 36308 18438 36350
rect 18562 36308 18609 36350
rect 18223 36268 18232 36308
rect 18394 36268 18396 36308
rect 18436 36268 18438 36308
rect 18600 36268 18609 36308
rect 18223 36226 18270 36268
rect 18394 36226 18438 36268
rect 18562 36226 18609 36268
rect 33343 36308 33390 36350
rect 33514 36308 33558 36350
rect 33682 36308 33729 36350
rect 33343 36268 33352 36308
rect 33514 36268 33516 36308
rect 33556 36268 33558 36308
rect 33720 36268 33729 36308
rect 33343 36226 33390 36268
rect 33514 36226 33558 36268
rect 33682 36226 33729 36268
rect 48463 36308 48510 36350
rect 48634 36308 48678 36350
rect 48802 36308 48849 36350
rect 48463 36268 48472 36308
rect 48634 36268 48636 36308
rect 48676 36268 48678 36308
rect 48840 36268 48849 36308
rect 48463 36226 48510 36268
rect 48634 36226 48678 36268
rect 48802 36226 48849 36268
rect 63583 36308 63630 36350
rect 63754 36308 63798 36350
rect 63922 36308 63969 36350
rect 63583 36268 63592 36308
rect 63754 36268 63756 36308
rect 63796 36268 63798 36308
rect 63960 36268 63969 36308
rect 63583 36226 63630 36268
rect 63754 36226 63798 36268
rect 63922 36226 63969 36268
rect 78703 36308 78750 36350
rect 78874 36308 78918 36350
rect 79042 36308 79089 36350
rect 78703 36268 78712 36308
rect 78874 36268 78876 36308
rect 78916 36268 78918 36308
rect 79080 36268 79089 36308
rect 78703 36226 78750 36268
rect 78874 36226 78918 36268
rect 79042 36226 79089 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 19463 35552 19510 35594
rect 19634 35552 19678 35594
rect 19802 35552 19849 35594
rect 19463 35512 19472 35552
rect 19634 35512 19636 35552
rect 19676 35512 19678 35552
rect 19840 35512 19849 35552
rect 19463 35470 19510 35512
rect 19634 35470 19678 35512
rect 19802 35470 19849 35512
rect 34583 35552 34630 35594
rect 34754 35552 34798 35594
rect 34922 35552 34969 35594
rect 34583 35512 34592 35552
rect 34754 35512 34756 35552
rect 34796 35512 34798 35552
rect 34960 35512 34969 35552
rect 34583 35470 34630 35512
rect 34754 35470 34798 35512
rect 34922 35470 34969 35512
rect 49703 35552 49750 35594
rect 49874 35552 49918 35594
rect 50042 35552 50089 35594
rect 49703 35512 49712 35552
rect 49874 35512 49876 35552
rect 49916 35512 49918 35552
rect 50080 35512 50089 35552
rect 49703 35470 49750 35512
rect 49874 35470 49918 35512
rect 50042 35470 50089 35512
rect 64823 35552 64870 35594
rect 64994 35552 65038 35594
rect 65162 35552 65209 35594
rect 64823 35512 64832 35552
rect 64994 35512 64996 35552
rect 65036 35512 65038 35552
rect 65200 35512 65209 35552
rect 64823 35470 64870 35512
rect 64994 35470 65038 35512
rect 65162 35470 65209 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 18223 34796 18270 34838
rect 18394 34796 18438 34838
rect 18562 34796 18609 34838
rect 18223 34756 18232 34796
rect 18394 34756 18396 34796
rect 18436 34756 18438 34796
rect 18600 34756 18609 34796
rect 18223 34714 18270 34756
rect 18394 34714 18438 34756
rect 18562 34714 18609 34756
rect 33343 34796 33390 34838
rect 33514 34796 33558 34838
rect 33682 34796 33729 34838
rect 33343 34756 33352 34796
rect 33514 34756 33516 34796
rect 33556 34756 33558 34796
rect 33720 34756 33729 34796
rect 33343 34714 33390 34756
rect 33514 34714 33558 34756
rect 33682 34714 33729 34756
rect 48463 34796 48510 34838
rect 48634 34796 48678 34838
rect 48802 34796 48849 34838
rect 48463 34756 48472 34796
rect 48634 34756 48636 34796
rect 48676 34756 48678 34796
rect 48840 34756 48849 34796
rect 48463 34714 48510 34756
rect 48634 34714 48678 34756
rect 48802 34714 48849 34756
rect 63583 34796 63630 34838
rect 63754 34796 63798 34838
rect 63922 34796 63969 34838
rect 63583 34756 63592 34796
rect 63754 34756 63756 34796
rect 63796 34756 63798 34796
rect 63960 34756 63969 34796
rect 63583 34714 63630 34756
rect 63754 34714 63798 34756
rect 63922 34714 63969 34756
rect 78703 34796 78750 34838
rect 78874 34796 78918 34838
rect 79042 34796 79089 34838
rect 78703 34756 78712 34796
rect 78874 34756 78876 34796
rect 78916 34756 78918 34796
rect 79080 34756 79089 34796
rect 78703 34714 78750 34756
rect 78874 34714 78918 34756
rect 79042 34714 79089 34756
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 19463 34040 19510 34082
rect 19634 34040 19678 34082
rect 19802 34040 19849 34082
rect 19463 34000 19472 34040
rect 19634 34000 19636 34040
rect 19676 34000 19678 34040
rect 19840 34000 19849 34040
rect 19463 33958 19510 34000
rect 19634 33958 19678 34000
rect 19802 33958 19849 34000
rect 34583 34040 34630 34082
rect 34754 34040 34798 34082
rect 34922 34040 34969 34082
rect 34583 34000 34592 34040
rect 34754 34000 34756 34040
rect 34796 34000 34798 34040
rect 34960 34000 34969 34040
rect 34583 33958 34630 34000
rect 34754 33958 34798 34000
rect 34922 33958 34969 34000
rect 49703 34040 49750 34082
rect 49874 34040 49918 34082
rect 50042 34040 50089 34082
rect 49703 34000 49712 34040
rect 49874 34000 49876 34040
rect 49916 34000 49918 34040
rect 50080 34000 50089 34040
rect 49703 33958 49750 34000
rect 49874 33958 49918 34000
rect 50042 33958 50089 34000
rect 64823 34040 64870 34082
rect 64994 34040 65038 34082
rect 65162 34040 65209 34082
rect 64823 34000 64832 34040
rect 64994 34000 64996 34040
rect 65036 34000 65038 34040
rect 65200 34000 65209 34040
rect 64823 33958 64870 34000
rect 64994 33958 65038 34000
rect 65162 33958 65209 34000
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 18223 33284 18270 33326
rect 18394 33284 18438 33326
rect 18562 33284 18609 33326
rect 18223 33244 18232 33284
rect 18394 33244 18396 33284
rect 18436 33244 18438 33284
rect 18600 33244 18609 33284
rect 18223 33202 18270 33244
rect 18394 33202 18438 33244
rect 18562 33202 18609 33244
rect 33343 33284 33390 33326
rect 33514 33284 33558 33326
rect 33682 33284 33729 33326
rect 33343 33244 33352 33284
rect 33514 33244 33516 33284
rect 33556 33244 33558 33284
rect 33720 33244 33729 33284
rect 33343 33202 33390 33244
rect 33514 33202 33558 33244
rect 33682 33202 33729 33244
rect 48463 33284 48510 33326
rect 48634 33284 48678 33326
rect 48802 33284 48849 33326
rect 48463 33244 48472 33284
rect 48634 33244 48636 33284
rect 48676 33244 48678 33284
rect 48840 33244 48849 33284
rect 48463 33202 48510 33244
rect 48634 33202 48678 33244
rect 48802 33202 48849 33244
rect 63583 33284 63630 33326
rect 63754 33284 63798 33326
rect 63922 33284 63969 33326
rect 63583 33244 63592 33284
rect 63754 33244 63756 33284
rect 63796 33244 63798 33284
rect 63960 33244 63969 33284
rect 63583 33202 63630 33244
rect 63754 33202 63798 33244
rect 63922 33202 63969 33244
rect 78703 33284 78750 33326
rect 78874 33284 78918 33326
rect 79042 33284 79089 33326
rect 78703 33244 78712 33284
rect 78874 33244 78876 33284
rect 78916 33244 78918 33284
rect 79080 33244 79089 33284
rect 78703 33202 78750 33244
rect 78874 33202 78918 33244
rect 79042 33202 79089 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 19463 32528 19510 32570
rect 19634 32528 19678 32570
rect 19802 32528 19849 32570
rect 19463 32488 19472 32528
rect 19634 32488 19636 32528
rect 19676 32488 19678 32528
rect 19840 32488 19849 32528
rect 19463 32446 19510 32488
rect 19634 32446 19678 32488
rect 19802 32446 19849 32488
rect 34583 32528 34630 32570
rect 34754 32528 34798 32570
rect 34922 32528 34969 32570
rect 34583 32488 34592 32528
rect 34754 32488 34756 32528
rect 34796 32488 34798 32528
rect 34960 32488 34969 32528
rect 34583 32446 34630 32488
rect 34754 32446 34798 32488
rect 34922 32446 34969 32488
rect 49703 32528 49750 32570
rect 49874 32528 49918 32570
rect 50042 32528 50089 32570
rect 49703 32488 49712 32528
rect 49874 32488 49876 32528
rect 49916 32488 49918 32528
rect 50080 32488 50089 32528
rect 49703 32446 49750 32488
rect 49874 32446 49918 32488
rect 50042 32446 50089 32488
rect 64823 32528 64870 32570
rect 64994 32528 65038 32570
rect 65162 32528 65209 32570
rect 64823 32488 64832 32528
rect 64994 32488 64996 32528
rect 65036 32488 65038 32528
rect 65200 32488 65209 32528
rect 64823 32446 64870 32488
rect 64994 32446 65038 32488
rect 65162 32446 65209 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 18223 31772 18270 31814
rect 18394 31772 18438 31814
rect 18562 31772 18609 31814
rect 18223 31732 18232 31772
rect 18394 31732 18396 31772
rect 18436 31732 18438 31772
rect 18600 31732 18609 31772
rect 18223 31690 18270 31732
rect 18394 31690 18438 31732
rect 18562 31690 18609 31732
rect 33343 31772 33390 31814
rect 33514 31772 33558 31814
rect 33682 31772 33729 31814
rect 33343 31732 33352 31772
rect 33514 31732 33516 31772
rect 33556 31732 33558 31772
rect 33720 31732 33729 31772
rect 33343 31690 33390 31732
rect 33514 31690 33558 31732
rect 33682 31690 33729 31732
rect 48463 31772 48510 31814
rect 48634 31772 48678 31814
rect 48802 31772 48849 31814
rect 48463 31732 48472 31772
rect 48634 31732 48636 31772
rect 48676 31732 48678 31772
rect 48840 31732 48849 31772
rect 48463 31690 48510 31732
rect 48634 31690 48678 31732
rect 48802 31690 48849 31732
rect 63583 31772 63630 31814
rect 63754 31772 63798 31814
rect 63922 31772 63969 31814
rect 63583 31732 63592 31772
rect 63754 31732 63756 31772
rect 63796 31732 63798 31772
rect 63960 31732 63969 31772
rect 63583 31690 63630 31732
rect 63754 31690 63798 31732
rect 63922 31690 63969 31732
rect 78703 31772 78750 31814
rect 78874 31772 78918 31814
rect 79042 31772 79089 31814
rect 78703 31732 78712 31772
rect 78874 31732 78876 31772
rect 78916 31732 78918 31772
rect 79080 31732 79089 31772
rect 78703 31690 78750 31732
rect 78874 31690 78918 31732
rect 79042 31690 79089 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 19463 31016 19510 31058
rect 19634 31016 19678 31058
rect 19802 31016 19849 31058
rect 19463 30976 19472 31016
rect 19634 30976 19636 31016
rect 19676 30976 19678 31016
rect 19840 30976 19849 31016
rect 19463 30934 19510 30976
rect 19634 30934 19678 30976
rect 19802 30934 19849 30976
rect 34583 31016 34630 31058
rect 34754 31016 34798 31058
rect 34922 31016 34969 31058
rect 34583 30976 34592 31016
rect 34754 30976 34756 31016
rect 34796 30976 34798 31016
rect 34960 30976 34969 31016
rect 34583 30934 34630 30976
rect 34754 30934 34798 30976
rect 34922 30934 34969 30976
rect 49703 31016 49750 31058
rect 49874 31016 49918 31058
rect 50042 31016 50089 31058
rect 49703 30976 49712 31016
rect 49874 30976 49876 31016
rect 49916 30976 49918 31016
rect 50080 30976 50089 31016
rect 49703 30934 49750 30976
rect 49874 30934 49918 30976
rect 50042 30934 50089 30976
rect 64823 31016 64870 31058
rect 64994 31016 65038 31058
rect 65162 31016 65209 31058
rect 64823 30976 64832 31016
rect 64994 30976 64996 31016
rect 65036 30976 65038 31016
rect 65200 30976 65209 31016
rect 64823 30934 64870 30976
rect 64994 30934 65038 30976
rect 65162 30934 65209 30976
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 18223 30260 18270 30302
rect 18394 30260 18438 30302
rect 18562 30260 18609 30302
rect 18223 30220 18232 30260
rect 18394 30220 18396 30260
rect 18436 30220 18438 30260
rect 18600 30220 18609 30260
rect 18223 30178 18270 30220
rect 18394 30178 18438 30220
rect 18562 30178 18609 30220
rect 33343 30260 33390 30302
rect 33514 30260 33558 30302
rect 33682 30260 33729 30302
rect 33343 30220 33352 30260
rect 33514 30220 33516 30260
rect 33556 30220 33558 30260
rect 33720 30220 33729 30260
rect 33343 30178 33390 30220
rect 33514 30178 33558 30220
rect 33682 30178 33729 30220
rect 48463 30260 48510 30302
rect 48634 30260 48678 30302
rect 48802 30260 48849 30302
rect 48463 30220 48472 30260
rect 48634 30220 48636 30260
rect 48676 30220 48678 30260
rect 48840 30220 48849 30260
rect 48463 30178 48510 30220
rect 48634 30178 48678 30220
rect 48802 30178 48849 30220
rect 63583 30260 63630 30302
rect 63754 30260 63798 30302
rect 63922 30260 63969 30302
rect 63583 30220 63592 30260
rect 63754 30220 63756 30260
rect 63796 30220 63798 30260
rect 63960 30220 63969 30260
rect 63583 30178 63630 30220
rect 63754 30178 63798 30220
rect 63922 30178 63969 30220
rect 78703 30260 78750 30302
rect 78874 30260 78918 30302
rect 79042 30260 79089 30302
rect 78703 30220 78712 30260
rect 78874 30220 78876 30260
rect 78916 30220 78918 30260
rect 79080 30220 79089 30260
rect 78703 30178 78750 30220
rect 78874 30178 78918 30220
rect 79042 30178 79089 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 19463 29504 19510 29546
rect 19634 29504 19678 29546
rect 19802 29504 19849 29546
rect 19463 29464 19472 29504
rect 19634 29464 19636 29504
rect 19676 29464 19678 29504
rect 19840 29464 19849 29504
rect 19463 29422 19510 29464
rect 19634 29422 19678 29464
rect 19802 29422 19849 29464
rect 34583 29504 34630 29546
rect 34754 29504 34798 29546
rect 34922 29504 34969 29546
rect 34583 29464 34592 29504
rect 34754 29464 34756 29504
rect 34796 29464 34798 29504
rect 34960 29464 34969 29504
rect 34583 29422 34630 29464
rect 34754 29422 34798 29464
rect 34922 29422 34969 29464
rect 49703 29504 49750 29546
rect 49874 29504 49918 29546
rect 50042 29504 50089 29546
rect 49703 29464 49712 29504
rect 49874 29464 49876 29504
rect 49916 29464 49918 29504
rect 50080 29464 50089 29504
rect 49703 29422 49750 29464
rect 49874 29422 49918 29464
rect 50042 29422 50089 29464
rect 64823 29504 64870 29546
rect 64994 29504 65038 29546
rect 65162 29504 65209 29546
rect 64823 29464 64832 29504
rect 64994 29464 64996 29504
rect 65036 29464 65038 29504
rect 65200 29464 65209 29504
rect 64823 29422 64870 29464
rect 64994 29422 65038 29464
rect 65162 29422 65209 29464
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 18223 28748 18270 28790
rect 18394 28748 18438 28790
rect 18562 28748 18609 28790
rect 18223 28708 18232 28748
rect 18394 28708 18396 28748
rect 18436 28708 18438 28748
rect 18600 28708 18609 28748
rect 18223 28666 18270 28708
rect 18394 28666 18438 28708
rect 18562 28666 18609 28708
rect 33343 28748 33390 28790
rect 33514 28748 33558 28790
rect 33682 28748 33729 28790
rect 33343 28708 33352 28748
rect 33514 28708 33516 28748
rect 33556 28708 33558 28748
rect 33720 28708 33729 28748
rect 33343 28666 33390 28708
rect 33514 28666 33558 28708
rect 33682 28666 33729 28708
rect 48463 28748 48510 28790
rect 48634 28748 48678 28790
rect 48802 28748 48849 28790
rect 48463 28708 48472 28748
rect 48634 28708 48636 28748
rect 48676 28708 48678 28748
rect 48840 28708 48849 28748
rect 48463 28666 48510 28708
rect 48634 28666 48678 28708
rect 48802 28666 48849 28708
rect 63583 28748 63630 28790
rect 63754 28748 63798 28790
rect 63922 28748 63969 28790
rect 63583 28708 63592 28748
rect 63754 28708 63756 28748
rect 63796 28708 63798 28748
rect 63960 28708 63969 28748
rect 63583 28666 63630 28708
rect 63754 28666 63798 28708
rect 63922 28666 63969 28708
rect 78703 28748 78750 28790
rect 78874 28748 78918 28790
rect 79042 28748 79089 28790
rect 78703 28708 78712 28748
rect 78874 28708 78876 28748
rect 78916 28708 78918 28748
rect 79080 28708 79089 28748
rect 78703 28666 78750 28708
rect 78874 28666 78918 28708
rect 79042 28666 79089 28708
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 19463 27992 19510 28034
rect 19634 27992 19678 28034
rect 19802 27992 19849 28034
rect 19463 27952 19472 27992
rect 19634 27952 19636 27992
rect 19676 27952 19678 27992
rect 19840 27952 19849 27992
rect 19463 27910 19510 27952
rect 19634 27910 19678 27952
rect 19802 27910 19849 27952
rect 34583 27992 34630 28034
rect 34754 27992 34798 28034
rect 34922 27992 34969 28034
rect 34583 27952 34592 27992
rect 34754 27952 34756 27992
rect 34796 27952 34798 27992
rect 34960 27952 34969 27992
rect 34583 27910 34630 27952
rect 34754 27910 34798 27952
rect 34922 27910 34969 27952
rect 49703 27992 49750 28034
rect 49874 27992 49918 28034
rect 50042 27992 50089 28034
rect 49703 27952 49712 27992
rect 49874 27952 49876 27992
rect 49916 27952 49918 27992
rect 50080 27952 50089 27992
rect 49703 27910 49750 27952
rect 49874 27910 49918 27952
rect 50042 27910 50089 27952
rect 64823 27992 64870 28034
rect 64994 27992 65038 28034
rect 65162 27992 65209 28034
rect 64823 27952 64832 27992
rect 64994 27952 64996 27992
rect 65036 27952 65038 27992
rect 65200 27952 65209 27992
rect 64823 27910 64870 27952
rect 64994 27910 65038 27952
rect 65162 27910 65209 27952
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 18223 27236 18270 27278
rect 18394 27236 18438 27278
rect 18562 27236 18609 27278
rect 18223 27196 18232 27236
rect 18394 27196 18396 27236
rect 18436 27196 18438 27236
rect 18600 27196 18609 27236
rect 18223 27154 18270 27196
rect 18394 27154 18438 27196
rect 18562 27154 18609 27196
rect 33343 27236 33390 27278
rect 33514 27236 33558 27278
rect 33682 27236 33729 27278
rect 33343 27196 33352 27236
rect 33514 27196 33516 27236
rect 33556 27196 33558 27236
rect 33720 27196 33729 27236
rect 33343 27154 33390 27196
rect 33514 27154 33558 27196
rect 33682 27154 33729 27196
rect 48463 27236 48510 27278
rect 48634 27236 48678 27278
rect 48802 27236 48849 27278
rect 48463 27196 48472 27236
rect 48634 27196 48636 27236
rect 48676 27196 48678 27236
rect 48840 27196 48849 27236
rect 48463 27154 48510 27196
rect 48634 27154 48678 27196
rect 48802 27154 48849 27196
rect 63583 27236 63630 27278
rect 63754 27236 63798 27278
rect 63922 27236 63969 27278
rect 63583 27196 63592 27236
rect 63754 27196 63756 27236
rect 63796 27196 63798 27236
rect 63960 27196 63969 27236
rect 63583 27154 63630 27196
rect 63754 27154 63798 27196
rect 63922 27154 63969 27196
rect 78703 27236 78750 27278
rect 78874 27236 78918 27278
rect 79042 27236 79089 27278
rect 78703 27196 78712 27236
rect 78874 27196 78876 27236
rect 78916 27196 78918 27236
rect 79080 27196 79089 27236
rect 78703 27154 78750 27196
rect 78874 27154 78918 27196
rect 79042 27154 79089 27196
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 19463 26480 19510 26522
rect 19634 26480 19678 26522
rect 19802 26480 19849 26522
rect 19463 26440 19472 26480
rect 19634 26440 19636 26480
rect 19676 26440 19678 26480
rect 19840 26440 19849 26480
rect 19463 26398 19510 26440
rect 19634 26398 19678 26440
rect 19802 26398 19849 26440
rect 34583 26480 34630 26522
rect 34754 26480 34798 26522
rect 34922 26480 34969 26522
rect 34583 26440 34592 26480
rect 34754 26440 34756 26480
rect 34796 26440 34798 26480
rect 34960 26440 34969 26480
rect 34583 26398 34630 26440
rect 34754 26398 34798 26440
rect 34922 26398 34969 26440
rect 49703 26480 49750 26522
rect 49874 26480 49918 26522
rect 50042 26480 50089 26522
rect 49703 26440 49712 26480
rect 49874 26440 49876 26480
rect 49916 26440 49918 26480
rect 50080 26440 50089 26480
rect 49703 26398 49750 26440
rect 49874 26398 49918 26440
rect 50042 26398 50089 26440
rect 64823 26480 64870 26522
rect 64994 26480 65038 26522
rect 65162 26480 65209 26522
rect 64823 26440 64832 26480
rect 64994 26440 64996 26480
rect 65036 26440 65038 26480
rect 65200 26440 65209 26480
rect 64823 26398 64870 26440
rect 64994 26398 65038 26440
rect 65162 26398 65209 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 18223 25724 18270 25766
rect 18394 25724 18438 25766
rect 18562 25724 18609 25766
rect 18223 25684 18232 25724
rect 18394 25684 18396 25724
rect 18436 25684 18438 25724
rect 18600 25684 18609 25724
rect 18223 25642 18270 25684
rect 18394 25642 18438 25684
rect 18562 25642 18609 25684
rect 33343 25724 33390 25766
rect 33514 25724 33558 25766
rect 33682 25724 33729 25766
rect 33343 25684 33352 25724
rect 33514 25684 33516 25724
rect 33556 25684 33558 25724
rect 33720 25684 33729 25724
rect 33343 25642 33390 25684
rect 33514 25642 33558 25684
rect 33682 25642 33729 25684
rect 48463 25724 48510 25766
rect 48634 25724 48678 25766
rect 48802 25724 48849 25766
rect 48463 25684 48472 25724
rect 48634 25684 48636 25724
rect 48676 25684 48678 25724
rect 48840 25684 48849 25724
rect 48463 25642 48510 25684
rect 48634 25642 48678 25684
rect 48802 25642 48849 25684
rect 63583 25724 63630 25766
rect 63754 25724 63798 25766
rect 63922 25724 63969 25766
rect 63583 25684 63592 25724
rect 63754 25684 63756 25724
rect 63796 25684 63798 25724
rect 63960 25684 63969 25724
rect 63583 25642 63630 25684
rect 63754 25642 63798 25684
rect 63922 25642 63969 25684
rect 78703 25724 78750 25766
rect 78874 25724 78918 25766
rect 79042 25724 79089 25766
rect 78703 25684 78712 25724
rect 78874 25684 78876 25724
rect 78916 25684 78918 25724
rect 79080 25684 79089 25724
rect 78703 25642 78750 25684
rect 78874 25642 78918 25684
rect 79042 25642 79089 25684
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 19463 24968 19510 25010
rect 19634 24968 19678 25010
rect 19802 24968 19849 25010
rect 19463 24928 19472 24968
rect 19634 24928 19636 24968
rect 19676 24928 19678 24968
rect 19840 24928 19849 24968
rect 19463 24886 19510 24928
rect 19634 24886 19678 24928
rect 19802 24886 19849 24928
rect 34583 24968 34630 25010
rect 34754 24968 34798 25010
rect 34922 24968 34969 25010
rect 34583 24928 34592 24968
rect 34754 24928 34756 24968
rect 34796 24928 34798 24968
rect 34960 24928 34969 24968
rect 34583 24886 34630 24928
rect 34754 24886 34798 24928
rect 34922 24886 34969 24928
rect 49703 24968 49750 25010
rect 49874 24968 49918 25010
rect 50042 24968 50089 25010
rect 49703 24928 49712 24968
rect 49874 24928 49876 24968
rect 49916 24928 49918 24968
rect 50080 24928 50089 24968
rect 49703 24886 49750 24928
rect 49874 24886 49918 24928
rect 50042 24886 50089 24928
rect 64823 24968 64870 25010
rect 64994 24968 65038 25010
rect 65162 24968 65209 25010
rect 64823 24928 64832 24968
rect 64994 24928 64996 24968
rect 65036 24928 65038 24968
rect 65200 24928 65209 24968
rect 64823 24886 64870 24928
rect 64994 24886 65038 24928
rect 65162 24886 65209 24928
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 18223 24212 18270 24254
rect 18394 24212 18438 24254
rect 18562 24212 18609 24254
rect 18223 24172 18232 24212
rect 18394 24172 18396 24212
rect 18436 24172 18438 24212
rect 18600 24172 18609 24212
rect 18223 24130 18270 24172
rect 18394 24130 18438 24172
rect 18562 24130 18609 24172
rect 33343 24212 33390 24254
rect 33514 24212 33558 24254
rect 33682 24212 33729 24254
rect 33343 24172 33352 24212
rect 33514 24172 33516 24212
rect 33556 24172 33558 24212
rect 33720 24172 33729 24212
rect 33343 24130 33390 24172
rect 33514 24130 33558 24172
rect 33682 24130 33729 24172
rect 48463 24212 48510 24254
rect 48634 24212 48678 24254
rect 48802 24212 48849 24254
rect 48463 24172 48472 24212
rect 48634 24172 48636 24212
rect 48676 24172 48678 24212
rect 48840 24172 48849 24212
rect 48463 24130 48510 24172
rect 48634 24130 48678 24172
rect 48802 24130 48849 24172
rect 40483 23836 40492 23876
rect 40532 23836 44044 23876
rect 44084 23836 61036 23876
rect 61076 23836 61085 23876
rect 52579 23752 52588 23792
rect 52628 23752 79084 23792
rect 79124 23752 79133 23792
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 19463 23456 19510 23498
rect 19634 23456 19678 23498
rect 19802 23456 19849 23498
rect 19463 23416 19472 23456
rect 19634 23416 19636 23456
rect 19676 23416 19678 23456
rect 19840 23416 19849 23456
rect 19463 23374 19510 23416
rect 19634 23374 19678 23416
rect 19802 23374 19849 23416
rect 34583 23456 34630 23498
rect 34754 23456 34798 23498
rect 34922 23456 34969 23498
rect 34583 23416 34592 23456
rect 34754 23416 34756 23456
rect 34796 23416 34798 23456
rect 34960 23416 34969 23456
rect 34583 23374 34630 23416
rect 34754 23374 34798 23416
rect 34922 23374 34969 23416
rect 49703 23456 49750 23498
rect 49874 23456 49918 23498
rect 50042 23456 50089 23498
rect 49703 23416 49712 23456
rect 49874 23416 49876 23456
rect 49916 23416 49918 23456
rect 50080 23416 50089 23456
rect 51811 23416 51820 23456
rect 51860 23416 56812 23456
rect 56852 23416 56861 23456
rect 49703 23374 49750 23416
rect 49874 23374 49918 23416
rect 50042 23374 50089 23416
rect 51043 23332 51052 23372
rect 51092 23332 56044 23372
rect 56084 23332 56093 23372
rect 51331 23248 51340 23288
rect 51380 23248 56428 23288
rect 56468 23248 56477 23288
rect 50851 23164 50860 23204
rect 50900 23164 55276 23204
rect 55316 23164 55325 23204
rect 52291 23080 52300 23120
rect 52340 23080 54796 23120
rect 54836 23080 54845 23120
rect 51907 22828 51916 22868
rect 51956 22828 58444 22868
rect 58484 22828 58828 22868
rect 58868 22828 58877 22868
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 18223 22700 18270 22742
rect 18394 22700 18438 22742
rect 18562 22700 18609 22742
rect 18223 22660 18232 22700
rect 18394 22660 18396 22700
rect 18436 22660 18438 22700
rect 18600 22660 18609 22700
rect 18223 22618 18270 22660
rect 18394 22618 18438 22660
rect 18562 22618 18609 22660
rect 33343 22700 33390 22742
rect 33514 22700 33558 22742
rect 33682 22700 33729 22742
rect 33343 22660 33352 22700
rect 33514 22660 33516 22700
rect 33556 22660 33558 22700
rect 33720 22660 33729 22700
rect 33343 22618 33390 22660
rect 33514 22618 33558 22660
rect 33682 22618 33729 22660
rect 48463 22700 48510 22742
rect 48634 22700 48678 22742
rect 48802 22700 48849 22742
rect 48463 22660 48472 22700
rect 48634 22660 48636 22700
rect 48676 22660 48678 22700
rect 48840 22660 48849 22700
rect 48463 22618 48510 22660
rect 48634 22618 48678 22660
rect 48802 22618 48849 22660
rect 64796 22541 65236 22652
rect 64796 22417 64870 22541
rect 64994 22417 65038 22541
rect 65162 22417 65236 22541
rect 64796 22373 65236 22417
rect 64796 22249 64870 22373
rect 64994 22249 65038 22373
rect 65162 22249 65236 22373
rect 64796 22205 65236 22249
rect 64796 22081 64870 22205
rect 64994 22081 65038 22205
rect 65162 22081 65236 22205
rect 64796 22037 65236 22081
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 19463 21944 19510 21986
rect 19634 21944 19678 21986
rect 19802 21944 19849 21986
rect 19463 21904 19472 21944
rect 19634 21904 19636 21944
rect 19676 21904 19678 21944
rect 19840 21904 19849 21944
rect 19463 21862 19510 21904
rect 19634 21862 19678 21904
rect 19802 21862 19849 21904
rect 34583 21944 34630 21986
rect 34754 21944 34798 21986
rect 34922 21944 34969 21986
rect 34583 21904 34592 21944
rect 34754 21904 34756 21944
rect 34796 21904 34798 21944
rect 34960 21904 34969 21944
rect 34583 21862 34630 21904
rect 34754 21862 34798 21904
rect 34922 21862 34969 21904
rect 49703 21944 49750 21986
rect 49874 21944 49918 21986
rect 50042 21944 50089 21986
rect 49703 21904 49712 21944
rect 49874 21904 49876 21944
rect 49916 21904 49918 21944
rect 50080 21904 50089 21944
rect 49703 21862 49750 21904
rect 49874 21862 49918 21904
rect 50042 21862 50089 21904
rect 64796 21913 64870 22037
rect 64994 21913 65038 22037
rect 65162 21913 65236 22037
rect 64796 21869 65236 21913
rect 64796 21745 64870 21869
rect 64994 21745 65038 21869
rect 65162 21745 65236 21869
rect 64796 21701 65236 21745
rect 64796 21577 64870 21701
rect 64994 21577 65038 21701
rect 65162 21577 65236 21701
rect 64796 21533 65236 21577
rect 64796 21409 64870 21533
rect 64994 21409 65038 21533
rect 65162 21409 65236 21533
rect 64796 21365 65236 21409
rect 64796 21241 64870 21365
rect 64994 21241 65038 21365
rect 65162 21241 65236 21365
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 18223 21188 18270 21230
rect 18394 21188 18438 21230
rect 18562 21188 18609 21230
rect 18223 21148 18232 21188
rect 18394 21148 18396 21188
rect 18436 21148 18438 21188
rect 18600 21148 18609 21188
rect 18223 21106 18270 21148
rect 18394 21106 18438 21148
rect 18562 21106 18609 21148
rect 33343 21188 33390 21230
rect 33514 21188 33558 21230
rect 33682 21188 33729 21230
rect 33343 21148 33352 21188
rect 33514 21148 33516 21188
rect 33556 21148 33558 21188
rect 33720 21148 33729 21188
rect 33343 21106 33390 21148
rect 33514 21106 33558 21148
rect 33682 21106 33729 21148
rect 48463 21188 48510 21230
rect 48634 21188 48678 21230
rect 48802 21188 48849 21230
rect 48463 21148 48472 21188
rect 48634 21148 48636 21188
rect 48676 21148 48678 21188
rect 48840 21148 48849 21188
rect 48463 21106 48510 21148
rect 48634 21106 48678 21148
rect 48802 21106 48849 21148
rect 64796 21197 65236 21241
rect 64796 21073 64870 21197
rect 64994 21073 65038 21197
rect 65162 21073 65236 21197
rect 64796 21029 65236 21073
rect 64796 20905 64870 21029
rect 64994 20905 65038 21029
rect 65162 20905 65236 21029
rect 64796 20861 65236 20905
rect 64796 20737 64870 20861
rect 64994 20737 65038 20861
rect 65162 20737 65236 20861
rect 64796 20693 65236 20737
rect 64796 20569 64870 20693
rect 64994 20569 65038 20693
rect 65162 20569 65236 20693
rect 64796 20525 65236 20569
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 19463 20432 19510 20474
rect 19634 20432 19678 20474
rect 19802 20432 19849 20474
rect 19463 20392 19472 20432
rect 19634 20392 19636 20432
rect 19676 20392 19678 20432
rect 19840 20392 19849 20432
rect 19463 20350 19510 20392
rect 19634 20350 19678 20392
rect 19802 20350 19849 20392
rect 34583 20432 34630 20474
rect 34754 20432 34798 20474
rect 34922 20432 34969 20474
rect 34583 20392 34592 20432
rect 34754 20392 34756 20432
rect 34796 20392 34798 20432
rect 34960 20392 34969 20432
rect 34583 20350 34630 20392
rect 34754 20350 34798 20392
rect 34922 20350 34969 20392
rect 49703 20432 49750 20474
rect 49874 20432 49918 20474
rect 50042 20432 50089 20474
rect 49703 20392 49712 20432
rect 49874 20392 49876 20432
rect 49916 20392 49918 20432
rect 50080 20392 50089 20432
rect 49703 20350 49750 20392
rect 49874 20350 49918 20392
rect 50042 20350 50089 20392
rect 64796 20401 64870 20525
rect 64994 20401 65038 20525
rect 65162 20401 65236 20525
rect 64796 20290 65236 20401
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 18223 19676 18270 19718
rect 18394 19676 18438 19718
rect 18562 19676 18609 19718
rect 18223 19636 18232 19676
rect 18394 19636 18396 19676
rect 18436 19636 18438 19676
rect 18600 19636 18609 19676
rect 18223 19594 18270 19636
rect 18394 19594 18438 19636
rect 18562 19594 18609 19636
rect 33343 19676 33390 19718
rect 33514 19676 33558 19718
rect 33682 19676 33729 19718
rect 33343 19636 33352 19676
rect 33514 19636 33516 19676
rect 33556 19636 33558 19676
rect 33720 19636 33729 19676
rect 33343 19594 33390 19636
rect 33514 19594 33558 19636
rect 33682 19594 33729 19636
rect 48463 19676 48510 19718
rect 48634 19676 48678 19718
rect 48802 19676 48849 19718
rect 48463 19636 48472 19676
rect 48634 19636 48636 19676
rect 48676 19636 48678 19676
rect 48840 19636 48849 19676
rect 48463 19594 48510 19636
rect 48634 19594 48678 19636
rect 48802 19594 48849 19636
rect 63556 19665 63996 19776
rect 63556 19541 63630 19665
rect 63754 19541 63798 19665
rect 63922 19541 63996 19665
rect 63556 19497 63996 19541
rect 63556 19373 63630 19497
rect 63754 19373 63798 19497
rect 63922 19373 63996 19497
rect 63556 19329 63996 19373
rect 63556 19205 63630 19329
rect 63754 19205 63798 19329
rect 63922 19205 63996 19329
rect 63556 19161 63996 19205
rect 63556 19037 63630 19161
rect 63754 19037 63798 19161
rect 63922 19037 63996 19161
rect 63556 18993 63996 19037
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 19463 18920 19510 18962
rect 19634 18920 19678 18962
rect 19802 18920 19849 18962
rect 19463 18880 19472 18920
rect 19634 18880 19636 18920
rect 19676 18880 19678 18920
rect 19840 18880 19849 18920
rect 19463 18838 19510 18880
rect 19634 18838 19678 18880
rect 19802 18838 19849 18880
rect 34583 18920 34630 18962
rect 34754 18920 34798 18962
rect 34922 18920 34969 18962
rect 34583 18880 34592 18920
rect 34754 18880 34756 18920
rect 34796 18880 34798 18920
rect 34960 18880 34969 18920
rect 34583 18838 34630 18880
rect 34754 18838 34798 18880
rect 34922 18838 34969 18880
rect 49703 18920 49750 18962
rect 49874 18920 49918 18962
rect 50042 18920 50089 18962
rect 49703 18880 49712 18920
rect 49874 18880 49876 18920
rect 49916 18880 49918 18920
rect 50080 18880 50089 18920
rect 49703 18838 49750 18880
rect 49874 18838 49918 18880
rect 50042 18838 50089 18880
rect 63556 18869 63630 18993
rect 63754 18869 63798 18993
rect 63922 18869 63996 18993
rect 63556 18825 63996 18869
rect 63556 18701 63630 18825
rect 63754 18701 63798 18825
rect 63922 18701 63996 18825
rect 63556 18657 63996 18701
rect 22339 18544 22348 18584
rect 22388 18544 27724 18584
rect 27764 18544 27773 18584
rect 63556 18533 63630 18657
rect 63754 18533 63798 18657
rect 63922 18533 63996 18657
rect 23683 18460 23692 18500
rect 23732 18460 28492 18500
rect 28532 18460 28541 18500
rect 63556 18489 63996 18533
rect 63556 18365 63630 18489
rect 63754 18365 63798 18489
rect 63922 18365 63996 18489
rect 63556 18321 63996 18365
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 18223 18164 18270 18206
rect 18394 18164 18438 18206
rect 18562 18164 18609 18206
rect 18223 18124 18232 18164
rect 18394 18124 18396 18164
rect 18436 18124 18438 18164
rect 18600 18124 18609 18164
rect 18223 18082 18270 18124
rect 18394 18082 18438 18124
rect 18562 18082 18609 18124
rect 33343 18164 33390 18206
rect 33514 18164 33558 18206
rect 33682 18164 33729 18206
rect 33343 18124 33352 18164
rect 33514 18124 33516 18164
rect 33556 18124 33558 18164
rect 33720 18124 33729 18164
rect 33343 18082 33390 18124
rect 33514 18082 33558 18124
rect 33682 18082 33729 18124
rect 48463 18164 48510 18206
rect 48634 18164 48678 18206
rect 48802 18164 48849 18206
rect 48463 18124 48472 18164
rect 48634 18124 48636 18164
rect 48676 18124 48678 18164
rect 48840 18124 48849 18164
rect 48463 18082 48510 18124
rect 48634 18082 48678 18124
rect 48802 18082 48849 18124
rect 63556 18197 63630 18321
rect 63754 18197 63798 18321
rect 63922 18197 63996 18321
rect 63556 18153 63996 18197
rect 63556 18029 63630 18153
rect 63754 18029 63798 18153
rect 63922 18029 63996 18153
rect 63556 17985 63996 18029
rect 63556 17861 63630 17985
rect 63754 17861 63798 17985
rect 63922 17861 63996 17985
rect 63556 17817 63996 17861
rect 63556 17693 63630 17817
rect 63754 17693 63798 17817
rect 63922 17693 63996 17817
rect 29539 17620 29548 17660
rect 29588 17620 49612 17660
rect 49652 17620 49661 17660
rect 63556 17649 63996 17693
rect 25795 17536 25804 17576
rect 25844 17536 51916 17576
rect 51956 17536 51965 17576
rect 63556 17525 63630 17649
rect 63754 17525 63798 17649
rect 63922 17525 63996 17649
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 19463 17408 19510 17450
rect 19634 17408 19678 17450
rect 19802 17408 19849 17450
rect 19463 17368 19472 17408
rect 19634 17368 19636 17408
rect 19676 17368 19678 17408
rect 19840 17368 19849 17408
rect 19463 17326 19510 17368
rect 19634 17326 19678 17368
rect 19802 17326 19849 17368
rect 34583 17408 34630 17450
rect 34754 17408 34798 17450
rect 34922 17408 34969 17450
rect 34583 17368 34592 17408
rect 34754 17368 34756 17408
rect 34796 17368 34798 17408
rect 34960 17368 34969 17408
rect 34583 17326 34630 17368
rect 34754 17326 34798 17368
rect 34922 17326 34969 17368
rect 49703 17408 49750 17450
rect 49874 17408 49918 17450
rect 50042 17408 50089 17450
rect 63556 17414 63996 17525
rect 78676 19665 79116 19776
rect 78676 19541 78750 19665
rect 78874 19541 78918 19665
rect 79042 19541 79116 19665
rect 78676 19497 79116 19541
rect 78676 19373 78750 19497
rect 78874 19373 78918 19497
rect 79042 19373 79116 19497
rect 78676 19329 79116 19373
rect 78676 19205 78750 19329
rect 78874 19205 78918 19329
rect 79042 19205 79116 19329
rect 78676 19161 79116 19205
rect 78676 19037 78750 19161
rect 78874 19037 78918 19161
rect 79042 19037 79116 19161
rect 78676 18993 79116 19037
rect 78676 18869 78750 18993
rect 78874 18869 78918 18993
rect 79042 18869 79116 18993
rect 78676 18825 79116 18869
rect 78676 18701 78750 18825
rect 78874 18701 78918 18825
rect 79042 18701 79116 18825
rect 78676 18657 79116 18701
rect 78676 18533 78750 18657
rect 78874 18533 78918 18657
rect 79042 18533 79116 18657
rect 78676 18489 79116 18533
rect 78676 18365 78750 18489
rect 78874 18365 78918 18489
rect 79042 18365 79116 18489
rect 78676 18321 79116 18365
rect 78676 18197 78750 18321
rect 78874 18197 78918 18321
rect 79042 18197 79116 18321
rect 78676 18153 79116 18197
rect 78676 18029 78750 18153
rect 78874 18029 78918 18153
rect 79042 18029 79116 18153
rect 78676 17985 79116 18029
rect 78676 17861 78750 17985
rect 78874 17861 78918 17985
rect 79042 17861 79116 17985
rect 78676 17817 79116 17861
rect 78676 17693 78750 17817
rect 78874 17693 78918 17817
rect 79042 17693 79116 17817
rect 78676 17649 79116 17693
rect 78676 17525 78750 17649
rect 78874 17525 78918 17649
rect 79042 17525 79116 17649
rect 78676 17414 79116 17525
rect 49703 17368 49712 17408
rect 49874 17368 49876 17408
rect 49916 17368 49918 17408
rect 50080 17368 50089 17408
rect 49703 17326 49750 17368
rect 49874 17326 49918 17368
rect 50042 17326 50089 17368
rect 51907 17200 51916 17240
rect 51956 17200 53932 17240
rect 53972 17200 53981 17240
rect 41155 17116 41164 17156
rect 41204 17116 48940 17156
rect 48980 17116 48989 17156
rect 50563 17116 50572 17156
rect 50612 17116 55084 17156
rect 55124 17116 55133 17156
rect 52579 17032 52588 17072
rect 52628 17032 78892 17072
rect 78932 17032 78941 17072
rect 32707 16948 32716 16988
rect 32756 16948 49036 16988
rect 49076 16948 49085 16988
rect 50371 16948 50380 16988
rect 50420 16948 55468 16988
rect 55508 16948 55517 16988
rect 39715 16864 39724 16904
rect 39764 16864 57868 16904
rect 57908 16864 57917 16904
rect 36643 16780 36652 16820
rect 36692 16780 53300 16820
rect 53260 16736 53300 16780
rect 53260 16696 58252 16736
rect 58292 16696 58301 16736
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 18223 16652 18270 16694
rect 18394 16652 18438 16694
rect 18562 16652 18609 16694
rect 18223 16612 18232 16652
rect 18394 16612 18396 16652
rect 18436 16612 18438 16652
rect 18600 16612 18609 16652
rect 18223 16570 18270 16612
rect 18394 16570 18438 16612
rect 18562 16570 18609 16612
rect 33343 16652 33390 16694
rect 33514 16652 33558 16694
rect 33682 16652 33729 16694
rect 33343 16612 33352 16652
rect 33514 16612 33516 16652
rect 33556 16612 33558 16652
rect 33720 16612 33729 16652
rect 33343 16570 33390 16612
rect 33514 16570 33558 16612
rect 33682 16570 33729 16612
rect 48463 16652 48510 16694
rect 48634 16652 48678 16694
rect 48802 16652 48849 16694
rect 48463 16612 48472 16652
rect 48634 16612 48636 16652
rect 48676 16612 48678 16652
rect 48840 16612 48849 16652
rect 49027 16612 49036 16652
rect 49076 16612 54700 16652
rect 54740 16612 54749 16652
rect 48463 16570 48510 16612
rect 48634 16570 48678 16612
rect 48802 16570 48849 16612
rect 48931 16528 48940 16568
rect 48980 16528 55660 16568
rect 55700 16528 55709 16568
rect 50467 16276 50476 16316
rect 50516 16276 61708 16316
rect 61748 16276 61757 16316
rect 51715 16192 51724 16232
rect 51764 16192 64972 16232
rect 65012 16192 65021 16232
rect 52675 16024 52684 16064
rect 52724 16024 53260 16064
rect 53300 16024 53309 16064
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 19463 15896 19510 15938
rect 19634 15896 19678 15938
rect 19802 15896 19849 15938
rect 19463 15856 19472 15896
rect 19634 15856 19636 15896
rect 19676 15856 19678 15896
rect 19840 15856 19849 15896
rect 19463 15814 19510 15856
rect 19634 15814 19678 15856
rect 19802 15814 19849 15856
rect 34583 15896 34630 15938
rect 34754 15896 34798 15938
rect 34922 15896 34969 15938
rect 34583 15856 34592 15896
rect 34754 15856 34756 15896
rect 34796 15856 34798 15896
rect 34960 15856 34969 15896
rect 34583 15814 34630 15856
rect 34754 15814 34798 15856
rect 34922 15814 34969 15856
rect 49703 15896 49750 15938
rect 49874 15896 49918 15938
rect 50042 15896 50089 15938
rect 49703 15856 49712 15896
rect 49874 15856 49876 15896
rect 49916 15856 49918 15896
rect 50080 15856 50089 15896
rect 49703 15814 49750 15856
rect 49874 15814 49918 15856
rect 50042 15814 50089 15856
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 18223 15140 18270 15182
rect 18394 15140 18438 15182
rect 18562 15140 18609 15182
rect 18223 15100 18232 15140
rect 18394 15100 18396 15140
rect 18436 15100 18438 15140
rect 18600 15100 18609 15140
rect 18223 15058 18270 15100
rect 18394 15058 18438 15100
rect 18562 15058 18609 15100
rect 33343 15140 33390 15182
rect 33514 15140 33558 15182
rect 33682 15140 33729 15182
rect 33343 15100 33352 15140
rect 33514 15100 33516 15140
rect 33556 15100 33558 15140
rect 33720 15100 33729 15140
rect 33343 15058 33390 15100
rect 33514 15058 33558 15100
rect 33682 15058 33729 15100
rect 48463 15140 48510 15182
rect 48634 15140 48678 15182
rect 48802 15140 48849 15182
rect 48463 15100 48472 15140
rect 48634 15100 48636 15140
rect 48676 15100 48678 15140
rect 48840 15100 48849 15140
rect 48463 15058 48510 15100
rect 48634 15058 48678 15100
rect 48802 15058 48849 15100
rect 63583 15140 63630 15182
rect 63754 15140 63798 15182
rect 63922 15140 63969 15182
rect 63583 15100 63592 15140
rect 63754 15100 63756 15140
rect 63796 15100 63798 15140
rect 63960 15100 63969 15140
rect 63583 15058 63630 15100
rect 63754 15058 63798 15100
rect 63922 15058 63969 15100
rect 78703 15140 78750 15182
rect 78874 15140 78918 15182
rect 79042 15140 79089 15182
rect 78703 15100 78712 15140
rect 78874 15100 78876 15140
rect 78916 15100 78918 15140
rect 79080 15100 79089 15140
rect 78703 15058 78750 15100
rect 78874 15058 78918 15100
rect 79042 15058 79089 15100
rect 51523 14848 51532 14888
rect 51572 14848 63340 14888
rect 63380 14848 63389 14888
rect 51235 14764 51244 14804
rect 51284 14764 58924 14804
rect 58964 14764 67180 14804
rect 67220 14764 67229 14804
rect 52483 14680 52492 14720
rect 52532 14680 54700 14720
rect 54740 14680 54749 14720
rect 32611 14512 32620 14552
rect 32660 14512 58540 14552
rect 58580 14512 58589 14552
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 19463 14384 19510 14426
rect 19634 14384 19678 14426
rect 19802 14384 19849 14426
rect 19463 14344 19472 14384
rect 19634 14344 19636 14384
rect 19676 14344 19678 14384
rect 19840 14344 19849 14384
rect 19463 14302 19510 14344
rect 19634 14302 19678 14344
rect 19802 14302 19849 14344
rect 34583 14384 34630 14426
rect 34754 14384 34798 14426
rect 34922 14384 34969 14426
rect 34583 14344 34592 14384
rect 34754 14344 34756 14384
rect 34796 14344 34798 14384
rect 34960 14344 34969 14384
rect 34583 14302 34630 14344
rect 34754 14302 34798 14344
rect 34922 14302 34969 14344
rect 49703 14384 49750 14426
rect 49874 14384 49918 14426
rect 50042 14384 50089 14426
rect 49703 14344 49712 14384
rect 49874 14344 49876 14384
rect 49916 14344 49918 14384
rect 50080 14344 50089 14384
rect 49703 14302 49750 14344
rect 49874 14302 49918 14344
rect 50042 14302 50089 14344
rect 64823 14384 64870 14426
rect 64994 14384 65038 14426
rect 65162 14384 65209 14426
rect 64823 14344 64832 14384
rect 64994 14344 64996 14384
rect 65036 14344 65038 14384
rect 65200 14344 65209 14384
rect 64823 14302 64870 14344
rect 64994 14302 65038 14344
rect 65162 14302 65209 14344
rect 57763 13924 57772 13964
rect 57812 13924 69196 13964
rect 69236 13924 69245 13964
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 18223 13628 18270 13670
rect 18394 13628 18438 13670
rect 18562 13628 18609 13670
rect 18223 13588 18232 13628
rect 18394 13588 18396 13628
rect 18436 13588 18438 13628
rect 18600 13588 18609 13628
rect 18223 13546 18270 13588
rect 18394 13546 18438 13588
rect 18562 13546 18609 13588
rect 33343 13628 33390 13670
rect 33514 13628 33558 13670
rect 33682 13628 33729 13670
rect 33343 13588 33352 13628
rect 33514 13588 33516 13628
rect 33556 13588 33558 13628
rect 33720 13588 33729 13628
rect 33343 13546 33390 13588
rect 33514 13546 33558 13588
rect 33682 13546 33729 13588
rect 48463 13628 48510 13670
rect 48634 13628 48678 13670
rect 48802 13628 48849 13670
rect 48463 13588 48472 13628
rect 48634 13588 48636 13628
rect 48676 13588 48678 13628
rect 48840 13588 48849 13628
rect 48463 13546 48510 13588
rect 48634 13546 48678 13588
rect 48802 13546 48849 13588
rect 63583 13628 63630 13670
rect 63754 13628 63798 13670
rect 63922 13628 63969 13670
rect 63583 13588 63592 13628
rect 63754 13588 63756 13628
rect 63796 13588 63798 13628
rect 63960 13588 63969 13628
rect 63583 13546 63630 13588
rect 63754 13546 63798 13588
rect 63922 13546 63969 13588
rect 78703 13628 78750 13670
rect 78874 13628 78918 13670
rect 79042 13628 79089 13670
rect 78703 13588 78712 13628
rect 78874 13588 78876 13628
rect 78916 13588 78918 13628
rect 79080 13588 79089 13628
rect 78703 13546 78750 13588
rect 78874 13546 78918 13588
rect 79042 13546 79089 13588
rect 51427 13000 51436 13040
rect 51476 13000 57772 13040
rect 57812 13000 57821 13040
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 19463 12872 19510 12914
rect 19634 12872 19678 12914
rect 19802 12872 19849 12914
rect 19463 12832 19472 12872
rect 19634 12832 19636 12872
rect 19676 12832 19678 12872
rect 19840 12832 19849 12872
rect 19463 12790 19510 12832
rect 19634 12790 19678 12832
rect 19802 12790 19849 12832
rect 34583 12872 34630 12914
rect 34754 12872 34798 12914
rect 34922 12872 34969 12914
rect 34583 12832 34592 12872
rect 34754 12832 34756 12872
rect 34796 12832 34798 12872
rect 34960 12832 34969 12872
rect 34583 12790 34630 12832
rect 34754 12790 34798 12832
rect 34922 12790 34969 12832
rect 49703 12872 49750 12914
rect 49874 12872 49918 12914
rect 50042 12872 50089 12914
rect 49703 12832 49712 12872
rect 49874 12832 49876 12872
rect 49916 12832 49918 12872
rect 50080 12832 50089 12872
rect 49703 12790 49750 12832
rect 49874 12790 49918 12832
rect 50042 12790 50089 12832
rect 64823 12872 64870 12914
rect 64994 12872 65038 12914
rect 65162 12872 65209 12914
rect 64823 12832 64832 12872
rect 64994 12832 64996 12872
rect 65036 12832 65038 12872
rect 65200 12832 65209 12872
rect 64823 12790 64870 12832
rect 64994 12790 65038 12832
rect 65162 12790 65209 12832
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 18223 12116 18270 12158
rect 18394 12116 18438 12158
rect 18562 12116 18609 12158
rect 18223 12076 18232 12116
rect 18394 12076 18396 12116
rect 18436 12076 18438 12116
rect 18600 12076 18609 12116
rect 18223 12034 18270 12076
rect 18394 12034 18438 12076
rect 18562 12034 18609 12076
rect 33343 12116 33390 12158
rect 33514 12116 33558 12158
rect 33682 12116 33729 12158
rect 33343 12076 33352 12116
rect 33514 12076 33516 12116
rect 33556 12076 33558 12116
rect 33720 12076 33729 12116
rect 33343 12034 33390 12076
rect 33514 12034 33558 12076
rect 33682 12034 33729 12076
rect 48463 12116 48510 12158
rect 48634 12116 48678 12158
rect 48802 12116 48849 12158
rect 48463 12076 48472 12116
rect 48634 12076 48636 12116
rect 48676 12076 48678 12116
rect 48840 12076 48849 12116
rect 48463 12034 48510 12076
rect 48634 12034 48678 12076
rect 48802 12034 48849 12076
rect 63583 12116 63630 12158
rect 63754 12116 63798 12158
rect 63922 12116 63969 12158
rect 63583 12076 63592 12116
rect 63754 12076 63756 12116
rect 63796 12076 63798 12116
rect 63960 12076 63969 12116
rect 63583 12034 63630 12076
rect 63754 12034 63798 12076
rect 63922 12034 63969 12076
rect 78703 12116 78750 12158
rect 78874 12116 78918 12158
rect 79042 12116 79089 12158
rect 78703 12076 78712 12116
rect 78874 12076 78876 12116
rect 78916 12076 78918 12116
rect 79080 12076 79089 12116
rect 78703 12034 78750 12076
rect 78874 12034 78918 12076
rect 79042 12034 79089 12076
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 19463 11360 19510 11402
rect 19634 11360 19678 11402
rect 19802 11360 19849 11402
rect 19463 11320 19472 11360
rect 19634 11320 19636 11360
rect 19676 11320 19678 11360
rect 19840 11320 19849 11360
rect 19463 11278 19510 11320
rect 19634 11278 19678 11320
rect 19802 11278 19849 11320
rect 34583 11360 34630 11402
rect 34754 11360 34798 11402
rect 34922 11360 34969 11402
rect 34583 11320 34592 11360
rect 34754 11320 34756 11360
rect 34796 11320 34798 11360
rect 34960 11320 34969 11360
rect 34583 11278 34630 11320
rect 34754 11278 34798 11320
rect 34922 11278 34969 11320
rect 49703 11360 49750 11402
rect 49874 11360 49918 11402
rect 50042 11360 50089 11402
rect 49703 11320 49712 11360
rect 49874 11320 49876 11360
rect 49916 11320 49918 11360
rect 50080 11320 50089 11360
rect 49703 11278 49750 11320
rect 49874 11278 49918 11320
rect 50042 11278 50089 11320
rect 64823 11360 64870 11402
rect 64994 11360 65038 11402
rect 65162 11360 65209 11402
rect 64823 11320 64832 11360
rect 64994 11320 64996 11360
rect 65036 11320 65038 11360
rect 65200 11320 65209 11360
rect 64823 11278 64870 11320
rect 64994 11278 65038 11320
rect 65162 11278 65209 11320
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 18223 10604 18270 10646
rect 18394 10604 18438 10646
rect 18562 10604 18609 10646
rect 18223 10564 18232 10604
rect 18394 10564 18396 10604
rect 18436 10564 18438 10604
rect 18600 10564 18609 10604
rect 18223 10522 18270 10564
rect 18394 10522 18438 10564
rect 18562 10522 18609 10564
rect 33343 10604 33390 10646
rect 33514 10604 33558 10646
rect 33682 10604 33729 10646
rect 33343 10564 33352 10604
rect 33514 10564 33516 10604
rect 33556 10564 33558 10604
rect 33720 10564 33729 10604
rect 33343 10522 33390 10564
rect 33514 10522 33558 10564
rect 33682 10522 33729 10564
rect 48463 10604 48510 10646
rect 48634 10604 48678 10646
rect 48802 10604 48849 10646
rect 48463 10564 48472 10604
rect 48634 10564 48636 10604
rect 48676 10564 48678 10604
rect 48840 10564 48849 10604
rect 48463 10522 48510 10564
rect 48634 10522 48678 10564
rect 48802 10522 48849 10564
rect 63583 10604 63630 10646
rect 63754 10604 63798 10646
rect 63922 10604 63969 10646
rect 63583 10564 63592 10604
rect 63754 10564 63756 10604
rect 63796 10564 63798 10604
rect 63960 10564 63969 10604
rect 63583 10522 63630 10564
rect 63754 10522 63798 10564
rect 63922 10522 63969 10564
rect 78703 10604 78750 10646
rect 78874 10604 78918 10646
rect 79042 10604 79089 10646
rect 78703 10564 78712 10604
rect 78874 10564 78876 10604
rect 78916 10564 78918 10604
rect 79080 10564 79089 10604
rect 78703 10522 78750 10564
rect 78874 10522 78918 10564
rect 79042 10522 79089 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 19463 9848 19510 9890
rect 19634 9848 19678 9890
rect 19802 9848 19849 9890
rect 19463 9808 19472 9848
rect 19634 9808 19636 9848
rect 19676 9808 19678 9848
rect 19840 9808 19849 9848
rect 19463 9766 19510 9808
rect 19634 9766 19678 9808
rect 19802 9766 19849 9808
rect 34583 9848 34630 9890
rect 34754 9848 34798 9890
rect 34922 9848 34969 9890
rect 34583 9808 34592 9848
rect 34754 9808 34756 9848
rect 34796 9808 34798 9848
rect 34960 9808 34969 9848
rect 34583 9766 34630 9808
rect 34754 9766 34798 9808
rect 34922 9766 34969 9808
rect 49703 9848 49750 9890
rect 49874 9848 49918 9890
rect 50042 9848 50089 9890
rect 49703 9808 49712 9848
rect 49874 9808 49876 9848
rect 49916 9808 49918 9848
rect 50080 9808 50089 9848
rect 49703 9766 49750 9808
rect 49874 9766 49918 9808
rect 50042 9766 50089 9808
rect 64823 9848 64870 9890
rect 64994 9848 65038 9890
rect 65162 9848 65209 9890
rect 64823 9808 64832 9848
rect 64994 9808 64996 9848
rect 65036 9808 65038 9848
rect 65200 9808 65209 9848
rect 64823 9766 64870 9808
rect 64994 9766 65038 9808
rect 65162 9766 65209 9808
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 18223 9092 18270 9134
rect 18394 9092 18438 9134
rect 18562 9092 18609 9134
rect 18223 9052 18232 9092
rect 18394 9052 18396 9092
rect 18436 9052 18438 9092
rect 18600 9052 18609 9092
rect 18223 9010 18270 9052
rect 18394 9010 18438 9052
rect 18562 9010 18609 9052
rect 33343 9092 33390 9134
rect 33514 9092 33558 9134
rect 33682 9092 33729 9134
rect 33343 9052 33352 9092
rect 33514 9052 33516 9092
rect 33556 9052 33558 9092
rect 33720 9052 33729 9092
rect 33343 9010 33390 9052
rect 33514 9010 33558 9052
rect 33682 9010 33729 9052
rect 48463 9092 48510 9134
rect 48634 9092 48678 9134
rect 48802 9092 48849 9134
rect 48463 9052 48472 9092
rect 48634 9052 48636 9092
rect 48676 9052 48678 9092
rect 48840 9052 48849 9092
rect 48463 9010 48510 9052
rect 48634 9010 48678 9052
rect 48802 9010 48849 9052
rect 63583 9092 63630 9134
rect 63754 9092 63798 9134
rect 63922 9092 63969 9134
rect 63583 9052 63592 9092
rect 63754 9052 63756 9092
rect 63796 9052 63798 9092
rect 63960 9052 63969 9092
rect 63583 9010 63630 9052
rect 63754 9010 63798 9052
rect 63922 9010 63969 9052
rect 78703 9092 78750 9134
rect 78874 9092 78918 9134
rect 79042 9092 79089 9134
rect 78703 9052 78712 9092
rect 78874 9052 78876 9092
rect 78916 9052 78918 9092
rect 79080 9052 79089 9092
rect 78703 9010 78750 9052
rect 78874 9010 78918 9052
rect 79042 9010 79089 9052
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 19463 8336 19510 8378
rect 19634 8336 19678 8378
rect 19802 8336 19849 8378
rect 19463 8296 19472 8336
rect 19634 8296 19636 8336
rect 19676 8296 19678 8336
rect 19840 8296 19849 8336
rect 19463 8254 19510 8296
rect 19634 8254 19678 8296
rect 19802 8254 19849 8296
rect 34583 8336 34630 8378
rect 34754 8336 34798 8378
rect 34922 8336 34969 8378
rect 34583 8296 34592 8336
rect 34754 8296 34756 8336
rect 34796 8296 34798 8336
rect 34960 8296 34969 8336
rect 34583 8254 34630 8296
rect 34754 8254 34798 8296
rect 34922 8254 34969 8296
rect 49703 8336 49750 8378
rect 49874 8336 49918 8378
rect 50042 8336 50089 8378
rect 49703 8296 49712 8336
rect 49874 8296 49876 8336
rect 49916 8296 49918 8336
rect 50080 8296 50089 8336
rect 49703 8254 49750 8296
rect 49874 8254 49918 8296
rect 50042 8254 50089 8296
rect 64823 8336 64870 8378
rect 64994 8336 65038 8378
rect 65162 8336 65209 8378
rect 64823 8296 64832 8336
rect 64994 8296 64996 8336
rect 65036 8296 65038 8336
rect 65200 8296 65209 8336
rect 64823 8254 64870 8296
rect 64994 8254 65038 8296
rect 65162 8254 65209 8296
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 18223 7580 18270 7622
rect 18394 7580 18438 7622
rect 18562 7580 18609 7622
rect 18223 7540 18232 7580
rect 18394 7540 18396 7580
rect 18436 7540 18438 7580
rect 18600 7540 18609 7580
rect 18223 7498 18270 7540
rect 18394 7498 18438 7540
rect 18562 7498 18609 7540
rect 33343 7580 33390 7622
rect 33514 7580 33558 7622
rect 33682 7580 33729 7622
rect 33343 7540 33352 7580
rect 33514 7540 33516 7580
rect 33556 7540 33558 7580
rect 33720 7540 33729 7580
rect 33343 7498 33390 7540
rect 33514 7498 33558 7540
rect 33682 7498 33729 7540
rect 48463 7580 48510 7622
rect 48634 7580 48678 7622
rect 48802 7580 48849 7622
rect 48463 7540 48472 7580
rect 48634 7540 48636 7580
rect 48676 7540 48678 7580
rect 48840 7540 48849 7580
rect 48463 7498 48510 7540
rect 48634 7498 48678 7540
rect 48802 7498 48849 7540
rect 63583 7580 63630 7622
rect 63754 7580 63798 7622
rect 63922 7580 63969 7622
rect 63583 7540 63592 7580
rect 63754 7540 63756 7580
rect 63796 7540 63798 7580
rect 63960 7540 63969 7580
rect 63583 7498 63630 7540
rect 63754 7498 63798 7540
rect 63922 7498 63969 7540
rect 78703 7580 78750 7622
rect 78874 7580 78918 7622
rect 79042 7580 79089 7622
rect 78703 7540 78712 7580
rect 78874 7540 78876 7580
rect 78916 7540 78918 7580
rect 79080 7540 79089 7580
rect 78703 7498 78750 7540
rect 78874 7498 78918 7540
rect 79042 7498 79089 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 19463 6824 19510 6866
rect 19634 6824 19678 6866
rect 19802 6824 19849 6866
rect 19463 6784 19472 6824
rect 19634 6784 19636 6824
rect 19676 6784 19678 6824
rect 19840 6784 19849 6824
rect 19463 6742 19510 6784
rect 19634 6742 19678 6784
rect 19802 6742 19849 6784
rect 34583 6824 34630 6866
rect 34754 6824 34798 6866
rect 34922 6824 34969 6866
rect 34583 6784 34592 6824
rect 34754 6784 34756 6824
rect 34796 6784 34798 6824
rect 34960 6784 34969 6824
rect 34583 6742 34630 6784
rect 34754 6742 34798 6784
rect 34922 6742 34969 6784
rect 49703 6824 49750 6866
rect 49874 6824 49918 6866
rect 50042 6824 50089 6866
rect 49703 6784 49712 6824
rect 49874 6784 49876 6824
rect 49916 6784 49918 6824
rect 50080 6784 50089 6824
rect 49703 6742 49750 6784
rect 49874 6742 49918 6784
rect 50042 6742 50089 6784
rect 64823 6824 64870 6866
rect 64994 6824 65038 6866
rect 65162 6824 65209 6866
rect 64823 6784 64832 6824
rect 64994 6784 64996 6824
rect 65036 6784 65038 6824
rect 65200 6784 65209 6824
rect 64823 6742 64870 6784
rect 64994 6742 65038 6784
rect 65162 6742 65209 6784
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 18223 6068 18270 6110
rect 18394 6068 18438 6110
rect 18562 6068 18609 6110
rect 18223 6028 18232 6068
rect 18394 6028 18396 6068
rect 18436 6028 18438 6068
rect 18600 6028 18609 6068
rect 18223 5986 18270 6028
rect 18394 5986 18438 6028
rect 18562 5986 18609 6028
rect 33343 6068 33390 6110
rect 33514 6068 33558 6110
rect 33682 6068 33729 6110
rect 33343 6028 33352 6068
rect 33514 6028 33516 6068
rect 33556 6028 33558 6068
rect 33720 6028 33729 6068
rect 33343 5986 33390 6028
rect 33514 5986 33558 6028
rect 33682 5986 33729 6028
rect 48463 6068 48510 6110
rect 48634 6068 48678 6110
rect 48802 6068 48849 6110
rect 48463 6028 48472 6068
rect 48634 6028 48636 6068
rect 48676 6028 48678 6068
rect 48840 6028 48849 6068
rect 48463 5986 48510 6028
rect 48634 5986 48678 6028
rect 48802 5986 48849 6028
rect 63583 6068 63630 6110
rect 63754 6068 63798 6110
rect 63922 6068 63969 6110
rect 63583 6028 63592 6068
rect 63754 6028 63756 6068
rect 63796 6028 63798 6068
rect 63960 6028 63969 6068
rect 63583 5986 63630 6028
rect 63754 5986 63798 6028
rect 63922 5986 63969 6028
rect 78703 6068 78750 6110
rect 78874 6068 78918 6110
rect 79042 6068 79089 6110
rect 78703 6028 78712 6068
rect 78874 6028 78876 6068
rect 78916 6028 78918 6068
rect 79080 6028 79089 6068
rect 78703 5986 78750 6028
rect 78874 5986 78918 6028
rect 79042 5986 79089 6028
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 19463 5312 19510 5354
rect 19634 5312 19678 5354
rect 19802 5312 19849 5354
rect 19463 5272 19472 5312
rect 19634 5272 19636 5312
rect 19676 5272 19678 5312
rect 19840 5272 19849 5312
rect 19463 5230 19510 5272
rect 19634 5230 19678 5272
rect 19802 5230 19849 5272
rect 34583 5312 34630 5354
rect 34754 5312 34798 5354
rect 34922 5312 34969 5354
rect 34583 5272 34592 5312
rect 34754 5272 34756 5312
rect 34796 5272 34798 5312
rect 34960 5272 34969 5312
rect 34583 5230 34630 5272
rect 34754 5230 34798 5272
rect 34922 5230 34969 5272
rect 49703 5312 49750 5354
rect 49874 5312 49918 5354
rect 50042 5312 50089 5354
rect 49703 5272 49712 5312
rect 49874 5272 49876 5312
rect 49916 5272 49918 5312
rect 50080 5272 50089 5312
rect 49703 5230 49750 5272
rect 49874 5230 49918 5272
rect 50042 5230 50089 5272
rect 64823 5312 64870 5354
rect 64994 5312 65038 5354
rect 65162 5312 65209 5354
rect 64823 5272 64832 5312
rect 64994 5272 64996 5312
rect 65036 5272 65038 5312
rect 65200 5272 65209 5312
rect 64823 5230 64870 5272
rect 64994 5230 65038 5272
rect 65162 5230 65209 5272
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 18223 4556 18270 4598
rect 18394 4556 18438 4598
rect 18562 4556 18609 4598
rect 18223 4516 18232 4556
rect 18394 4516 18396 4556
rect 18436 4516 18438 4556
rect 18600 4516 18609 4556
rect 18223 4474 18270 4516
rect 18394 4474 18438 4516
rect 18562 4474 18609 4516
rect 33343 4556 33390 4598
rect 33514 4556 33558 4598
rect 33682 4556 33729 4598
rect 33343 4516 33352 4556
rect 33514 4516 33516 4556
rect 33556 4516 33558 4556
rect 33720 4516 33729 4556
rect 33343 4474 33390 4516
rect 33514 4474 33558 4516
rect 33682 4474 33729 4516
rect 48463 4556 48510 4598
rect 48634 4556 48678 4598
rect 48802 4556 48849 4598
rect 48463 4516 48472 4556
rect 48634 4516 48636 4556
rect 48676 4516 48678 4556
rect 48840 4516 48849 4556
rect 48463 4474 48510 4516
rect 48634 4474 48678 4516
rect 48802 4474 48849 4516
rect 63583 4556 63630 4598
rect 63754 4556 63798 4598
rect 63922 4556 63969 4598
rect 63583 4516 63592 4556
rect 63754 4516 63756 4556
rect 63796 4516 63798 4556
rect 63960 4516 63969 4556
rect 63583 4474 63630 4516
rect 63754 4474 63798 4516
rect 63922 4474 63969 4516
rect 78703 4556 78750 4598
rect 78874 4556 78918 4598
rect 79042 4556 79089 4598
rect 78703 4516 78712 4556
rect 78874 4516 78876 4556
rect 78916 4516 78918 4556
rect 79080 4516 79089 4556
rect 78703 4474 78750 4516
rect 78874 4474 78918 4516
rect 79042 4474 79089 4516
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 19463 3800 19510 3842
rect 19634 3800 19678 3842
rect 19802 3800 19849 3842
rect 19463 3760 19472 3800
rect 19634 3760 19636 3800
rect 19676 3760 19678 3800
rect 19840 3760 19849 3800
rect 19463 3718 19510 3760
rect 19634 3718 19678 3760
rect 19802 3718 19849 3760
rect 34583 3800 34630 3842
rect 34754 3800 34798 3842
rect 34922 3800 34969 3842
rect 34583 3760 34592 3800
rect 34754 3760 34756 3800
rect 34796 3760 34798 3800
rect 34960 3760 34969 3800
rect 34583 3718 34630 3760
rect 34754 3718 34798 3760
rect 34922 3718 34969 3760
rect 49703 3800 49750 3842
rect 49874 3800 49918 3842
rect 50042 3800 50089 3842
rect 49703 3760 49712 3800
rect 49874 3760 49876 3800
rect 49916 3760 49918 3800
rect 50080 3760 50089 3800
rect 49703 3718 49750 3760
rect 49874 3718 49918 3760
rect 50042 3718 50089 3760
rect 64823 3800 64870 3842
rect 64994 3800 65038 3842
rect 65162 3800 65209 3842
rect 64823 3760 64832 3800
rect 64994 3760 64996 3800
rect 65036 3760 65038 3800
rect 65200 3760 65209 3800
rect 64823 3718 64870 3760
rect 64994 3718 65038 3760
rect 65162 3718 65209 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 18223 3044 18270 3086
rect 18394 3044 18438 3086
rect 18562 3044 18609 3086
rect 18223 3004 18232 3044
rect 18394 3004 18396 3044
rect 18436 3004 18438 3044
rect 18600 3004 18609 3044
rect 18223 2962 18270 3004
rect 18394 2962 18438 3004
rect 18562 2962 18609 3004
rect 33343 3044 33390 3086
rect 33514 3044 33558 3086
rect 33682 3044 33729 3086
rect 33343 3004 33352 3044
rect 33514 3004 33516 3044
rect 33556 3004 33558 3044
rect 33720 3004 33729 3044
rect 33343 2962 33390 3004
rect 33514 2962 33558 3004
rect 33682 2962 33729 3004
rect 48463 3044 48510 3086
rect 48634 3044 48678 3086
rect 48802 3044 48849 3086
rect 48463 3004 48472 3044
rect 48634 3004 48636 3044
rect 48676 3004 48678 3044
rect 48840 3004 48849 3044
rect 48463 2962 48510 3004
rect 48634 2962 48678 3004
rect 48802 2962 48849 3004
rect 63583 3044 63630 3086
rect 63754 3044 63798 3086
rect 63922 3044 63969 3086
rect 63583 3004 63592 3044
rect 63754 3004 63756 3044
rect 63796 3004 63798 3044
rect 63960 3004 63969 3044
rect 63583 2962 63630 3004
rect 63754 2962 63798 3004
rect 63922 2962 63969 3004
rect 78703 3044 78750 3086
rect 78874 3044 78918 3086
rect 79042 3044 79089 3086
rect 78703 3004 78712 3044
rect 78874 3004 78876 3044
rect 78916 3004 78918 3044
rect 79080 3004 79089 3044
rect 78703 2962 78750 3004
rect 78874 2962 78918 3004
rect 79042 2962 79089 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 19463 2288 19510 2330
rect 19634 2288 19678 2330
rect 19802 2288 19849 2330
rect 19463 2248 19472 2288
rect 19634 2248 19636 2288
rect 19676 2248 19678 2288
rect 19840 2248 19849 2288
rect 19463 2206 19510 2248
rect 19634 2206 19678 2248
rect 19802 2206 19849 2248
rect 34583 2288 34630 2330
rect 34754 2288 34798 2330
rect 34922 2288 34969 2330
rect 34583 2248 34592 2288
rect 34754 2248 34756 2288
rect 34796 2248 34798 2288
rect 34960 2248 34969 2288
rect 34583 2206 34630 2248
rect 34754 2206 34798 2248
rect 34922 2206 34969 2248
rect 49703 2288 49750 2330
rect 49874 2288 49918 2330
rect 50042 2288 50089 2330
rect 49703 2248 49712 2288
rect 49874 2248 49876 2288
rect 49916 2248 49918 2288
rect 50080 2248 50089 2288
rect 49703 2206 49750 2248
rect 49874 2206 49918 2248
rect 50042 2206 50089 2248
rect 64823 2288 64870 2330
rect 64994 2288 65038 2330
rect 65162 2288 65209 2330
rect 64823 2248 64832 2288
rect 64994 2248 64996 2288
rect 65036 2248 65038 2288
rect 65200 2248 65209 2288
rect 64823 2206 64870 2248
rect 64994 2206 65038 2248
rect 65162 2206 65209 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 18223 1532 18270 1574
rect 18394 1532 18438 1574
rect 18562 1532 18609 1574
rect 18223 1492 18232 1532
rect 18394 1492 18396 1532
rect 18436 1492 18438 1532
rect 18600 1492 18609 1532
rect 18223 1450 18270 1492
rect 18394 1450 18438 1492
rect 18562 1450 18609 1492
rect 33343 1532 33390 1574
rect 33514 1532 33558 1574
rect 33682 1532 33729 1574
rect 33343 1492 33352 1532
rect 33514 1492 33516 1532
rect 33556 1492 33558 1532
rect 33720 1492 33729 1532
rect 33343 1450 33390 1492
rect 33514 1450 33558 1492
rect 33682 1450 33729 1492
rect 48463 1532 48510 1574
rect 48634 1532 48678 1574
rect 48802 1532 48849 1574
rect 48463 1492 48472 1532
rect 48634 1492 48636 1532
rect 48676 1492 48678 1532
rect 48840 1492 48849 1532
rect 48463 1450 48510 1492
rect 48634 1450 48678 1492
rect 48802 1450 48849 1492
rect 63583 1532 63630 1574
rect 63754 1532 63798 1574
rect 63922 1532 63969 1574
rect 63583 1492 63592 1532
rect 63754 1492 63756 1532
rect 63796 1492 63798 1532
rect 63960 1492 63969 1532
rect 63583 1450 63630 1492
rect 63754 1450 63798 1492
rect 63922 1450 63969 1492
rect 78703 1532 78750 1574
rect 78874 1532 78918 1574
rect 79042 1532 79089 1574
rect 78703 1492 78712 1532
rect 78874 1492 78876 1532
rect 78916 1492 78918 1532
rect 79080 1492 79089 1532
rect 78703 1450 78750 1492
rect 78874 1450 78918 1492
rect 79042 1450 79089 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 19463 776 19510 818
rect 19634 776 19678 818
rect 19802 776 19849 818
rect 19463 736 19472 776
rect 19634 736 19636 776
rect 19676 736 19678 776
rect 19840 736 19849 776
rect 19463 694 19510 736
rect 19634 694 19678 736
rect 19802 694 19849 736
rect 34583 776 34630 818
rect 34754 776 34798 818
rect 34922 776 34969 818
rect 34583 736 34592 776
rect 34754 736 34756 776
rect 34796 736 34798 776
rect 34960 736 34969 776
rect 34583 694 34630 736
rect 34754 694 34798 736
rect 34922 694 34969 736
rect 49703 776 49750 818
rect 49874 776 49918 818
rect 50042 776 50089 818
rect 49703 736 49712 776
rect 49874 736 49876 776
rect 49916 736 49918 776
rect 50080 736 50089 776
rect 49703 694 49750 736
rect 49874 694 49918 736
rect 50042 694 50089 736
rect 64823 776 64870 818
rect 64994 776 65038 818
rect 65162 776 65209 818
rect 64823 736 64832 776
rect 64994 736 64996 776
rect 65036 736 65038 776
rect 65200 736 65209 776
rect 64823 694 64870 736
rect 64994 694 65038 736
rect 65162 694 65209 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 19510 38576 19634 38618
rect 19678 38576 19802 38618
rect 19510 38536 19512 38576
rect 19512 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19634 38576
rect 19678 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19800 38576
rect 19800 38536 19802 38576
rect 19510 38494 19634 38536
rect 19678 38494 19802 38536
rect 34630 38576 34754 38618
rect 34798 38576 34922 38618
rect 34630 38536 34632 38576
rect 34632 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34754 38576
rect 34798 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34920 38576
rect 34920 38536 34922 38576
rect 34630 38494 34754 38536
rect 34798 38494 34922 38536
rect 49750 38576 49874 38618
rect 49918 38576 50042 38618
rect 49750 38536 49752 38576
rect 49752 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49874 38576
rect 49918 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50040 38576
rect 50040 38536 50042 38576
rect 49750 38494 49874 38536
rect 49918 38494 50042 38536
rect 64870 38576 64994 38618
rect 65038 38576 65162 38618
rect 64870 38536 64872 38576
rect 64872 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64994 38576
rect 65038 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65160 38576
rect 65160 38536 65162 38576
rect 64870 38494 64994 38536
rect 65038 38494 65162 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 18270 37820 18394 37862
rect 18438 37820 18562 37862
rect 18270 37780 18272 37820
rect 18272 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18394 37820
rect 18438 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18560 37820
rect 18560 37780 18562 37820
rect 18270 37738 18394 37780
rect 18438 37738 18562 37780
rect 33390 37820 33514 37862
rect 33558 37820 33682 37862
rect 33390 37780 33392 37820
rect 33392 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33514 37820
rect 33558 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33680 37820
rect 33680 37780 33682 37820
rect 33390 37738 33514 37780
rect 33558 37738 33682 37780
rect 48510 37820 48634 37862
rect 48678 37820 48802 37862
rect 48510 37780 48512 37820
rect 48512 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48634 37820
rect 48678 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48800 37820
rect 48800 37780 48802 37820
rect 48510 37738 48634 37780
rect 48678 37738 48802 37780
rect 63630 37820 63754 37862
rect 63798 37820 63922 37862
rect 63630 37780 63632 37820
rect 63632 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63754 37820
rect 63798 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63920 37820
rect 63920 37780 63922 37820
rect 63630 37738 63754 37780
rect 63798 37738 63922 37780
rect 78750 37820 78874 37862
rect 78918 37820 79042 37862
rect 78750 37780 78752 37820
rect 78752 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78874 37820
rect 78918 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79040 37820
rect 79040 37780 79042 37820
rect 78750 37738 78874 37780
rect 78918 37738 79042 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 19510 37064 19634 37106
rect 19678 37064 19802 37106
rect 19510 37024 19512 37064
rect 19512 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19634 37064
rect 19678 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19800 37064
rect 19800 37024 19802 37064
rect 19510 36982 19634 37024
rect 19678 36982 19802 37024
rect 34630 37064 34754 37106
rect 34798 37064 34922 37106
rect 34630 37024 34632 37064
rect 34632 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34754 37064
rect 34798 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34920 37064
rect 34920 37024 34922 37064
rect 34630 36982 34754 37024
rect 34798 36982 34922 37024
rect 49750 37064 49874 37106
rect 49918 37064 50042 37106
rect 49750 37024 49752 37064
rect 49752 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49874 37064
rect 49918 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50040 37064
rect 50040 37024 50042 37064
rect 49750 36982 49874 37024
rect 49918 36982 50042 37024
rect 64870 37064 64994 37106
rect 65038 37064 65162 37106
rect 64870 37024 64872 37064
rect 64872 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64994 37064
rect 65038 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65160 37064
rect 65160 37024 65162 37064
rect 64870 36982 64994 37024
rect 65038 36982 65162 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 18270 36308 18394 36350
rect 18438 36308 18562 36350
rect 18270 36268 18272 36308
rect 18272 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18394 36308
rect 18438 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18560 36308
rect 18560 36268 18562 36308
rect 18270 36226 18394 36268
rect 18438 36226 18562 36268
rect 33390 36308 33514 36350
rect 33558 36308 33682 36350
rect 33390 36268 33392 36308
rect 33392 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33514 36308
rect 33558 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33680 36308
rect 33680 36268 33682 36308
rect 33390 36226 33514 36268
rect 33558 36226 33682 36268
rect 48510 36308 48634 36350
rect 48678 36308 48802 36350
rect 48510 36268 48512 36308
rect 48512 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48634 36308
rect 48678 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48800 36308
rect 48800 36268 48802 36308
rect 48510 36226 48634 36268
rect 48678 36226 48802 36268
rect 63630 36308 63754 36350
rect 63798 36308 63922 36350
rect 63630 36268 63632 36308
rect 63632 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63754 36308
rect 63798 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63920 36308
rect 63920 36268 63922 36308
rect 63630 36226 63754 36268
rect 63798 36226 63922 36268
rect 78750 36308 78874 36350
rect 78918 36308 79042 36350
rect 78750 36268 78752 36308
rect 78752 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78874 36308
rect 78918 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79040 36308
rect 79040 36268 79042 36308
rect 78750 36226 78874 36268
rect 78918 36226 79042 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 19510 35552 19634 35594
rect 19678 35552 19802 35594
rect 19510 35512 19512 35552
rect 19512 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19634 35552
rect 19678 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19800 35552
rect 19800 35512 19802 35552
rect 19510 35470 19634 35512
rect 19678 35470 19802 35512
rect 34630 35552 34754 35594
rect 34798 35552 34922 35594
rect 34630 35512 34632 35552
rect 34632 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34754 35552
rect 34798 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34920 35552
rect 34920 35512 34922 35552
rect 34630 35470 34754 35512
rect 34798 35470 34922 35512
rect 49750 35552 49874 35594
rect 49918 35552 50042 35594
rect 49750 35512 49752 35552
rect 49752 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49874 35552
rect 49918 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50040 35552
rect 50040 35512 50042 35552
rect 49750 35470 49874 35512
rect 49918 35470 50042 35512
rect 64870 35552 64994 35594
rect 65038 35552 65162 35594
rect 64870 35512 64872 35552
rect 64872 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64994 35552
rect 65038 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65160 35552
rect 65160 35512 65162 35552
rect 64870 35470 64994 35512
rect 65038 35470 65162 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 18270 34796 18394 34838
rect 18438 34796 18562 34838
rect 18270 34756 18272 34796
rect 18272 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18394 34796
rect 18438 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18560 34796
rect 18560 34756 18562 34796
rect 18270 34714 18394 34756
rect 18438 34714 18562 34756
rect 33390 34796 33514 34838
rect 33558 34796 33682 34838
rect 33390 34756 33392 34796
rect 33392 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33514 34796
rect 33558 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33680 34796
rect 33680 34756 33682 34796
rect 33390 34714 33514 34756
rect 33558 34714 33682 34756
rect 48510 34796 48634 34838
rect 48678 34796 48802 34838
rect 48510 34756 48512 34796
rect 48512 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48634 34796
rect 48678 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48800 34796
rect 48800 34756 48802 34796
rect 48510 34714 48634 34756
rect 48678 34714 48802 34756
rect 63630 34796 63754 34838
rect 63798 34796 63922 34838
rect 63630 34756 63632 34796
rect 63632 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63754 34796
rect 63798 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63920 34796
rect 63920 34756 63922 34796
rect 63630 34714 63754 34756
rect 63798 34714 63922 34756
rect 78750 34796 78874 34838
rect 78918 34796 79042 34838
rect 78750 34756 78752 34796
rect 78752 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78874 34796
rect 78918 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79040 34796
rect 79040 34756 79042 34796
rect 78750 34714 78874 34756
rect 78918 34714 79042 34756
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 19510 34040 19634 34082
rect 19678 34040 19802 34082
rect 19510 34000 19512 34040
rect 19512 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19634 34040
rect 19678 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19800 34040
rect 19800 34000 19802 34040
rect 19510 33958 19634 34000
rect 19678 33958 19802 34000
rect 34630 34040 34754 34082
rect 34798 34040 34922 34082
rect 34630 34000 34632 34040
rect 34632 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34754 34040
rect 34798 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34920 34040
rect 34920 34000 34922 34040
rect 34630 33958 34754 34000
rect 34798 33958 34922 34000
rect 49750 34040 49874 34082
rect 49918 34040 50042 34082
rect 49750 34000 49752 34040
rect 49752 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49874 34040
rect 49918 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50040 34040
rect 50040 34000 50042 34040
rect 49750 33958 49874 34000
rect 49918 33958 50042 34000
rect 64870 34040 64994 34082
rect 65038 34040 65162 34082
rect 64870 34000 64872 34040
rect 64872 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64994 34040
rect 65038 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65160 34040
rect 65160 34000 65162 34040
rect 64870 33958 64994 34000
rect 65038 33958 65162 34000
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 18270 33284 18394 33326
rect 18438 33284 18562 33326
rect 18270 33244 18272 33284
rect 18272 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18394 33284
rect 18438 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18560 33284
rect 18560 33244 18562 33284
rect 18270 33202 18394 33244
rect 18438 33202 18562 33244
rect 33390 33284 33514 33326
rect 33558 33284 33682 33326
rect 33390 33244 33392 33284
rect 33392 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33514 33284
rect 33558 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33680 33284
rect 33680 33244 33682 33284
rect 33390 33202 33514 33244
rect 33558 33202 33682 33244
rect 48510 33284 48634 33326
rect 48678 33284 48802 33326
rect 48510 33244 48512 33284
rect 48512 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48634 33284
rect 48678 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48800 33284
rect 48800 33244 48802 33284
rect 48510 33202 48634 33244
rect 48678 33202 48802 33244
rect 63630 33284 63754 33326
rect 63798 33284 63922 33326
rect 63630 33244 63632 33284
rect 63632 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63754 33284
rect 63798 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63920 33284
rect 63920 33244 63922 33284
rect 63630 33202 63754 33244
rect 63798 33202 63922 33244
rect 78750 33284 78874 33326
rect 78918 33284 79042 33326
rect 78750 33244 78752 33284
rect 78752 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78874 33284
rect 78918 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79040 33284
rect 79040 33244 79042 33284
rect 78750 33202 78874 33244
rect 78918 33202 79042 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 19510 32528 19634 32570
rect 19678 32528 19802 32570
rect 19510 32488 19512 32528
rect 19512 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19634 32528
rect 19678 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19800 32528
rect 19800 32488 19802 32528
rect 19510 32446 19634 32488
rect 19678 32446 19802 32488
rect 34630 32528 34754 32570
rect 34798 32528 34922 32570
rect 34630 32488 34632 32528
rect 34632 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34754 32528
rect 34798 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34920 32528
rect 34920 32488 34922 32528
rect 34630 32446 34754 32488
rect 34798 32446 34922 32488
rect 49750 32528 49874 32570
rect 49918 32528 50042 32570
rect 49750 32488 49752 32528
rect 49752 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49874 32528
rect 49918 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50040 32528
rect 50040 32488 50042 32528
rect 49750 32446 49874 32488
rect 49918 32446 50042 32488
rect 64870 32528 64994 32570
rect 65038 32528 65162 32570
rect 64870 32488 64872 32528
rect 64872 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64994 32528
rect 65038 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65160 32528
rect 65160 32488 65162 32528
rect 64870 32446 64994 32488
rect 65038 32446 65162 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 18270 31772 18394 31814
rect 18438 31772 18562 31814
rect 18270 31732 18272 31772
rect 18272 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18394 31772
rect 18438 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18560 31772
rect 18560 31732 18562 31772
rect 18270 31690 18394 31732
rect 18438 31690 18562 31732
rect 33390 31772 33514 31814
rect 33558 31772 33682 31814
rect 33390 31732 33392 31772
rect 33392 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33514 31772
rect 33558 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33680 31772
rect 33680 31732 33682 31772
rect 33390 31690 33514 31732
rect 33558 31690 33682 31732
rect 48510 31772 48634 31814
rect 48678 31772 48802 31814
rect 48510 31732 48512 31772
rect 48512 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48634 31772
rect 48678 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48800 31772
rect 48800 31732 48802 31772
rect 48510 31690 48634 31732
rect 48678 31690 48802 31732
rect 63630 31772 63754 31814
rect 63798 31772 63922 31814
rect 63630 31732 63632 31772
rect 63632 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63754 31772
rect 63798 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63920 31772
rect 63920 31732 63922 31772
rect 63630 31690 63754 31732
rect 63798 31690 63922 31732
rect 78750 31772 78874 31814
rect 78918 31772 79042 31814
rect 78750 31732 78752 31772
rect 78752 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78874 31772
rect 78918 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79040 31772
rect 79040 31732 79042 31772
rect 78750 31690 78874 31732
rect 78918 31690 79042 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 19510 31016 19634 31058
rect 19678 31016 19802 31058
rect 19510 30976 19512 31016
rect 19512 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19634 31016
rect 19678 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19800 31016
rect 19800 30976 19802 31016
rect 19510 30934 19634 30976
rect 19678 30934 19802 30976
rect 34630 31016 34754 31058
rect 34798 31016 34922 31058
rect 34630 30976 34632 31016
rect 34632 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34754 31016
rect 34798 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34920 31016
rect 34920 30976 34922 31016
rect 34630 30934 34754 30976
rect 34798 30934 34922 30976
rect 49750 31016 49874 31058
rect 49918 31016 50042 31058
rect 49750 30976 49752 31016
rect 49752 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49874 31016
rect 49918 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50040 31016
rect 50040 30976 50042 31016
rect 49750 30934 49874 30976
rect 49918 30934 50042 30976
rect 64870 31016 64994 31058
rect 65038 31016 65162 31058
rect 64870 30976 64872 31016
rect 64872 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64994 31016
rect 65038 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65160 31016
rect 65160 30976 65162 31016
rect 64870 30934 64994 30976
rect 65038 30934 65162 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 18270 30260 18394 30302
rect 18438 30260 18562 30302
rect 18270 30220 18272 30260
rect 18272 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18394 30260
rect 18438 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18560 30260
rect 18560 30220 18562 30260
rect 18270 30178 18394 30220
rect 18438 30178 18562 30220
rect 33390 30260 33514 30302
rect 33558 30260 33682 30302
rect 33390 30220 33392 30260
rect 33392 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33514 30260
rect 33558 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33680 30260
rect 33680 30220 33682 30260
rect 33390 30178 33514 30220
rect 33558 30178 33682 30220
rect 48510 30260 48634 30302
rect 48678 30260 48802 30302
rect 48510 30220 48512 30260
rect 48512 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48634 30260
rect 48678 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48800 30260
rect 48800 30220 48802 30260
rect 48510 30178 48634 30220
rect 48678 30178 48802 30220
rect 63630 30260 63754 30302
rect 63798 30260 63922 30302
rect 63630 30220 63632 30260
rect 63632 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63754 30260
rect 63798 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63920 30260
rect 63920 30220 63922 30260
rect 63630 30178 63754 30220
rect 63798 30178 63922 30220
rect 78750 30260 78874 30302
rect 78918 30260 79042 30302
rect 78750 30220 78752 30260
rect 78752 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78874 30260
rect 78918 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79040 30260
rect 79040 30220 79042 30260
rect 78750 30178 78874 30220
rect 78918 30178 79042 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 19510 29504 19634 29546
rect 19678 29504 19802 29546
rect 19510 29464 19512 29504
rect 19512 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19634 29504
rect 19678 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19800 29504
rect 19800 29464 19802 29504
rect 19510 29422 19634 29464
rect 19678 29422 19802 29464
rect 34630 29504 34754 29546
rect 34798 29504 34922 29546
rect 34630 29464 34632 29504
rect 34632 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34754 29504
rect 34798 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34920 29504
rect 34920 29464 34922 29504
rect 34630 29422 34754 29464
rect 34798 29422 34922 29464
rect 49750 29504 49874 29546
rect 49918 29504 50042 29546
rect 49750 29464 49752 29504
rect 49752 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49874 29504
rect 49918 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50040 29504
rect 50040 29464 50042 29504
rect 49750 29422 49874 29464
rect 49918 29422 50042 29464
rect 64870 29504 64994 29546
rect 65038 29504 65162 29546
rect 64870 29464 64872 29504
rect 64872 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64994 29504
rect 65038 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65160 29504
rect 65160 29464 65162 29504
rect 64870 29422 64994 29464
rect 65038 29422 65162 29464
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 18270 28748 18394 28790
rect 18438 28748 18562 28790
rect 18270 28708 18272 28748
rect 18272 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18394 28748
rect 18438 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18560 28748
rect 18560 28708 18562 28748
rect 18270 28666 18394 28708
rect 18438 28666 18562 28708
rect 33390 28748 33514 28790
rect 33558 28748 33682 28790
rect 33390 28708 33392 28748
rect 33392 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33514 28748
rect 33558 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33680 28748
rect 33680 28708 33682 28748
rect 33390 28666 33514 28708
rect 33558 28666 33682 28708
rect 48510 28748 48634 28790
rect 48678 28748 48802 28790
rect 48510 28708 48512 28748
rect 48512 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48634 28748
rect 48678 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48800 28748
rect 48800 28708 48802 28748
rect 48510 28666 48634 28708
rect 48678 28666 48802 28708
rect 63630 28748 63754 28790
rect 63798 28748 63922 28790
rect 63630 28708 63632 28748
rect 63632 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63754 28748
rect 63798 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63920 28748
rect 63920 28708 63922 28748
rect 63630 28666 63754 28708
rect 63798 28666 63922 28708
rect 78750 28748 78874 28790
rect 78918 28748 79042 28790
rect 78750 28708 78752 28748
rect 78752 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78874 28748
rect 78918 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79040 28748
rect 79040 28708 79042 28748
rect 78750 28666 78874 28708
rect 78918 28666 79042 28708
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 19510 27992 19634 28034
rect 19678 27992 19802 28034
rect 19510 27952 19512 27992
rect 19512 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19634 27992
rect 19678 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19800 27992
rect 19800 27952 19802 27992
rect 19510 27910 19634 27952
rect 19678 27910 19802 27952
rect 34630 27992 34754 28034
rect 34798 27992 34922 28034
rect 34630 27952 34632 27992
rect 34632 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34754 27992
rect 34798 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34920 27992
rect 34920 27952 34922 27992
rect 34630 27910 34754 27952
rect 34798 27910 34922 27952
rect 49750 27992 49874 28034
rect 49918 27992 50042 28034
rect 49750 27952 49752 27992
rect 49752 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49874 27992
rect 49918 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50040 27992
rect 50040 27952 50042 27992
rect 49750 27910 49874 27952
rect 49918 27910 50042 27952
rect 64870 27992 64994 28034
rect 65038 27992 65162 28034
rect 64870 27952 64872 27992
rect 64872 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64994 27992
rect 65038 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65160 27992
rect 65160 27952 65162 27992
rect 64870 27910 64994 27952
rect 65038 27910 65162 27952
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 18270 27236 18394 27278
rect 18438 27236 18562 27278
rect 18270 27196 18272 27236
rect 18272 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18394 27236
rect 18438 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18560 27236
rect 18560 27196 18562 27236
rect 18270 27154 18394 27196
rect 18438 27154 18562 27196
rect 33390 27236 33514 27278
rect 33558 27236 33682 27278
rect 33390 27196 33392 27236
rect 33392 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33514 27236
rect 33558 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33680 27236
rect 33680 27196 33682 27236
rect 33390 27154 33514 27196
rect 33558 27154 33682 27196
rect 48510 27236 48634 27278
rect 48678 27236 48802 27278
rect 48510 27196 48512 27236
rect 48512 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48634 27236
rect 48678 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48800 27236
rect 48800 27196 48802 27236
rect 48510 27154 48634 27196
rect 48678 27154 48802 27196
rect 63630 27236 63754 27278
rect 63798 27236 63922 27278
rect 63630 27196 63632 27236
rect 63632 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63754 27236
rect 63798 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63920 27236
rect 63920 27196 63922 27236
rect 63630 27154 63754 27196
rect 63798 27154 63922 27196
rect 78750 27236 78874 27278
rect 78918 27236 79042 27278
rect 78750 27196 78752 27236
rect 78752 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78874 27236
rect 78918 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79040 27236
rect 79040 27196 79042 27236
rect 78750 27154 78874 27196
rect 78918 27154 79042 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 19510 26480 19634 26522
rect 19678 26480 19802 26522
rect 19510 26440 19512 26480
rect 19512 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19634 26480
rect 19678 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19800 26480
rect 19800 26440 19802 26480
rect 19510 26398 19634 26440
rect 19678 26398 19802 26440
rect 34630 26480 34754 26522
rect 34798 26480 34922 26522
rect 34630 26440 34632 26480
rect 34632 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34754 26480
rect 34798 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34920 26480
rect 34920 26440 34922 26480
rect 34630 26398 34754 26440
rect 34798 26398 34922 26440
rect 49750 26480 49874 26522
rect 49918 26480 50042 26522
rect 49750 26440 49752 26480
rect 49752 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49874 26480
rect 49918 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50040 26480
rect 50040 26440 50042 26480
rect 49750 26398 49874 26440
rect 49918 26398 50042 26440
rect 64870 26480 64994 26522
rect 65038 26480 65162 26522
rect 64870 26440 64872 26480
rect 64872 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64994 26480
rect 65038 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65160 26480
rect 65160 26440 65162 26480
rect 64870 26398 64994 26440
rect 65038 26398 65162 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 18270 25724 18394 25766
rect 18438 25724 18562 25766
rect 18270 25684 18272 25724
rect 18272 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18394 25724
rect 18438 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18560 25724
rect 18560 25684 18562 25724
rect 18270 25642 18394 25684
rect 18438 25642 18562 25684
rect 33390 25724 33514 25766
rect 33558 25724 33682 25766
rect 33390 25684 33392 25724
rect 33392 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33514 25724
rect 33558 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33680 25724
rect 33680 25684 33682 25724
rect 33390 25642 33514 25684
rect 33558 25642 33682 25684
rect 48510 25724 48634 25766
rect 48678 25724 48802 25766
rect 48510 25684 48512 25724
rect 48512 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48634 25724
rect 48678 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48800 25724
rect 48800 25684 48802 25724
rect 48510 25642 48634 25684
rect 48678 25642 48802 25684
rect 63630 25724 63754 25766
rect 63798 25724 63922 25766
rect 63630 25684 63632 25724
rect 63632 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63754 25724
rect 63798 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63920 25724
rect 63920 25684 63922 25724
rect 63630 25642 63754 25684
rect 63798 25642 63922 25684
rect 78750 25724 78874 25766
rect 78918 25724 79042 25766
rect 78750 25684 78752 25724
rect 78752 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78874 25724
rect 78918 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79040 25724
rect 79040 25684 79042 25724
rect 78750 25642 78874 25684
rect 78918 25642 79042 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 19510 24968 19634 25010
rect 19678 24968 19802 25010
rect 19510 24928 19512 24968
rect 19512 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19634 24968
rect 19678 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19800 24968
rect 19800 24928 19802 24968
rect 19510 24886 19634 24928
rect 19678 24886 19802 24928
rect 34630 24968 34754 25010
rect 34798 24968 34922 25010
rect 34630 24928 34632 24968
rect 34632 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34754 24968
rect 34798 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34920 24968
rect 34920 24928 34922 24968
rect 34630 24886 34754 24928
rect 34798 24886 34922 24928
rect 49750 24968 49874 25010
rect 49918 24968 50042 25010
rect 49750 24928 49752 24968
rect 49752 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49874 24968
rect 49918 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50040 24968
rect 50040 24928 50042 24968
rect 49750 24886 49874 24928
rect 49918 24886 50042 24928
rect 64870 24968 64994 25010
rect 65038 24968 65162 25010
rect 64870 24928 64872 24968
rect 64872 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64994 24968
rect 65038 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65160 24968
rect 65160 24928 65162 24968
rect 64870 24886 64994 24928
rect 65038 24886 65162 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 18270 24212 18394 24254
rect 18438 24212 18562 24254
rect 18270 24172 18272 24212
rect 18272 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18394 24212
rect 18438 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18560 24212
rect 18560 24172 18562 24212
rect 18270 24130 18394 24172
rect 18438 24130 18562 24172
rect 33390 24212 33514 24254
rect 33558 24212 33682 24254
rect 33390 24172 33392 24212
rect 33392 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33514 24212
rect 33558 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33680 24212
rect 33680 24172 33682 24212
rect 33390 24130 33514 24172
rect 33558 24130 33682 24172
rect 48510 24212 48634 24254
rect 48678 24212 48802 24254
rect 48510 24172 48512 24212
rect 48512 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48634 24212
rect 48678 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48800 24212
rect 48800 24172 48802 24212
rect 48510 24130 48634 24172
rect 48678 24130 48802 24172
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 19510 23456 19634 23498
rect 19678 23456 19802 23498
rect 19510 23416 19512 23456
rect 19512 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19634 23456
rect 19678 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19800 23456
rect 19800 23416 19802 23456
rect 19510 23374 19634 23416
rect 19678 23374 19802 23416
rect 34630 23456 34754 23498
rect 34798 23456 34922 23498
rect 34630 23416 34632 23456
rect 34632 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34754 23456
rect 34798 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34920 23456
rect 34920 23416 34922 23456
rect 34630 23374 34754 23416
rect 34798 23374 34922 23416
rect 49750 23456 49874 23498
rect 49918 23456 50042 23498
rect 49750 23416 49752 23456
rect 49752 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49874 23456
rect 49918 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50040 23456
rect 50040 23416 50042 23456
rect 49750 23374 49874 23416
rect 49918 23374 50042 23416
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 18270 22700 18394 22742
rect 18438 22700 18562 22742
rect 18270 22660 18272 22700
rect 18272 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18394 22700
rect 18438 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18560 22700
rect 18560 22660 18562 22700
rect 18270 22618 18394 22660
rect 18438 22618 18562 22660
rect 33390 22700 33514 22742
rect 33558 22700 33682 22742
rect 33390 22660 33392 22700
rect 33392 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33514 22700
rect 33558 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33680 22700
rect 33680 22660 33682 22700
rect 33390 22618 33514 22660
rect 33558 22618 33682 22660
rect 48510 22700 48634 22742
rect 48678 22700 48802 22742
rect 48510 22660 48512 22700
rect 48512 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48634 22700
rect 48678 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48800 22700
rect 48800 22660 48802 22700
rect 48510 22618 48634 22660
rect 48678 22618 48802 22660
rect 64870 22417 64994 22541
rect 65038 22417 65162 22541
rect 64870 22249 64994 22373
rect 65038 22249 65162 22373
rect 64870 22081 64994 22205
rect 65038 22081 65162 22205
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 19510 21944 19634 21986
rect 19678 21944 19802 21986
rect 19510 21904 19512 21944
rect 19512 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19634 21944
rect 19678 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19800 21944
rect 19800 21904 19802 21944
rect 19510 21862 19634 21904
rect 19678 21862 19802 21904
rect 34630 21944 34754 21986
rect 34798 21944 34922 21986
rect 34630 21904 34632 21944
rect 34632 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34754 21944
rect 34798 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34920 21944
rect 34920 21904 34922 21944
rect 34630 21862 34754 21904
rect 34798 21862 34922 21904
rect 49750 21944 49874 21986
rect 49918 21944 50042 21986
rect 49750 21904 49752 21944
rect 49752 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49874 21944
rect 49918 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50040 21944
rect 50040 21904 50042 21944
rect 49750 21862 49874 21904
rect 49918 21862 50042 21904
rect 64870 21913 64994 22037
rect 65038 21913 65162 22037
rect 64870 21745 64994 21869
rect 65038 21745 65162 21869
rect 64870 21577 64994 21701
rect 65038 21577 65162 21701
rect 64870 21409 64994 21533
rect 65038 21409 65162 21533
rect 64870 21241 64994 21365
rect 65038 21241 65162 21365
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 18270 21188 18394 21230
rect 18438 21188 18562 21230
rect 18270 21148 18272 21188
rect 18272 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18394 21188
rect 18438 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18560 21188
rect 18560 21148 18562 21188
rect 18270 21106 18394 21148
rect 18438 21106 18562 21148
rect 33390 21188 33514 21230
rect 33558 21188 33682 21230
rect 33390 21148 33392 21188
rect 33392 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33514 21188
rect 33558 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33680 21188
rect 33680 21148 33682 21188
rect 33390 21106 33514 21148
rect 33558 21106 33682 21148
rect 48510 21188 48634 21230
rect 48678 21188 48802 21230
rect 48510 21148 48512 21188
rect 48512 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48634 21188
rect 48678 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48800 21188
rect 48800 21148 48802 21188
rect 48510 21106 48634 21148
rect 48678 21106 48802 21148
rect 64870 21073 64994 21197
rect 65038 21073 65162 21197
rect 64870 20905 64994 21029
rect 65038 20905 65162 21029
rect 64870 20737 64994 20861
rect 65038 20737 65162 20861
rect 64870 20569 64994 20693
rect 65038 20569 65162 20693
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 19510 20432 19634 20474
rect 19678 20432 19802 20474
rect 19510 20392 19512 20432
rect 19512 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19634 20432
rect 19678 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19800 20432
rect 19800 20392 19802 20432
rect 19510 20350 19634 20392
rect 19678 20350 19802 20392
rect 34630 20432 34754 20474
rect 34798 20432 34922 20474
rect 34630 20392 34632 20432
rect 34632 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34754 20432
rect 34798 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34920 20432
rect 34920 20392 34922 20432
rect 34630 20350 34754 20392
rect 34798 20350 34922 20392
rect 49750 20432 49874 20474
rect 49918 20432 50042 20474
rect 49750 20392 49752 20432
rect 49752 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49874 20432
rect 49918 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50040 20432
rect 50040 20392 50042 20432
rect 49750 20350 49874 20392
rect 49918 20350 50042 20392
rect 64870 20401 64994 20525
rect 65038 20401 65162 20525
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 18270 19676 18394 19718
rect 18438 19676 18562 19718
rect 18270 19636 18272 19676
rect 18272 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18394 19676
rect 18438 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18560 19676
rect 18560 19636 18562 19676
rect 18270 19594 18394 19636
rect 18438 19594 18562 19636
rect 33390 19676 33514 19718
rect 33558 19676 33682 19718
rect 33390 19636 33392 19676
rect 33392 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33514 19676
rect 33558 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33680 19676
rect 33680 19636 33682 19676
rect 33390 19594 33514 19636
rect 33558 19594 33682 19636
rect 48510 19676 48634 19718
rect 48678 19676 48802 19718
rect 48510 19636 48512 19676
rect 48512 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48634 19676
rect 48678 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48800 19676
rect 48800 19636 48802 19676
rect 48510 19594 48634 19636
rect 48678 19594 48802 19636
rect 63630 19541 63754 19665
rect 63798 19541 63922 19665
rect 63630 19373 63754 19497
rect 63798 19373 63922 19497
rect 63630 19205 63754 19329
rect 63798 19205 63922 19329
rect 63630 19037 63754 19161
rect 63798 19037 63922 19161
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 19510 18920 19634 18962
rect 19678 18920 19802 18962
rect 19510 18880 19512 18920
rect 19512 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19634 18920
rect 19678 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19800 18920
rect 19800 18880 19802 18920
rect 19510 18838 19634 18880
rect 19678 18838 19802 18880
rect 34630 18920 34754 18962
rect 34798 18920 34922 18962
rect 34630 18880 34632 18920
rect 34632 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34754 18920
rect 34798 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34920 18920
rect 34920 18880 34922 18920
rect 34630 18838 34754 18880
rect 34798 18838 34922 18880
rect 49750 18920 49874 18962
rect 49918 18920 50042 18962
rect 49750 18880 49752 18920
rect 49752 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49874 18920
rect 49918 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50040 18920
rect 50040 18880 50042 18920
rect 49750 18838 49874 18880
rect 49918 18838 50042 18880
rect 63630 18869 63754 18993
rect 63798 18869 63922 18993
rect 63630 18701 63754 18825
rect 63798 18701 63922 18825
rect 63630 18533 63754 18657
rect 63798 18533 63922 18657
rect 63630 18365 63754 18489
rect 63798 18365 63922 18489
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 18270 18164 18394 18206
rect 18438 18164 18562 18206
rect 18270 18124 18272 18164
rect 18272 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18394 18164
rect 18438 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18560 18164
rect 18560 18124 18562 18164
rect 18270 18082 18394 18124
rect 18438 18082 18562 18124
rect 33390 18164 33514 18206
rect 33558 18164 33682 18206
rect 33390 18124 33392 18164
rect 33392 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33514 18164
rect 33558 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33680 18164
rect 33680 18124 33682 18164
rect 33390 18082 33514 18124
rect 33558 18082 33682 18124
rect 48510 18164 48634 18206
rect 48678 18164 48802 18206
rect 48510 18124 48512 18164
rect 48512 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48634 18164
rect 48678 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48800 18164
rect 48800 18124 48802 18164
rect 48510 18082 48634 18124
rect 48678 18082 48802 18124
rect 63630 18197 63754 18321
rect 63798 18197 63922 18321
rect 63630 18029 63754 18153
rect 63798 18029 63922 18153
rect 63630 17861 63754 17985
rect 63798 17861 63922 17985
rect 63630 17693 63754 17817
rect 63798 17693 63922 17817
rect 63630 17525 63754 17649
rect 63798 17525 63922 17649
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 19510 17408 19634 17450
rect 19678 17408 19802 17450
rect 19510 17368 19512 17408
rect 19512 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19634 17408
rect 19678 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19800 17408
rect 19800 17368 19802 17408
rect 19510 17326 19634 17368
rect 19678 17326 19802 17368
rect 34630 17408 34754 17450
rect 34798 17408 34922 17450
rect 34630 17368 34632 17408
rect 34632 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34754 17408
rect 34798 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34920 17408
rect 34920 17368 34922 17408
rect 34630 17326 34754 17368
rect 34798 17326 34922 17368
rect 49750 17408 49874 17450
rect 49918 17408 50042 17450
rect 78750 19541 78874 19665
rect 78918 19541 79042 19665
rect 78750 19373 78874 19497
rect 78918 19373 79042 19497
rect 78750 19205 78874 19329
rect 78918 19205 79042 19329
rect 78750 19037 78874 19161
rect 78918 19037 79042 19161
rect 78750 18869 78874 18993
rect 78918 18869 79042 18993
rect 78750 18701 78874 18825
rect 78918 18701 79042 18825
rect 78750 18533 78874 18657
rect 78918 18533 79042 18657
rect 78750 18365 78874 18489
rect 78918 18365 79042 18489
rect 78750 18197 78874 18321
rect 78918 18197 79042 18321
rect 78750 18029 78874 18153
rect 78918 18029 79042 18153
rect 78750 17861 78874 17985
rect 78918 17861 79042 17985
rect 78750 17693 78874 17817
rect 78918 17693 79042 17817
rect 78750 17525 78874 17649
rect 78918 17525 79042 17649
rect 49750 17368 49752 17408
rect 49752 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49874 17408
rect 49918 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50040 17408
rect 50040 17368 50042 17408
rect 49750 17326 49874 17368
rect 49918 17326 50042 17368
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 18270 16652 18394 16694
rect 18438 16652 18562 16694
rect 18270 16612 18272 16652
rect 18272 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18394 16652
rect 18438 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18560 16652
rect 18560 16612 18562 16652
rect 18270 16570 18394 16612
rect 18438 16570 18562 16612
rect 33390 16652 33514 16694
rect 33558 16652 33682 16694
rect 33390 16612 33392 16652
rect 33392 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33514 16652
rect 33558 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33680 16652
rect 33680 16612 33682 16652
rect 33390 16570 33514 16612
rect 33558 16570 33682 16612
rect 48510 16652 48634 16694
rect 48678 16652 48802 16694
rect 48510 16612 48512 16652
rect 48512 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48634 16652
rect 48678 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48800 16652
rect 48800 16612 48802 16652
rect 48510 16570 48634 16612
rect 48678 16570 48802 16612
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 19510 15896 19634 15938
rect 19678 15896 19802 15938
rect 19510 15856 19512 15896
rect 19512 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19634 15896
rect 19678 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19800 15896
rect 19800 15856 19802 15896
rect 19510 15814 19634 15856
rect 19678 15814 19802 15856
rect 34630 15896 34754 15938
rect 34798 15896 34922 15938
rect 34630 15856 34632 15896
rect 34632 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34754 15896
rect 34798 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34920 15896
rect 34920 15856 34922 15896
rect 34630 15814 34754 15856
rect 34798 15814 34922 15856
rect 49750 15896 49874 15938
rect 49918 15896 50042 15938
rect 49750 15856 49752 15896
rect 49752 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49874 15896
rect 49918 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50040 15896
rect 50040 15856 50042 15896
rect 49750 15814 49874 15856
rect 49918 15814 50042 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 18270 15140 18394 15182
rect 18438 15140 18562 15182
rect 18270 15100 18272 15140
rect 18272 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18394 15140
rect 18438 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18560 15140
rect 18560 15100 18562 15140
rect 18270 15058 18394 15100
rect 18438 15058 18562 15100
rect 33390 15140 33514 15182
rect 33558 15140 33682 15182
rect 33390 15100 33392 15140
rect 33392 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33514 15140
rect 33558 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33680 15140
rect 33680 15100 33682 15140
rect 33390 15058 33514 15100
rect 33558 15058 33682 15100
rect 48510 15140 48634 15182
rect 48678 15140 48802 15182
rect 48510 15100 48512 15140
rect 48512 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48634 15140
rect 48678 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48800 15140
rect 48800 15100 48802 15140
rect 48510 15058 48634 15100
rect 48678 15058 48802 15100
rect 63630 15140 63754 15182
rect 63798 15140 63922 15182
rect 63630 15100 63632 15140
rect 63632 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63754 15140
rect 63798 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63920 15140
rect 63920 15100 63922 15140
rect 63630 15058 63754 15100
rect 63798 15058 63922 15100
rect 78750 15140 78874 15182
rect 78918 15140 79042 15182
rect 78750 15100 78752 15140
rect 78752 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78874 15140
rect 78918 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79040 15140
rect 79040 15100 79042 15140
rect 78750 15058 78874 15100
rect 78918 15058 79042 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 19510 14384 19634 14426
rect 19678 14384 19802 14426
rect 19510 14344 19512 14384
rect 19512 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19634 14384
rect 19678 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19800 14384
rect 19800 14344 19802 14384
rect 19510 14302 19634 14344
rect 19678 14302 19802 14344
rect 34630 14384 34754 14426
rect 34798 14384 34922 14426
rect 34630 14344 34632 14384
rect 34632 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34754 14384
rect 34798 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34920 14384
rect 34920 14344 34922 14384
rect 34630 14302 34754 14344
rect 34798 14302 34922 14344
rect 49750 14384 49874 14426
rect 49918 14384 50042 14426
rect 49750 14344 49752 14384
rect 49752 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49874 14384
rect 49918 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50040 14384
rect 50040 14344 50042 14384
rect 49750 14302 49874 14344
rect 49918 14302 50042 14344
rect 64870 14384 64994 14426
rect 65038 14384 65162 14426
rect 64870 14344 64872 14384
rect 64872 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64994 14384
rect 65038 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65160 14384
rect 65160 14344 65162 14384
rect 64870 14302 64994 14344
rect 65038 14302 65162 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 18270 13628 18394 13670
rect 18438 13628 18562 13670
rect 18270 13588 18272 13628
rect 18272 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18394 13628
rect 18438 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18560 13628
rect 18560 13588 18562 13628
rect 18270 13546 18394 13588
rect 18438 13546 18562 13588
rect 33390 13628 33514 13670
rect 33558 13628 33682 13670
rect 33390 13588 33392 13628
rect 33392 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33514 13628
rect 33558 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33680 13628
rect 33680 13588 33682 13628
rect 33390 13546 33514 13588
rect 33558 13546 33682 13588
rect 48510 13628 48634 13670
rect 48678 13628 48802 13670
rect 48510 13588 48512 13628
rect 48512 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48634 13628
rect 48678 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48800 13628
rect 48800 13588 48802 13628
rect 48510 13546 48634 13588
rect 48678 13546 48802 13588
rect 63630 13628 63754 13670
rect 63798 13628 63922 13670
rect 63630 13588 63632 13628
rect 63632 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63754 13628
rect 63798 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63920 13628
rect 63920 13588 63922 13628
rect 63630 13546 63754 13588
rect 63798 13546 63922 13588
rect 78750 13628 78874 13670
rect 78918 13628 79042 13670
rect 78750 13588 78752 13628
rect 78752 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78874 13628
rect 78918 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79040 13628
rect 79040 13588 79042 13628
rect 78750 13546 78874 13588
rect 78918 13546 79042 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 19510 12872 19634 12914
rect 19678 12872 19802 12914
rect 19510 12832 19512 12872
rect 19512 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19634 12872
rect 19678 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19800 12872
rect 19800 12832 19802 12872
rect 19510 12790 19634 12832
rect 19678 12790 19802 12832
rect 34630 12872 34754 12914
rect 34798 12872 34922 12914
rect 34630 12832 34632 12872
rect 34632 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34754 12872
rect 34798 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34920 12872
rect 34920 12832 34922 12872
rect 34630 12790 34754 12832
rect 34798 12790 34922 12832
rect 49750 12872 49874 12914
rect 49918 12872 50042 12914
rect 49750 12832 49752 12872
rect 49752 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49874 12872
rect 49918 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50040 12872
rect 50040 12832 50042 12872
rect 49750 12790 49874 12832
rect 49918 12790 50042 12832
rect 64870 12872 64994 12914
rect 65038 12872 65162 12914
rect 64870 12832 64872 12872
rect 64872 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64994 12872
rect 65038 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65160 12872
rect 65160 12832 65162 12872
rect 64870 12790 64994 12832
rect 65038 12790 65162 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 18270 12116 18394 12158
rect 18438 12116 18562 12158
rect 18270 12076 18272 12116
rect 18272 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18394 12116
rect 18438 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18560 12116
rect 18560 12076 18562 12116
rect 18270 12034 18394 12076
rect 18438 12034 18562 12076
rect 33390 12116 33514 12158
rect 33558 12116 33682 12158
rect 33390 12076 33392 12116
rect 33392 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33514 12116
rect 33558 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33680 12116
rect 33680 12076 33682 12116
rect 33390 12034 33514 12076
rect 33558 12034 33682 12076
rect 48510 12116 48634 12158
rect 48678 12116 48802 12158
rect 48510 12076 48512 12116
rect 48512 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48634 12116
rect 48678 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48800 12116
rect 48800 12076 48802 12116
rect 48510 12034 48634 12076
rect 48678 12034 48802 12076
rect 63630 12116 63754 12158
rect 63798 12116 63922 12158
rect 63630 12076 63632 12116
rect 63632 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63754 12116
rect 63798 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63920 12116
rect 63920 12076 63922 12116
rect 63630 12034 63754 12076
rect 63798 12034 63922 12076
rect 78750 12116 78874 12158
rect 78918 12116 79042 12158
rect 78750 12076 78752 12116
rect 78752 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78874 12116
rect 78918 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79040 12116
rect 79040 12076 79042 12116
rect 78750 12034 78874 12076
rect 78918 12034 79042 12076
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 19510 11360 19634 11402
rect 19678 11360 19802 11402
rect 19510 11320 19512 11360
rect 19512 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19634 11360
rect 19678 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19800 11360
rect 19800 11320 19802 11360
rect 19510 11278 19634 11320
rect 19678 11278 19802 11320
rect 34630 11360 34754 11402
rect 34798 11360 34922 11402
rect 34630 11320 34632 11360
rect 34632 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34754 11360
rect 34798 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34920 11360
rect 34920 11320 34922 11360
rect 34630 11278 34754 11320
rect 34798 11278 34922 11320
rect 49750 11360 49874 11402
rect 49918 11360 50042 11402
rect 49750 11320 49752 11360
rect 49752 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49874 11360
rect 49918 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50040 11360
rect 50040 11320 50042 11360
rect 49750 11278 49874 11320
rect 49918 11278 50042 11320
rect 64870 11360 64994 11402
rect 65038 11360 65162 11402
rect 64870 11320 64872 11360
rect 64872 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64994 11360
rect 65038 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65160 11360
rect 65160 11320 65162 11360
rect 64870 11278 64994 11320
rect 65038 11278 65162 11320
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 18270 10604 18394 10646
rect 18438 10604 18562 10646
rect 18270 10564 18272 10604
rect 18272 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18394 10604
rect 18438 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18560 10604
rect 18560 10564 18562 10604
rect 18270 10522 18394 10564
rect 18438 10522 18562 10564
rect 33390 10604 33514 10646
rect 33558 10604 33682 10646
rect 33390 10564 33392 10604
rect 33392 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33514 10604
rect 33558 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33680 10604
rect 33680 10564 33682 10604
rect 33390 10522 33514 10564
rect 33558 10522 33682 10564
rect 48510 10604 48634 10646
rect 48678 10604 48802 10646
rect 48510 10564 48512 10604
rect 48512 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48634 10604
rect 48678 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48800 10604
rect 48800 10564 48802 10604
rect 48510 10522 48634 10564
rect 48678 10522 48802 10564
rect 63630 10604 63754 10646
rect 63798 10604 63922 10646
rect 63630 10564 63632 10604
rect 63632 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63754 10604
rect 63798 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63920 10604
rect 63920 10564 63922 10604
rect 63630 10522 63754 10564
rect 63798 10522 63922 10564
rect 78750 10604 78874 10646
rect 78918 10604 79042 10646
rect 78750 10564 78752 10604
rect 78752 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78874 10604
rect 78918 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79040 10604
rect 79040 10564 79042 10604
rect 78750 10522 78874 10564
rect 78918 10522 79042 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 19510 9848 19634 9890
rect 19678 9848 19802 9890
rect 19510 9808 19512 9848
rect 19512 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19634 9848
rect 19678 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19800 9848
rect 19800 9808 19802 9848
rect 19510 9766 19634 9808
rect 19678 9766 19802 9808
rect 34630 9848 34754 9890
rect 34798 9848 34922 9890
rect 34630 9808 34632 9848
rect 34632 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34754 9848
rect 34798 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34920 9848
rect 34920 9808 34922 9848
rect 34630 9766 34754 9808
rect 34798 9766 34922 9808
rect 49750 9848 49874 9890
rect 49918 9848 50042 9890
rect 49750 9808 49752 9848
rect 49752 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49874 9848
rect 49918 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50040 9848
rect 50040 9808 50042 9848
rect 49750 9766 49874 9808
rect 49918 9766 50042 9808
rect 64870 9848 64994 9890
rect 65038 9848 65162 9890
rect 64870 9808 64872 9848
rect 64872 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64994 9848
rect 65038 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65160 9848
rect 65160 9808 65162 9848
rect 64870 9766 64994 9808
rect 65038 9766 65162 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 18270 9092 18394 9134
rect 18438 9092 18562 9134
rect 18270 9052 18272 9092
rect 18272 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18394 9092
rect 18438 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18560 9092
rect 18560 9052 18562 9092
rect 18270 9010 18394 9052
rect 18438 9010 18562 9052
rect 33390 9092 33514 9134
rect 33558 9092 33682 9134
rect 33390 9052 33392 9092
rect 33392 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33514 9092
rect 33558 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33680 9092
rect 33680 9052 33682 9092
rect 33390 9010 33514 9052
rect 33558 9010 33682 9052
rect 48510 9092 48634 9134
rect 48678 9092 48802 9134
rect 48510 9052 48512 9092
rect 48512 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48634 9092
rect 48678 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48800 9092
rect 48800 9052 48802 9092
rect 48510 9010 48634 9052
rect 48678 9010 48802 9052
rect 63630 9092 63754 9134
rect 63798 9092 63922 9134
rect 63630 9052 63632 9092
rect 63632 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63754 9092
rect 63798 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63920 9092
rect 63920 9052 63922 9092
rect 63630 9010 63754 9052
rect 63798 9010 63922 9052
rect 78750 9092 78874 9134
rect 78918 9092 79042 9134
rect 78750 9052 78752 9092
rect 78752 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78874 9092
rect 78918 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79040 9092
rect 79040 9052 79042 9092
rect 78750 9010 78874 9052
rect 78918 9010 79042 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 19510 8336 19634 8378
rect 19678 8336 19802 8378
rect 19510 8296 19512 8336
rect 19512 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19634 8336
rect 19678 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19800 8336
rect 19800 8296 19802 8336
rect 19510 8254 19634 8296
rect 19678 8254 19802 8296
rect 34630 8336 34754 8378
rect 34798 8336 34922 8378
rect 34630 8296 34632 8336
rect 34632 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34754 8336
rect 34798 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34920 8336
rect 34920 8296 34922 8336
rect 34630 8254 34754 8296
rect 34798 8254 34922 8296
rect 49750 8336 49874 8378
rect 49918 8336 50042 8378
rect 49750 8296 49752 8336
rect 49752 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49874 8336
rect 49918 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50040 8336
rect 50040 8296 50042 8336
rect 49750 8254 49874 8296
rect 49918 8254 50042 8296
rect 64870 8336 64994 8378
rect 65038 8336 65162 8378
rect 64870 8296 64872 8336
rect 64872 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64994 8336
rect 65038 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65160 8336
rect 65160 8296 65162 8336
rect 64870 8254 64994 8296
rect 65038 8254 65162 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 18270 7580 18394 7622
rect 18438 7580 18562 7622
rect 18270 7540 18272 7580
rect 18272 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18394 7580
rect 18438 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18560 7580
rect 18560 7540 18562 7580
rect 18270 7498 18394 7540
rect 18438 7498 18562 7540
rect 33390 7580 33514 7622
rect 33558 7580 33682 7622
rect 33390 7540 33392 7580
rect 33392 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33514 7580
rect 33558 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33680 7580
rect 33680 7540 33682 7580
rect 33390 7498 33514 7540
rect 33558 7498 33682 7540
rect 48510 7580 48634 7622
rect 48678 7580 48802 7622
rect 48510 7540 48512 7580
rect 48512 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48634 7580
rect 48678 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48800 7580
rect 48800 7540 48802 7580
rect 48510 7498 48634 7540
rect 48678 7498 48802 7540
rect 63630 7580 63754 7622
rect 63798 7580 63922 7622
rect 63630 7540 63632 7580
rect 63632 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63754 7580
rect 63798 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63920 7580
rect 63920 7540 63922 7580
rect 63630 7498 63754 7540
rect 63798 7498 63922 7540
rect 78750 7580 78874 7622
rect 78918 7580 79042 7622
rect 78750 7540 78752 7580
rect 78752 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78874 7580
rect 78918 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79040 7580
rect 79040 7540 79042 7580
rect 78750 7498 78874 7540
rect 78918 7498 79042 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 19510 6824 19634 6866
rect 19678 6824 19802 6866
rect 19510 6784 19512 6824
rect 19512 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19634 6824
rect 19678 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19800 6824
rect 19800 6784 19802 6824
rect 19510 6742 19634 6784
rect 19678 6742 19802 6784
rect 34630 6824 34754 6866
rect 34798 6824 34922 6866
rect 34630 6784 34632 6824
rect 34632 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34754 6824
rect 34798 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34920 6824
rect 34920 6784 34922 6824
rect 34630 6742 34754 6784
rect 34798 6742 34922 6784
rect 49750 6824 49874 6866
rect 49918 6824 50042 6866
rect 49750 6784 49752 6824
rect 49752 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49874 6824
rect 49918 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50040 6824
rect 50040 6784 50042 6824
rect 49750 6742 49874 6784
rect 49918 6742 50042 6784
rect 64870 6824 64994 6866
rect 65038 6824 65162 6866
rect 64870 6784 64872 6824
rect 64872 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64994 6824
rect 65038 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65160 6824
rect 65160 6784 65162 6824
rect 64870 6742 64994 6784
rect 65038 6742 65162 6784
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 18270 6068 18394 6110
rect 18438 6068 18562 6110
rect 18270 6028 18272 6068
rect 18272 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18394 6068
rect 18438 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18560 6068
rect 18560 6028 18562 6068
rect 18270 5986 18394 6028
rect 18438 5986 18562 6028
rect 33390 6068 33514 6110
rect 33558 6068 33682 6110
rect 33390 6028 33392 6068
rect 33392 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33514 6068
rect 33558 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33680 6068
rect 33680 6028 33682 6068
rect 33390 5986 33514 6028
rect 33558 5986 33682 6028
rect 48510 6068 48634 6110
rect 48678 6068 48802 6110
rect 48510 6028 48512 6068
rect 48512 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48634 6068
rect 48678 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48800 6068
rect 48800 6028 48802 6068
rect 48510 5986 48634 6028
rect 48678 5986 48802 6028
rect 63630 6068 63754 6110
rect 63798 6068 63922 6110
rect 63630 6028 63632 6068
rect 63632 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63754 6068
rect 63798 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63920 6068
rect 63920 6028 63922 6068
rect 63630 5986 63754 6028
rect 63798 5986 63922 6028
rect 78750 6068 78874 6110
rect 78918 6068 79042 6110
rect 78750 6028 78752 6068
rect 78752 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78874 6068
rect 78918 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79040 6068
rect 79040 6028 79042 6068
rect 78750 5986 78874 6028
rect 78918 5986 79042 6028
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 19510 5312 19634 5354
rect 19678 5312 19802 5354
rect 19510 5272 19512 5312
rect 19512 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19634 5312
rect 19678 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19800 5312
rect 19800 5272 19802 5312
rect 19510 5230 19634 5272
rect 19678 5230 19802 5272
rect 34630 5312 34754 5354
rect 34798 5312 34922 5354
rect 34630 5272 34632 5312
rect 34632 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34754 5312
rect 34798 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34920 5312
rect 34920 5272 34922 5312
rect 34630 5230 34754 5272
rect 34798 5230 34922 5272
rect 49750 5312 49874 5354
rect 49918 5312 50042 5354
rect 49750 5272 49752 5312
rect 49752 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49874 5312
rect 49918 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50040 5312
rect 50040 5272 50042 5312
rect 49750 5230 49874 5272
rect 49918 5230 50042 5272
rect 64870 5312 64994 5354
rect 65038 5312 65162 5354
rect 64870 5272 64872 5312
rect 64872 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64994 5312
rect 65038 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65160 5312
rect 65160 5272 65162 5312
rect 64870 5230 64994 5272
rect 65038 5230 65162 5272
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 18270 4556 18394 4598
rect 18438 4556 18562 4598
rect 18270 4516 18272 4556
rect 18272 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18394 4556
rect 18438 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18560 4556
rect 18560 4516 18562 4556
rect 18270 4474 18394 4516
rect 18438 4474 18562 4516
rect 33390 4556 33514 4598
rect 33558 4556 33682 4598
rect 33390 4516 33392 4556
rect 33392 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33514 4556
rect 33558 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33680 4556
rect 33680 4516 33682 4556
rect 33390 4474 33514 4516
rect 33558 4474 33682 4516
rect 48510 4556 48634 4598
rect 48678 4556 48802 4598
rect 48510 4516 48512 4556
rect 48512 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48634 4556
rect 48678 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48800 4556
rect 48800 4516 48802 4556
rect 48510 4474 48634 4516
rect 48678 4474 48802 4516
rect 63630 4556 63754 4598
rect 63798 4556 63922 4598
rect 63630 4516 63632 4556
rect 63632 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63754 4556
rect 63798 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63920 4556
rect 63920 4516 63922 4556
rect 63630 4474 63754 4516
rect 63798 4474 63922 4516
rect 78750 4556 78874 4598
rect 78918 4556 79042 4598
rect 78750 4516 78752 4556
rect 78752 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78874 4556
rect 78918 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79040 4556
rect 79040 4516 79042 4556
rect 78750 4474 78874 4516
rect 78918 4474 79042 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 19510 3800 19634 3842
rect 19678 3800 19802 3842
rect 19510 3760 19512 3800
rect 19512 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19634 3800
rect 19678 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19800 3800
rect 19800 3760 19802 3800
rect 19510 3718 19634 3760
rect 19678 3718 19802 3760
rect 34630 3800 34754 3842
rect 34798 3800 34922 3842
rect 34630 3760 34632 3800
rect 34632 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34754 3800
rect 34798 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34920 3800
rect 34920 3760 34922 3800
rect 34630 3718 34754 3760
rect 34798 3718 34922 3760
rect 49750 3800 49874 3842
rect 49918 3800 50042 3842
rect 49750 3760 49752 3800
rect 49752 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49874 3800
rect 49918 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50040 3800
rect 50040 3760 50042 3800
rect 49750 3718 49874 3760
rect 49918 3718 50042 3760
rect 64870 3800 64994 3842
rect 65038 3800 65162 3842
rect 64870 3760 64872 3800
rect 64872 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64994 3800
rect 65038 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65160 3800
rect 65160 3760 65162 3800
rect 64870 3718 64994 3760
rect 65038 3718 65162 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 18270 3044 18394 3086
rect 18438 3044 18562 3086
rect 18270 3004 18272 3044
rect 18272 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18394 3044
rect 18438 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18560 3044
rect 18560 3004 18562 3044
rect 18270 2962 18394 3004
rect 18438 2962 18562 3004
rect 33390 3044 33514 3086
rect 33558 3044 33682 3086
rect 33390 3004 33392 3044
rect 33392 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33514 3044
rect 33558 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33680 3044
rect 33680 3004 33682 3044
rect 33390 2962 33514 3004
rect 33558 2962 33682 3004
rect 48510 3044 48634 3086
rect 48678 3044 48802 3086
rect 48510 3004 48512 3044
rect 48512 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48634 3044
rect 48678 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48800 3044
rect 48800 3004 48802 3044
rect 48510 2962 48634 3004
rect 48678 2962 48802 3004
rect 63630 3044 63754 3086
rect 63798 3044 63922 3086
rect 63630 3004 63632 3044
rect 63632 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63754 3044
rect 63798 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63920 3044
rect 63920 3004 63922 3044
rect 63630 2962 63754 3004
rect 63798 2962 63922 3004
rect 78750 3044 78874 3086
rect 78918 3044 79042 3086
rect 78750 3004 78752 3044
rect 78752 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78874 3044
rect 78918 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79040 3044
rect 79040 3004 79042 3044
rect 78750 2962 78874 3004
rect 78918 2962 79042 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 19510 2288 19634 2330
rect 19678 2288 19802 2330
rect 19510 2248 19512 2288
rect 19512 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19634 2288
rect 19678 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19800 2288
rect 19800 2248 19802 2288
rect 19510 2206 19634 2248
rect 19678 2206 19802 2248
rect 34630 2288 34754 2330
rect 34798 2288 34922 2330
rect 34630 2248 34632 2288
rect 34632 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34754 2288
rect 34798 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34920 2288
rect 34920 2248 34922 2288
rect 34630 2206 34754 2248
rect 34798 2206 34922 2248
rect 49750 2288 49874 2330
rect 49918 2288 50042 2330
rect 49750 2248 49752 2288
rect 49752 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49874 2288
rect 49918 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50040 2288
rect 50040 2248 50042 2288
rect 49750 2206 49874 2248
rect 49918 2206 50042 2248
rect 64870 2288 64994 2330
rect 65038 2288 65162 2330
rect 64870 2248 64872 2288
rect 64872 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64994 2288
rect 65038 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65160 2288
rect 65160 2248 65162 2288
rect 64870 2206 64994 2248
rect 65038 2206 65162 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 18270 1532 18394 1574
rect 18438 1532 18562 1574
rect 18270 1492 18272 1532
rect 18272 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18394 1532
rect 18438 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18560 1532
rect 18560 1492 18562 1532
rect 18270 1450 18394 1492
rect 18438 1450 18562 1492
rect 33390 1532 33514 1574
rect 33558 1532 33682 1574
rect 33390 1492 33392 1532
rect 33392 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33514 1532
rect 33558 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33680 1532
rect 33680 1492 33682 1532
rect 33390 1450 33514 1492
rect 33558 1450 33682 1492
rect 48510 1532 48634 1574
rect 48678 1532 48802 1574
rect 48510 1492 48512 1532
rect 48512 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48634 1532
rect 48678 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48800 1532
rect 48800 1492 48802 1532
rect 48510 1450 48634 1492
rect 48678 1450 48802 1492
rect 63630 1532 63754 1574
rect 63798 1532 63922 1574
rect 63630 1492 63632 1532
rect 63632 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63754 1532
rect 63798 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63920 1532
rect 63920 1492 63922 1532
rect 63630 1450 63754 1492
rect 63798 1450 63922 1492
rect 78750 1532 78874 1574
rect 78918 1532 79042 1574
rect 78750 1492 78752 1532
rect 78752 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78874 1532
rect 78918 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79040 1532
rect 79040 1492 79042 1532
rect 78750 1450 78874 1492
rect 78918 1450 79042 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 19510 776 19634 818
rect 19678 776 19802 818
rect 19510 736 19512 776
rect 19512 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19634 776
rect 19678 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19800 776
rect 19800 736 19802 776
rect 19510 694 19634 736
rect 19678 694 19802 736
rect 34630 776 34754 818
rect 34798 776 34922 818
rect 34630 736 34632 776
rect 34632 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34754 776
rect 34798 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34920 776
rect 34920 736 34922 776
rect 34630 694 34754 736
rect 34798 694 34922 736
rect 49750 776 49874 818
rect 49918 776 50042 818
rect 49750 736 49752 776
rect 49752 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49874 776
rect 49918 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50040 776
rect 50040 736 50042 776
rect 49750 694 49874 736
rect 49918 694 50042 736
rect 64870 776 64994 818
rect 65038 776 65162 818
rect 64870 736 64872 776
rect 64872 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64994 776
rect 65038 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65160 776
rect 65160 736 65162 776
rect 64870 694 64994 736
rect 65038 694 65162 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 19436 38618 19876 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 18196 37862 18636 38600
rect 18196 37738 18270 37862
rect 18394 37738 18438 37862
rect 18562 37738 18636 37862
rect 18196 36350 18636 37738
rect 18196 36226 18270 36350
rect 18394 36226 18438 36350
rect 18562 36226 18636 36350
rect 18196 34838 18636 36226
rect 18196 34714 18270 34838
rect 18394 34714 18438 34838
rect 18562 34714 18636 34838
rect 18196 33326 18636 34714
rect 18196 33202 18270 33326
rect 18394 33202 18438 33326
rect 18562 33202 18636 33326
rect 18196 31814 18636 33202
rect 18196 31690 18270 31814
rect 18394 31690 18438 31814
rect 18562 31690 18636 31814
rect 18196 30302 18636 31690
rect 18196 30178 18270 30302
rect 18394 30178 18438 30302
rect 18562 30178 18636 30302
rect 18196 28790 18636 30178
rect 18196 28666 18270 28790
rect 18394 28666 18438 28790
rect 18562 28666 18636 28790
rect 18196 27278 18636 28666
rect 18196 27154 18270 27278
rect 18394 27154 18438 27278
rect 18562 27154 18636 27278
rect 18196 25766 18636 27154
rect 18196 25642 18270 25766
rect 18394 25642 18438 25766
rect 18562 25642 18636 25766
rect 18196 24254 18636 25642
rect 18196 24130 18270 24254
rect 18394 24130 18438 24254
rect 18562 24130 18636 24254
rect 18196 22742 18636 24130
rect 18196 22618 18270 22742
rect 18394 22618 18438 22742
rect 18562 22618 18636 22742
rect 18196 21230 18636 22618
rect 18196 21106 18270 21230
rect 18394 21106 18438 21230
rect 18562 21106 18636 21230
rect 18196 19718 18636 21106
rect 18196 19594 18270 19718
rect 18394 19594 18438 19718
rect 18562 19594 18636 19718
rect 18196 18206 18636 19594
rect 18196 18082 18270 18206
rect 18394 18082 18438 18206
rect 18562 18082 18636 18206
rect 18196 16694 18636 18082
rect 18196 16570 18270 16694
rect 18394 16570 18438 16694
rect 18562 16570 18636 16694
rect 18196 15182 18636 16570
rect 18196 15058 18270 15182
rect 18394 15058 18438 15182
rect 18562 15058 18636 15182
rect 18196 13670 18636 15058
rect 18196 13546 18270 13670
rect 18394 13546 18438 13670
rect 18562 13546 18636 13670
rect 18196 12158 18636 13546
rect 18196 12034 18270 12158
rect 18394 12034 18438 12158
rect 18562 12034 18636 12158
rect 18196 10646 18636 12034
rect 18196 10522 18270 10646
rect 18394 10522 18438 10646
rect 18562 10522 18636 10646
rect 18196 9134 18636 10522
rect 18196 9010 18270 9134
rect 18394 9010 18438 9134
rect 18562 9010 18636 9134
rect 18196 7622 18636 9010
rect 18196 7498 18270 7622
rect 18394 7498 18438 7622
rect 18562 7498 18636 7622
rect 18196 6110 18636 7498
rect 18196 5986 18270 6110
rect 18394 5986 18438 6110
rect 18562 5986 18636 6110
rect 18196 4598 18636 5986
rect 18196 4474 18270 4598
rect 18394 4474 18438 4598
rect 18562 4474 18636 4598
rect 18196 3086 18636 4474
rect 18196 2962 18270 3086
rect 18394 2962 18438 3086
rect 18562 2962 18636 3086
rect 18196 1574 18636 2962
rect 18196 1450 18270 1574
rect 18394 1450 18438 1574
rect 18562 1450 18636 1574
rect 18196 712 18636 1450
rect 19436 38494 19510 38618
rect 19634 38494 19678 38618
rect 19802 38494 19876 38618
rect 34556 38618 34996 38682
rect 19436 37106 19876 38494
rect 19436 36982 19510 37106
rect 19634 36982 19678 37106
rect 19802 36982 19876 37106
rect 19436 35594 19876 36982
rect 19436 35470 19510 35594
rect 19634 35470 19678 35594
rect 19802 35470 19876 35594
rect 19436 34082 19876 35470
rect 19436 33958 19510 34082
rect 19634 33958 19678 34082
rect 19802 33958 19876 34082
rect 19436 32570 19876 33958
rect 19436 32446 19510 32570
rect 19634 32446 19678 32570
rect 19802 32446 19876 32570
rect 19436 31058 19876 32446
rect 19436 30934 19510 31058
rect 19634 30934 19678 31058
rect 19802 30934 19876 31058
rect 19436 29546 19876 30934
rect 19436 29422 19510 29546
rect 19634 29422 19678 29546
rect 19802 29422 19876 29546
rect 19436 28034 19876 29422
rect 19436 27910 19510 28034
rect 19634 27910 19678 28034
rect 19802 27910 19876 28034
rect 19436 26522 19876 27910
rect 19436 26398 19510 26522
rect 19634 26398 19678 26522
rect 19802 26398 19876 26522
rect 19436 25010 19876 26398
rect 19436 24886 19510 25010
rect 19634 24886 19678 25010
rect 19802 24886 19876 25010
rect 19436 23498 19876 24886
rect 19436 23374 19510 23498
rect 19634 23374 19678 23498
rect 19802 23374 19876 23498
rect 19436 21986 19876 23374
rect 19436 21862 19510 21986
rect 19634 21862 19678 21986
rect 19802 21862 19876 21986
rect 19436 20474 19876 21862
rect 19436 20350 19510 20474
rect 19634 20350 19678 20474
rect 19802 20350 19876 20474
rect 19436 18962 19876 20350
rect 19436 18838 19510 18962
rect 19634 18838 19678 18962
rect 19802 18838 19876 18962
rect 19436 17450 19876 18838
rect 19436 17326 19510 17450
rect 19634 17326 19678 17450
rect 19802 17326 19876 17450
rect 19436 15938 19876 17326
rect 19436 15814 19510 15938
rect 19634 15814 19678 15938
rect 19802 15814 19876 15938
rect 19436 14426 19876 15814
rect 19436 14302 19510 14426
rect 19634 14302 19678 14426
rect 19802 14302 19876 14426
rect 19436 12914 19876 14302
rect 19436 12790 19510 12914
rect 19634 12790 19678 12914
rect 19802 12790 19876 12914
rect 19436 11402 19876 12790
rect 19436 11278 19510 11402
rect 19634 11278 19678 11402
rect 19802 11278 19876 11402
rect 19436 9890 19876 11278
rect 19436 9766 19510 9890
rect 19634 9766 19678 9890
rect 19802 9766 19876 9890
rect 19436 8378 19876 9766
rect 19436 8254 19510 8378
rect 19634 8254 19678 8378
rect 19802 8254 19876 8378
rect 19436 6866 19876 8254
rect 19436 6742 19510 6866
rect 19634 6742 19678 6866
rect 19802 6742 19876 6866
rect 19436 5354 19876 6742
rect 19436 5230 19510 5354
rect 19634 5230 19678 5354
rect 19802 5230 19876 5354
rect 19436 3842 19876 5230
rect 19436 3718 19510 3842
rect 19634 3718 19678 3842
rect 19802 3718 19876 3842
rect 19436 2330 19876 3718
rect 19436 2206 19510 2330
rect 19634 2206 19678 2330
rect 19802 2206 19876 2330
rect 19436 818 19876 2206
rect 4316 630 4756 694
rect 19436 694 19510 818
rect 19634 694 19678 818
rect 19802 694 19876 818
rect 33316 37862 33756 38600
rect 33316 37738 33390 37862
rect 33514 37738 33558 37862
rect 33682 37738 33756 37862
rect 33316 36350 33756 37738
rect 33316 36226 33390 36350
rect 33514 36226 33558 36350
rect 33682 36226 33756 36350
rect 33316 34838 33756 36226
rect 33316 34714 33390 34838
rect 33514 34714 33558 34838
rect 33682 34714 33756 34838
rect 33316 33326 33756 34714
rect 33316 33202 33390 33326
rect 33514 33202 33558 33326
rect 33682 33202 33756 33326
rect 33316 31814 33756 33202
rect 33316 31690 33390 31814
rect 33514 31690 33558 31814
rect 33682 31690 33756 31814
rect 33316 30302 33756 31690
rect 33316 30178 33390 30302
rect 33514 30178 33558 30302
rect 33682 30178 33756 30302
rect 33316 28790 33756 30178
rect 33316 28666 33390 28790
rect 33514 28666 33558 28790
rect 33682 28666 33756 28790
rect 33316 27278 33756 28666
rect 33316 27154 33390 27278
rect 33514 27154 33558 27278
rect 33682 27154 33756 27278
rect 33316 25766 33756 27154
rect 33316 25642 33390 25766
rect 33514 25642 33558 25766
rect 33682 25642 33756 25766
rect 33316 24254 33756 25642
rect 33316 24130 33390 24254
rect 33514 24130 33558 24254
rect 33682 24130 33756 24254
rect 33316 22742 33756 24130
rect 33316 22618 33390 22742
rect 33514 22618 33558 22742
rect 33682 22618 33756 22742
rect 33316 21230 33756 22618
rect 33316 21106 33390 21230
rect 33514 21106 33558 21230
rect 33682 21106 33756 21230
rect 33316 19718 33756 21106
rect 33316 19594 33390 19718
rect 33514 19594 33558 19718
rect 33682 19594 33756 19718
rect 33316 18206 33756 19594
rect 33316 18082 33390 18206
rect 33514 18082 33558 18206
rect 33682 18082 33756 18206
rect 33316 16694 33756 18082
rect 33316 16570 33390 16694
rect 33514 16570 33558 16694
rect 33682 16570 33756 16694
rect 33316 15182 33756 16570
rect 33316 15058 33390 15182
rect 33514 15058 33558 15182
rect 33682 15058 33756 15182
rect 33316 13670 33756 15058
rect 33316 13546 33390 13670
rect 33514 13546 33558 13670
rect 33682 13546 33756 13670
rect 33316 12158 33756 13546
rect 33316 12034 33390 12158
rect 33514 12034 33558 12158
rect 33682 12034 33756 12158
rect 33316 10646 33756 12034
rect 33316 10522 33390 10646
rect 33514 10522 33558 10646
rect 33682 10522 33756 10646
rect 33316 9134 33756 10522
rect 33316 9010 33390 9134
rect 33514 9010 33558 9134
rect 33682 9010 33756 9134
rect 33316 7622 33756 9010
rect 33316 7498 33390 7622
rect 33514 7498 33558 7622
rect 33682 7498 33756 7622
rect 33316 6110 33756 7498
rect 33316 5986 33390 6110
rect 33514 5986 33558 6110
rect 33682 5986 33756 6110
rect 33316 4598 33756 5986
rect 33316 4474 33390 4598
rect 33514 4474 33558 4598
rect 33682 4474 33756 4598
rect 33316 3086 33756 4474
rect 33316 2962 33390 3086
rect 33514 2962 33558 3086
rect 33682 2962 33756 3086
rect 33316 1574 33756 2962
rect 33316 1450 33390 1574
rect 33514 1450 33558 1574
rect 33682 1450 33756 1574
rect 33316 712 33756 1450
rect 34556 38494 34630 38618
rect 34754 38494 34798 38618
rect 34922 38494 34996 38618
rect 49676 38618 50116 38682
rect 34556 37106 34996 38494
rect 34556 36982 34630 37106
rect 34754 36982 34798 37106
rect 34922 36982 34996 37106
rect 34556 35594 34996 36982
rect 34556 35470 34630 35594
rect 34754 35470 34798 35594
rect 34922 35470 34996 35594
rect 34556 34082 34996 35470
rect 34556 33958 34630 34082
rect 34754 33958 34798 34082
rect 34922 33958 34996 34082
rect 34556 32570 34996 33958
rect 34556 32446 34630 32570
rect 34754 32446 34798 32570
rect 34922 32446 34996 32570
rect 34556 31058 34996 32446
rect 34556 30934 34630 31058
rect 34754 30934 34798 31058
rect 34922 30934 34996 31058
rect 34556 29546 34996 30934
rect 34556 29422 34630 29546
rect 34754 29422 34798 29546
rect 34922 29422 34996 29546
rect 34556 28034 34996 29422
rect 34556 27910 34630 28034
rect 34754 27910 34798 28034
rect 34922 27910 34996 28034
rect 34556 26522 34996 27910
rect 34556 26398 34630 26522
rect 34754 26398 34798 26522
rect 34922 26398 34996 26522
rect 34556 25010 34996 26398
rect 34556 24886 34630 25010
rect 34754 24886 34798 25010
rect 34922 24886 34996 25010
rect 34556 23498 34996 24886
rect 34556 23374 34630 23498
rect 34754 23374 34798 23498
rect 34922 23374 34996 23498
rect 34556 21986 34996 23374
rect 34556 21862 34630 21986
rect 34754 21862 34798 21986
rect 34922 21862 34996 21986
rect 34556 20474 34996 21862
rect 34556 20350 34630 20474
rect 34754 20350 34798 20474
rect 34922 20350 34996 20474
rect 34556 18962 34996 20350
rect 34556 18838 34630 18962
rect 34754 18838 34798 18962
rect 34922 18838 34996 18962
rect 34556 17450 34996 18838
rect 34556 17326 34630 17450
rect 34754 17326 34798 17450
rect 34922 17326 34996 17450
rect 34556 15938 34996 17326
rect 34556 15814 34630 15938
rect 34754 15814 34798 15938
rect 34922 15814 34996 15938
rect 34556 14426 34996 15814
rect 34556 14302 34630 14426
rect 34754 14302 34798 14426
rect 34922 14302 34996 14426
rect 34556 12914 34996 14302
rect 34556 12790 34630 12914
rect 34754 12790 34798 12914
rect 34922 12790 34996 12914
rect 34556 11402 34996 12790
rect 34556 11278 34630 11402
rect 34754 11278 34798 11402
rect 34922 11278 34996 11402
rect 34556 9890 34996 11278
rect 34556 9766 34630 9890
rect 34754 9766 34798 9890
rect 34922 9766 34996 9890
rect 34556 8378 34996 9766
rect 34556 8254 34630 8378
rect 34754 8254 34798 8378
rect 34922 8254 34996 8378
rect 34556 6866 34996 8254
rect 34556 6742 34630 6866
rect 34754 6742 34798 6866
rect 34922 6742 34996 6866
rect 34556 5354 34996 6742
rect 34556 5230 34630 5354
rect 34754 5230 34798 5354
rect 34922 5230 34996 5354
rect 34556 3842 34996 5230
rect 34556 3718 34630 3842
rect 34754 3718 34798 3842
rect 34922 3718 34996 3842
rect 34556 2330 34996 3718
rect 34556 2206 34630 2330
rect 34754 2206 34798 2330
rect 34922 2206 34996 2330
rect 34556 818 34996 2206
rect 19436 630 19876 694
rect 34556 694 34630 818
rect 34754 694 34798 818
rect 34922 694 34996 818
rect 48436 37862 48876 38600
rect 48436 37738 48510 37862
rect 48634 37738 48678 37862
rect 48802 37738 48876 37862
rect 48436 36350 48876 37738
rect 48436 36226 48510 36350
rect 48634 36226 48678 36350
rect 48802 36226 48876 36350
rect 48436 34838 48876 36226
rect 48436 34714 48510 34838
rect 48634 34714 48678 34838
rect 48802 34714 48876 34838
rect 48436 33326 48876 34714
rect 48436 33202 48510 33326
rect 48634 33202 48678 33326
rect 48802 33202 48876 33326
rect 48436 31814 48876 33202
rect 48436 31690 48510 31814
rect 48634 31690 48678 31814
rect 48802 31690 48876 31814
rect 48436 30302 48876 31690
rect 48436 30178 48510 30302
rect 48634 30178 48678 30302
rect 48802 30178 48876 30302
rect 48436 28790 48876 30178
rect 48436 28666 48510 28790
rect 48634 28666 48678 28790
rect 48802 28666 48876 28790
rect 48436 27278 48876 28666
rect 48436 27154 48510 27278
rect 48634 27154 48678 27278
rect 48802 27154 48876 27278
rect 48436 25766 48876 27154
rect 48436 25642 48510 25766
rect 48634 25642 48678 25766
rect 48802 25642 48876 25766
rect 48436 24254 48876 25642
rect 48436 24130 48510 24254
rect 48634 24130 48678 24254
rect 48802 24130 48876 24254
rect 48436 22742 48876 24130
rect 48436 22618 48510 22742
rect 48634 22618 48678 22742
rect 48802 22618 48876 22742
rect 48436 21230 48876 22618
rect 48436 21106 48510 21230
rect 48634 21106 48678 21230
rect 48802 21106 48876 21230
rect 48436 19718 48876 21106
rect 48436 19594 48510 19718
rect 48634 19594 48678 19718
rect 48802 19594 48876 19718
rect 48436 18206 48876 19594
rect 48436 18082 48510 18206
rect 48634 18082 48678 18206
rect 48802 18082 48876 18206
rect 48436 16694 48876 18082
rect 48436 16570 48510 16694
rect 48634 16570 48678 16694
rect 48802 16570 48876 16694
rect 48436 15182 48876 16570
rect 48436 15058 48510 15182
rect 48634 15058 48678 15182
rect 48802 15058 48876 15182
rect 48436 13670 48876 15058
rect 48436 13546 48510 13670
rect 48634 13546 48678 13670
rect 48802 13546 48876 13670
rect 48436 12158 48876 13546
rect 48436 12034 48510 12158
rect 48634 12034 48678 12158
rect 48802 12034 48876 12158
rect 48436 10646 48876 12034
rect 48436 10522 48510 10646
rect 48634 10522 48678 10646
rect 48802 10522 48876 10646
rect 48436 9134 48876 10522
rect 48436 9010 48510 9134
rect 48634 9010 48678 9134
rect 48802 9010 48876 9134
rect 48436 7622 48876 9010
rect 48436 7498 48510 7622
rect 48634 7498 48678 7622
rect 48802 7498 48876 7622
rect 48436 6110 48876 7498
rect 48436 5986 48510 6110
rect 48634 5986 48678 6110
rect 48802 5986 48876 6110
rect 48436 4598 48876 5986
rect 48436 4474 48510 4598
rect 48634 4474 48678 4598
rect 48802 4474 48876 4598
rect 48436 3086 48876 4474
rect 48436 2962 48510 3086
rect 48634 2962 48678 3086
rect 48802 2962 48876 3086
rect 48436 1574 48876 2962
rect 48436 1450 48510 1574
rect 48634 1450 48678 1574
rect 48802 1450 48876 1574
rect 48436 712 48876 1450
rect 49676 38494 49750 38618
rect 49874 38494 49918 38618
rect 50042 38494 50116 38618
rect 64796 38618 65236 38682
rect 49676 37106 50116 38494
rect 49676 36982 49750 37106
rect 49874 36982 49918 37106
rect 50042 36982 50116 37106
rect 49676 35594 50116 36982
rect 49676 35470 49750 35594
rect 49874 35470 49918 35594
rect 50042 35470 50116 35594
rect 49676 34082 50116 35470
rect 49676 33958 49750 34082
rect 49874 33958 49918 34082
rect 50042 33958 50116 34082
rect 49676 32570 50116 33958
rect 49676 32446 49750 32570
rect 49874 32446 49918 32570
rect 50042 32446 50116 32570
rect 49676 31058 50116 32446
rect 49676 30934 49750 31058
rect 49874 30934 49918 31058
rect 50042 30934 50116 31058
rect 49676 29546 50116 30934
rect 49676 29422 49750 29546
rect 49874 29422 49918 29546
rect 50042 29422 50116 29546
rect 49676 28034 50116 29422
rect 49676 27910 49750 28034
rect 49874 27910 49918 28034
rect 50042 27910 50116 28034
rect 49676 26522 50116 27910
rect 49676 26398 49750 26522
rect 49874 26398 49918 26522
rect 50042 26398 50116 26522
rect 49676 25010 50116 26398
rect 49676 24886 49750 25010
rect 49874 24886 49918 25010
rect 50042 24886 50116 25010
rect 49676 23498 50116 24886
rect 49676 23374 49750 23498
rect 49874 23374 49918 23498
rect 50042 23374 50116 23498
rect 49676 21986 50116 23374
rect 49676 21862 49750 21986
rect 49874 21862 49918 21986
rect 50042 21862 50116 21986
rect 49676 20474 50116 21862
rect 49676 20350 49750 20474
rect 49874 20350 49918 20474
rect 50042 20350 50116 20474
rect 49676 18962 50116 20350
rect 49676 18838 49750 18962
rect 49874 18838 49918 18962
rect 50042 18838 50116 18962
rect 49676 17450 50116 18838
rect 49676 17326 49750 17450
rect 49874 17326 49918 17450
rect 50042 17326 50116 17450
rect 49676 15938 50116 17326
rect 49676 15814 49750 15938
rect 49874 15814 49918 15938
rect 50042 15814 50116 15938
rect 49676 14426 50116 15814
rect 49676 14302 49750 14426
rect 49874 14302 49918 14426
rect 50042 14302 50116 14426
rect 49676 12914 50116 14302
rect 49676 12790 49750 12914
rect 49874 12790 49918 12914
rect 50042 12790 50116 12914
rect 49676 11402 50116 12790
rect 49676 11278 49750 11402
rect 49874 11278 49918 11402
rect 50042 11278 50116 11402
rect 49676 9890 50116 11278
rect 49676 9766 49750 9890
rect 49874 9766 49918 9890
rect 50042 9766 50116 9890
rect 49676 8378 50116 9766
rect 49676 8254 49750 8378
rect 49874 8254 49918 8378
rect 50042 8254 50116 8378
rect 49676 6866 50116 8254
rect 49676 6742 49750 6866
rect 49874 6742 49918 6866
rect 50042 6742 50116 6866
rect 49676 5354 50116 6742
rect 49676 5230 49750 5354
rect 49874 5230 49918 5354
rect 50042 5230 50116 5354
rect 49676 3842 50116 5230
rect 49676 3718 49750 3842
rect 49874 3718 49918 3842
rect 50042 3718 50116 3842
rect 49676 2330 50116 3718
rect 49676 2206 49750 2330
rect 49874 2206 49918 2330
rect 50042 2206 50116 2330
rect 49676 818 50116 2206
rect 34556 630 34996 694
rect 49676 694 49750 818
rect 49874 694 49918 818
rect 50042 694 50116 818
rect 63556 37862 63996 38600
rect 63556 37738 63630 37862
rect 63754 37738 63798 37862
rect 63922 37738 63996 37862
rect 63556 36350 63996 37738
rect 63556 36226 63630 36350
rect 63754 36226 63798 36350
rect 63922 36226 63996 36350
rect 63556 34838 63996 36226
rect 63556 34714 63630 34838
rect 63754 34714 63798 34838
rect 63922 34714 63996 34838
rect 63556 33326 63996 34714
rect 63556 33202 63630 33326
rect 63754 33202 63798 33326
rect 63922 33202 63996 33326
rect 63556 31814 63996 33202
rect 63556 31690 63630 31814
rect 63754 31690 63798 31814
rect 63922 31690 63996 31814
rect 63556 30302 63996 31690
rect 63556 30178 63630 30302
rect 63754 30178 63798 30302
rect 63922 30178 63996 30302
rect 63556 28790 63996 30178
rect 63556 28666 63630 28790
rect 63754 28666 63798 28790
rect 63922 28666 63996 28790
rect 63556 27278 63996 28666
rect 63556 27154 63630 27278
rect 63754 27154 63798 27278
rect 63922 27154 63996 27278
rect 63556 25766 63996 27154
rect 63556 25642 63630 25766
rect 63754 25642 63798 25766
rect 63922 25642 63996 25766
rect 63556 19665 63996 25642
rect 63556 19541 63630 19665
rect 63754 19541 63798 19665
rect 63922 19541 63996 19665
rect 63556 19497 63996 19541
rect 63556 19373 63630 19497
rect 63754 19373 63798 19497
rect 63922 19373 63996 19497
rect 63556 19329 63996 19373
rect 63556 19205 63630 19329
rect 63754 19205 63798 19329
rect 63922 19205 63996 19329
rect 63556 19161 63996 19205
rect 63556 19037 63630 19161
rect 63754 19037 63798 19161
rect 63922 19037 63996 19161
rect 63556 18993 63996 19037
rect 63556 18869 63630 18993
rect 63754 18869 63798 18993
rect 63922 18869 63996 18993
rect 63556 18825 63996 18869
rect 63556 18701 63630 18825
rect 63754 18701 63798 18825
rect 63922 18701 63996 18825
rect 63556 18657 63996 18701
rect 63556 18533 63630 18657
rect 63754 18533 63798 18657
rect 63922 18533 63996 18657
rect 63556 18489 63996 18533
rect 63556 18365 63630 18489
rect 63754 18365 63798 18489
rect 63922 18365 63996 18489
rect 63556 18321 63996 18365
rect 63556 18197 63630 18321
rect 63754 18197 63798 18321
rect 63922 18197 63996 18321
rect 63556 18153 63996 18197
rect 63556 18029 63630 18153
rect 63754 18029 63798 18153
rect 63922 18029 63996 18153
rect 63556 17985 63996 18029
rect 63556 17861 63630 17985
rect 63754 17861 63798 17985
rect 63922 17861 63996 17985
rect 63556 17817 63996 17861
rect 63556 17693 63630 17817
rect 63754 17693 63798 17817
rect 63922 17693 63996 17817
rect 63556 17649 63996 17693
rect 63556 17525 63630 17649
rect 63754 17525 63798 17649
rect 63922 17525 63996 17649
rect 63556 15182 63996 17525
rect 63556 15058 63630 15182
rect 63754 15058 63798 15182
rect 63922 15058 63996 15182
rect 63556 13670 63996 15058
rect 63556 13546 63630 13670
rect 63754 13546 63798 13670
rect 63922 13546 63996 13670
rect 63556 12158 63996 13546
rect 63556 12034 63630 12158
rect 63754 12034 63798 12158
rect 63922 12034 63996 12158
rect 63556 10646 63996 12034
rect 63556 10522 63630 10646
rect 63754 10522 63798 10646
rect 63922 10522 63996 10646
rect 63556 9134 63996 10522
rect 63556 9010 63630 9134
rect 63754 9010 63798 9134
rect 63922 9010 63996 9134
rect 63556 7622 63996 9010
rect 63556 7498 63630 7622
rect 63754 7498 63798 7622
rect 63922 7498 63996 7622
rect 63556 6110 63996 7498
rect 63556 5986 63630 6110
rect 63754 5986 63798 6110
rect 63922 5986 63996 6110
rect 63556 4598 63996 5986
rect 63556 4474 63630 4598
rect 63754 4474 63798 4598
rect 63922 4474 63996 4598
rect 63556 3086 63996 4474
rect 63556 2962 63630 3086
rect 63754 2962 63798 3086
rect 63922 2962 63996 3086
rect 63556 1574 63996 2962
rect 63556 1450 63630 1574
rect 63754 1450 63798 1574
rect 63922 1450 63996 1574
rect 63556 712 63996 1450
rect 64796 38494 64870 38618
rect 64994 38494 65038 38618
rect 65162 38494 65236 38618
rect 64796 37106 65236 38494
rect 64796 36982 64870 37106
rect 64994 36982 65038 37106
rect 65162 36982 65236 37106
rect 64796 35594 65236 36982
rect 64796 35470 64870 35594
rect 64994 35470 65038 35594
rect 65162 35470 65236 35594
rect 64796 34082 65236 35470
rect 64796 33958 64870 34082
rect 64994 33958 65038 34082
rect 65162 33958 65236 34082
rect 64796 32570 65236 33958
rect 64796 32446 64870 32570
rect 64994 32446 65038 32570
rect 65162 32446 65236 32570
rect 64796 31058 65236 32446
rect 64796 30934 64870 31058
rect 64994 30934 65038 31058
rect 65162 30934 65236 31058
rect 64796 29546 65236 30934
rect 64796 29422 64870 29546
rect 64994 29422 65038 29546
rect 65162 29422 65236 29546
rect 64796 28034 65236 29422
rect 64796 27910 64870 28034
rect 64994 27910 65038 28034
rect 65162 27910 65236 28034
rect 64796 26522 65236 27910
rect 64796 26398 64870 26522
rect 64994 26398 65038 26522
rect 65162 26398 65236 26522
rect 64796 25010 65236 26398
rect 64796 24886 64870 25010
rect 64994 24886 65038 25010
rect 65162 24886 65236 25010
rect 64796 22541 65236 24886
rect 64796 22417 64870 22541
rect 64994 22417 65038 22541
rect 65162 22417 65236 22541
rect 64796 22373 65236 22417
rect 64796 22249 64870 22373
rect 64994 22249 65038 22373
rect 65162 22249 65236 22373
rect 64796 22205 65236 22249
rect 64796 22081 64870 22205
rect 64994 22081 65038 22205
rect 65162 22081 65236 22205
rect 64796 22037 65236 22081
rect 64796 21913 64870 22037
rect 64994 21913 65038 22037
rect 65162 21913 65236 22037
rect 64796 21869 65236 21913
rect 64796 21745 64870 21869
rect 64994 21745 65038 21869
rect 65162 21745 65236 21869
rect 64796 21701 65236 21745
rect 64796 21577 64870 21701
rect 64994 21577 65038 21701
rect 65162 21577 65236 21701
rect 64796 21533 65236 21577
rect 64796 21409 64870 21533
rect 64994 21409 65038 21533
rect 65162 21409 65236 21533
rect 64796 21365 65236 21409
rect 64796 21241 64870 21365
rect 64994 21241 65038 21365
rect 65162 21241 65236 21365
rect 64796 21197 65236 21241
rect 64796 21073 64870 21197
rect 64994 21073 65038 21197
rect 65162 21073 65236 21197
rect 64796 21029 65236 21073
rect 64796 20905 64870 21029
rect 64994 20905 65038 21029
rect 65162 20905 65236 21029
rect 64796 20861 65236 20905
rect 64796 20737 64870 20861
rect 64994 20737 65038 20861
rect 65162 20737 65236 20861
rect 64796 20693 65236 20737
rect 64796 20569 64870 20693
rect 64994 20569 65038 20693
rect 65162 20569 65236 20693
rect 64796 20525 65236 20569
rect 64796 20401 64870 20525
rect 64994 20401 65038 20525
rect 65162 20401 65236 20525
rect 64796 14426 65236 20401
rect 64796 14302 64870 14426
rect 64994 14302 65038 14426
rect 65162 14302 65236 14426
rect 64796 12914 65236 14302
rect 64796 12790 64870 12914
rect 64994 12790 65038 12914
rect 65162 12790 65236 12914
rect 64796 11402 65236 12790
rect 64796 11278 64870 11402
rect 64994 11278 65038 11402
rect 65162 11278 65236 11402
rect 64796 9890 65236 11278
rect 64796 9766 64870 9890
rect 64994 9766 65038 9890
rect 65162 9766 65236 9890
rect 64796 8378 65236 9766
rect 64796 8254 64870 8378
rect 64994 8254 65038 8378
rect 65162 8254 65236 8378
rect 64796 6866 65236 8254
rect 64796 6742 64870 6866
rect 64994 6742 65038 6866
rect 65162 6742 65236 6866
rect 64796 5354 65236 6742
rect 64796 5230 64870 5354
rect 64994 5230 65038 5354
rect 65162 5230 65236 5354
rect 64796 3842 65236 5230
rect 64796 3718 64870 3842
rect 64994 3718 65038 3842
rect 65162 3718 65236 3842
rect 64796 2330 65236 3718
rect 64796 2206 64870 2330
rect 64994 2206 65038 2330
rect 65162 2206 65236 2330
rect 64796 818 65236 2206
rect 49676 630 50116 694
rect 64796 694 64870 818
rect 64994 694 65038 818
rect 65162 694 65236 818
rect 78676 37862 79116 38600
rect 78676 37738 78750 37862
rect 78874 37738 78918 37862
rect 79042 37738 79116 37862
rect 78676 36350 79116 37738
rect 78676 36226 78750 36350
rect 78874 36226 78918 36350
rect 79042 36226 79116 36350
rect 78676 34838 79116 36226
rect 78676 34714 78750 34838
rect 78874 34714 78918 34838
rect 79042 34714 79116 34838
rect 78676 33326 79116 34714
rect 78676 33202 78750 33326
rect 78874 33202 78918 33326
rect 79042 33202 79116 33326
rect 78676 31814 79116 33202
rect 78676 31690 78750 31814
rect 78874 31690 78918 31814
rect 79042 31690 79116 31814
rect 78676 30302 79116 31690
rect 78676 30178 78750 30302
rect 78874 30178 78918 30302
rect 79042 30178 79116 30302
rect 78676 28790 79116 30178
rect 78676 28666 78750 28790
rect 78874 28666 78918 28790
rect 79042 28666 79116 28790
rect 78676 27278 79116 28666
rect 78676 27154 78750 27278
rect 78874 27154 78918 27278
rect 79042 27154 79116 27278
rect 78676 25766 79116 27154
rect 78676 25642 78750 25766
rect 78874 25642 78918 25766
rect 79042 25642 79116 25766
rect 78676 19665 79116 25642
rect 78676 19541 78750 19665
rect 78874 19541 78918 19665
rect 79042 19541 79116 19665
rect 78676 19497 79116 19541
rect 78676 19373 78750 19497
rect 78874 19373 78918 19497
rect 79042 19373 79116 19497
rect 78676 19329 79116 19373
rect 78676 19205 78750 19329
rect 78874 19205 78918 19329
rect 79042 19205 79116 19329
rect 78676 19161 79116 19205
rect 78676 19037 78750 19161
rect 78874 19037 78918 19161
rect 79042 19037 79116 19161
rect 78676 18993 79116 19037
rect 78676 18869 78750 18993
rect 78874 18869 78918 18993
rect 79042 18869 79116 18993
rect 78676 18825 79116 18869
rect 78676 18701 78750 18825
rect 78874 18701 78918 18825
rect 79042 18701 79116 18825
rect 78676 18657 79116 18701
rect 78676 18533 78750 18657
rect 78874 18533 78918 18657
rect 79042 18533 79116 18657
rect 78676 18489 79116 18533
rect 78676 18365 78750 18489
rect 78874 18365 78918 18489
rect 79042 18365 79116 18489
rect 78676 18321 79116 18365
rect 78676 18197 78750 18321
rect 78874 18197 78918 18321
rect 79042 18197 79116 18321
rect 78676 18153 79116 18197
rect 78676 18029 78750 18153
rect 78874 18029 78918 18153
rect 79042 18029 79116 18153
rect 78676 17985 79116 18029
rect 78676 17861 78750 17985
rect 78874 17861 78918 17985
rect 79042 17861 79116 17985
rect 78676 17817 79116 17861
rect 78676 17693 78750 17817
rect 78874 17693 78918 17817
rect 79042 17693 79116 17817
rect 78676 17649 79116 17693
rect 78676 17525 78750 17649
rect 78874 17525 78918 17649
rect 79042 17525 79116 17649
rect 78676 15182 79116 17525
rect 78676 15058 78750 15182
rect 78874 15058 78918 15182
rect 79042 15058 79116 15182
rect 78676 13670 79116 15058
rect 78676 13546 78750 13670
rect 78874 13546 78918 13670
rect 79042 13546 79116 13670
rect 78676 12158 79116 13546
rect 78676 12034 78750 12158
rect 78874 12034 78918 12158
rect 79042 12034 79116 12158
rect 78676 10646 79116 12034
rect 78676 10522 78750 10646
rect 78874 10522 78918 10646
rect 79042 10522 79116 10646
rect 78676 9134 79116 10522
rect 78676 9010 78750 9134
rect 78874 9010 78918 9134
rect 79042 9010 79116 9134
rect 78676 7622 79116 9010
rect 78676 7498 78750 7622
rect 78874 7498 78918 7622
rect 79042 7498 79116 7622
rect 78676 6110 79116 7498
rect 78676 5986 78750 6110
rect 78874 5986 78918 6110
rect 79042 5986 79116 6110
rect 78676 4598 79116 5986
rect 78676 4474 78750 4598
rect 78874 4474 78918 4598
rect 79042 4474 79116 4598
rect 78676 3086 79116 4474
rect 78676 2962 78750 3086
rect 78874 2962 78918 3086
rect 79042 2962 79116 3086
rect 78676 1574 79116 2962
rect 78676 1450 78750 1574
rect 78874 1450 78918 1574
rect 79042 1450 79116 1574
rect 78676 712 79116 1450
rect 64796 630 65236 694
use sg13g2_inv_1  _1284_
timestamp 1676382929
transform 1 0 52224 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1285_
timestamp 1676382929
transform -1 0 4416 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1286_
timestamp 1676382929
transform 1 0 52512 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1287_
timestamp 1676382929
transform 1 0 52224 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1288_
timestamp 1676382929
transform 1 0 54720 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1289_
timestamp 1676382929
transform 1 0 55104 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1290_
timestamp 1676382929
transform -1 0 56256 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1291_
timestamp 1676382929
transform -1 0 56544 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1292_
timestamp 1676382929
transform 1 0 56544 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1293_
timestamp 1676382929
transform 1 0 56832 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1294_
timestamp 1676382929
transform 1 0 57216 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1295_
timestamp 1676382929
transform 1 0 57600 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1296_
timestamp 1676382929
transform 1 0 57984 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1297_
timestamp 1676382929
transform 1 0 58368 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1298_
timestamp 1676382929
transform 1 0 58752 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1299_
timestamp 1676382929
transform 1 0 59232 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1300_
timestamp 1676382929
transform 1 0 59616 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1301_
timestamp 1676382929
transform 1 0 60000 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1302_
timestamp 1676382929
transform 1 0 60384 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1303_
timestamp 1676382929
transform 1 0 60768 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1304_
timestamp 1676382929
transform 1 0 61248 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1305_
timestamp 1676382929
transform 1 0 61632 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1306_
timestamp 1676382929
transform 1 0 62016 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1307_
timestamp 1676382929
transform 1 0 62400 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1308_
timestamp 1676382929
transform 1 0 62784 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1309_
timestamp 1676382929
transform 1 0 63168 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1310_
timestamp 1676382929
transform 1 0 63552 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1311_
timestamp 1676382929
transform 1 0 64032 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1312_
timestamp 1676382929
transform 1 0 64416 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1313_
timestamp 1676382929
transform 1 0 64800 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1314_
timestamp 1676382929
transform 1 0 65184 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1315_
timestamp 1676382929
transform 1 0 65664 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1316_
timestamp 1676382929
transform 1 0 66048 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1317_
timestamp 1676382929
transform 1 0 66432 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1318_
timestamp 1676382929
transform 1 0 66816 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1319_
timestamp 1676382929
transform 1 0 67200 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1320_
timestamp 1676382929
transform 1 0 67584 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1321_
timestamp 1676382929
transform 1 0 68064 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1322_
timestamp 1676382929
transform 1 0 68448 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1323_
timestamp 1676382929
transform 1 0 68832 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1324_
timestamp 1676382929
transform 1 0 69216 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1325_
timestamp 1676382929
transform 1 0 69600 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1326_
timestamp 1676382929
transform 1 0 70080 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1327_
timestamp 1676382929
transform 1 0 70464 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1328_
timestamp 1676382929
transform 1 0 70848 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1329_
timestamp 1676382929
transform 1 0 71232 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1330_
timestamp 1676382929
transform 1 0 71616 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1331_
timestamp 1676382929
transform 1 0 72000 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1332_
timestamp 1676382929
transform 1 0 72384 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1333_
timestamp 1676382929
transform 1 0 72768 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1334_
timestamp 1676382929
transform 1 0 73248 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1335_
timestamp 1676382929
transform 1 0 73632 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1336_
timestamp 1676382929
transform 1 0 74016 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1337_
timestamp 1676382929
transform 1 0 74400 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1338_
timestamp 1676382929
transform 1 0 74784 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1339_
timestamp 1676382929
transform 1 0 75168 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1340_
timestamp 1676382929
transform 1 0 75552 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1341_
timestamp 1676382929
transform 1 0 76032 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1342_
timestamp 1676382929
transform -1 0 77088 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1343_
timestamp 1676382929
transform -1 0 77376 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1344_
timestamp 1676382929
transform -1 0 77664 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1345_
timestamp 1676382929
transform 1 0 77664 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1346_
timestamp 1676382929
transform 1 0 78048 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1347_
timestamp 1676382929
transform 1 0 78432 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1348_
timestamp 1676382929
transform 1 0 78720 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1349_
timestamp 1676382929
transform 1 0 79104 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1350_
timestamp 1676382929
transform 1 0 78528 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1351_
timestamp 1676382929
transform 1 0 78144 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1352_
timestamp 1676382929
transform 1 0 77856 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1353_
timestamp 1676382929
transform 1 0 77472 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1354_
timestamp 1676382929
transform 1 0 77088 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1355_
timestamp 1676382929
transform -1 0 77088 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1356_
timestamp 1676382929
transform -1 0 76704 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1357_
timestamp 1676382929
transform 1 0 75648 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1358_
timestamp 1676382929
transform 1 0 75264 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1359_
timestamp 1676382929
transform 1 0 74880 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1360_
timestamp 1676382929
transform 1 0 74496 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1361_
timestamp 1676382929
transform 1 0 74112 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1362_
timestamp 1676382929
transform 1 0 73632 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1363_
timestamp 1676382929
transform 1 0 73248 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1364_
timestamp 1676382929
transform 1 0 72864 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1365_
timestamp 1676382929
transform 1 0 72480 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1366_
timestamp 1676382929
transform 1 0 72096 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1367_
timestamp 1676382929
transform 1 0 71712 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1368_
timestamp 1676382929
transform 1 0 71232 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1369_
timestamp 1676382929
transform 1 0 70848 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1370_
timestamp 1676382929
transform 1 0 70464 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1371_
timestamp 1676382929
transform 1 0 70080 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1372_
timestamp 1676382929
transform 1 0 69696 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1373_
timestamp 1676382929
transform 1 0 69312 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1374_
timestamp 1676382929
transform 1 0 68832 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1375_
timestamp 1676382929
transform 1 0 68448 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1376_
timestamp 1676382929
transform 1 0 68064 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1377_
timestamp 1676382929
transform 1 0 67680 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1378_
timestamp 1676382929
transform 1 0 67296 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1379_
timestamp 1676382929
transform 1 0 66912 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1380_
timestamp 1676382929
transform 1 0 66432 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1381_
timestamp 1676382929
transform 1 0 66048 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1382_
timestamp 1676382929
transform 1 0 65664 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1383_
timestamp 1676382929
transform 1 0 65280 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1384_
timestamp 1676382929
transform 1 0 64896 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1385_
timestamp 1676382929
transform 1 0 64416 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1386_
timestamp 1676382929
transform 1 0 64032 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1387_
timestamp 1676382929
transform 1 0 63648 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1388_
timestamp 1676382929
transform 1 0 63264 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1389_
timestamp 1676382929
transform 1 0 62880 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1390_
timestamp 1676382929
transform 1 0 62592 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1391_
timestamp 1676382929
transform 1 0 62304 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1392_
timestamp 1676382929
transform 1 0 62016 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1393_
timestamp 1676382929
transform 1 0 61344 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1394_
timestamp 1676382929
transform 1 0 60672 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1395_
timestamp 1676382929
transform 1 0 60384 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1396_
timestamp 1676382929
transform 1 0 60000 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1397_
timestamp 1676382929
transform 1 0 59616 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1398_
timestamp 1676382929
transform 1 0 59232 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1399_
timestamp 1676382929
transform 1 0 58848 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1400_
timestamp 1676382929
transform 1 0 58464 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1401_
timestamp 1676382929
transform 1 0 58176 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1402_
timestamp 1676382929
transform 1 0 57888 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1403_
timestamp 1676382929
transform 1 0 57216 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1404_
timestamp 1676382929
transform 1 0 56832 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1405_
timestamp 1676382929
transform 1 0 56448 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1406_
timestamp 1676382929
transform 1 0 55968 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1407_
timestamp 1676382929
transform 1 0 55584 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1408_
timestamp 1676382929
transform 1 0 55200 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1409_
timestamp 1676382929
transform 1 0 54912 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1410_
timestamp 1676382929
transform 1 0 54624 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1411_
timestamp 1676382929
transform 1 0 52224 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1412_
timestamp 1676382929
transform 1 0 52224 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1413_
timestamp 1676382929
transform -1 0 4800 0 -1 20412
box -48 -56 336 834
use sg13g2_mux2_1  _1414_
timestamp 1677247768
transform -1 0 23616 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1415_
timestamp 1676557249
transform 1 0 22464 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1416_
timestamp 1676627187
transform -1 0 2208 0 -1 23436
box -48 -56 432 834
use sg13g2_or2_1  _1417_
timestamp 1684236171
transform 1 0 1344 0 -1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _1418_
timestamp 1683973020
transform -1 0 3936 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1419_
timestamp 1685175443
transform -1 0 22560 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1420_
timestamp 1683973020
transform 1 0 22464 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1421_
timestamp 1677247768
transform 1 0 26688 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1422_
timestamp 1676557249
transform 1 0 27648 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1423_
timestamp 1683973020
transform -1 0 25632 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1424_
timestamp 1685175443
transform -1 0 26112 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1425_
timestamp 1683973020
transform 1 0 26112 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1426_
timestamp 1677247768
transform -1 0 30912 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1427_
timestamp 1676557249
transform -1 0 29952 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1428_
timestamp 1683973020
transform -1 0 29088 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1429_
timestamp 1685175443
transform -1 0 30336 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1430_
timestamp 1683973020
transform -1 0 29184 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1431_
timestamp 1677247768
transform 1 0 32736 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1432_
timestamp 1676557249
transform 1 0 33696 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1433_
timestamp 1683973020
transform -1 0 32256 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1434_
timestamp 1685175443
transform -1 0 33024 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1435_
timestamp 1683973020
transform -1 0 32544 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1436_
timestamp 1677247768
transform -1 0 36960 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1437_
timestamp 1676557249
transform -1 0 36000 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1438_
timestamp 1683973020
transform -1 0 35232 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1439_
timestamp 1685175443
transform -1 0 36384 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1440_
timestamp 1683973020
transform -1 0 35904 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1441_
timestamp 1677247768
transform -1 0 39936 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1442_
timestamp 1676557249
transform -1 0 38592 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1443_
timestamp 1683973020
transform -1 0 38208 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1444_
timestamp 1685175443
transform -1 0 39360 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1445_
timestamp 1683973020
transform -1 0 38592 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _1446_
timestamp 1677247768
transform 1 0 42624 0 1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1447_
timestamp 1676557249
transform 1 0 43488 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1448_
timestamp 1683973020
transform -1 0 41376 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1449_
timestamp 1685175443
transform -1 0 42720 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1450_
timestamp 1683973020
transform -1 0 42336 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1451_
timestamp 1677247768
transform 1 0 42048 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1452_
timestamp 1676557249
transform 1 0 43872 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1453_
timestamp 1683973020
transform 1 0 42336 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1454_
timestamp 1685175443
transform -1 0 42048 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1455_
timestamp 1683973020
transform 1 0 41856 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1456_
timestamp 1677247768
transform -1 0 43776 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1457_
timestamp 1676557249
transform -1 0 43008 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1458_
timestamp 1683973020
transform 1 0 41760 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1459_
timestamp 1685175443
transform 1 0 41088 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1460_
timestamp 1683973020
transform 1 0 41376 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1461_
timestamp 1677247768
transform -1 0 40320 0 -1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1462_
timestamp 1676557249
transform 1 0 38976 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1463_
timestamp 1683973020
transform -1 0 40224 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1464_
timestamp 1685175443
transform 1 0 39072 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1465_
timestamp 1683973020
transform 1 0 39936 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1466_
timestamp 1677247768
transform 1 0 36672 0 1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1467_
timestamp 1676557249
transform -1 0 38592 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1468_
timestamp 1683973020
transform 1 0 38400 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1469_
timestamp 1685175443
transform 1 0 36192 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1470_
timestamp 1683973020
transform 1 0 36672 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1471_
timestamp 1677247768
transform 1 0 33600 0 1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1472_
timestamp 1676557249
transform 1 0 34560 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1473_
timestamp 1683973020
transform 1 0 34848 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1474_
timestamp 1685175443
transform 1 0 33312 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1475_
timestamp 1683973020
transform 1 0 33792 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1476_
timestamp 1677247768
transform 1 0 32064 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1477_
timestamp 1676557249
transform -1 0 33120 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1478_
timestamp 1683973020
transform 1 0 33120 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1479_
timestamp 1685175443
transform -1 0 32064 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1480_
timestamp 1683973020
transform 1 0 32736 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1481_
timestamp 1677247768
transform -1 0 37344 0 -1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1482_
timestamp 1676557249
transform -1 0 36480 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1483_
timestamp 1683973020
transform -1 0 35328 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1484_
timestamp 1685175443
transform -1 0 35712 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1485_
timestamp 1683973020
transform 1 0 34752 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1486_
timestamp 1677247768
transform 1 0 38400 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1487_
timestamp 1676557249
transform -1 0 39744 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1488_
timestamp 1683973020
transform -1 0 36864 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1489_
timestamp 1685175443
transform -1 0 37824 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1490_
timestamp 1683973020
transform -1 0 37344 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1491_
timestamp 1677247768
transform 1 0 41376 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1492_
timestamp 1676557249
transform 1 0 42816 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1493_
timestamp 1683973020
transform -1 0 39648 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1494_
timestamp 1685175443
transform -1 0 41088 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1495_
timestamp 1683973020
transform -1 0 40416 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1496_
timestamp 1677247768
transform -1 0 44448 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1497_
timestamp 1676557249
transform 1 0 43872 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1498_
timestamp 1683973020
transform -1 0 42144 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1499_
timestamp 1685175443
transform -1 0 43200 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1500_
timestamp 1683973020
transform -1 0 42624 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1501_
timestamp 1677247768
transform -1 0 47232 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1502_
timestamp 1676557249
transform 1 0 46656 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1503_
timestamp 1683973020
transform -1 0 44544 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1504_
timestamp 1685175443
transform -1 0 45792 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1505_
timestamp 1683973020
transform -1 0 45120 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1506_
timestamp 1677247768
transform 1 0 47808 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1507_
timestamp 1676557249
transform -1 0 48768 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1508_
timestamp 1683973020
transform -1 0 47136 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1509_
timestamp 1685175443
transform -1 0 47616 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1510_
timestamp 1683973020
transform -1 0 47616 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1511_
timestamp 1677247768
transform 1 0 48000 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1512_
timestamp 1676557249
transform -1 0 48768 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1513_
timestamp 1683973020
transform 1 0 47616 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1514_
timestamp 1685175443
transform -1 0 47808 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1515_
timestamp 1683973020
transform 1 0 47136 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1516_
timestamp 1677247768
transform 1 0 51552 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1517_
timestamp 1676557249
transform 1 0 52416 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1518_
timestamp 1683973020
transform -1 0 49248 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1519_
timestamp 1685175443
transform -1 0 51072 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1520_
timestamp 1683973020
transform -1 0 50496 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1521_
timestamp 1677247768
transform 1 0 53664 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1522_
timestamp 1676557249
transform -1 0 54528 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1523_
timestamp 1683973020
transform -1 0 52416 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1524_
timestamp 1685175443
transform -1 0 53184 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1525_
timestamp 1683973020
transform -1 0 52704 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1526_
timestamp 1677247768
transform 1 0 52992 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1527_
timestamp 1676557249
transform -1 0 53952 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1528_
timestamp 1683973020
transform 1 0 53184 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1529_
timestamp 1685175443
transform -1 0 53472 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1530_
timestamp 1683973020
transform 1 0 52704 0 1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _1531_
timestamp 1677247768
transform 1 0 52608 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1532_
timestamp 1676557249
transform 1 0 53568 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1533_
timestamp 1683973020
transform 1 0 52608 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1534_
timestamp 1685175443
transform 1 0 52128 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1535_
timestamp 1683973020
transform 1 0 52416 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1536_
timestamp 1677247768
transform 1 0 50688 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1537_
timestamp 1676557249
transform 1 0 52128 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1538_
timestamp 1683973020
transform 1 0 51360 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1539_
timestamp 1685175443
transform 1 0 50688 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1540_
timestamp 1683973020
transform 1 0 51168 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1541_
timestamp 1677247768
transform 1 0 47808 0 -1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1542_
timestamp 1676557249
transform -1 0 48864 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1543_
timestamp 1683973020
transform 1 0 49152 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1544_
timestamp 1685175443
transform 1 0 47712 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1545_
timestamp 1683973020
transform 1 0 48192 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1546_
timestamp 1677247768
transform 1 0 46848 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1547_
timestamp 1676557249
transform -1 0 47808 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1548_
timestamp 1683973020
transform 1 0 47808 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1549_
timestamp 1685175443
transform -1 0 46080 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1550_
timestamp 1683973020
transform 1 0 46080 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1551_
timestamp 1677247768
transform 1 0 45216 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1552_
timestamp 1676557249
transform 1 0 47040 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1553_
timestamp 1683973020
transform -1 0 46464 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1554_
timestamp 1685175443
transform 1 0 45408 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1555_
timestamp 1683973020
transform 1 0 45888 0 -1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _1556_
timestamp 1677247768
transform 1 0 48192 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _1557_
timestamp 1676557249
transform -1 0 49536 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1558_
timestamp 1683973020
transform -1 0 46560 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1559_
timestamp 1685175443
transform -1 0 47808 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1560_
timestamp 1683973020
transform -1 0 47136 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1561_
timestamp 1677247768
transform 1 0 50208 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2_1  _1562_
timestamp 1676557249
transform 1 0 51552 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1563_
timestamp 1683973020
transform -1 0 49056 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1564_
timestamp 1685175443
transform -1 0 50112 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1565_
timestamp 1683973020
transform -1 0 49536 0 -1 17388
box -48 -56 528 834
use sg13g2_mux2_1  _1566_
timestamp 1677247768
transform -1 0 52992 0 1 15876
box -48 -56 1008 834
use sg13g2_nand2_1  _1567_
timestamp 1676557249
transform 1 0 52416 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1568_
timestamp 1683973020
transform -1 0 51168 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1569_
timestamp 1685175443
transform -1 0 51936 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1570_
timestamp 1683973020
transform -1 0 51552 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1571_
timestamp 1677247768
transform 1 0 55872 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1572_
timestamp 1676557249
transform -1 0 56736 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1573_
timestamp 1683973020
transform -1 0 53664 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1574_
timestamp 1685175443
transform -1 0 55488 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1575_
timestamp 1683973020
transform -1 0 54816 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1576_
timestamp 1677247768
transform 1 0 57600 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1577_
timestamp 1676557249
transform -1 0 58464 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1578_
timestamp 1683973020
transform -1 0 56448 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1579_
timestamp 1685175443
transform -1 0 56928 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1580_
timestamp 1683973020
transform 1 0 56448 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1581_
timestamp 1677247768
transform -1 0 60000 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1582_
timestamp 1676557249
transform 1 0 59040 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1583_
timestamp 1683973020
transform 1 0 57600 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1584_
timestamp 1685175443
transform -1 0 58560 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1585_
timestamp 1683973020
transform -1 0 58176 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1586_
timestamp 1677247768
transform 1 0 58176 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1587_
timestamp 1676557249
transform -1 0 58944 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1588_
timestamp 1683973020
transform 1 0 58176 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1589_
timestamp 1685175443
transform -1 0 58176 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1590_
timestamp 1683973020
transform 1 0 57696 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1591_
timestamp 1677247768
transform 1 0 59520 0 1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1592_
timestamp 1676557249
transform -1 0 60480 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1593_
timestamp 1683973020
transform -1 0 58944 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1594_
timestamp 1685175443
transform -1 0 58944 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1595_
timestamp 1683973020
transform 1 0 57984 0 -1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _1596_
timestamp 1677247768
transform 1 0 60672 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1597_
timestamp 1676557249
transform 1 0 62112 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1598_
timestamp 1683973020
transform -1 0 59616 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1599_
timestamp 1685175443
transform 1 0 58944 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1600_
timestamp 1683973020
transform 1 0 59136 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1601_
timestamp 1677247768
transform 1 0 56064 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1602_
timestamp 1676557249
transform -1 0 57024 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1603_
timestamp 1683973020
transform 1 0 57888 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1604_
timestamp 1685175443
transform -1 0 56064 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1605_
timestamp 1683973020
transform 1 0 57024 0 1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1606_
timestamp 1677247768
transform -1 0 56832 0 1 756
box -48 -56 1008 834
use sg13g2_nand2_1  _1607_
timestamp 1676557249
transform 1 0 56064 0 -1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1608_
timestamp 1683973020
transform 1 0 55680 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1609_
timestamp 1685175443
transform -1 0 55680 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1610_
timestamp 1683973020
transform 1 0 55296 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1611_
timestamp 1677247768
transform 1 0 59232 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1612_
timestamp 1676557249
transform 1 0 60192 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1613_
timestamp 1683973020
transform -1 0 57600 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _1614_
timestamp 1685175443
transform -1 0 58944 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1615_
timestamp 1683973020
transform 1 0 58944 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1616_
timestamp 1677247768
transform 1 0 63552 0 1 756
box -48 -56 1008 834
use sg13g2_nand2_1  _1617_
timestamp 1676557249
transform 1 0 64512 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _1618_
timestamp 1683973020
transform -1 0 62112 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _1619_
timestamp 1685175443
transform -1 0 63168 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1620_
timestamp 1683973020
transform -1 0 62688 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1621_
timestamp 1677247768
transform 1 0 65376 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1622_
timestamp 1676557249
transform -1 0 66528 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1623_
timestamp 1683973020
transform -1 0 64128 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1624_
timestamp 1685175443
transform -1 0 64704 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1625_
timestamp 1683973020
transform -1 0 64224 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1626_
timestamp 1677247768
transform 1 0 65568 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1627_
timestamp 1676557249
transform -1 0 66528 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1628_
timestamp 1683973020
transform 1 0 65664 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1629_
timestamp 1685175443
transform -1 0 65472 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1630_
timestamp 1683973020
transform 1 0 64512 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1631_
timestamp 1677247768
transform 1 0 64512 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1632_
timestamp 1676557249
transform -1 0 65568 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1633_
timestamp 1683973020
transform 1 0 64704 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1634_
timestamp 1685175443
transform -1 0 64512 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1635_
timestamp 1683973020
transform 1 0 63552 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1636_
timestamp 1677247768
transform -1 0 65088 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1637_
timestamp 1676557249
transform 1 0 64416 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1638_
timestamp 1683973020
transform 1 0 64224 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1639_
timestamp 1685175443
transform 1 0 63744 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1640_
timestamp 1683973020
transform 1 0 64704 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1641_
timestamp 1677247768
transform 1 0 63168 0 -1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1642_
timestamp 1676557249
transform -1 0 64128 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1643_
timestamp 1683973020
transform 1 0 63360 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1644_
timestamp 1685175443
transform 1 0 62688 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1645_
timestamp 1683973020
transform 1 0 63168 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1646_
timestamp 1677247768
transform 1 0 60960 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1647_
timestamp 1676557249
transform 1 0 61728 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1648_
timestamp 1683973020
transform 1 0 61920 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1649_
timestamp 1685175443
transform -1 0 61728 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1650_
timestamp 1683973020
transform -1 0 61248 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1651_
timestamp 1677247768
transform -1 0 65088 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1652_
timestamp 1676557249
transform -1 0 64128 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1653_
timestamp 1683973020
transform -1 0 64224 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1654_
timestamp 1685175443
transform -1 0 65088 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1655_
timestamp 1683973020
transform -1 0 64608 0 1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1656_
timestamp 1677247768
transform 1 0 69504 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1657_
timestamp 1676557249
transform -1 0 70368 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1658_
timestamp 1683973020
transform -1 0 67680 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1659_
timestamp 1685175443
transform -1 0 68928 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1660_
timestamp 1683973020
transform -1 0 68448 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1661_
timestamp 1677247768
transform 1 0 69312 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1662_
timestamp 1676557249
transform -1 0 69984 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1663_
timestamp 1683973020
transform -1 0 69408 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1664_
timestamp 1685175443
transform -1 0 68928 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1665_
timestamp 1683973020
transform 1 0 68832 0 1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1666_
timestamp 1677247768
transform 1 0 69120 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1667_
timestamp 1676557249
transform -1 0 70080 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1668_
timestamp 1683973020
transform 1 0 68832 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1669_
timestamp 1685175443
transform -1 0 68640 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1670_
timestamp 1683973020
transform 1 0 68640 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1671_
timestamp 1677247768
transform 1 0 70656 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1672_
timestamp 1676557249
transform -1 0 71616 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1673_
timestamp 1683973020
transform -1 0 69888 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1674_
timestamp 1685175443
transform -1 0 69984 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1675_
timestamp 1683973020
transform 1 0 69216 0 1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1676_
timestamp 1677247768
transform -1 0 72000 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2_1  _1677_
timestamp 1676557249
transform 1 0 71136 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1678_
timestamp 1683973020
transform 1 0 69984 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1679_
timestamp 1685175443
transform 1 0 69216 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1680_
timestamp 1683973020
transform 1 0 69696 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1681_
timestamp 1677247768
transform 1 0 67776 0 -1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1682_
timestamp 1676557249
transform 1 0 68544 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1683_
timestamp 1683973020
transform 1 0 68832 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1684_
timestamp 1685175443
transform -1 0 68544 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1685_
timestamp 1683973020
transform 1 0 67296 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1686_
timestamp 1677247768
transform 1 0 71040 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1687_
timestamp 1676557249
transform -1 0 71904 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1688_
timestamp 1683973020
transform -1 0 69024 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1689_
timestamp 1685175443
transform -1 0 70176 0 -1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1690_
timestamp 1683973020
transform -1 0 69600 0 -1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1691_
timestamp 1677247768
transform 1 0 72096 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1692_
timestamp 1676557249
transform 1 0 75072 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1693_
timestamp 1683973020
transform -1 0 72480 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1694_
timestamp 1685175443
transform -1 0 72096 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1695_
timestamp 1683973020
transform 1 0 72384 0 1 756
box -48 -56 528 834
use sg13g2_mux2_1  _1696_
timestamp 1677247768
transform 1 0 76608 0 1 2268
box -48 -56 1008 834
use sg13g2_nand2_1  _1697_
timestamp 1676557249
transform 1 0 77568 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1698_
timestamp 1683973020
transform -1 0 74976 0 -1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1699_
timestamp 1685175443
transform -1 0 76320 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _1700_
timestamp 1683973020
transform -1 0 75552 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _1701_
timestamp 1677247768
transform 1 0 76032 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _1702_
timestamp 1676557249
transform 1 0 76896 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1703_
timestamp 1683973020
transform 1 0 76320 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1704_
timestamp 1685175443
transform -1 0 76032 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1705_
timestamp 1683973020
transform 1 0 75072 0 1 3780
box -48 -56 528 834
use sg13g2_mux2_1  _1706_
timestamp 1677247768
transform 1 0 76032 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _1707_
timestamp 1676557249
transform 1 0 76800 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1708_
timestamp 1683973020
transform -1 0 76320 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1709_
timestamp 1685175443
transform -1 0 76032 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1710_
timestamp 1683973020
transform 1 0 76128 0 1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _1711_
timestamp 1677247768
transform 1 0 76032 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _1712_
timestamp 1676557249
transform -1 0 77760 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1713_
timestamp 1683973020
transform 1 0 75840 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1714_
timestamp 1685175443
transform 1 0 75360 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1715_
timestamp 1683973020
transform 1 0 76128 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _1716_
timestamp 1677247768
transform 1 0 76032 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2_1  _1717_
timestamp 1676557249
transform 1 0 76992 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1718_
timestamp 1683973020
transform -1 0 76032 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1719_
timestamp 1685175443
transform -1 0 75936 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1720_
timestamp 1683973020
transform 1 0 75936 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _1721_
timestamp 1677247768
transform 1 0 75168 0 1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _1722_
timestamp 1676557249
transform 1 0 76032 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1723_
timestamp 1683973020
transform 1 0 75552 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1724_
timestamp 1685175443
transform -1 0 75072 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1725_
timestamp 1683973020
transform 1 0 75072 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _1726_
timestamp 1677247768
transform 1 0 75264 0 1 12852
box -48 -56 1008 834
use sg13g2_nand2_1  _1727_
timestamp 1676557249
transform -1 0 76320 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1728_
timestamp 1683973020
transform 1 0 74688 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1729_
timestamp 1685175443
transform -1 0 75264 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1730_
timestamp 1683973020
transform 1 0 74208 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _1731_
timestamp 1677247768
transform 1 0 74496 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _1732_
timestamp 1676557249
transform -1 0 75456 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1733_
timestamp 1683973020
transform 1 0 74688 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1734_
timestamp 1685175443
transform -1 0 74496 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1735_
timestamp 1683973020
transform 1 0 73536 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _1736_
timestamp 1677247768
transform 1 0 75264 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1737_
timestamp 1676557249
transform -1 0 76128 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1738_
timestamp 1683973020
transform 1 0 74208 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1739_
timestamp 1685175443
transform -1 0 75072 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1740_
timestamp 1683973020
transform -1 0 74592 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1741_
timestamp 1677247768
transform 1 0 76032 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1742_
timestamp 1676557249
transform -1 0 77088 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1743_
timestamp 1683973020
transform 1 0 75072 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1744_
timestamp 1685175443
transform -1 0 76032 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1745_
timestamp 1683973020
transform 1 0 74784 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1746_
timestamp 1677247768
transform 1 0 75936 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1747_
timestamp 1676557249
transform -1 0 76800 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1748_
timestamp 1683973020
transform 1 0 75360 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1749_
timestamp 1685175443
transform -1 0 75648 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1750_
timestamp 1683973020
transform 1 0 75168 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1751_
timestamp 1677247768
transform 1 0 76032 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1752_
timestamp 1676557249
transform 1 0 76896 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1753_
timestamp 1683973020
transform 1 0 75648 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1754_
timestamp 1685175443
transform -1 0 75264 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1755_
timestamp 1683973020
transform 1 0 75264 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1756_
timestamp 1677247768
transform 1 0 77280 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1757_
timestamp 1676557249
transform -1 0 78624 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1758_
timestamp 1683973020
transform 1 0 75744 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1759_
timestamp 1685175443
transform -1 0 76608 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1760_
timestamp 1683973020
transform -1 0 76128 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1761_
timestamp 1677247768
transform 1 0 76416 0 1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1762_
timestamp 1676557249
transform -1 0 77376 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1763_
timestamp 1683973020
transform 1 0 76608 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1764_
timestamp 1685175443
transform -1 0 75936 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1765_
timestamp 1683973020
transform 1 0 75936 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1766_
timestamp 1677247768
transform 1 0 76800 0 -1 38556
box -48 -56 1008 834
use sg13g2_nand2_1  _1767_
timestamp 1676557249
transform -1 0 77760 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1768_
timestamp 1683973020
transform 1 0 76128 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1769_
timestamp 1685175443
transform 1 0 74880 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1770_
timestamp 1683973020
transform 1 0 76032 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1771_
timestamp 1677247768
transform 1 0 72672 0 1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1772_
timestamp 1676557249
transform -1 0 73632 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1773_
timestamp 1683973020
transform 1 0 74208 0 1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1774_
timestamp 1685175443
transform 1 0 72768 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1775_
timestamp 1683973020
transform 1 0 73728 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1776_
timestamp 1677247768
transform 1 0 70752 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1777_
timestamp 1676557249
transform 1 0 71424 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1778_
timestamp 1683973020
transform 1 0 71808 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1779_
timestamp 1685175443
transform 1 0 70272 0 -1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1780_
timestamp 1683973020
transform 1 0 71712 0 -1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _1781_
timestamp 1677247768
transform 1 0 68064 0 -1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1782_
timestamp 1676557249
transform 1 0 70944 0 -1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _1783_
timestamp 1683973020
transform 1 0 69600 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1784_
timestamp 1685175443
transform -1 0 68352 0 -1 38556
box -48 -56 538 834
use sg13g2_a21oi_1  _1785_
timestamp 1683973020
transform 1 0 67392 0 -1 38556
box -48 -56 528 834
use sg13g2_mux2_1  _1786_
timestamp 1677247768
transform -1 0 67200 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1787_
timestamp 1676557249
transform -1 0 66240 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1788_
timestamp 1683973020
transform 1 0 67104 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1789_
timestamp 1685175443
transform 1 0 66912 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1790_
timestamp 1683973020
transform 1 0 66432 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1791_
timestamp 1677247768
transform 1 0 65664 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1792_
timestamp 1676557249
transform -1 0 66912 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1793_
timestamp 1683973020
transform 1 0 66048 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1794_
timestamp 1685175443
transform -1 0 66240 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1795_
timestamp 1683973020
transform 1 0 66048 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1796_
timestamp 1677247768
transform 1 0 71520 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1797_
timestamp 1676557249
transform 1 0 72384 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1798_
timestamp 1683973020
transform -1 0 69312 0 1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1799_
timestamp 1685175443
transform -1 0 70656 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1800_
timestamp 1683973020
transform -1 0 70176 0 -1 32508
box -48 -56 528 834
use sg13g2_mux2_1  _1801_
timestamp 1677247768
transform -1 0 71616 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1802_
timestamp 1676557249
transform 1 0 70944 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1803_
timestamp 1683973020
transform 1 0 70656 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1804_
timestamp 1685175443
transform -1 0 71232 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1805_
timestamp 1683973020
transform 1 0 70464 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1806_
timestamp 1677247768
transform 1 0 70176 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1807_
timestamp 1676557249
transform -1 0 70944 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1808_
timestamp 1683973020
transform 1 0 69408 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1809_
timestamp 1685175443
transform -1 0 70752 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1810_
timestamp 1683973020
transform -1 0 70368 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1811_
timestamp 1677247768
transform 1 0 70752 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1812_
timestamp 1676557249
transform 1 0 71712 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1813_
timestamp 1683973020
transform 1 0 69984 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1814_
timestamp 1685175443
transform 1 0 69216 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1815_
timestamp 1683973020
transform 1 0 69504 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1816_
timestamp 1677247768
transform 1 0 66912 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1817_
timestamp 1676557249
transform -1 0 68448 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1818_
timestamp 1683973020
transform 1 0 68256 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1819_
timestamp 1685175443
transform 1 0 67104 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1820_
timestamp 1683973020
transform 1 0 67584 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1821_
timestamp 1677247768
transform 1 0 62976 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1822_
timestamp 1676557249
transform 1 0 64704 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1823_
timestamp 1683973020
transform 1 0 65376 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1824_
timestamp 1685175443
transform 1 0 64128 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1825_
timestamp 1683973020
transform 1 0 64608 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1826_
timestamp 1677247768
transform 1 0 64416 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1827_
timestamp 1676557249
transform -1 0 65280 0 -1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1828_
timestamp 1683973020
transform 1 0 63744 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1829_
timestamp 1685175443
transform 1 0 63744 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1830_
timestamp 1683973020
transform -1 0 64224 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1831_
timestamp 1677247768
transform 1 0 64992 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1832_
timestamp 1676557249
transform -1 0 65952 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1833_
timestamp 1683973020
transform 1 0 63264 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1834_
timestamp 1685175443
transform -1 0 63552 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1835_
timestamp 1683973020
transform 1 0 63552 0 1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1836_
timestamp 1677247768
transform -1 0 63840 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1837_
timestamp 1676557249
transform 1 0 62784 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1838_
timestamp 1683973020
transform 1 0 62976 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1839_
timestamp 1685175443
transform -1 0 62784 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1840_
timestamp 1683973020
transform 1 0 62400 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1841_
timestamp 1677247768
transform -1 0 63360 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1842_
timestamp 1676557249
transform 1 0 62592 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1843_
timestamp 1683973020
transform 1 0 62112 0 -1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1844_
timestamp 1685175443
transform -1 0 61920 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1845_
timestamp 1683973020
transform 1 0 61920 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1846_
timestamp 1677247768
transform 1 0 62784 0 -1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1847_
timestamp 1676557249
transform 1 0 63744 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _1848_
timestamp 1683973020
transform -1 0 62400 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1849_
timestamp 1685175443
transform 1 0 61632 0 -1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1850_
timestamp 1683973020
transform 1 0 62112 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1851_
timestamp 1677247768
transform -1 0 59040 0 -1 37044
box -48 -56 1008 834
use sg13g2_nand2_1  _1852_
timestamp 1676557249
transform 1 0 58464 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1853_
timestamp 1683973020
transform 1 0 60096 0 1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1854_
timestamp 1685175443
transform 1 0 58752 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _1855_
timestamp 1683973020
transform 1 0 59232 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1856_
timestamp 1677247768
transform 1 0 55680 0 1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1857_
timestamp 1676557249
transform -1 0 56832 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1858_
timestamp 1683973020
transform 1 0 57216 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _1859_
timestamp 1685175443
transform -1 0 56448 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _1860_
timestamp 1683973020
transform 1 0 55680 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _1861_
timestamp 1677247768
transform 1 0 58176 0 -1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1862_
timestamp 1676557249
transform 1 0 59136 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1863_
timestamp 1683973020
transform 1 0 57696 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _1864_
timestamp 1685175443
transform -1 0 58752 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1865_
timestamp 1683973020
transform -1 0 57888 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1866_
timestamp 1677247768
transform 1 0 59520 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1867_
timestamp 1676557249
transform 1 0 60672 0 -1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1868_
timestamp 1683973020
transform -1 0 60000 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1869_
timestamp 1685175443
transform 1 0 59520 0 1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1870_
timestamp 1683973020
transform 1 0 60480 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1871_
timestamp 1677247768
transform -1 0 60288 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1872_
timestamp 1676557249
transform 1 0 59616 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1873_
timestamp 1683973020
transform 1 0 59424 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1874_
timestamp 1685175443
transform -1 0 60096 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1875_
timestamp 1683973020
transform 1 0 59136 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1876_
timestamp 1677247768
transform -1 0 60096 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1877_
timestamp 1676557249
transform -1 0 59712 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1878_
timestamp 1683973020
transform 1 0 58752 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1879_
timestamp 1685175443
transform 1 0 57984 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1880_
timestamp 1683973020
transform 1 0 58272 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1881_
timestamp 1677247768
transform 1 0 55296 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1882_
timestamp 1676557249
transform 1 0 56064 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1883_
timestamp 1683973020
transform 1 0 56736 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1884_
timestamp 1685175443
transform 1 0 55584 0 -1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1885_
timestamp 1683973020
transform 1 0 56256 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1886_
timestamp 1677247768
transform -1 0 56160 0 1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1887_
timestamp 1676557249
transform 1 0 55392 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1888_
timestamp 1683973020
transform 1 0 55104 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1889_
timestamp 1685175443
transform -1 0 55968 0 -1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1890_
timestamp 1683973020
transform 1 0 54624 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1891_
timestamp 1677247768
transform 1 0 55008 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1892_
timestamp 1676557249
transform -1 0 55968 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1893_
timestamp 1683973020
transform 1 0 54816 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _1894_
timestamp 1685175443
transform -1 0 55104 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1895_
timestamp 1683973020
transform 1 0 54528 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1896_
timestamp 1677247768
transform 1 0 54144 0 -1 34020
box -48 -56 1008 834
use sg13g2_nand2_1  _1897_
timestamp 1676557249
transform -1 0 55488 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _1898_
timestamp 1683973020
transform 1 0 54144 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _1899_
timestamp 1685175443
transform 1 0 53376 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1900_
timestamp 1683973020
transform 1 0 53760 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1901_
timestamp 1677247768
transform -1 0 52032 0 -1 35532
box -48 -56 1008 834
use sg13g2_nand2_1  _1902_
timestamp 1676557249
transform 1 0 51264 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _1903_
timestamp 1683973020
transform 1 0 52128 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1904_
timestamp 1685175443
transform 1 0 50400 0 1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1905_
timestamp 1683973020
transform 1 0 50880 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1906_
timestamp 1677247768
transform 1 0 46272 0 1 32508
box -48 -56 1008 834
use sg13g2_nand2_1  _1907_
timestamp 1676557249
transform -1 0 48000 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1908_
timestamp 1683973020
transform 1 0 49152 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _1909_
timestamp 1685175443
transform -1 0 47136 0 -1 34020
box -48 -56 538 834
use sg13g2_a21oi_1  _1910_
timestamp 1683973020
transform -1 0 46560 0 1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1911_
timestamp 1677247768
transform -1 0 51072 0 1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1912_
timestamp 1676557249
transform 1 0 50304 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1913_
timestamp 1683973020
transform -1 0 49344 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1914_
timestamp 1685175443
transform -1 0 49056 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1915_
timestamp 1683973020
transform 1 0 49152 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _1916_
timestamp 1677247768
transform 1 0 49920 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1917_
timestamp 1676557249
transform -1 0 50880 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _1918_
timestamp 1683973020
transform 1 0 49632 0 1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1919_
timestamp 1685175443
transform -1 0 50016 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1920_
timestamp 1683973020
transform 1 0 49440 0 -1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1921_
timestamp 1677247768
transform 1 0 51072 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1922_
timestamp 1676557249
transform -1 0 52032 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1923_
timestamp 1683973020
transform 1 0 49344 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1924_
timestamp 1685175443
transform -1 0 50784 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _1925_
timestamp 1683973020
transform -1 0 50304 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1926_
timestamp 1677247768
transform 1 0 51264 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1927_
timestamp 1676557249
transform -1 0 52320 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1928_
timestamp 1683973020
transform 1 0 50016 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1929_
timestamp 1685175443
transform 1 0 50496 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1930_
timestamp 1683973020
transform -1 0 50976 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1931_
timestamp 1677247768
transform 1 0 50208 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1932_
timestamp 1676557249
transform -1 0 51168 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1933_
timestamp 1683973020
transform 1 0 50304 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1934_
timestamp 1685175443
transform 1 0 49728 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1935_
timestamp 1683973020
transform 1 0 50592 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1936_
timestamp 1677247768
transform -1 0 50784 0 -1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _1937_
timestamp 1676557249
transform -1 0 49824 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _1938_
timestamp 1683973020
transform 1 0 49344 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1939_
timestamp 1685175443
transform 1 0 48480 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1940_
timestamp 1683973020
transform 1 0 48768 0 -1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1941_
timestamp 1677247768
transform -1 0 45888 0 -1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _1942_
timestamp 1676557249
transform -1 0 45120 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _1943_
timestamp 1683973020
transform 1 0 46272 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1944_
timestamp 1685175443
transform 1 0 44736 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1945_
timestamp 1683973020
transform 1 0 45120 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1946_
timestamp 1677247768
transform 1 0 44832 0 1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1947_
timestamp 1676557249
transform 1 0 45792 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1948_
timestamp 1683973020
transform 1 0 44544 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1949_
timestamp 1685175443
transform -1 0 44352 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1950_
timestamp 1683973020
transform 1 0 44352 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1951_
timestamp 1677247768
transform 1 0 45984 0 1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1952_
timestamp 1676557249
transform -1 0 46944 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1953_
timestamp 1683973020
transform 1 0 44832 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1954_
timestamp 1685175443
transform -1 0 45696 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1955_
timestamp 1683973020
transform -1 0 45216 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _1956_
timestamp 1677247768
transform -1 0 47040 0 -1 27972
box -48 -56 1008 834
use sg13g2_nand2_1  _1957_
timestamp 1676557249
transform 1 0 46176 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1958_
timestamp 1683973020
transform -1 0 45984 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1959_
timestamp 1685175443
transform 1 0 45024 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1960_
timestamp 1683973020
transform 1 0 45408 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1961_
timestamp 1677247768
transform -1 0 46944 0 1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1962_
timestamp 1676557249
transform 1 0 45888 0 -1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1963_
timestamp 1683973020
transform -1 0 45408 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1964_
timestamp 1685175443
transform 1 0 44544 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _1965_
timestamp 1683973020
transform 1 0 44832 0 -1 29484
box -48 -56 528 834
use sg13g2_mux2_1  _1966_
timestamp 1677247768
transform -1 0 43680 0 1 30996
box -48 -56 1008 834
use sg13g2_nand2_1  _1967_
timestamp 1676557249
transform 1 0 42816 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _1968_
timestamp 1683973020
transform 1 0 43680 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1969_
timestamp 1685175443
transform 1 0 42240 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _1970_
timestamp 1683973020
transform 1 0 42624 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _1971_
timestamp 1677247768
transform 1 0 40896 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2_1  _1972_
timestamp 1676557249
transform -1 0 41664 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _1973_
timestamp 1683973020
transform 1 0 41376 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _1974_
timestamp 1685175443
transform 1 0 40512 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _1975_
timestamp 1683973020
transform 1 0 40800 0 1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1976_
timestamp 1677247768
transform 1 0 40224 0 1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1977_
timestamp 1676557249
transform -1 0 41280 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1978_
timestamp 1683973020
transform 1 0 40128 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _1979_
timestamp 1685175443
transform -1 0 40224 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1980_
timestamp 1683973020
transform 1 0 40224 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _1981_
timestamp 1677247768
transform 1 0 39456 0 -1 24948
box -48 -56 1008 834
use sg13g2_nand2_1  _1982_
timestamp 1676557249
transform -1 0 40416 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1983_
timestamp 1683973020
transform 1 0 39744 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1984_
timestamp 1685175443
transform 1 0 39744 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1985_
timestamp 1683973020
transform 1 0 39264 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1986_
timestamp 1677247768
transform -1 0 41952 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1987_
timestamp 1676557249
transform -1 0 41184 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1988_
timestamp 1683973020
transform 1 0 39168 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1989_
timestamp 1685175443
transform 1 0 38688 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1990_
timestamp 1683973020
transform 1 0 38976 0 1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _1991_
timestamp 1677247768
transform 1 0 36096 0 -1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _1992_
timestamp 1676557249
transform 1 0 37056 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1993_
timestamp 1683973020
transform 1 0 37728 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1994_
timestamp 1685175443
transform 1 0 36000 0 1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1995_
timestamp 1683973020
transform 1 0 36480 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _1996_
timestamp 1677247768
transform 1 0 34752 0 -1 26460
box -48 -56 1008 834
use sg13g2_nand2_1  _1997_
timestamp 1676557249
transform -1 0 35520 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1998_
timestamp 1683973020
transform 1 0 35616 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1999_
timestamp 1685175443
transform 1 0 34368 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _2000_
timestamp 1683973020
transform 1 0 34848 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _2001_
timestamp 1677247768
transform 1 0 31680 0 1 23436
box -48 -56 1008 834
use sg13g2_nand2_1  _2002_
timestamp 1676557249
transform -1 0 32448 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2003_
timestamp 1683973020
transform 1 0 33024 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _2004_
timestamp 1685175443
transform 1 0 31584 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _2005_
timestamp 1683973020
transform 1 0 32064 0 -1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _2006_
timestamp 1677247768
transform 1 0 31008 0 1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _2007_
timestamp 1676557249
transform -1 0 32064 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2008_
timestamp 1683973020
transform 1 0 31200 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _2009_
timestamp 1685175443
transform 1 0 30528 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _2010_
timestamp 1683973020
transform 1 0 30912 0 -1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _2011_
timestamp 1677247768
transform 1 0 28032 0 -1 21924
box -48 -56 1008 834
use sg13g2_nand2_1  _2012_
timestamp 1676557249
transform -1 0 28800 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2013_
timestamp 1683973020
transform 1 0 29472 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _2014_
timestamp 1685175443
transform 1 0 27744 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _2015_
timestamp 1683973020
transform 1 0 28224 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _2016_
timestamp 1677247768
transform 1 0 10464 0 -1 18900
box -48 -56 1008 834
use sg13g2_nand2_1  _2017_
timestamp 1676557249
transform 1 0 11424 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2018_
timestamp 1683973020
transform 1 0 26400 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _2019_
timestamp 1685175443
transform 1 0 10848 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _2020_
timestamp 1683973020
transform 1 0 11328 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _2021_
timestamp 1677247768
transform 1 0 3360 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2_1  _2022_
timestamp 1676557249
transform 1 0 4128 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2023_
timestamp 1683973020
transform 1 0 2784 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _2024_
timestamp 1685175443
transform 1 0 2016 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _2025_
timestamp 1683973020
transform 1 0 2304 0 1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _2026_
timestamp 1677247768
transform -1 0 4704 0 -1 6804
box -48 -56 1008 834
use sg13g2_nand2_1  _2027_
timestamp 1676557249
transform 1 0 3648 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2028_
timestamp 1683973020
transform 1 0 2496 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _2029_
timestamp 1685175443
transform 1 0 1632 0 -1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _2030_
timestamp 1683973020
transform 1 0 2112 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _2031_
timestamp 1677247768
transform 1 0 3168 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _2032_
timestamp 1676557249
transform 1 0 3936 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2033_
timestamp 1683973020
transform 1 0 2592 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _2034_
timestamp 1685175443
transform 1 0 1920 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _2035_
timestamp 1683973020
transform 1 0 2112 0 -1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _2036_
timestamp 1677247768
transform 1 0 2592 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2_1  _2037_
timestamp 1676557249
transform 1 0 3552 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2038_
timestamp 1683973020
transform 1 0 2496 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _2039_
timestamp 1685175443
transform 1 0 1632 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _2040_
timestamp 1683973020
transform 1 0 2112 0 1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _2041_
timestamp 1677247768
transform 1 0 2976 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2_1  _2042_
timestamp 1676557249
transform 1 0 3840 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2043_
timestamp 1683973020
transform 1 0 2496 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _2044_
timestamp 1685175443
transform 1 0 1728 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _2045_
timestamp 1683973020
transform 1 0 2208 0 -1 11340
box -48 -56 528 834
use sg13g2_mux2_1  _2046_
timestamp 1677247768
transform 1 0 3072 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _2047_
timestamp 1676557249
transform 1 0 3936 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2048_
timestamp 1683973020
transform 1 0 2688 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _2049_
timestamp 1685175443
transform 1 0 2016 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _2050_
timestamp 1683973020
transform 1 0 2208 0 -1 12852
box -48 -56 528 834
use sg13g2_mux2_1  _2051_
timestamp 1677247768
transform 1 0 2784 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2_1  _2052_
timestamp 1676557249
transform 1 0 3648 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2053_
timestamp 1683973020
transform -1 0 3072 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _2054_
timestamp 1685175443
transform 1 0 2304 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _2055_
timestamp 1683973020
transform 1 0 2688 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2056_
timestamp 1676557249
transform 1 0 23520 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2057_
timestamp 1683973020
transform -1 0 23328 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2058_
timestamp 1676557249
transform -1 0 27552 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2059_
timestamp 1683973020
transform 1 0 26592 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2060_
timestamp 1676557249
transform -1 0 30720 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2061_
timestamp 1683973020
transform 1 0 29760 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2062_
timestamp 1676557249
transform -1 0 33600 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2063_
timestamp 1683973020
transform 1 0 32352 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2064_
timestamp 1676557249
transform -1 0 36768 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2065_
timestamp 1683973020
transform 1 0 35616 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2066_
timestamp 1676557249
transform -1 0 38976 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _2067_
timestamp 1683973020
transform 1 0 38496 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2068_
timestamp 1676557249
transform -1 0 44736 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2069_
timestamp 1683973020
transform 1 0 43872 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2070_
timestamp 1676557249
transform -1 0 43296 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2071_
timestamp 1683973020
transform 1 0 42528 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2072_
timestamp 1676557249
transform -1 0 43488 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2073_
timestamp 1683973020
transform 1 0 42624 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2074_
timestamp 1676557249
transform 1 0 39744 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2075_
timestamp 1683973020
transform 1 0 40320 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2076_
timestamp 1676557249
transform -1 0 37248 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2077_
timestamp 1683973020
transform -1 0 38112 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2078_
timestamp 1676557249
transform -1 0 33696 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2079_
timestamp 1683973020
transform -1 0 34176 0 -1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2080_
timestamp 1676557249
transform -1 0 32352 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2081_
timestamp 1683973020
transform 1 0 31488 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2082_
timestamp 1676557249
transform -1 0 36864 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2083_
timestamp 1683973020
transform -1 0 36960 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2084_
timestamp 1676557249
transform -1 0 39648 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2085_
timestamp 1683973020
transform 1 0 38784 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2086_
timestamp 1676557249
transform -1 0 42720 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2087_
timestamp 1683973020
transform -1 0 42336 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2088_
timestamp 1676557249
transform 1 0 43872 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2089_
timestamp 1683973020
transform -1 0 44928 0 1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2090_
timestamp 1676557249
transform -1 0 47232 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2091_
timestamp 1683973020
transform 1 0 46272 0 1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2092_
timestamp 1676557249
transform 1 0 48768 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2093_
timestamp 1683973020
transform 1 0 48768 0 1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2094_
timestamp 1676557249
transform -1 0 50208 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2095_
timestamp 1683973020
transform 1 0 48960 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2096_
timestamp 1676557249
transform -1 0 52896 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2097_
timestamp 1683973020
transform -1 0 51936 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2098_
timestamp 1676557249
transform 1 0 54624 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2099_
timestamp 1683973020
transform 1 0 54048 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2100_
timestamp 1676557249
transform 1 0 54048 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2101_
timestamp 1683973020
transform 1 0 53856 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2102_
timestamp 1676557249
transform 1 0 52992 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2103_
timestamp 1683973020
transform -1 0 53856 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2104_
timestamp 1676557249
transform 1 0 51840 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2105_
timestamp 1683973020
transform 1 0 51648 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2106_
timestamp 1676557249
transform -1 0 49632 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2107_
timestamp 1683973020
transform 1 0 48768 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2108_
timestamp 1676557249
transform -1 0 48192 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2109_
timestamp 1683973020
transform 1 0 47520 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2110_
timestamp 1676557249
transform 1 0 45696 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2111_
timestamp 1683973020
transform -1 0 46368 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2112_
timestamp 1676557249
transform 1 0 49056 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _2113_
timestamp 1683973020
transform 1 0 48864 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2114_
timestamp 1676557249
transform 1 0 49344 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2115_
timestamp 1683973020
transform -1 0 50208 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _2116_
timestamp 1676557249
transform -1 0 53856 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2117_
timestamp 1683973020
transform 1 0 52992 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2118_
timestamp 1676557249
transform -1 0 57696 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2119_
timestamp 1683973020
transform 1 0 56832 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2120_
timestamp 1676557249
transform -1 0 58080 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2121_
timestamp 1683973020
transform -1 0 59040 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2122_
timestamp 1676557249
transform -1 0 59616 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2123_
timestamp 1683973020
transform 1 0 58752 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2124_
timestamp 1676557249
transform -1 0 59808 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2125_
timestamp 1683973020
transform 1 0 58944 0 1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2126_
timestamp 1676557249
transform -1 0 60768 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2127_
timestamp 1683973020
transform -1 0 60960 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2128_
timestamp 1676557249
transform -1 0 61728 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2129_
timestamp 1683973020
transform 1 0 60768 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2130_
timestamp 1676557249
transform -1 0 56544 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2131_
timestamp 1683973020
transform 1 0 55584 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2132_
timestamp 1676557249
transform -1 0 57024 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2133_
timestamp 1683973020
transform 1 0 56160 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2134_
timestamp 1676557249
transform -1 0 59616 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2135_
timestamp 1683973020
transform -1 0 59232 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2136_
timestamp 1676557249
transform -1 0 64992 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2137_
timestamp 1683973020
transform 1 0 64128 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2138_
timestamp 1676557249
transform -1 0 66912 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2139_
timestamp 1683973020
transform 1 0 66048 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2140_
timestamp 1676557249
transform -1 0 67008 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2141_
timestamp 1683973020
transform 1 0 66336 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2142_
timestamp 1676557249
transform -1 0 66336 0 -1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _2143_
timestamp 1683973020
transform 1 0 65472 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2144_
timestamp 1676557249
transform -1 0 65568 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2145_
timestamp 1683973020
transform 1 0 64800 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2146_
timestamp 1676557249
transform 1 0 64320 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2147_
timestamp 1683973020
transform 1 0 64128 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2148_
timestamp 1676557249
transform -1 0 62688 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2149_
timestamp 1683973020
transform 1 0 60480 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2150_
timestamp 1676557249
transform 1 0 64800 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2151_
timestamp 1683973020
transform -1 0 65568 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2152_
timestamp 1676557249
transform -1 0 71232 0 -1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _2153_
timestamp 1683973020
transform -1 0 70464 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _2154_
timestamp 1676557249
transform -1 0 70752 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2155_
timestamp 1683973020
transform -1 0 70368 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2156_
timestamp 1676557249
transform -1 0 71136 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2157_
timestamp 1683973020
transform 1 0 69888 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2158_
timestamp 1676557249
transform -1 0 72000 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2159_
timestamp 1683973020
transform 1 0 71328 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2160_
timestamp 1676557249
transform -1 0 72384 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2161_
timestamp 1683973020
transform 1 0 71520 0 1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _2162_
timestamp 1676557249
transform -1 0 69312 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2163_
timestamp 1683973020
transform -1 0 69024 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _2164_
timestamp 1676557249
transform -1 0 72384 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2165_
timestamp 1683973020
transform 1 0 71520 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2166_
timestamp 1676557249
transform 1 0 74304 0 1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2167_
timestamp 1683973020
transform 1 0 73920 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2168_
timestamp 1676557249
transform -1 0 79008 0 -1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _2169_
timestamp 1683973020
transform 1 0 78144 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _2170_
timestamp 1676557249
transform -1 0 77760 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2171_
timestamp 1683973020
transform 1 0 77088 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2172_
timestamp 1676557249
transform -1 0 77856 0 1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _2173_
timestamp 1683973020
transform 1 0 76992 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _2174_
timestamp 1676557249
transform -1 0 77664 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2175_
timestamp 1683973020
transform 1 0 76896 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2176_
timestamp 1676557249
transform -1 0 77856 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2177_
timestamp 1683973020
transform 1 0 76992 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2178_
timestamp 1676557249
transform -1 0 77280 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2179_
timestamp 1683973020
transform 1 0 76416 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2180_
timestamp 1676557249
transform -1 0 77280 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2181_
timestamp 1683973020
transform 1 0 76416 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _2182_
timestamp 1676557249
transform -1 0 76128 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _2183_
timestamp 1683973020
transform 1 0 75456 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2184_
timestamp 1676557249
transform -1 0 76704 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2185_
timestamp 1683973020
transform -1 0 76608 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2186_
timestamp 1676557249
transform -1 0 77472 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2187_
timestamp 1683973020
transform 1 0 76800 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2188_
timestamp 1676557249
transform -1 0 77472 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2189_
timestamp 1683973020
transform 1 0 76608 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2190_
timestamp 1676557249
transform -1 0 77760 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2191_
timestamp 1683973020
transform 1 0 76992 0 1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2192_
timestamp 1676557249
transform -1 0 78144 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2193_
timestamp 1683973020
transform 1 0 77184 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2194_
timestamp 1676557249
transform -1 0 78240 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2195_
timestamp 1683973020
transform 1 0 77376 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2196_
timestamp 1676557249
transform -1 0 78336 0 1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2197_
timestamp 1683973020
transform 1 0 76512 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2198_
timestamp 1676557249
transform -1 0 74016 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2199_
timestamp 1683973020
transform 1 0 73248 0 1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2200_
timestamp 1676557249
transform -1 0 71904 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2201_
timestamp 1683973020
transform -1 0 72000 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2202_
timestamp 1676557249
transform 1 0 69504 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2203_
timestamp 1683973020
transform 1 0 69024 0 -1 37044
box -48 -56 528 834
use sg13g2_nand2_1  _2204_
timestamp 1676557249
transform -1 0 67680 0 1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2205_
timestamp 1683973020
transform 1 0 66816 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2206_
timestamp 1676557249
transform -1 0 67104 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2207_
timestamp 1683973020
transform 1 0 66240 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2208_
timestamp 1676557249
transform -1 0 72864 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2209_
timestamp 1683973020
transform 1 0 71904 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2210_
timestamp 1676557249
transform -1 0 72384 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _2211_
timestamp 1683973020
transform 1 0 71328 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2212_
timestamp 1676557249
transform -1 0 71616 0 -1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _2213_
timestamp 1683973020
transform 1 0 70944 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2214_
timestamp 1676557249
transform -1 0 71520 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2215_
timestamp 1683973020
transform 1 0 70656 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2216_
timestamp 1676557249
transform -1 0 68448 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2217_
timestamp 1683973020
transform 1 0 67584 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2218_
timestamp 1676557249
transform -1 0 64704 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2219_
timestamp 1683973020
transform 1 0 63840 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2220_
timestamp 1676557249
transform -1 0 65952 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2221_
timestamp 1683973020
transform 1 0 65088 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2222_
timestamp 1676557249
transform -1 0 66336 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2223_
timestamp 1683973020
transform 1 0 65568 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2224_
timestamp 1676557249
transform -1 0 64704 0 -1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2225_
timestamp 1683973020
transform 1 0 63840 0 -1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2226_
timestamp 1676557249
transform -1 0 63360 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2227_
timestamp 1683973020
transform 1 0 62592 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _2228_
timestamp 1676557249
transform -1 0 64512 0 -1 37044
box -48 -56 432 834
use sg13g2_a21oi_1  _2229_
timestamp 1683973020
transform 1 0 63264 0 -1 38556
box -48 -56 528 834
use sg13g2_nand2_1  _2230_
timestamp 1676557249
transform -1 0 59712 0 1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2231_
timestamp 1683973020
transform 1 0 58848 0 1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _2232_
timestamp 1676557249
transform -1 0 55104 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2233_
timestamp 1683973020
transform -1 0 55968 0 1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _2234_
timestamp 1676557249
transform -1 0 59136 0 -1 34020
box -48 -56 432 834
use sg13g2_a21oi_1  _2235_
timestamp 1683973020
transform 1 0 57984 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2236_
timestamp 1676557249
transform -1 0 61344 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2237_
timestamp 1683973020
transform -1 0 60672 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2238_
timestamp 1676557249
transform -1 0 60864 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2239_
timestamp 1683973020
transform 1 0 60000 0 1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2240_
timestamp 1676557249
transform -1 0 60480 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2241_
timestamp 1683973020
transform -1 0 60192 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2242_
timestamp 1676557249
transform -1 0 55968 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2243_
timestamp 1683973020
transform 1 0 55200 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2244_
timestamp 1676557249
transform -1 0 56544 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2245_
timestamp 1683973020
transform 1 0 55776 0 1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2246_
timestamp 1676557249
transform -1 0 56352 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2247_
timestamp 1683973020
transform 1 0 55584 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2248_
timestamp 1676557249
transform -1 0 54720 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2249_
timestamp 1683973020
transform -1 0 55200 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2250_
timestamp 1676557249
transform -1 0 52896 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _2251_
timestamp 1683973020
transform 1 0 52032 0 -1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _2252_
timestamp 1676557249
transform -1 0 46944 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2253_
timestamp 1683973020
transform 1 0 45792 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _2254_
timestamp 1676557249
transform 1 0 50976 0 1 32508
box -48 -56 432 834
use sg13g2_a21oi_1  _2255_
timestamp 1683973020
transform -1 0 51552 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2256_
timestamp 1676557249
transform 1 0 50880 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2257_
timestamp 1683973020
transform -1 0 51168 0 1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2258_
timestamp 1676557249
transform -1 0 52416 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2259_
timestamp 1683973020
transform 1 0 51552 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2260_
timestamp 1676557249
transform -1 0 52704 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2261_
timestamp 1683973020
transform 1 0 52032 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2262_
timestamp 1676557249
transform -1 0 51552 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2263_
timestamp 1683973020
transform -1 0 51552 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2264_
timestamp 1676557249
transform 1 0 50496 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2265_
timestamp 1683973020
transform -1 0 51264 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2266_
timestamp 1676557249
transform 1 0 45600 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2267_
timestamp 1683973020
transform 1 0 45408 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _2268_
timestamp 1676557249
transform 1 0 45408 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _2269_
timestamp 1683973020
transform -1 0 46272 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2270_
timestamp 1676557249
transform -1 0 48288 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2271_
timestamp 1683973020
transform 1 0 46656 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2272_
timestamp 1676557249
transform -1 0 47904 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2273_
timestamp 1683973020
transform 1 0 47040 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _2274_
timestamp 1676557249
transform -1 0 47328 0 1 29484
box -48 -56 432 834
use sg13g2_a21oi_1  _2275_
timestamp 1683973020
transform 1 0 45984 0 -1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2276_
timestamp 1676557249
transform 1 0 43104 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _2277_
timestamp 1683973020
transform -1 0 44160 0 1 30996
box -48 -56 528 834
use sg13g2_nand2_1  _2278_
timestamp 1676557249
transform 1 0 41280 0 1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _2279_
timestamp 1683973020
transform -1 0 42336 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2_1  _2280_
timestamp 1676557249
transform -1 0 41568 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2281_
timestamp 1683973020
transform -1 0 41568 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2282_
timestamp 1676557249
transform -1 0 41280 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2283_
timestamp 1683973020
transform 1 0 40416 0 -1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _2284_
timestamp 1676557249
transform -1 0 41472 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2285_
timestamp 1683973020
transform -1 0 41088 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2286_
timestamp 1676557249
transform -1 0 36864 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2287_
timestamp 1683973020
transform 1 0 36000 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2288_
timestamp 1676557249
transform -1 0 36576 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2289_
timestamp 1683973020
transform 1 0 35712 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _2290_
timestamp 1676557249
transform 1 0 32640 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _2291_
timestamp 1683973020
transform 1 0 32448 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _2292_
timestamp 1676557249
transform 1 0 32256 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2293_
timestamp 1683973020
transform 1 0 32064 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _2294_
timestamp 1676557249
transform -1 0 29184 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2295_
timestamp 1683973020
transform -1 0 29184 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _2296_
timestamp 1676557249
transform -1 0 12384 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _2297_
timestamp 1683973020
transform 1 0 11712 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _2298_
timestamp 1676557249
transform -1 0 5376 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _2299_
timestamp 1683973020
transform 1 0 4512 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2300_
timestamp 1676557249
transform -1 0 5184 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2301_
timestamp 1683973020
transform 1 0 4512 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _2302_
timestamp 1676557249
transform -1 0 5088 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _2303_
timestamp 1683973020
transform 1 0 4224 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _2304_
timestamp 1676557249
transform -1 0 5184 0 -1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _2305_
timestamp 1683973020
transform 1 0 4320 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _2306_
timestamp 1676557249
transform -1 0 5184 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _2307_
timestamp 1683973020
transform 1 0 4416 0 1 11340
box -48 -56 528 834
use sg13g2_nand2_1  _2308_
timestamp 1676557249
transform 1 0 4128 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _2309_
timestamp 1683973020
transform -1 0 4800 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _2310_
timestamp 1676557249
transform 1 0 4128 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _2311_
timestamp 1683973020
transform -1 0 4704 0 -1 15876
box -48 -56 528 834
use sg13g2_tiehi  _2312__328
timestamp 1680000651
transform -1 0 23424 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2312_
timestamp 1746535128
transform 1 0 22560 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2313__327
timestamp 1680000651
transform -1 0 27264 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2313_
timestamp 1746535128
transform 1 0 26112 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2314__325
timestamp 1680000651
transform 1 0 29472 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2314_
timestamp 1746535128
transform 1 0 29184 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2315__323
timestamp 1680000651
transform -1 0 33024 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2315_
timestamp 1746535128
transform 1 0 32160 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2316__321
timestamp 1680000651
transform -1 0 36000 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2316_
timestamp 1746535128
transform 1 0 35232 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2317__319
timestamp 1680000651
transform -1 0 39744 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2317_
timestamp 1746535128
transform 1 0 38592 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2318__317
timestamp 1680000651
transform -1 0 42240 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2318_
timestamp 1746535128
transform 1 0 41376 0 -1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2319__315
timestamp 1680000651
transform 1 0 38112 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2319_
timestamp 1746535128
transform 1 0 39744 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2320_
timestamp 1746535128
transform 1 0 40224 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2320__313
timestamp 1680000651
transform -1 0 41088 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2321__311
timestamp 1680000651
transform 1 0 37824 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2321_
timestamp 1746535128
transform -1 0 39936 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2322__309
timestamp 1680000651
transform 1 0 35424 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2322_
timestamp 1746535128
transform -1 0 37344 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2323__307
timestamp 1680000651
transform -1 0 31872 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2323_
timestamp 1746535128
transform 1 0 31008 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2324_
timestamp 1746535128
transform 1 0 33024 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2324__305
timestamp 1680000651
transform -1 0 33888 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2325_
timestamp 1746535128
transform 1 0 33792 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2325__303
timestamp 1680000651
transform -1 0 34656 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2326__301
timestamp 1680000651
transform -1 0 37344 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2326_
timestamp 1746535128
transform 1 0 36384 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2327__299
timestamp 1680000651
transform -1 0 40320 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2327_
timestamp 1746535128
transform 1 0 39360 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2328__297
timestamp 1680000651
transform 1 0 41280 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2328_
timestamp 1746535128
transform 1 0 41472 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2329__295
timestamp 1680000651
transform -1 0 44928 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2329_
timestamp 1746535128
transform 1 0 44064 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2330__293
timestamp 1680000651
transform -1 0 46272 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2330_
timestamp 1746535128
transform 1 0 45312 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2331__291
timestamp 1680000651
transform -1 0 46656 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2331_
timestamp 1746535128
transform 1 0 45792 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2332__289
timestamp 1680000651
transform -1 0 50496 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2332_
timestamp 1746535128
transform 1 0 49536 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2333__287
timestamp 1680000651
transform -1 0 52224 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2333_
timestamp 1746535128
transform 1 0 51360 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2334__285
timestamp 1680000651
transform -1 0 51264 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2334_
timestamp 1746535128
transform 1 0 50400 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2335_
timestamp 1746535128
transform 1 0 49728 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2335__283
timestamp 1680000651
transform -1 0 50688 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2336_
timestamp 1746535128
transform -1 0 50688 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2336__281
timestamp 1680000651
transform 1 0 48672 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2337_
timestamp 1746535128
transform 1 0 45216 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2337__279
timestamp 1680000651
transform -1 0 46080 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2338__277
timestamp 1680000651
transform -1 0 45408 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2338_
timestamp 1746535128
transform 1 0 44544 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2339__275
timestamp 1680000651
transform -1 0 44160 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2339_
timestamp 1746535128
transform 1 0 43296 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2340__273
timestamp 1680000651
transform -1 0 47040 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2340_
timestamp 1746535128
transform 1 0 46176 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2341__271
timestamp 1680000651
transform -1 0 49440 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2341_
timestamp 1746535128
transform 1 0 48576 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2342_
timestamp 1746535128
transform 1 0 50688 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2342__269
timestamp 1680000651
transform -1 0 51936 0 -1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2343__267
timestamp 1680000651
transform -1 0 54624 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2343_
timestamp 1746535128
transform 1 0 53664 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2344_
timestamp 1746535128
transform 1 0 54720 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2344__265
timestamp 1680000651
transform -1 0 55584 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2345__263
timestamp 1680000651
transform 1 0 56064 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2345_
timestamp 1746535128
transform 1 0 56448 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2346__261
timestamp 1680000651
transform -1 0 56736 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2346_
timestamp 1746535128
transform 1 0 55872 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2347_
timestamp 1746535128
transform 1 0 56832 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2347__259
timestamp 1680000651
transform -1 0 57696 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2348__257
timestamp 1680000651
transform -1 0 60000 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2348_
timestamp 1746535128
transform 1 0 58848 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2349__255
timestamp 1680000651
transform 1 0 54912 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2349_
timestamp 1746535128
transform -1 0 56448 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2350__253
timestamp 1680000651
transform -1 0 54336 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2350_
timestamp 1746535128
transform 1 0 53472 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2351__251
timestamp 1680000651
transform -1 0 61056 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2351_
timestamp 1746535128
transform 1 0 59040 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2352__249
timestamp 1680000651
transform -1 0 62496 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2352_
timestamp 1746535128
transform 1 0 61632 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2353_
timestamp 1746535128
transform 1 0 62784 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2353__247
timestamp 1680000651
transform -1 0 63648 0 -1 3780
box -48 -56 432 834
use sg13g2_tiehi  _2354__245
timestamp 1680000651
transform -1 0 63936 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2354_
timestamp 1746535128
transform 1 0 63072 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2355__243
timestamp 1680000651
transform -1 0 63360 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2355_
timestamp 1746535128
transform 1 0 62112 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2356__241
timestamp 1680000651
transform 1 0 62112 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2356_
timestamp 1746535128
transform 1 0 62112 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2357__239
timestamp 1680000651
transform 1 0 61824 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2357_
timestamp 1746535128
transform -1 0 63456 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2358_
timestamp 1746535128
transform 1 0 61152 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2358__237
timestamp 1680000651
transform -1 0 62496 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2359_
timestamp 1746535128
transform 1 0 64512 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2359__235
timestamp 1680000651
transform -1 0 65472 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2360__233
timestamp 1680000651
transform -1 0 68352 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2360_
timestamp 1746535128
transform 1 0 67488 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2361_
timestamp 1746535128
transform 1 0 67296 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2361__231
timestamp 1680000651
transform 1 0 67200 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2362__229
timestamp 1680000651
transform -1 0 68160 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2362_
timestamp 1746535128
transform 1 0 66816 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2363__227
timestamp 1680000651
transform -1 0 70464 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2363_
timestamp 1746535128
transform 1 0 68256 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2364__225
timestamp 1680000651
transform 1 0 69120 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2364_
timestamp 1746535128
transform 1 0 69216 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2365__223
timestamp 1680000651
transform -1 0 66816 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2365_
timestamp 1746535128
transform 1 0 65952 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2366__221
timestamp 1680000651
transform -1 0 69696 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2366_
timestamp 1746535128
transform 1 0 68928 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2367__219
timestamp 1680000651
transform 1 0 71232 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2367_
timestamp 1746535128
transform 1 0 71328 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2368__217
timestamp 1680000651
transform -1 0 76416 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2368_
timestamp 1746535128
transform 1 0 75552 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2369__215
timestamp 1680000651
transform -1 0 74592 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2369_
timestamp 1746535128
transform 1 0 73728 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2370__213
timestamp 1680000651
transform -1 0 74784 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2370_
timestamp 1746535128
transform 1 0 73536 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2371__211
timestamp 1680000651
transform -1 0 74592 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2371_
timestamp 1746535128
transform 1 0 73536 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2372_
timestamp 1746535128
transform 1 0 73440 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2372__209
timestamp 1680000651
transform -1 0 74304 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2373__207
timestamp 1680000651
transform -1 0 73344 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2373_
timestamp 1746535128
transform 1 0 72480 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2374__205
timestamp 1680000651
transform 1 0 71808 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2374_
timestamp 1746535128
transform 1 0 72192 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2375__203
timestamp 1680000651
transform -1 0 72960 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2375_
timestamp 1746535128
transform 1 0 72096 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2376__457
timestamp 1680000651
transform 1 0 73152 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2376_
timestamp 1746535128
transform 1 0 73152 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2377__455
timestamp 1680000651
transform -1 0 73824 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2377_
timestamp 1746535128
transform 1 0 72960 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2378__453
timestamp 1680000651
transform -1 0 74208 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2378_
timestamp 1746535128
transform 1 0 73344 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2379__451
timestamp 1680000651
transform -1 0 74400 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2379_
timestamp 1746535128
transform 1 0 73536 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2380__449
timestamp 1680000651
transform 1 0 74880 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2380_
timestamp 1746535128
transform 1 0 74688 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2381_
timestamp 1746535128
transform 1 0 74112 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2381__447
timestamp 1680000651
transform -1 0 74976 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  _2382__445
timestamp 1680000651
transform -1 0 76224 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2382_
timestamp 1746535128
transform 1 0 75360 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2383__443
timestamp 1680000651
transform 1 0 71712 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2383_
timestamp 1746535128
transform -1 0 73440 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2384__441
timestamp 1680000651
transform 1 0 69216 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2384_
timestamp 1746535128
transform -1 0 71328 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2385__439
timestamp 1680000651
transform 1 0 66240 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2385_
timestamp 1746535128
transform 1 0 66240 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2386_
timestamp 1746535128
transform 1 0 64320 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2386__437
timestamp 1680000651
transform -1 0 65184 0 -1 35532
box -48 -56 432 834
use sg13g2_tiehi  _2387__435
timestamp 1680000651
transform -1 0 67296 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2387_
timestamp 1746535128
transform 1 0 66240 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2388__433
timestamp 1680000651
transform -1 0 70176 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2388_
timestamp 1746535128
transform 1 0 69312 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2389__431
timestamp 1680000651
transform -1 0 69024 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2389_
timestamp 1746535128
transform 1 0 68160 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2390_
timestamp 1746535128
transform 1 0 67680 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2390__429
timestamp 1680000651
transform -1 0 68640 0 1 27972
box -48 -56 432 834
use sg13g2_tiehi  _2391__427
timestamp 1680000651
transform 1 0 69120 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2391_
timestamp 1746535128
transform 1 0 69024 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2392_
timestamp 1746535128
transform -1 0 68256 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2392__425
timestamp 1680000651
transform 1 0 66144 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2393__423
timestamp 1680000651
transform -1 0 62400 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2393_
timestamp 1746535128
transform 1 0 61536 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2394__421
timestamp 1680000651
transform -1 0 62688 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2394_
timestamp 1746535128
transform 1 0 61824 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2395__419
timestamp 1680000651
transform -1 0 63840 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2395_
timestamp 1746535128
transform 1 0 62976 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2396__417
timestamp 1680000651
transform -1 0 61440 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2396_
timestamp 1746535128
transform 1 0 60288 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2397__415
timestamp 1680000651
transform -1 0 60672 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2397_
timestamp 1746535128
transform 1 0 59808 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2398__413
timestamp 1680000651
transform -1 0 61920 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2398_
timestamp 1746535128
transform 1 0 61056 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2399__411
timestamp 1680000651
transform 1 0 56640 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2399_
timestamp 1746535128
transform -1 0 58752 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2400__409
timestamp 1680000651
transform -1 0 55488 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2400_
timestamp 1746535128
transform 1 0 54624 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2401__407
timestamp 1680000651
transform -1 0 58752 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2401_
timestamp 1746535128
transform 1 0 57888 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2402_
timestamp 1746535128
transform -1 0 60480 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2402__405
timestamp 1680000651
transform 1 0 58368 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2403_
timestamp 1746535128
transform 1 0 57024 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2403__403
timestamp 1680000651
transform -1 0 57888 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2404_
timestamp 1746535128
transform 1 0 57312 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2404__401
timestamp 1680000651
transform -1 0 58176 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2405_
timestamp 1746535128
transform -1 0 56736 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2405__399
timestamp 1680000651
transform 1 0 54624 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2406_
timestamp 1746535128
transform 1 0 52896 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2406__397
timestamp 1680000651
transform -1 0 53760 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2407__395
timestamp 1680000651
transform -1 0 53664 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2407_
timestamp 1746535128
transform 1 0 52800 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2408__393
timestamp 1680000651
transform 1 0 51744 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2408_
timestamp 1746535128
transform 1 0 51552 0 -1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2409__391
timestamp 1680000651
transform 1 0 48960 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2409_
timestamp 1746535128
transform -1 0 51072 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2410__389
timestamp 1680000651
transform -1 0 47424 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2410_
timestamp 1746535128
transform 1 0 46560 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2411__387
timestamp 1680000651
transform -1 0 49152 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2411_
timestamp 1746535128
transform 1 0 48384 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2412__385
timestamp 1680000651
transform -1 0 48576 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2412_
timestamp 1746535128
transform 1 0 47712 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2413__383
timestamp 1680000651
transform 1 0 48960 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2413_
timestamp 1746535128
transform 1 0 48768 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2414__381
timestamp 1680000651
transform 1 0 48288 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2414_
timestamp 1746535128
transform 1 0 48672 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2415__379
timestamp 1680000651
transform -1 0 48864 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2415_
timestamp 1746535128
transform 1 0 48000 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2416__377
timestamp 1680000651
transform -1 0 48480 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2416_
timestamp 1746535128
transform 1 0 47616 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2417__375
timestamp 1680000651
transform -1 0 43200 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2417_
timestamp 1746535128
transform 1 0 42336 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2418_
timestamp 1746535128
transform 1 0 42240 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2418__373
timestamp 1680000651
transform -1 0 43104 0 1 23436
box -48 -56 432 834
use sg13g2_tiehi  _2419__371
timestamp 1680000651
transform -1 0 44448 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2419_
timestamp 1746535128
transform 1 0 43584 0 -1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2420__369
timestamp 1680000651
transform -1 0 44640 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2420_
timestamp 1746535128
transform 1 0 43488 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2421__367
timestamp 1680000651
transform -1 0 44544 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2421_
timestamp 1746535128
transform 1 0 43392 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2422__365
timestamp 1680000651
transform -1 0 40992 0 -1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2422_
timestamp 1746535128
transform 1 0 40128 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2423__363
timestamp 1680000651
transform -1 0 39168 0 1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2423_
timestamp 1746535128
transform 1 0 38304 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2424__361
timestamp 1680000651
transform -1 0 38496 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2424_
timestamp 1746535128
transform 1 0 37632 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2425_
timestamp 1746535128
transform 1 0 37152 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2425__359
timestamp 1680000651
transform -1 0 38016 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2426_
timestamp 1746535128
transform 1 0 38400 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2426__357
timestamp 1680000651
transform 1 0 38592 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2427_
timestamp 1746535128
transform 1 0 34848 0 -1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2427__355
timestamp 1680000651
transform -1 0 35808 0 1 23436
box -48 -56 432 834
use sg13g2_tiehi  _2428__353
timestamp 1680000651
transform 1 0 32736 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2428_
timestamp 1746535128
transform -1 0 34752 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2429_
timestamp 1746535128
transform 1 0 29664 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2429__351
timestamp 1680000651
transform -1 0 30528 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2430__349
timestamp 1680000651
transform -1 0 29184 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2430_
timestamp 1746535128
transform 1 0 28320 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2431__347
timestamp 1680000651
transform 1 0 25920 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2431_
timestamp 1746535128
transform -1 0 28032 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2432__345
timestamp 1680000651
transform 1 0 9312 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2432_
timestamp 1746535128
transform -1 0 11424 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2433__343
timestamp 1680000651
transform 1 0 1632 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2433_
timestamp 1746535128
transform 1 0 1344 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2434_
timestamp 1746535128
transform 1 0 1152 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2434__341
timestamp 1680000651
transform -1 0 2016 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2435__339
timestamp 1680000651
transform 1 0 1056 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2435_
timestamp 1746535128
transform 1 0 1248 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2436_
timestamp 1746535128
transform 1 0 960 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2436__337
timestamp 1680000651
transform 1 0 1248 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2437__335
timestamp 1680000651
transform -1 0 2208 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2437_
timestamp 1746535128
transform 1 0 1248 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2438__333
timestamp 1680000651
transform 1 0 1632 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2438_
timestamp 1746535128
transform 1 0 1344 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2439_
timestamp 1746535128
transform -1 0 3648 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2439__331
timestamp 1680000651
transform 1 0 1536 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2440_
timestamp 1746535128
transform 1 0 23328 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2440__329
timestamp 1680000651
transform -1 0 24288 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2441_
timestamp 1746535128
transform 1 0 27072 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2441__326
timestamp 1680000651
transform -1 0 27936 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2442_
timestamp 1746535128
transform 1 0 30240 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2442__322
timestamp 1680000651
transform -1 0 31104 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2443__318
timestamp 1680000651
transform -1 0 33696 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2443_
timestamp 1746535128
transform 1 0 32832 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2444__314
timestamp 1680000651
transform -1 0 37344 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2444_
timestamp 1746535128
transform 1 0 36096 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2445_
timestamp 1746535128
transform 1 0 38688 0 -1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2445__310
timestamp 1680000651
transform -1 0 39744 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2446__306
timestamp 1680000651
transform -1 0 45024 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2446_
timestamp 1746535128
transform 1 0 43584 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2447_
timestamp 1746535128
transform 1 0 43008 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2447__302
timestamp 1680000651
transform -1 0 43872 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2448__298
timestamp 1680000651
transform -1 0 44160 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2448_
timestamp 1746535128
transform 1 0 43008 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2449_
timestamp 1746535128
transform 1 0 40128 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2449__294
timestamp 1680000651
transform -1 0 41184 0 -1 15876
box -48 -56 432 834
use sg13g2_tiehi  _2450__290
timestamp 1680000651
transform -1 0 38208 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2450_
timestamp 1746535128
transform 1 0 37248 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2451__286
timestamp 1680000651
transform -1 0 35136 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2451_
timestamp 1746535128
transform 1 0 34176 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2452_
timestamp 1746535128
transform 1 0 30144 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2452__282
timestamp 1680000651
transform -1 0 31008 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2453_
timestamp 1746535128
transform 1 0 36864 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2453__278
timestamp 1680000651
transform -1 0 37728 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2454_
timestamp 1746535128
transform 1 0 39072 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2454__274
timestamp 1680000651
transform -1 0 40032 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2455__270
timestamp 1680000651
transform -1 0 43200 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2455_
timestamp 1746535128
transform 1 0 42336 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2456__266
timestamp 1680000651
transform -1 0 45312 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2456_
timestamp 1746535128
transform 1 0 44256 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2457_
timestamp 1746535128
transform 1 0 46752 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2457__262
timestamp 1680000651
transform -1 0 47616 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2458__258
timestamp 1680000651
transform -1 0 49632 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2458_
timestamp 1746535128
transform 1 0 48672 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2459__254
timestamp 1680000651
transform -1 0 49824 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2459_
timestamp 1746535128
transform 1 0 48768 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2460__250
timestamp 1680000651
transform -1 0 53184 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2460_
timestamp 1746535128
transform 1 0 52320 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2461__246
timestamp 1680000651
transform -1 0 55584 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2461_
timestamp 1746535128
transform 1 0 54528 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2462__242
timestamp 1680000651
transform -1 0 55104 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2462_
timestamp 1746535128
transform 1 0 54240 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2463_
timestamp 1746535128
transform 1 0 53856 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _2463__238
timestamp 1680000651
transform -1 0 54720 0 1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2464__234
timestamp 1680000651
transform -1 0 52800 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2464_
timestamp 1746535128
transform 1 0 51936 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2465_
timestamp 1746535128
transform 1 0 49152 0 1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2465__230
timestamp 1680000651
transform -1 0 50016 0 -1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2466__226
timestamp 1680000651
transform -1 0 48768 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2466_
timestamp 1746535128
transform 1 0 47904 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2467_
timestamp 1746535128
transform 1 0 46176 0 -1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2467__222
timestamp 1680000651
transform -1 0 47040 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  _2468__218
timestamp 1680000651
transform -1 0 50400 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2468_
timestamp 1746535128
transform 1 0 49536 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2469__214
timestamp 1680000651
transform -1 0 51072 0 -1 18900
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2469_
timestamp 1746535128
transform 1 0 50208 0 1 17388
box -48 -56 2640 834
use sg13g2_tiehi  _2470__210
timestamp 1680000651
transform -1 0 54240 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2470_
timestamp 1746535128
transform 1 0 52992 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2471__206
timestamp 1680000651
transform -1 0 57888 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2471_
timestamp 1746535128
transform 1 0 57024 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2472__202
timestamp 1680000651
transform -1 0 58944 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2472_
timestamp 1746535128
transform 1 0 58080 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2473__454
timestamp 1680000651
transform -1 0 60096 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2473_
timestamp 1746535128
transform 1 0 59232 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2474_
timestamp 1746535128
transform 1 0 59520 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2474__450
timestamp 1680000651
transform -1 0 60384 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2475_
timestamp 1746535128
transform 1 0 60384 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2475__446
timestamp 1680000651
transform -1 0 61344 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2476_
timestamp 1746535128
transform 1 0 61248 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2476__442
timestamp 1680000651
transform -1 0 62112 0 -1 5292
box -48 -56 432 834
use sg13g2_tiehi  _2477__438
timestamp 1680000651
transform -1 0 56928 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2477_
timestamp 1746535128
transform 1 0 56064 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2478__434
timestamp 1680000651
transform -1 0 57408 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2478_
timestamp 1746535128
transform 1 0 56448 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2479__430
timestamp 1680000651
transform -1 0 60480 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2479_
timestamp 1746535128
transform 1 0 59616 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2480__426
timestamp 1680000651
transform -1 0 65280 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2480_
timestamp 1746535128
transform 1 0 64416 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2481__422
timestamp 1680000651
transform -1 0 67200 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2481_
timestamp 1746535128
transform 1 0 66336 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2482_
timestamp 1746535128
transform 1 0 66624 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2482__418
timestamp 1680000651
transform -1 0 67488 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2483_
timestamp 1746535128
transform 1 0 65952 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2483__414
timestamp 1680000651
transform -1 0 66816 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2484__410
timestamp 1680000651
transform -1 0 66048 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2484_
timestamp 1746535128
transform 1 0 65184 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2485_
timestamp 1746535128
transform 1 0 64704 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2485__406
timestamp 1680000651
transform -1 0 65568 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2486_
timestamp 1746535128
transform 1 0 60480 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2486__402
timestamp 1680000651
transform -1 0 61344 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2487_
timestamp 1746535128
transform 1 0 65376 0 -1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2487__398
timestamp 1680000651
transform -1 0 66240 0 1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2488__394
timestamp 1680000651
transform -1 0 71616 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2488_
timestamp 1746535128
transform 1 0 70272 0 1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2489__390
timestamp 1680000651
transform -1 0 71232 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2489_
timestamp 1746535128
transform 1 0 70368 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2490__386
timestamp 1680000651
transform -1 0 71616 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2490_
timestamp 1746535128
transform 1 0 70464 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2491__382
timestamp 1680000651
transform -1 0 72480 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2491_
timestamp 1746535128
transform 1 0 71616 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2492__378
timestamp 1680000651
transform -1 0 72672 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2492_
timestamp 1746535128
transform 1 0 71808 0 -1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _2493__374
timestamp 1680000651
transform -1 0 69600 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2493_
timestamp 1746535128
transform 1 0 68736 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _2494__370
timestamp 1680000651
transform -1 0 72768 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2494_
timestamp 1746535128
transform 1 0 71904 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2495__366
timestamp 1680000651
transform 1 0 74688 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2495_
timestamp 1746535128
transform -1 0 75744 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2496__362
timestamp 1680000651
transform 1 0 77952 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2496_
timestamp 1746535128
transform -1 0 79584 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _2497__358
timestamp 1680000651
transform -1 0 78144 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2497_
timestamp 1746535128
transform 1 0 76992 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2498__354
timestamp 1680000651
transform -1 0 78144 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2498_
timestamp 1746535128
transform 1 0 76992 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2499_
timestamp 1746535128
transform 1 0 76992 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _2499__350
timestamp 1680000651
transform -1 0 78144 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2500__346
timestamp 1680000651
transform -1 0 77952 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2500_
timestamp 1746535128
transform 1 0 76992 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2501_
timestamp 1746535128
transform 1 0 76800 0 -1 12852
box -48 -56 2640 834
use sg13g2_tiehi  _2501__342
timestamp 1680000651
transform -1 0 77664 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2502_
timestamp 1746535128
transform 1 0 76896 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2502__338
timestamp 1680000651
transform -1 0 77760 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _2503__334
timestamp 1680000651
transform -1 0 76992 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2503_
timestamp 1746535128
transform 1 0 76128 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2504_
timestamp 1746535128
transform 1 0 76608 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2504__330
timestamp 1680000651
transform -1 0 77472 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2505__324
timestamp 1680000651
transform -1 0 77856 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2505_
timestamp 1746535128
transform 1 0 76992 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2506_
timestamp 1746535128
transform 1 0 76992 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2506__316
timestamp 1680000651
transform -1 0 77856 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2507_
timestamp 1746535128
transform 1 0 76992 0 -1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2507__308
timestamp 1680000651
transform -1 0 77952 0 1 29484
box -48 -56 432 834
use sg13g2_tiehi  _2508__300
timestamp 1680000651
transform -1 0 78144 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2508_
timestamp 1746535128
transform 1 0 76992 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2509__292
timestamp 1680000651
transform -1 0 78144 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2509_
timestamp 1746535128
transform 1 0 76992 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2510__284
timestamp 1680000651
transform -1 0 78720 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2510_
timestamp 1746535128
transform 1 0 76992 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2511__276
timestamp 1680000651
transform -1 0 74400 0 1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2511_
timestamp 1746535128
transform 1 0 73440 0 -1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2512__268
timestamp 1680000651
transform -1 0 72864 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2512_
timestamp 1746535128
transform 1 0 72000 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2513__260
timestamp 1680000651
transform -1 0 71712 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2513_
timestamp 1746535128
transform 1 0 69120 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2514_
timestamp 1746535128
transform 1 0 67200 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2514__252
timestamp 1680000651
transform -1 0 68064 0 1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2515_
timestamp 1746535128
transform 1 0 66624 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2515__244
timestamp 1680000651
transform -1 0 67488 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  _2516__236
timestamp 1680000651
transform -1 0 73152 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2516_
timestamp 1746535128
transform 1 0 72096 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2517__228
timestamp 1680000651
transform -1 0 72576 0 1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2517_
timestamp 1746535128
transform 1 0 71616 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2518_
timestamp 1746535128
transform 1 0 71328 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2518__220
timestamp 1680000651
transform -1 0 72192 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2519_
timestamp 1746535128
transform 1 0 70560 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2519__212
timestamp 1680000651
transform -1 0 71904 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2520_
timestamp 1746535128
transform 1 0 67872 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2520__204
timestamp 1680000651
transform -1 0 68832 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2521_
timestamp 1746535128
transform 1 0 63936 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2521__452
timestamp 1680000651
transform -1 0 65472 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2522_
timestamp 1746535128
transform 1 0 65664 0 1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2522__444
timestamp 1680000651
transform -1 0 66528 0 -1 27972
box -48 -56 432 834
use sg13g2_tiehi  _2523__436
timestamp 1680000651
transform -1 0 66816 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2523_
timestamp 1746535128
transform 1 0 65952 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2524__428
timestamp 1680000651
transform -1 0 64032 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2524_
timestamp 1746535128
transform 1 0 63168 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2525__420
timestamp 1680000651
transform -1 0 63936 0 -1 35532
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2525_
timestamp 1746535128
transform 1 0 63072 0 1 34020
box -48 -56 2640 834
use sg13g2_tiehi  _2526__412
timestamp 1680000651
transform -1 0 64512 0 -1 38556
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2526_
timestamp 1746535128
transform 1 0 63648 0 1 37044
box -48 -56 2640 834
use sg13g2_tiehi  _2527__404
timestamp 1680000651
transform -1 0 60096 0 1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2527_
timestamp 1746535128
transform 1 0 59040 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2528_
timestamp 1746535128
transform 1 0 55104 0 -1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2528__396
timestamp 1680000651
transform 1 0 55296 0 1 34020
box -48 -56 432 834
use sg13g2_tiehi  _2529__388
timestamp 1680000651
transform -1 0 59520 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2529_
timestamp 1746535128
transform 1 0 58464 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2530__380
timestamp 1680000651
transform -1 0 61728 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2530_
timestamp 1746535128
transform 1 0 60480 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2531_
timestamp 1746535128
transform 1 0 60384 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2531__372
timestamp 1680000651
transform -1 0 61440 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2532_
timestamp 1746535128
transform 1 0 60192 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2532__364
timestamp 1680000651
transform -1 0 61248 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2533__356
timestamp 1680000651
transform -1 0 56064 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2533_
timestamp 1746535128
transform 1 0 54816 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2534_
timestamp 1746535128
transform 1 0 56256 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2534__348
timestamp 1680000651
transform -1 0 57120 0 1 27972
box -48 -56 432 834
use sg13g2_tiehi  _2535__340
timestamp 1680000651
transform -1 0 56928 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2535_
timestamp 1746535128
transform 1 0 56064 0 1 30996
box -48 -56 2640 834
use sg13g2_tiehi  _2536__332
timestamp 1680000651
transform -1 0 56160 0 -1 34020
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2536_
timestamp 1746535128
transform 1 0 55200 0 1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2537__320
timestamp 1680000651
transform -1 0 52800 0 -1 37044
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2537_
timestamp 1746535128
transform 1 0 51936 0 1 35532
box -48 -56 2640 834
use sg13g2_tiehi  _2538__304
timestamp 1680000651
transform -1 0 47616 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2538_
timestamp 1746535128
transform 1 0 45984 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2539_
timestamp 1746535128
transform 1 0 51072 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2539__288
timestamp 1680000651
transform -1 0 51936 0 1 30996
box -48 -56 432 834
use sg13g2_tiehi  _2540__272
timestamp 1680000651
transform -1 0 52032 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2540_
timestamp 1746535128
transform 1 0 51168 0 1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2541__256
timestamp 1680000651
transform -1 0 52800 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2541_
timestamp 1746535128
transform 1 0 52032 0 -1 27972
box -48 -56 2640 834
use sg13g2_tiehi  _2542__240
timestamp 1680000651
transform -1 0 53088 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2542_
timestamp 1746535128
transform 1 0 52224 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2543__224
timestamp 1680000651
transform -1 0 52896 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2543_
timestamp 1746535128
transform 1 0 51648 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2544__208
timestamp 1680000651
transform -1 0 51648 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2544_
timestamp 1746535128
transform 1 0 50208 0 1 20412
box -48 -56 2640 834
use sg13g2_tiehi  _2545__448
timestamp 1680000651
transform -1 0 46752 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2545_
timestamp 1746535128
transform 1 0 45888 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2546__432
timestamp 1680000651
transform -1 0 47232 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2546_
timestamp 1746535128
transform 1 0 46272 0 -1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2547__416
timestamp 1680000651
transform -1 0 47904 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2547_
timestamp 1746535128
transform 1 0 46944 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2548__400
timestamp 1680000651
transform -1 0 47808 0 1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2548_
timestamp 1746535128
transform 1 0 46944 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2549__384
timestamp 1680000651
transform -1 0 47136 0 -1 30996
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2549_
timestamp 1746535128
transform 1 0 46272 0 -1 29484
box -48 -56 2640 834
use sg13g2_tiehi  _2550__368
timestamp 1680000651
transform -1 0 44160 0 1 32508
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2550_
timestamp 1746535128
transform 1 0 43296 0 -1 32508
box -48 -56 2640 834
use sg13g2_tiehi  _2551__352
timestamp 1680000651
transform -1 0 42720 0 -1 29484
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2551_
timestamp 1746535128
transform 1 0 41664 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2552_
timestamp 1746535128
transform 1 0 41568 0 1 26460
box -48 -56 2640 834
use sg13g2_tiehi  _2552__336
timestamp 1680000651
transform -1 0 42432 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2553_
timestamp 1746535128
transform 1 0 40800 0 1 24948
box -48 -56 2640 834
use sg13g2_tiehi  _2553__312
timestamp 1680000651
transform -1 0 41664 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2554__280
timestamp 1680000651
transform -1 0 42336 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2554_
timestamp 1746535128
transform 1 0 41088 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2555__248
timestamp 1680000651
transform 1 0 35712 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2555_
timestamp 1746535128
transform 1 0 35616 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2556__216
timestamp 1680000651
transform -1 0 36768 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2556_
timestamp 1746535128
transform 1 0 35904 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2557_
timestamp 1746535128
transform 1 0 32832 0 1 23436
box -48 -56 2640 834
use sg13g2_tiehi  _2557__440
timestamp 1680000651
transform -1 0 33696 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2558_
timestamp 1746535128
transform 1 0 32736 0 1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2558__408
timestamp 1680000651
transform -1 0 33600 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2559_
timestamp 1746535128
transform 1 0 29280 0 -1 21924
box -48 -56 2640 834
use sg13g2_tiehi  _2559__376
timestamp 1680000651
transform -1 0 30144 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  _2560__344
timestamp 1680000651
transform -1 0 13056 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2560_
timestamp 1746535128
transform 1 0 12192 0 1 18900
box -48 -56 2640 834
use sg13g2_tiehi  _2561__296
timestamp 1680000651
transform -1 0 5856 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2561_
timestamp 1746535128
transform 1 0 4992 0 1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _2562__232
timestamp 1680000651
transform -1 0 5760 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2562_
timestamp 1746535128
transform 1 0 4896 0 1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _2563__424
timestamp 1680000651
transform -1 0 5568 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2563_
timestamp 1746535128
transform 1 0 4704 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2564_
timestamp 1746535128
transform 1 0 4704 0 1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _2564__360
timestamp 1680000651
transform -1 0 5568 0 -1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2565__264
timestamp 1680000651
transform -1 0 6144 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2565_
timestamp 1746535128
transform 1 0 4896 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2566_
timestamp 1746535128
transform 1 0 4800 0 -1 14364
box -48 -56 2640 834
use sg13g2_tiehi  _2566__392
timestamp 1680000651
transform -1 0 5856 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _2567_
timestamp 1746535128
transform 1 0 4512 0 1 15876
box -48 -56 2640 834
use sg13g2_tiehi  _2567__456
timestamp 1680000651
transform -1 0 5376 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2832_
timestamp 1676381911
transform -1 0 1824 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _2833_
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _2834_
timestamp 1676381911
transform -1 0 1728 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _2835_
timestamp 1676381911
transform -1 0 1248 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _2836_
timestamp 1676381911
transform -1 0 1440 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2837_
timestamp 1676381911
transform -1 0 1344 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2838_
timestamp 1676381911
transform -1 0 1632 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _2839_
timestamp 1676381911
transform -1 0 1824 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _2840_
timestamp 1676381911
transform -1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _2841_
timestamp 1676381911
transform -1 0 1344 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _2842_
timestamp 1676381911
transform -1 0 1632 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _2843_
timestamp 1676381911
transform -1 0 1152 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _2844_
timestamp 1676381911
transform -1 0 1824 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _2845_
timestamp 1676381911
transform -1 0 1824 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _2846_
timestamp 1676381911
transform -1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2847_
timestamp 1676381911
transform -1 0 1440 0 1 14364
box -48 -56 432 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform -1 0 41376 0 -1 20412
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_0__f_clk
timestamp 1676553496
transform -1 0 42816 0 -1 11340
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_1__f_clk
timestamp 1676553496
transform 1 0 29184 0 -1 12852
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_2__f_clk
timestamp 1676553496
transform -1 0 55680 0 1 14364
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_3__f_clk
timestamp 1676553496
transform -1 0 55200 0 1 27972
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_leaf_0_clk
timestamp 1676451365
transform 1 0 4512 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_1_clk
timestamp 1676451365
transform 1 0 30912 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_2_clk
timestamp 1676451365
transform -1 0 34368 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_3_clk
timestamp 1676451365
transform -1 0 47520 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_4_clk
timestamp 1676451365
transform -1 0 50304 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_5_clk
timestamp 1676451365
transform -1 0 52800 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_6_clk
timestamp 1676451365
transform -1 0 69600 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_7_clk
timestamp 1676451365
transform 1 0 74112 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_8_clk
timestamp 1676451365
transform -1 0 70944 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_9_clk
timestamp 1676451365
transform -1 0 52800 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_10_clk
timestamp 1676451365
transform 1 0 51552 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_11_clk
timestamp 1676451365
transform -1 0 72384 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_12_clk
timestamp 1676451365
transform -1 0 71136 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_13_clk
timestamp 1676451365
transform 1 0 73056 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_14_clk
timestamp 1676451365
transform 1 0 59424 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_15_clk
timestamp 1676451365
transform 1 0 49152 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_16_clk
timestamp 1676451365
transform 1 0 46560 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_17_clk
timestamp 1676451365
transform 1 0 37152 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_18_clk
timestamp 1676451365
transform -1 0 5280 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkload0
timestamp 1676451365
transform 1 0 51648 0 -1 29484
box -48 -56 1296 834
use sg13g2_inv_1  clkload1
timestamp 1676382929
transform 1 0 45696 0 1 24948
box -48 -56 336 834
use sg13g2_inv_2  clkload2
timestamp 1676382947
transform 1 0 51168 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_2  clkload3
timestamp 1676382947
transform 1 0 48288 0 1 6804
box -48 -56 432 834
use sg13g2_inv_2  clkload4
timestamp 1676382947
transform 1 0 47136 0 -1 14364
box -48 -56 432 834
use sg13g2_inv_8  clkload5
timestamp 1676383150
transform 1 0 4512 0 1 12852
box -48 -56 1008 834
use sg13g2_inv_1  clkload6
timestamp 1676382929
transform 1 0 32736 0 1 24948
box -48 -56 336 834
use sg13g2_inv_4  clkload7
timestamp 1676383058
transform 1 0 37152 0 -1 15876
box -48 -56 624 834
use sg13g2_inv_8  clkload8
timestamp 1676383150
transform 1 0 3936 0 1 5292
box -48 -56 1008 834
use sg13g2_inv_2  clkload9
timestamp 1676382947
transform 1 0 51552 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  clkload10
timestamp 1676382929
transform -1 0 69888 0 1 756
box -48 -56 336 834
use sg13g2_inv_2  clkload11
timestamp 1676382947
transform 1 0 48480 0 1 30996
box -48 -56 432 834
use dac128module  dac
timestamp 0
transform 1 0 53240 0 1 17400
box 0 0 1 1
use sg13g2_inv_1  digitalen.g\[0\].u.inv1
timestamp 1676382929
transform 1 0 52512 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[0\].u.inv2
timestamp 1676382929
transform -1 0 52800 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv1
timestamp 1676382929
transform 1 0 78816 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv2
timestamp 1676382929
transform 1 0 79296 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv1
timestamp 1676382929
transform 1 0 79008 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv2
timestamp 1676382929
transform 1 0 79296 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv1
timestamp 1676382929
transform 1 0 52512 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv2
timestamp 1676382929
transform -1 0 52224 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform 1 0 22272 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform 1 0 27648 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 2304 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform 1 0 40800 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform -1 0 47616 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform 1 0 49728 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform 1 0 40128 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform -1 0 39456 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 39744 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 49920 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform -1 0 49536 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform 1 0 38880 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 57312 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform -1 0 57600 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform -1 0 69696 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 68640 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 60000 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform 1 0 58176 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform -1 0 70176 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform -1 0 67680 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 57408 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform 1 0 2688 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform -1 0 25824 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform 1 0 26304 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout47
timestamp 1676381911
transform 1 0 27072 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform -1 0 3744 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 41856 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout50
timestamp 1676381911
transform -1 0 50400 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform 1 0 50304 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout52
timestamp 1676381911
transform 1 0 41472 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform 1 0 38976 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 50304 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform 1 0 49344 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform 1 0 38592 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform 1 0 57312 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform -1 0 59040 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout59
timestamp 1676381911
transform 1 0 68832 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout60
timestamp 1676381911
transform 1 0 67104 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout61
timestamp 1676381911
transform -1 0 59136 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout62
timestamp 1676381911
transform 1 0 69024 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout63
timestamp 1676381911
transform 1 0 68352 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout64
timestamp 1676381911
transform 1 0 58752 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout65
timestamp 1676381911
transform 1 0 58368 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout66
timestamp 1676381911
transform 1 0 2976 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout67
timestamp 1676381911
transform -1 0 23520 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout68
timestamp 1676381911
transform -1 0 34464 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform 1 0 24384 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform 1 0 3744 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform -1 0 45792 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform 1 0 44832 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform 1 0 51552 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform -1 0 50592 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform 1 0 43968 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform 1 0 41184 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform -1 0 51648 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform 1 0 50112 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 40416 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform -1 0 60384 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform -1 0 70464 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform 1 0 70464 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 60480 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform 1 0 60192 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 61440 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 71808 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 70368 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform 1 0 60960 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform -1 0 4512 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform -1 0 3360 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform -1 0 4896 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout92
timestamp 1676381911
transform 1 0 31680 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout93
timestamp 1676381911
transform 1 0 36768 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout94
timestamp 1676381911
transform 1 0 24768 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout95
timestamp 1676381911
transform 1 0 30816 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout96
timestamp 1676381911
transform 1 0 35520 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout97
timestamp 1676381911
transform 1 0 26688 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout98
timestamp 1676381911
transform -1 0 4128 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout99
timestamp 1676381911
transform 1 0 42048 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform -1 0 46944 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout101
timestamp 1676381911
transform -1 0 40896 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout102
timestamp 1676381911
transform -1 0 43200 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout103
timestamp 1676381911
transform 1 0 54816 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform -1 0 52032 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform -1 0 51456 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout106
timestamp 1676381911
transform 1 0 42816 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform 1 0 44640 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout108
timestamp 1676381911
transform 1 0 39360 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform -1 0 40512 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout110
timestamp 1676381911
transform 1 0 52032 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout111
timestamp 1676381911
transform 1 0 54432 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout112
timestamp 1676381911
transform -1 0 51264 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout113
timestamp 1676381911
transform 1 0 50976 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout114
timestamp 1676381911
transform -1 0 40992 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout115
timestamp 1676381911
transform 1 0 64704 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout116
timestamp 1676381911
transform -1 0 59808 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout117
timestamp 1676381911
transform -1 0 62304 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout118
timestamp 1676381911
transform -1 0 71232 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout119
timestamp 1676381911
transform 1 0 76416 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout120
timestamp 1676381911
transform 1 0 76416 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout121
timestamp 1676381911
transform 1 0 70464 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout122
timestamp 1676381911
transform 1 0 70848 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout123
timestamp 1676381911
transform 1 0 61632 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout124
timestamp 1676381911
transform 1 0 59040 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout125
timestamp 1676381911
transform -1 0 59520 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout126
timestamp 1676381911
transform -1 0 61056 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout127
timestamp 1676381911
transform -1 0 68928 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout128
timestamp 1676381911
transform -1 0 72000 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout129
timestamp 1676381911
transform -1 0 75168 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout130
timestamp 1676381911
transform 1 0 71232 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout131
timestamp 1676381911
transform 1 0 60864 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout132
timestamp 1676381911
transform 1 0 4128 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout133
timestamp 1676381911
transform 1 0 21888 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout134
timestamp 1676381911
transform -1 0 23328 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout135
timestamp 1676381911
transform 1 0 2304 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout136
timestamp 1676381911
transform -1 0 23808 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout137
timestamp 1676381911
transform -1 0 43584 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout138
timestamp 1676381911
transform 1 0 44448 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout139
timestamp 1676381911
transform -1 0 51264 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout140
timestamp 1676381911
transform 1 0 51168 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout141
timestamp 1676381911
transform 1 0 43584 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout142
timestamp 1676381911
transform 1 0 39360 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout143
timestamp 1676381911
transform 1 0 51456 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout144
timestamp 1676381911
transform 1 0 50112 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout145
timestamp 1676381911
transform -1 0 41664 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout146
timestamp 1676381911
transform -1 0 60000 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout147
timestamp 1676381911
transform 1 0 60768 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout148
timestamp 1676381911
transform -1 0 70080 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout149
timestamp 1676381911
transform -1 0 69984 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout150
timestamp 1676381911
transform -1 0 60480 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout151
timestamp 1676381911
transform 1 0 58752 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout152
timestamp 1676381911
transform -1 0 59136 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout153
timestamp 1676381911
transform -1 0 71136 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout154
timestamp 1676381911
transform 1 0 71616 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout155
timestamp 1676381911
transform 1 0 60576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout156
timestamp 1676381911
transform 1 0 3072 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout157
timestamp 1676381911
transform 1 0 3360 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout158
timestamp 1676381911
transform 1 0 24000 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout159
timestamp 1676381911
transform 1 0 23616 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout160
timestamp 1676381911
transform -1 0 1920 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout161
timestamp 1676381911
transform -1 0 45408 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout162
timestamp 1676381911
transform -1 0 44640 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout163
timestamp 1676381911
transform 1 0 51456 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout164
timestamp 1676381911
transform -1 0 44736 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout165
timestamp 1676381911
transform -1 0 40704 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout166
timestamp 1676381911
transform 1 0 51168 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout167
timestamp 1676381911
transform 1 0 51264 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout168
timestamp 1676381911
transform 1 0 40416 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout169
timestamp 1676381911
transform -1 0 59520 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout170
timestamp 1676381911
transform -1 0 63072 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout171
timestamp 1676381911
transform 1 0 70368 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout172
timestamp 1676381911
transform -1 0 70848 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout173
timestamp 1676381911
transform 1 0 60576 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout174
timestamp 1676381911
transform -1 0 60864 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout175
timestamp 1676381911
transform -1 0 72000 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout176
timestamp 1676381911
transform -1 0 72384 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout177
timestamp 1676381911
transform 1 0 60288 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout178
timestamp 1676381911
transform 1 0 1920 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout179
timestamp 1676381911
transform -1 0 2304 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout180
timestamp 1676381911
transform 1 0 21696 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout181
timestamp 1676381911
transform 1 0 28032 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout182
timestamp 1676381911
transform -1 0 5184 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout183
timestamp 1676381911
transform -1 0 41568 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout184
timestamp 1676381911
transform -1 0 48000 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout185
timestamp 1676381911
transform 1 0 49920 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout186
timestamp 1676381911
transform -1 0 43392 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout187
timestamp 1676381911
transform -1 0 40128 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout188
timestamp 1676381911
transform 1 0 42240 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout189
timestamp 1676381911
transform -1 0 57216 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout190
timestamp 1676381911
transform -1 0 51072 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout191
timestamp 1676381911
transform 1 0 42624 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout192
timestamp 1676381911
transform 1 0 58176 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout193
timestamp 1676381911
transform 1 0 57696 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout194
timestamp 1676381911
transform 1 0 70080 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout195
timestamp 1676381911
transform -1 0 69312 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout196
timestamp 1676381911
transform -1 0 59040 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout197
timestamp 1676381911
transform -1 0 59424 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout198
timestamp 1676381911
transform 1 0 67680 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout199
timestamp 1676381911
transform 1 0 67008 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout200
timestamp 1676381911
transform 1 0 58272 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout201
timestamp 1676381911
transform 1 0 4992 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_567
timestamp 1677580104
transform 1 0 55008 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_569
timestamp 1677579658
transform 1 0 55200 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_575
timestamp 1677579658
transform 1 0 55776 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_586
timestamp 1677580104
transform 1 0 56832 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_588
timestamp 1677579658
transform 1 0 57024 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_594
timestamp 1679581782
transform 1 0 57600 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_601
timestamp 1677580104
transform 1 0 58272 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_630
timestamp 1679577901
transform 1 0 61056 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_634
timestamp 1677580104
transform 1 0 61440 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_641
timestamp 1677579658
transform 1 0 62112 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_652
timestamp 1679577901
transform 1 0 63168 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_674
timestamp 1679581782
transform 1 0 65280 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_713
timestamp 1677580104
transform 1 0 69024 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_753
timestamp 1677580104
transform 1 0 72864 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_755
timestamp 1677579658
transform 1 0 73056 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_783
timestamp 1677579658
transform 1 0 75744 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_789
timestamp 1679581782
transform 1 0 76320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_546
timestamp 1679577901
transform 1 0 52992 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_550
timestamp 1677579658
transform 1 0 53376 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_663
timestamp 1677580104
transform 1 0 64224 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_692
timestamp 1677580104
transform 1 0 67008 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_694
timestamp 1677579658
transform 1 0 67200 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_769
timestamp 1677579658
transform 1 0 74400 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_775
timestamp 1677579658
transform 1 0 74976 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_817
timestamp 1679577901
transform 1 0 79008 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_821
timestamp 1677580104
transform 1 0 79392 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_4
timestamp 1679577901
transform 1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_8
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_13
timestamp 1679577901
transform 1 0 1824 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_17
timestamp 1677579658
transform 1 0 2208 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 3936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 4608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 5952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 6624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 7968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 8640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 9984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 14016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 14688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 16704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 18720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679581782
transform 1 0 19392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679581782
transform 1 0 20064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679581782
transform 1 0 20736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679581782
transform 1 0 21408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 22080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679581782
transform 1 0 22752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679581782
transform 1 0 23424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679581782
transform 1 0 24096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1679581782
transform 1 0 24768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1679581782
transform 1 0 25440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1679581782
transform 1 0 26112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1679581782
transform 1 0 26784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1679581782
transform 1 0 27456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1679581782
transform 1 0 28128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1679581782
transform 1 0 28800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1679581782
transform 1 0 29472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1679581782
transform 1 0 30144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_315
timestamp 1679581782
transform 1 0 30816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_322
timestamp 1679581782
transform 1 0 31488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_329
timestamp 1679581782
transform 1 0 32160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679581782
transform 1 0 32832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679581782
transform 1 0 33504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_350
timestamp 1679581782
transform 1 0 34176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_357
timestamp 1679581782
transform 1 0 34848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_364
timestamp 1679581782
transform 1 0 35520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_371
timestamp 1679581782
transform 1 0 36192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_378
timestamp 1679581782
transform 1 0 36864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_385
timestamp 1679581782
transform 1 0 37536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_392
timestamp 1679581782
transform 1 0 38208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_399
timestamp 1679581782
transform 1 0 38880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_406
timestamp 1679581782
transform 1 0 39552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_413
timestamp 1679581782
transform 1 0 40224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_420
timestamp 1679581782
transform 1 0 40896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_427
timestamp 1679581782
transform 1 0 41568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_434
timestamp 1679581782
transform 1 0 42240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_441
timestamp 1679581782
transform 1 0 42912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_448
timestamp 1679581782
transform 1 0 43584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_455
timestamp 1679581782
transform 1 0 44256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_462
timestamp 1679581782
transform 1 0 44928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_469
timestamp 1679581782
transform 1 0 45600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_476
timestamp 1679581782
transform 1 0 46272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_483
timestamp 1679581782
transform 1 0 46944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_490
timestamp 1679581782
transform 1 0 47616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_497
timestamp 1679581782
transform 1 0 48288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_504
timestamp 1679581782
transform 1 0 48960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_511
timestamp 1679581782
transform 1 0 49632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_518
timestamp 1679581782
transform 1 0 50304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_525
timestamp 1679581782
transform 1 0 50976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_532
timestamp 1679581782
transform 1 0 51648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_539
timestamp 1679581782
transform 1 0 52320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_546
timestamp 1679581782
transform 1 0 52992 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_553
timestamp 1677580104
transform 1 0 53664 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_555
timestamp 1677579658
transform 1 0 53856 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_560
timestamp 1679581782
transform 1 0 54336 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_567
timestamp 1677580104
transform 1 0 55008 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_625
timestamp 1679581782
transform 1 0 60576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_632
timestamp 1679581782
transform 1 0 61248 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_639
timestamp 1677580104
transform 1 0 61920 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_645
timestamp 1679581782
transform 1 0 62496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_652
timestamp 1679577901
transform 1 0 63168 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_656
timestamp 1677579658
transform 1 0 63552 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_671
timestamp 1679581782
transform 1 0 64992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_678
timestamp 1679581782
transform 1 0 65664 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_685
timestamp 1677579658
transform 1 0 66336 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_697
timestamp 1679577901
transform 1 0 67488 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_701
timestamp 1677580104
transform 1 0 67872 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_730
timestamp 1679577901
transform 1 0 70656 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_734
timestamp 1677580104
transform 1 0 71040 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_780
timestamp 1679577901
transform 1 0 75456 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_784
timestamp 1677580104
transform 1 0 75840 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_790
timestamp 1677580104
transform 1 0 76416 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_810
timestamp 1679581782
transform 1 0 78336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_817
timestamp 1679577901
transform 1 0 79008 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_821
timestamp 1677580104
transform 1 0 79392 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_35
timestamp 1677580104
transform 1 0 3936 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_50
timestamp 1679581782
transform 1 0 5376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_57
timestamp 1679581782
transform 1 0 6048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_64
timestamp 1679581782
transform 1 0 6720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_71
timestamp 1679581782
transform 1 0 7392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_78
timestamp 1679581782
transform 1 0 8064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_85
timestamp 1679581782
transform 1 0 8736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_92
timestamp 1679581782
transform 1 0 9408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_99
timestamp 1679581782
transform 1 0 10080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_106
timestamp 1679581782
transform 1 0 10752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_113
timestamp 1679581782
transform 1 0 11424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_120
timestamp 1679581782
transform 1 0 12096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_127
timestamp 1679581782
transform 1 0 12768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_134
timestamp 1679581782
transform 1 0 13440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_141
timestamp 1679581782
transform 1 0 14112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_148
timestamp 1679581782
transform 1 0 14784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_155
timestamp 1679581782
transform 1 0 15456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_162
timestamp 1679581782
transform 1 0 16128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_169
timestamp 1679581782
transform 1 0 16800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_176
timestamp 1679581782
transform 1 0 17472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_183
timestamp 1679581782
transform 1 0 18144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_190
timestamp 1679581782
transform 1 0 18816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_197
timestamp 1679581782
transform 1 0 19488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_204
timestamp 1679581782
transform 1 0 20160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_211
timestamp 1679581782
transform 1 0 20832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_218
timestamp 1679581782
transform 1 0 21504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_225
timestamp 1679581782
transform 1 0 22176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_232
timestamp 1679581782
transform 1 0 22848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_239
timestamp 1679581782
transform 1 0 23520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_246
timestamp 1679581782
transform 1 0 24192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_253
timestamp 1679581782
transform 1 0 24864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_260
timestamp 1679581782
transform 1 0 25536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_267
timestamp 1679581782
transform 1 0 26208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_274
timestamp 1679581782
transform 1 0 26880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_281
timestamp 1679581782
transform 1 0 27552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_288
timestamp 1679581782
transform 1 0 28224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_295
timestamp 1679581782
transform 1 0 28896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_302
timestamp 1679581782
transform 1 0 29568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_309
timestamp 1679581782
transform 1 0 30240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_316
timestamp 1679581782
transform 1 0 30912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_323
timestamp 1679581782
transform 1 0 31584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_330
timestamp 1679581782
transform 1 0 32256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_337
timestamp 1679581782
transform 1 0 32928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_344
timestamp 1679581782
transform 1 0 33600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_351
timestamp 1679581782
transform 1 0 34272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_358
timestamp 1679581782
transform 1 0 34944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_365
timestamp 1679581782
transform 1 0 35616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_372
timestamp 1679581782
transform 1 0 36288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_379
timestamp 1679581782
transform 1 0 36960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_386
timestamp 1679581782
transform 1 0 37632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_393
timestamp 1679581782
transform 1 0 38304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_400
timestamp 1679581782
transform 1 0 38976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_407
timestamp 1679581782
transform 1 0 39648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_414
timestamp 1679581782
transform 1 0 40320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_421
timestamp 1679581782
transform 1 0 40992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_428
timestamp 1679581782
transform 1 0 41664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_435
timestamp 1679581782
transform 1 0 42336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_442
timestamp 1679581782
transform 1 0 43008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_449
timestamp 1679581782
transform 1 0 43680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_456
timestamp 1679581782
transform 1 0 44352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_463
timestamp 1679581782
transform 1 0 45024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_470
timestamp 1679581782
transform 1 0 45696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_477
timestamp 1679581782
transform 1 0 46368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_484
timestamp 1679581782
transform 1 0 47040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_491
timestamp 1679581782
transform 1 0 47712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_498
timestamp 1679581782
transform 1 0 48384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_505
timestamp 1679581782
transform 1 0 49056 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_512
timestamp 1677580104
transform 1 0 49728 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_514
timestamp 1677579658
transform 1 0 49920 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_520
timestamp 1677579658
transform 1 0 50496 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_526
timestamp 1679577901
transform 1 0 51072 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_530
timestamp 1677579658
transform 1 0 51456 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_545
timestamp 1679581782
transform 1 0 52896 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_552
timestamp 1677580104
transform 1 0 53568 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_554
timestamp 1677579658
transform 1 0 53760 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_582
timestamp 1677580104
transform 1 0 56448 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_588
timestamp 1679581782
transform 1 0 57024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_595
timestamp 1679581782
transform 1 0 57696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_602
timestamp 1679581782
transform 1 0 58368 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_609
timestamp 1677580104
transform 1 0 59040 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_642
timestamp 1679581782
transform 1 0 62208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_649
timestamp 1679577901
transform 1 0 62880 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_657
timestamp 1677579658
transform 1 0 63648 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_668
timestamp 1679581782
transform 1 0 64704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_675
timestamp 1679581782
transform 1 0 65376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_691
timestamp 1679581782
transform 1 0 66912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_698
timestamp 1679581782
transform 1 0 67584 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_705
timestamp 1677580104
transform 1 0 68256 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_707
timestamp 1677579658
transform 1 0 68448 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_713
timestamp 1677579658
transform 1 0 69024 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_719
timestamp 1677579658
transform 1 0 69600 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_732
timestamp 1677580104
transform 1 0 70848 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_749
timestamp 1679581782
transform 1 0 72480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_756
timestamp 1679577901
transform 1 0 73152 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_760
timestamp 1677580104
transform 1 0 73536 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_794
timestamp 1677580104
transform 1 0 76800 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_796
timestamp 1677579658
transform 1 0 76992 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_8
timestamp 1677580104
transform 1 0 1344 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_10
timestamp 1677579658
transform 1 0 1536 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_25
timestamp 1679577901
transform 1 0 2976 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_39
timestamp 1677580104
transform 1 0 4320 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_73
timestamp 1679581782
transform 1 0 7584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_80
timestamp 1679581782
transform 1 0 8256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_87
timestamp 1679581782
transform 1 0 8928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_94
timestamp 1679581782
transform 1 0 9600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_101
timestamp 1679581782
transform 1 0 10272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_108
timestamp 1679581782
transform 1 0 10944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_115
timestamp 1679581782
transform 1 0 11616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_122
timestamp 1679581782
transform 1 0 12288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_129
timestamp 1679581782
transform 1 0 12960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_136
timestamp 1679581782
transform 1 0 13632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_143
timestamp 1679581782
transform 1 0 14304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_150
timestamp 1679581782
transform 1 0 14976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_157
timestamp 1679581782
transform 1 0 15648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_164
timestamp 1679581782
transform 1 0 16320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_171
timestamp 1679581782
transform 1 0 16992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_178
timestamp 1679581782
transform 1 0 17664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_185
timestamp 1679581782
transform 1 0 18336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_192
timestamp 1679581782
transform 1 0 19008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_199
timestamp 1679581782
transform 1 0 19680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_206
timestamp 1679581782
transform 1 0 20352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_213
timestamp 1679581782
transform 1 0 21024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_220
timestamp 1679581782
transform 1 0 21696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_227
timestamp 1679581782
transform 1 0 22368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_234
timestamp 1679581782
transform 1 0 23040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_241
timestamp 1679581782
transform 1 0 23712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_248
timestamp 1679581782
transform 1 0 24384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_255
timestamp 1679581782
transform 1 0 25056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_262
timestamp 1679581782
transform 1 0 25728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_269
timestamp 1679581782
transform 1 0 26400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_276
timestamp 1679581782
transform 1 0 27072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_283
timestamp 1679581782
transform 1 0 27744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_290
timestamp 1679581782
transform 1 0 28416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_297
timestamp 1679581782
transform 1 0 29088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_304
timestamp 1679581782
transform 1 0 29760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_311
timestamp 1679581782
transform 1 0 30432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_318
timestamp 1679581782
transform 1 0 31104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_325
timestamp 1679581782
transform 1 0 31776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_332
timestamp 1679581782
transform 1 0 32448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679581782
transform 1 0 33120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_346
timestamp 1679581782
transform 1 0 33792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_353
timestamp 1679581782
transform 1 0 34464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679581782
transform 1 0 35136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679581782
transform 1 0 35808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_374
timestamp 1679581782
transform 1 0 36480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_381
timestamp 1679581782
transform 1 0 37152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679581782
transform 1 0 37824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_395
timestamp 1679581782
transform 1 0 38496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679581782
transform 1 0 39168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_409
timestamp 1679581782
transform 1 0 39840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_416
timestamp 1679581782
transform 1 0 40512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_423
timestamp 1679581782
transform 1 0 41184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_430
timestamp 1679581782
transform 1 0 41856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_437
timestamp 1679581782
transform 1 0 42528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_444
timestamp 1679581782
transform 1 0 43200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_451
timestamp 1679581782
transform 1 0 43872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_458
timestamp 1679581782
transform 1 0 44544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_465
timestamp 1679581782
transform 1 0 45216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_472
timestamp 1679581782
transform 1 0 45888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_479
timestamp 1679581782
transform 1 0 46560 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_486
timestamp 1677579658
transform 1 0 47232 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_492
timestamp 1679581782
transform 1 0 47808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_499
timestamp 1679581782
transform 1 0 48480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_506
timestamp 1679577901
transform 1 0 49152 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_537
timestamp 1677580104
transform 1 0 52128 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_570
timestamp 1677580104
transform 1 0 55296 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_572
timestamp 1677579658
transform 1 0 55488 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_593
timestamp 1679577901
transform 1 0 57504 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_602
timestamp 1679577901
transform 1 0 58368 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_606
timestamp 1677580104
transform 1 0 58752 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_624
timestamp 1677580104
transform 1 0 60480 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_636
timestamp 1679581782
transform 1 0 61632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_643
timestamp 1679577901
transform 1 0 62304 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_647
timestamp 1677579658
transform 1 0 62688 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_770
timestamp 1679577901
transform 1 0 74496 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_774
timestamp 1677580104
transform 1 0 74880 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_4
timestamp 1677580104
transform 1 0 960 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_6
timestamp 1677579658
transform 1 0 1152 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 2592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_28
timestamp 1679577901
transform 1 0 3264 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_49
timestamp 1677580104
transform 1 0 5280 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_55
timestamp 1679581782
transform 1 0 5856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_62
timestamp 1679581782
transform 1 0 6528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_69
timestamp 1679581782
transform 1 0 7200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_76
timestamp 1679581782
transform 1 0 7872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_83
timestamp 1679581782
transform 1 0 8544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_90
timestamp 1679581782
transform 1 0 9216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_97
timestamp 1679581782
transform 1 0 9888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_104
timestamp 1679581782
transform 1 0 10560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_111
timestamp 1679581782
transform 1 0 11232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_118
timestamp 1679581782
transform 1 0 11904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_125
timestamp 1679581782
transform 1 0 12576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_132
timestamp 1679581782
transform 1 0 13248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_139
timestamp 1679581782
transform 1 0 13920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_146
timestamp 1679581782
transform 1 0 14592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_153
timestamp 1679581782
transform 1 0 15264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_160
timestamp 1679581782
transform 1 0 15936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_167
timestamp 1679581782
transform 1 0 16608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_174
timestamp 1679581782
transform 1 0 17280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_181
timestamp 1679581782
transform 1 0 17952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_188
timestamp 1679581782
transform 1 0 18624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_195
timestamp 1679581782
transform 1 0 19296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_202
timestamp 1679581782
transform 1 0 19968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_209
timestamp 1679581782
transform 1 0 20640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_216
timestamp 1679581782
transform 1 0 21312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_223
timestamp 1679581782
transform 1 0 21984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_230
timestamp 1679581782
transform 1 0 22656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_237
timestamp 1679581782
transform 1 0 23328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_244
timestamp 1679581782
transform 1 0 24000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_251
timestamp 1679581782
transform 1 0 24672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_258
timestamp 1679581782
transform 1 0 25344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_265
timestamp 1679581782
transform 1 0 26016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_272
timestamp 1679581782
transform 1 0 26688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_279
timestamp 1679581782
transform 1 0 27360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_286
timestamp 1679581782
transform 1 0 28032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_293
timestamp 1679581782
transform 1 0 28704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_300
timestamp 1679581782
transform 1 0 29376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_307
timestamp 1679581782
transform 1 0 30048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_314
timestamp 1679581782
transform 1 0 30720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_321
timestamp 1679581782
transform 1 0 31392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_328
timestamp 1679581782
transform 1 0 32064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_335
timestamp 1679581782
transform 1 0 32736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_342
timestamp 1679581782
transform 1 0 33408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_349
timestamp 1679581782
transform 1 0 34080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_356
timestamp 1679581782
transform 1 0 34752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_363
timestamp 1679581782
transform 1 0 35424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_370
timestamp 1679581782
transform 1 0 36096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_377
timestamp 1679581782
transform 1 0 36768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_384
timestamp 1679581782
transform 1 0 37440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_391
timestamp 1679581782
transform 1 0 38112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_398
timestamp 1679581782
transform 1 0 38784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_405
timestamp 1679581782
transform 1 0 39456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_412
timestamp 1679581782
transform 1 0 40128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_419
timestamp 1679581782
transform 1 0 40800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_426
timestamp 1679581782
transform 1 0 41472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_433
timestamp 1679581782
transform 1 0 42144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_440
timestamp 1679581782
transform 1 0 42816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_447
timestamp 1679581782
transform 1 0 43488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_454
timestamp 1679581782
transform 1 0 44160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_461
timestamp 1679581782
transform 1 0 44832 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_468
timestamp 1677580104
transform 1 0 45504 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_470
timestamp 1677579658
transform 1 0 45696 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_507
timestamp 1679581782
transform 1 0 49248 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_514
timestamp 1677580104
transform 1 0 49920 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_520
timestamp 1679581782
transform 1 0 50496 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_527
timestamp 1677580104
transform 1 0 51168 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_529
timestamp 1677579658
transform 1 0 51360 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_548
timestamp 1679581782
transform 1 0 53184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_555
timestamp 1679581782
transform 1 0 53856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_562
timestamp 1679581782
transform 1 0 54528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_569
timestamp 1679577901
transform 1 0 55200 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_605
timestamp 1677580104
transform 1 0 58656 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_634
timestamp 1677580104
transform 1 0 61440 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_636
timestamp 1677579658
transform 1 0 61632 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_645
timestamp 1679577901
transform 1 0 62496 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_649
timestamp 1677580104
transform 1 0 62880 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_687
timestamp 1677580104
transform 1 0 66528 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_689
timestamp 1677579658
transform 1 0 66720 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_694
timestamp 1679581782
transform 1 0 67200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_701
timestamp 1679581782
transform 1 0 67872 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_708
timestamp 1677580104
transform 1 0 68544 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_710
timestamp 1677579658
transform 1 0 68736 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_720
timestamp 1679581782
transform 1 0 69696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_727
timestamp 1679581782
transform 1 0 70368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_734
timestamp 1679577901
transform 1 0 71040 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_738
timestamp 1677579658
transform 1 0 71424 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_752
timestamp 1679581782
transform 1 0 72768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_759
timestamp 1679581782
transform 1 0 73440 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_766
timestamp 1677579658
transform 1 0 74112 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_771
timestamp 1679581782
transform 1 0 74592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_778
timestamp 1679577901
transform 1 0 75264 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_782
timestamp 1677580104
transform 1 0 75648 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_789
timestamp 1679577901
transform 1 0 76320 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_793
timestamp 1677580104
transform 1 0 76704 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_799
timestamp 1677579658
transform 1 0 77280 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679581782
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679581782
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_822
timestamp 1677579658
transform 1 0 79488 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 576 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_33
timestamp 1677580104
transform 1 0 3744 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_72
timestamp 1679581782
transform 1 0 7488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_79
timestamp 1679581782
transform 1 0 8160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_86
timestamp 1679581782
transform 1 0 8832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_93
timestamp 1679581782
transform 1 0 9504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_100
timestamp 1679581782
transform 1 0 10176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_107
timestamp 1679581782
transform 1 0 10848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_114
timestamp 1679581782
transform 1 0 11520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_121
timestamp 1679581782
transform 1 0 12192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_128
timestamp 1679581782
transform 1 0 12864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_135
timestamp 1679581782
transform 1 0 13536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_142
timestamp 1679581782
transform 1 0 14208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_149
timestamp 1679581782
transform 1 0 14880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_156
timestamp 1679581782
transform 1 0 15552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_163
timestamp 1679581782
transform 1 0 16224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_170
timestamp 1679581782
transform 1 0 16896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_177
timestamp 1679581782
transform 1 0 17568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_184
timestamp 1679581782
transform 1 0 18240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_191
timestamp 1679581782
transform 1 0 18912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_198
timestamp 1679581782
transform 1 0 19584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_205
timestamp 1679581782
transform 1 0 20256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_212
timestamp 1679581782
transform 1 0 20928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_219
timestamp 1679581782
transform 1 0 21600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_226
timestamp 1679581782
transform 1 0 22272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_233
timestamp 1679581782
transform 1 0 22944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_240
timestamp 1679581782
transform 1 0 23616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_247
timestamp 1679581782
transform 1 0 24288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_254
timestamp 1679581782
transform 1 0 24960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_261
timestamp 1679581782
transform 1 0 25632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_268
timestamp 1679581782
transform 1 0 26304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_275
timestamp 1679581782
transform 1 0 26976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_282
timestamp 1679581782
transform 1 0 27648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_289
timestamp 1679581782
transform 1 0 28320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_296
timestamp 1679581782
transform 1 0 28992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_303
timestamp 1679581782
transform 1 0 29664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_310
timestamp 1679581782
transform 1 0 30336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_317
timestamp 1679581782
transform 1 0 31008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_324
timestamp 1679581782
transform 1 0 31680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_331
timestamp 1679581782
transform 1 0 32352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_338
timestamp 1679581782
transform 1 0 33024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_345
timestamp 1679581782
transform 1 0 33696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_352
timestamp 1679581782
transform 1 0 34368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_359
timestamp 1679581782
transform 1 0 35040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_366
timestamp 1679581782
transform 1 0 35712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_373
timestamp 1679581782
transform 1 0 36384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_380
timestamp 1679581782
transform 1 0 37056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_387
timestamp 1679581782
transform 1 0 37728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_394
timestamp 1679581782
transform 1 0 38400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_401
timestamp 1679581782
transform 1 0 39072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_408
timestamp 1679581782
transform 1 0 39744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_415
timestamp 1679581782
transform 1 0 40416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_422
timestamp 1679581782
transform 1 0 41088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_429
timestamp 1679581782
transform 1 0 41760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_436
timestamp 1679581782
transform 1 0 42432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_443
timestamp 1679581782
transform 1 0 43104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_450
timestamp 1679581782
transform 1 0 43776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_457
timestamp 1679581782
transform 1 0 44448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_464
timestamp 1679581782
transform 1 0 45120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_471
timestamp 1679577901
transform 1 0 45792 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_475
timestamp 1677579658
transform 1 0 46176 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_480
timestamp 1679577901
transform 1 0 46656 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_484
timestamp 1677579658
transform 1 0 47040 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_490
timestamp 1679577901
transform 1 0 47616 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_517
timestamp 1679581782
transform 1 0 50208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_524
timestamp 1679581782
transform 1 0 50880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_531
timestamp 1679581782
transform 1 0 51552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_548
timestamp 1679577901
transform 1 0 53184 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_552
timestamp 1677579658
transform 1 0 53568 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_567
timestamp 1679581782
transform 1 0 55008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_574
timestamp 1679577901
transform 1 0 55680 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_578
timestamp 1677579658
transform 1 0 56064 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_587
timestamp 1679581782
transform 1 0 56928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_594
timestamp 1679581782
transform 1 0 57600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_601
timestamp 1679581782
transform 1 0 58272 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_608
timestamp 1677580104
transform 1 0 58944 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_619
timestamp 1679581782
transform 1 0 60000 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_626
timestamp 1677579658
transform 1 0 60672 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_659
timestamp 1679581782
transform 1 0 63840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679581782
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_683
timestamp 1677580104
transform 1 0 66144 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_690
timestamp 1677580104
transform 1 0 66816 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_692
timestamp 1677579658
transform 1 0 67008 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679581782
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679581782
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_711
timestamp 1679577901
transform 1 0 68832 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679581782
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_732
timestamp 1677580104
transform 1 0 70848 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_748
timestamp 1679581782
transform 1 0 72384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_755
timestamp 1679577901
transform 1 0 73056 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_759
timestamp 1677579658
transform 1 0 73440 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_792
timestamp 1679577901
transform 1 0 76608 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_805
timestamp 1679581782
transform 1 0 77856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_812
timestamp 1679581782
transform 1 0 78528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_819
timestamp 1679577901
transform 1 0 79200 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_4
timestamp 1679581782
transform 1 0 960 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_15
timestamp 1677579658
transform 1 0 2016 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_26
timestamp 1679581782
transform 1 0 3072 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_43
timestamp 1677579658
transform 1 0 4704 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_48
timestamp 1677580104
transform 1 0 5184 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_54
timestamp 1679581782
transform 1 0 5760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_61
timestamp 1679581782
transform 1 0 6432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_68
timestamp 1679581782
transform 1 0 7104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_75
timestamp 1679581782
transform 1 0 7776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_82
timestamp 1679581782
transform 1 0 8448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_89
timestamp 1679581782
transform 1 0 9120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679581782
transform 1 0 9792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_103
timestamp 1679581782
transform 1 0 10464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_110
timestamp 1679581782
transform 1 0 11136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_117
timestamp 1679581782
transform 1 0 11808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_124
timestamp 1679581782
transform 1 0 12480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_131
timestamp 1679581782
transform 1 0 13152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_138
timestamp 1679581782
transform 1 0 13824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_145
timestamp 1679581782
transform 1 0 14496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_152
timestamp 1679581782
transform 1 0 15168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_159
timestamp 1679581782
transform 1 0 15840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_166
timestamp 1679581782
transform 1 0 16512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_173
timestamp 1679581782
transform 1 0 17184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_180
timestamp 1679581782
transform 1 0 17856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_187
timestamp 1679581782
transform 1 0 18528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_194
timestamp 1679581782
transform 1 0 19200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_201
timestamp 1679581782
transform 1 0 19872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_208
timestamp 1679581782
transform 1 0 20544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_215
timestamp 1679581782
transform 1 0 21216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_222
timestamp 1679581782
transform 1 0 21888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_229
timestamp 1679581782
transform 1 0 22560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_236
timestamp 1679581782
transform 1 0 23232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_243
timestamp 1679581782
transform 1 0 23904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_250
timestamp 1679581782
transform 1 0 24576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_257
timestamp 1679581782
transform 1 0 25248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_264
timestamp 1679581782
transform 1 0 25920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_271
timestamp 1679581782
transform 1 0 26592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_278
timestamp 1679581782
transform 1 0 27264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_285
timestamp 1679581782
transform 1 0 27936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_292
timestamp 1679581782
transform 1 0 28608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_299
timestamp 1679581782
transform 1 0 29280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_306
timestamp 1679581782
transform 1 0 29952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_313
timestamp 1679581782
transform 1 0 30624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_320
timestamp 1679581782
transform 1 0 31296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_327
timestamp 1679581782
transform 1 0 31968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_334
timestamp 1679581782
transform 1 0 32640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_341
timestamp 1679581782
transform 1 0 33312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_348
timestamp 1679581782
transform 1 0 33984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_355
timestamp 1679581782
transform 1 0 34656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_362
timestamp 1679581782
transform 1 0 35328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_369
timestamp 1679581782
transform 1 0 36000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_376
timestamp 1679581782
transform 1 0 36672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_383
timestamp 1679581782
transform 1 0 37344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_390
timestamp 1679581782
transform 1 0 38016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_397
timestamp 1679581782
transform 1 0 38688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_404
timestamp 1679581782
transform 1 0 39360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_411
timestamp 1679581782
transform 1 0 40032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_418
timestamp 1679581782
transform 1 0 40704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_425
timestamp 1679581782
transform 1 0 41376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_432
timestamp 1679581782
transform 1 0 42048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_439
timestamp 1679581782
transform 1 0 42720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_446
timestamp 1679581782
transform 1 0 43392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_453
timestamp 1679581782
transform 1 0 44064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_460
timestamp 1679581782
transform 1 0 44736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_467
timestamp 1679581782
transform 1 0 45408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_474
timestamp 1679581782
transform 1 0 46080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_481
timestamp 1679577901
transform 1 0 46752 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_495
timestamp 1679581782
transform 1 0 48096 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_556
timestamp 1677579658
transform 1 0 53952 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_589
timestamp 1677580104
transform 1 0 57120 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_595
timestamp 1677580104
transform 1 0 57696 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_597
timestamp 1677579658
transform 1 0 57888 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_608
timestamp 1677580104
transform 1 0 58944 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_615
timestamp 1679577901
transform 1 0 59616 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_619
timestamp 1677579658
transform 1 0 60000 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_624
timestamp 1679581782
transform 1 0 60480 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_631
timestamp 1677580104
transform 1 0 61152 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_637
timestamp 1679581782
transform 1 0 61728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_644
timestamp 1679581782
transform 1 0 62400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_651
timestamp 1679577901
transform 1 0 63072 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_655
timestamp 1677579658
transform 1 0 63456 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_660
timestamp 1679581782
transform 1 0 63936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_667
timestamp 1679581782
transform 1 0 64608 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_674
timestamp 1677580104
transform 1 0 65280 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_676
timestamp 1677579658
transform 1 0 65472 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_687
timestamp 1677579658
transform 1 0 66528 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_773
timestamp 1679581782
transform 1 0 74784 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_780
timestamp 1677579658
transform 1 0 75456 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_4
timestamp 1677580104
transform 1 0 960 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_6
timestamp 1677579658
transform 1 0 1152 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_34
timestamp 1677579658
transform 1 0 3840 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_39
timestamp 1679577901
transform 1 0 4320 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_47
timestamp 1679581782
transform 1 0 5088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_54
timestamp 1679581782
transform 1 0 5760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_61
timestamp 1679581782
transform 1 0 6432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_68
timestamp 1679581782
transform 1 0 7104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_75
timestamp 1679581782
transform 1 0 7776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_82
timestamp 1679581782
transform 1 0 8448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_89
timestamp 1679581782
transform 1 0 9120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_96
timestamp 1679581782
transform 1 0 9792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_103
timestamp 1679581782
transform 1 0 10464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_110
timestamp 1679581782
transform 1 0 11136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_117
timestamp 1679581782
transform 1 0 11808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_124
timestamp 1679581782
transform 1 0 12480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_131
timestamp 1679581782
transform 1 0 13152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_138
timestamp 1679581782
transform 1 0 13824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_145
timestamp 1679581782
transform 1 0 14496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_152
timestamp 1679581782
transform 1 0 15168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_159
timestamp 1679581782
transform 1 0 15840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_166
timestamp 1679581782
transform 1 0 16512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_173
timestamp 1679581782
transform 1 0 17184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_180
timestamp 1679581782
transform 1 0 17856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_187
timestamp 1679581782
transform 1 0 18528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_194
timestamp 1679581782
transform 1 0 19200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_201
timestamp 1679581782
transform 1 0 19872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_208
timestamp 1679581782
transform 1 0 20544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_215
timestamp 1679581782
transform 1 0 21216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_222
timestamp 1679581782
transform 1 0 21888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_229
timestamp 1679581782
transform 1 0 22560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_236
timestamp 1679581782
transform 1 0 23232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_243
timestamp 1679581782
transform 1 0 23904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_250
timestamp 1679581782
transform 1 0 24576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_257
timestamp 1679581782
transform 1 0 25248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_264
timestamp 1679581782
transform 1 0 25920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_271
timestamp 1679581782
transform 1 0 26592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_278
timestamp 1679581782
transform 1 0 27264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_285
timestamp 1679581782
transform 1 0 27936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_292
timestamp 1679581782
transform 1 0 28608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_299
timestamp 1679581782
transform 1 0 29280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_306
timestamp 1679581782
transform 1 0 29952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_313
timestamp 1679581782
transform 1 0 30624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_320
timestamp 1679581782
transform 1 0 31296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_327
timestamp 1679581782
transform 1 0 31968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_334
timestamp 1679581782
transform 1 0 32640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_341
timestamp 1679581782
transform 1 0 33312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_348
timestamp 1679581782
transform 1 0 33984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_355
timestamp 1679581782
transform 1 0 34656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_362
timestamp 1679581782
transform 1 0 35328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_369
timestamp 1679581782
transform 1 0 36000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_376
timestamp 1679581782
transform 1 0 36672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_383
timestamp 1679581782
transform 1 0 37344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_390
timestamp 1679581782
transform 1 0 38016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_397
timestamp 1679581782
transform 1 0 38688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_404
timestamp 1679581782
transform 1 0 39360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_411
timestamp 1679581782
transform 1 0 40032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_418
timestamp 1679581782
transform 1 0 40704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_425
timestamp 1679581782
transform 1 0 41376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_432
timestamp 1679581782
transform 1 0 42048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_439
timestamp 1679581782
transform 1 0 42720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_446
timestamp 1679581782
transform 1 0 43392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_453
timestamp 1679581782
transform 1 0 44064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_460
timestamp 1679577901
transform 1 0 44736 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_464
timestamp 1677580104
transform 1 0 45120 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_493
timestamp 1679577901
transform 1 0 47904 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_528
timestamp 1679577901
transform 1 0 51264 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_532
timestamp 1677580104
transform 1 0 51648 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_538
timestamp 1679577901
transform 1 0 52224 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_542
timestamp 1677579658
transform 1 0 52608 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_553
timestamp 1679577901
transform 1 0 53664 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_557
timestamp 1677579658
transform 1 0 54048 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_562
timestamp 1677580104
transform 1 0 54528 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_564
timestamp 1677579658
transform 1 0 54720 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_573
timestamp 1679581782
transform 1 0 55584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_580
timestamp 1679577901
transform 1 0 56256 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_584
timestamp 1677580104
transform 1 0 56640 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_613
timestamp 1677579658
transform 1 0 59424 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_633
timestamp 1679581782
transform 1 0 61344 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_640
timestamp 1677579658
transform 1 0 62016 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_677
timestamp 1679577901
transform 1 0 65568 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_681
timestamp 1677580104
transform 1 0 65952 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_687
timestamp 1677579658
transform 1 0 66528 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_692
timestamp 1679581782
transform 1 0 67008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_699
timestamp 1679581782
transform 1 0 67680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_706
timestamp 1679581782
transform 1 0 68352 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_713
timestamp 1677579658
transform 1 0 69024 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 70464 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_744
timestamp 1677580104
transform 1 0 72000 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_746
timestamp 1677579658
transform 1 0 72192 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_751
timestamp 1679581782
transform 1 0 72672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_758
timestamp 1679581782
transform 1 0 73344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_765
timestamp 1679581782
transform 1 0 74016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_772
timestamp 1679581782
transform 1 0 74688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_789
timestamp 1679577901
transform 1 0 76320 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_793
timestamp 1677579658
transform 1 0 76704 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_798
timestamp 1677579658
transform 1 0 77184 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_803
timestamp 1677579658
transform 1 0 77664 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_808
timestamp 1679581782
transform 1 0 78144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_815
timestamp 1679581782
transform 1 0 78816 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_822
timestamp 1677579658
transform 1 0 79488 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_4
timestamp 1677579658
transform 1 0 960 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_13
timestamp 1677579658
transform 1 0 1824 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_19
timestamp 1677579658
transform 1 0 2400 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_25
timestamp 1677580104
transform 1 0 2976 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_37
timestamp 1677579658
transform 1 0 4128 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 7968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 8640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 9984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 10656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 12672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 14688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 16704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 18720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 20736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 21408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 22080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 22752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 23424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 24768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 25440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679581782
transform 1 0 26112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679581782
transform 1 0 26784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679581782
transform 1 0 27456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679581782
transform 1 0 28128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679581782
transform 1 0 28800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679581782
transform 1 0 29472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679581782
transform 1 0 30144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679581782
transform 1 0 30816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679581782
transform 1 0 31488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679581782
transform 1 0 32160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679581782
transform 1 0 32832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679581782
transform 1 0 33504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679581782
transform 1 0 34176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679581782
transform 1 0 34848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 35520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679581782
transform 1 0 36192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679581782
transform 1 0 36864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679581782
transform 1 0 37536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679581782
transform 1 0 38208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679581782
transform 1 0 38880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679581782
transform 1 0 39552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679581782
transform 1 0 40224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679581782
transform 1 0 40896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679581782
transform 1 0 41568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679581782
transform 1 0 42240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679581782
transform 1 0 42912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_448
timestamp 1679577901
transform 1 0 43584 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_452
timestamp 1677579658
transform 1 0 43968 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_458
timestamp 1677579658
transform 1 0 44544 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_464
timestamp 1677580104
transform 1 0 45120 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_471
timestamp 1677579658
transform 1 0 45792 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_476
timestamp 1679577901
transform 1 0 46272 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_490
timestamp 1677580104
transform 1 0 47616 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_551
timestamp 1679577901
transform 1 0 53472 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_560
timestamp 1679581782
transform 1 0 54336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_567
timestamp 1679581782
transform 1 0 55008 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_574
timestamp 1677580104
transform 1 0 55680 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_608
timestamp 1679581782
transform 1 0 58944 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_654
timestamp 1677580104
transform 1 0 63360 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_685
timestamp 1677579658
transform 1 0 66336 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_690
timestamp 1679581782
transform 1 0 66816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_697
timestamp 1679581782
transform 1 0 67488 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_704
timestamp 1677579658
transform 1 0 68160 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_732
timestamp 1679577901
transform 1 0 70848 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_736
timestamp 1677579658
transform 1 0 71232 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679581782
transform 1 0 71808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679581782
transform 1 0 72480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_756
timestamp 1679577901
transform 1 0 73152 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_792
timestamp 1677580104
transform 1 0 76608 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_794
timestamp 1677579658
transform 1 0 76800 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_808
timestamp 1679581782
transform 1 0 78144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_815
timestamp 1679581782
transform 1 0 78816 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_822
timestamp 1677579658
transform 1 0 79488 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_4
timestamp 1677580104
transform 1 0 960 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_6
timestamp 1677579658
transform 1 0 1152 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_31
timestamp 1679581782
transform 1 0 3552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_38
timestamp 1679581782
transform 1 0 4224 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_45
timestamp 1677580104
transform 1 0 4896 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_47
timestamp 1677579658
transform 1 0 5088 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_52
timestamp 1679581782
transform 1 0 5568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_59
timestamp 1679581782
transform 1 0 6240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_66
timestamp 1679581782
transform 1 0 6912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_73
timestamp 1679581782
transform 1 0 7584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_80
timestamp 1679581782
transform 1 0 8256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_87
timestamp 1679581782
transform 1 0 8928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_94
timestamp 1679581782
transform 1 0 9600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_101
timestamp 1679581782
transform 1 0 10272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_108
timestamp 1679581782
transform 1 0 10944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_115
timestamp 1679581782
transform 1 0 11616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_122
timestamp 1679581782
transform 1 0 12288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_129
timestamp 1679581782
transform 1 0 12960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_136
timestamp 1679581782
transform 1 0 13632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_143
timestamp 1679581782
transform 1 0 14304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_150
timestamp 1679581782
transform 1 0 14976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_157
timestamp 1679581782
transform 1 0 15648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_164
timestamp 1679581782
transform 1 0 16320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_171
timestamp 1679581782
transform 1 0 16992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_178
timestamp 1679581782
transform 1 0 17664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_185
timestamp 1679581782
transform 1 0 18336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_192
timestamp 1679581782
transform 1 0 19008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_199
timestamp 1679581782
transform 1 0 19680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_206
timestamp 1679581782
transform 1 0 20352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_213
timestamp 1679581782
transform 1 0 21024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_220
timestamp 1679581782
transform 1 0 21696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_227
timestamp 1679581782
transform 1 0 22368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_234
timestamp 1679581782
transform 1 0 23040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_241
timestamp 1679581782
transform 1 0 23712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_248
timestamp 1679581782
transform 1 0 24384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_255
timestamp 1679581782
transform 1 0 25056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_262
timestamp 1679581782
transform 1 0 25728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_269
timestamp 1679581782
transform 1 0 26400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_276
timestamp 1679581782
transform 1 0 27072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_283
timestamp 1679581782
transform 1 0 27744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_290
timestamp 1679581782
transform 1 0 28416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_297
timestamp 1679581782
transform 1 0 29088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_304
timestamp 1679581782
transform 1 0 29760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_311
timestamp 1679581782
transform 1 0 30432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_318
timestamp 1679581782
transform 1 0 31104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_325
timestamp 1679581782
transform 1 0 31776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_332
timestamp 1679581782
transform 1 0 32448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_339
timestamp 1679581782
transform 1 0 33120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_346
timestamp 1679581782
transform 1 0 33792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_353
timestamp 1679581782
transform 1 0 34464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_360
timestamp 1679581782
transform 1 0 35136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_367
timestamp 1679581782
transform 1 0 35808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_374
timestamp 1679581782
transform 1 0 36480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_381
timestamp 1679581782
transform 1 0 37152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_388
timestamp 1679581782
transform 1 0 37824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_395
timestamp 1679581782
transform 1 0 38496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_402
timestamp 1679581782
transform 1 0 39168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_409
timestamp 1679581782
transform 1 0 39840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_416
timestamp 1679581782
transform 1 0 40512 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_423
timestamp 1677580104
transform 1 0 41184 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_425
timestamp 1677579658
transform 1 0 41376 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_484
timestamp 1679581782
transform 1 0 47040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_491
timestamp 1679581782
transform 1 0 47712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_511
timestamp 1679581782
transform 1 0 49632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_518
timestamp 1679577901
transform 1 0 50304 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_522
timestamp 1677580104
transform 1 0 50688 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_528
timestamp 1679581782
transform 1 0 51264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_535
timestamp 1679581782
transform 1 0 51936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_542
timestamp 1679577901
transform 1 0 52608 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_556
timestamp 1677580104
transform 1 0 53952 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_558
timestamp 1677579658
transform 1 0 54144 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_586
timestamp 1679581782
transform 1 0 56832 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_593
timestamp 1677580104
transform 1 0 57504 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_617
timestamp 1677580104
transform 1 0 59808 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679581782
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679581782
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679581782
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679581782
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_655
timestamp 1677580104
transform 1 0 63456 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_657
timestamp 1677579658
transform 1 0 63648 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_672
timestamp 1679581782
transform 1 0 65088 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_679
timestamp 1677580104
transform 1 0 65760 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_708
timestamp 1677580104
transform 1 0 68544 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_710
timestamp 1677579658
transform 1 0 68736 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_728
timestamp 1677580104
transform 1 0 70464 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_771
timestamp 1679581782
transform 1 0 74592 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_778
timestamp 1677580104
transform 1 0 75264 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_780
timestamp 1677579658
transform 1 0 75456 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_35
timestamp 1679577901
transform 1 0 3936 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_52
timestamp 1679581782
transform 1 0 5568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_59
timestamp 1679581782
transform 1 0 6240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_66
timestamp 1679581782
transform 1 0 6912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_73
timestamp 1679581782
transform 1 0 7584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_80
timestamp 1679581782
transform 1 0 8256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_87
timestamp 1679581782
transform 1 0 8928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_94
timestamp 1679581782
transform 1 0 9600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_101
timestamp 1679581782
transform 1 0 10272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_108
timestamp 1679581782
transform 1 0 10944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_115
timestamp 1679581782
transform 1 0 11616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_122
timestamp 1679581782
transform 1 0 12288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_129
timestamp 1679581782
transform 1 0 12960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_136
timestamp 1679581782
transform 1 0 13632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_143
timestamp 1679581782
transform 1 0 14304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_150
timestamp 1679581782
transform 1 0 14976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_157
timestamp 1679581782
transform 1 0 15648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_164
timestamp 1679581782
transform 1 0 16320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_171
timestamp 1679581782
transform 1 0 16992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_178
timestamp 1679581782
transform 1 0 17664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_185
timestamp 1679581782
transform 1 0 18336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_192
timestamp 1679581782
transform 1 0 19008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_199
timestamp 1679581782
transform 1 0 19680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_206
timestamp 1679581782
transform 1 0 20352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_213
timestamp 1679581782
transform 1 0 21024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_220
timestamp 1679581782
transform 1 0 21696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_227
timestamp 1679581782
transform 1 0 22368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_234
timestamp 1679581782
transform 1 0 23040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_241
timestamp 1679581782
transform 1 0 23712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_248
timestamp 1679581782
transform 1 0 24384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_255
timestamp 1679581782
transform 1 0 25056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_262
timestamp 1679581782
transform 1 0 25728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_269
timestamp 1679581782
transform 1 0 26400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_276
timestamp 1679581782
transform 1 0 27072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_283
timestamp 1679581782
transform 1 0 27744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_290
timestamp 1679581782
transform 1 0 28416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_297
timestamp 1679581782
transform 1 0 29088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_304
timestamp 1679581782
transform 1 0 29760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_311
timestamp 1679581782
transform 1 0 30432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_318
timestamp 1679581782
transform 1 0 31104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_325
timestamp 1679581782
transform 1 0 31776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_332
timestamp 1679581782
transform 1 0 32448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_339
timestamp 1679581782
transform 1 0 33120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_346
timestamp 1679581782
transform 1 0 33792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_353
timestamp 1679581782
transform 1 0 34464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_360
timestamp 1679581782
transform 1 0 35136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_367
timestamp 1679581782
transform 1 0 35808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_374
timestamp 1679581782
transform 1 0 36480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_381
timestamp 1679581782
transform 1 0 37152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_388
timestamp 1679581782
transform 1 0 37824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_395
timestamp 1679581782
transform 1 0 38496 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_407
timestamp 1677580104
transform 1 0 39648 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_409
timestamp 1677579658
transform 1 0 39840 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_415
timestamp 1677580104
transform 1 0 40416 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_422
timestamp 1677580104
transform 1 0 41088 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_438
timestamp 1677579658
transform 1 0 42624 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_444
timestamp 1679581782
transform 1 0 43200 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_455
timestamp 1677580104
transform 1 0 44256 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_457
timestamp 1677579658
transform 1 0 44448 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_462
timestamp 1679581782
transform 1 0 44928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_469
timestamp 1679581782
transform 1 0 45600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_490
timestamp 1679581782
transform 1 0 47616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_497
timestamp 1679581782
transform 1 0 48288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679581782
transform 1 0 48960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679581782
transform 1 0 49632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_522
timestamp 1679581782
transform 1 0 50688 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_534
timestamp 1677580104
transform 1 0 51840 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_536
timestamp 1677579658
transform 1 0 52032 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_547
timestamp 1679577901
transform 1 0 53088 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_551
timestamp 1677579658
transform 1 0 53472 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_556
timestamp 1677579658
transform 1 0 53952 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_561
timestamp 1677580104
transform 1 0 54432 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_563
timestamp 1677579658
transform 1 0 54624 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_568
timestamp 1679581782
transform 1 0 55104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_575
timestamp 1679577901
transform 1 0 55776 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_579
timestamp 1677580104
transform 1 0 56160 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_585
timestamp 1679577901
transform 1 0 56736 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_589
timestamp 1677580104
transform 1 0 57120 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_677
timestamp 1679581782
transform 1 0 65568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_684
timestamp 1679577901
transform 1 0 66240 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_688
timestamp 1677580104
transform 1 0 66624 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_735
timestamp 1677579658
transform 1 0 71136 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_744
timestamp 1677579658
transform 1 0 72000 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679581782
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679581782
transform 1 0 73152 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_763
timestamp 1677579658
transform 1 0 73824 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_768
timestamp 1679581782
transform 1 0 74304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_775
timestamp 1679577901
transform 1 0 74976 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_779
timestamp 1677579658
transform 1 0 75360 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_794
timestamp 1677580104
transform 1 0 76800 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_805
timestamp 1679581782
transform 1 0 77856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_812
timestamp 1679581782
transform 1 0 78528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_819
timestamp 1679577901
transform 1 0 79200 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_4  FILLER_12_4
timestamp 1679577901
transform 1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_8
timestamp 1677579658
transform 1 0 1344 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_13
timestamp 1679581782
transform 1 0 1824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_29
timestamp 1679581782
transform 1 0 3360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_36
timestamp 1679581782
transform 1 0 4032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_70
timestamp 1679581782
transform 1 0 7296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_77
timestamp 1679581782
transform 1 0 7968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_84
timestamp 1679581782
transform 1 0 8640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_91
timestamp 1679581782
transform 1 0 9312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_98
timestamp 1679581782
transform 1 0 9984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_105
timestamp 1679581782
transform 1 0 10656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_112
timestamp 1679581782
transform 1 0 11328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_119
timestamp 1679581782
transform 1 0 12000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_126
timestamp 1679581782
transform 1 0 12672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_133
timestamp 1679581782
transform 1 0 13344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_140
timestamp 1679581782
transform 1 0 14016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_147
timestamp 1679581782
transform 1 0 14688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_154
timestamp 1679581782
transform 1 0 15360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_161
timestamp 1679581782
transform 1 0 16032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_168
timestamp 1679581782
transform 1 0 16704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_175
timestamp 1679581782
transform 1 0 17376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_182
timestamp 1679581782
transform 1 0 18048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_189
timestamp 1679581782
transform 1 0 18720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_196
timestamp 1679581782
transform 1 0 19392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_203
timestamp 1679581782
transform 1 0 20064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_210
timestamp 1679581782
transform 1 0 20736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_217
timestamp 1679581782
transform 1 0 21408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_224
timestamp 1679581782
transform 1 0 22080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_231
timestamp 1679581782
transform 1 0 22752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_238
timestamp 1679581782
transform 1 0 23424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_245
timestamp 1679581782
transform 1 0 24096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_252
timestamp 1679581782
transform 1 0 24768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_259
timestamp 1679581782
transform 1 0 25440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_266
timestamp 1679581782
transform 1 0 26112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_273
timestamp 1679581782
transform 1 0 26784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_280
timestamp 1679581782
transform 1 0 27456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_287
timestamp 1679581782
transform 1 0 28128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_294
timestamp 1679581782
transform 1 0 28800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1679581782
transform 1 0 29472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_308
timestamp 1679581782
transform 1 0 30144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_315
timestamp 1679581782
transform 1 0 30816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_322
timestamp 1679581782
transform 1 0 31488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_329
timestamp 1679581782
transform 1 0 32160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_336
timestamp 1679581782
transform 1 0 32832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_343
timestamp 1679581782
transform 1 0 33504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_350
timestamp 1679581782
transform 1 0 34176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_357
timestamp 1679581782
transform 1 0 34848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_364
timestamp 1679581782
transform 1 0 35520 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_371
timestamp 1677580104
transform 1 0 36192 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_400
timestamp 1679577901
transform 1 0 38976 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_431
timestamp 1677579658
transform 1 0 41952 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_436
timestamp 1679581782
transform 1 0 42432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_443
timestamp 1679577901
transform 1 0 43104 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_462
timestamp 1679581782
transform 1 0 44928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_469
timestamp 1679581782
transform 1 0 45600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_508
timestamp 1679577901
transform 1 0 49344 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_539
timestamp 1677580104
transform 1 0 52320 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_541
timestamp 1677579658
transform 1 0 52512 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_556
timestamp 1679577901
transform 1 0 53952 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_564
timestamp 1679581782
transform 1 0 54720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_571
timestamp 1679581782
transform 1 0 55392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_578
timestamp 1679581782
transform 1 0 56064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_585
timestamp 1679577901
transform 1 0 56736 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_589
timestamp 1677580104
transform 1 0 57120 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_617
timestamp 1679581782
transform 1 0 59808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_624
timestamp 1679581782
transform 1 0 60480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_631
timestamp 1679581782
transform 1 0 61152 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_638
timestamp 1677580104
transform 1 0 61824 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_640
timestamp 1677579658
transform 1 0 62016 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_645
timestamp 1679581782
transform 1 0 62496 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_652
timestamp 1677580104
transform 1 0 63168 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_659
timestamp 1677580104
transform 1 0 63840 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_661
timestamp 1677579658
transform 1 0 64032 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_672
timestamp 1677579658
transform 1 0 65088 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_755
timestamp 1679577901
transform 1 0 73056 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_22
timestamp 1677580104
transform 1 0 2688 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_24
timestamp 1677579658
transform 1 0 2880 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_35
timestamp 1679581782
transform 1 0 3936 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_42
timestamp 1677580104
transform 1 0 4608 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_48
timestamp 1679581782
transform 1 0 5184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_55
timestamp 1679581782
transform 1 0 5856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_62
timestamp 1679581782
transform 1 0 6528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_69
timestamp 1679581782
transform 1 0 7200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_76
timestamp 1679581782
transform 1 0 7872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_83
timestamp 1679581782
transform 1 0 8544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_90
timestamp 1679581782
transform 1 0 9216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_97
timestamp 1679581782
transform 1 0 9888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_104
timestamp 1679581782
transform 1 0 10560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_111
timestamp 1679581782
transform 1 0 11232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_118
timestamp 1679581782
transform 1 0 11904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_125
timestamp 1679581782
transform 1 0 12576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_132
timestamp 1679581782
transform 1 0 13248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_139
timestamp 1679581782
transform 1 0 13920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_146
timestamp 1679581782
transform 1 0 14592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_153
timestamp 1679581782
transform 1 0 15264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_160
timestamp 1679581782
transform 1 0 15936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_167
timestamp 1679581782
transform 1 0 16608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_174
timestamp 1679581782
transform 1 0 17280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_181
timestamp 1679581782
transform 1 0 17952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_188
timestamp 1679581782
transform 1 0 18624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_195
timestamp 1679581782
transform 1 0 19296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_202
timestamp 1679581782
transform 1 0 19968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_209
timestamp 1679581782
transform 1 0 20640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_216
timestamp 1679581782
transform 1 0 21312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_223
timestamp 1679581782
transform 1 0 21984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_230
timestamp 1679581782
transform 1 0 22656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_237
timestamp 1679581782
transform 1 0 23328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_244
timestamp 1679581782
transform 1 0 24000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_251
timestamp 1679581782
transform 1 0 24672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_258
timestamp 1679581782
transform 1 0 25344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_265
timestamp 1679581782
transform 1 0 26016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_272
timestamp 1679581782
transform 1 0 26688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_279
timestamp 1679581782
transform 1 0 27360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_286
timestamp 1679581782
transform 1 0 28032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_293
timestamp 1679581782
transform 1 0 28704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_300
timestamp 1679581782
transform 1 0 29376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_307
timestamp 1679581782
transform 1 0 30048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_314
timestamp 1679581782
transform 1 0 30720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_321
timestamp 1679581782
transform 1 0 31392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_328
timestamp 1679581782
transform 1 0 32064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_335
timestamp 1679581782
transform 1 0 32736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_342
timestamp 1679581782
transform 1 0 33408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_349
timestamp 1679581782
transform 1 0 34080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_356
timestamp 1679581782
transform 1 0 34752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_363
timestamp 1679581782
transform 1 0 35424 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_370
timestamp 1677580104
transform 1 0 36096 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_372
timestamp 1677579658
transform 1 0 36288 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_388
timestamp 1679577901
transform 1 0 37824 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_392
timestamp 1677580104
transform 1 0 38208 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_408
timestamp 1677580104
transform 1 0 39744 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_414
timestamp 1677579658
transform 1 0 40320 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_444
timestamp 1679581782
transform 1 0 43200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_486
timestamp 1679581782
transform 1 0 47232 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_493
timestamp 1677580104
transform 1 0 47904 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_536
timestamp 1679577901
transform 1 0 52032 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_545
timestamp 1677579658
transform 1 0 52896 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_619
timestamp 1679581782
transform 1 0 60000 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_626
timestamp 1677580104
transform 1 0 60672 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_655
timestamp 1679581782
transform 1 0 63456 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_662
timestamp 1677580104
transform 1 0 64128 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_664
timestamp 1677579658
transform 1 0 64320 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_674
timestamp 1679577901
transform 1 0 65280 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_682
timestamp 1679581782
transform 1 0 66048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_689
timestamp 1679581782
transform 1 0 66720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_696
timestamp 1679581782
transform 1 0 67392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_703
timestamp 1679581782
transform 1 0 68064 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_710
timestamp 1677579658
transform 1 0 68736 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_740
timestamp 1679581782
transform 1 0 71616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_747
timestamp 1679581782
transform 1 0 72288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_758
timestamp 1679581782
transform 1 0 73344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_765
timestamp 1679577901
transform 1 0 74016 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_769
timestamp 1677580104
transform 1 0 74400 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_794
timestamp 1677580104
transform 1 0 76800 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_800
timestamp 1677580104
transform 1 0 77376 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_806
timestamp 1679581782
transform 1 0 77952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_813
timestamp 1679581782
transform 1 0 78624 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_820
timestamp 1677580104
transform 1 0 79296 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_822
timestamp 1677579658
transform 1 0 79488 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1677580104
transform 1 0 576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_2
timestamp 1677579658
transform 1 0 768 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_38
timestamp 1677580104
transform 1 0 4224 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_72
timestamp 1679581782
transform 1 0 7488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_79
timestamp 1679581782
transform 1 0 8160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_86
timestamp 1679581782
transform 1 0 8832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_93
timestamp 1679581782
transform 1 0 9504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_100
timestamp 1679581782
transform 1 0 10176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_107
timestamp 1679581782
transform 1 0 10848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_114
timestamp 1679581782
transform 1 0 11520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_121
timestamp 1679581782
transform 1 0 12192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_128
timestamp 1679581782
transform 1 0 12864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_135
timestamp 1679581782
transform 1 0 13536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_142
timestamp 1679581782
transform 1 0 14208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_149
timestamp 1679581782
transform 1 0 14880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_156
timestamp 1679581782
transform 1 0 15552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_163
timestamp 1679581782
transform 1 0 16224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_170
timestamp 1679581782
transform 1 0 16896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_177
timestamp 1679581782
transform 1 0 17568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_184
timestamp 1679581782
transform 1 0 18240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_191
timestamp 1679581782
transform 1 0 18912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_198
timestamp 1679581782
transform 1 0 19584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_205
timestamp 1679581782
transform 1 0 20256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_212
timestamp 1679581782
transform 1 0 20928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_219
timestamp 1679581782
transform 1 0 21600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_226
timestamp 1679581782
transform 1 0 22272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_233
timestamp 1679581782
transform 1 0 22944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_240
timestamp 1679581782
transform 1 0 23616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_247
timestamp 1679581782
transform 1 0 24288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_254
timestamp 1679581782
transform 1 0 24960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_261
timestamp 1679581782
transform 1 0 25632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_268
timestamp 1679581782
transform 1 0 26304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_275
timestamp 1679581782
transform 1 0 26976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_282
timestamp 1679581782
transform 1 0 27648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_289
timestamp 1679581782
transform 1 0 28320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_296
timestamp 1679581782
transform 1 0 28992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_303
timestamp 1679581782
transform 1 0 29664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_310
timestamp 1679581782
transform 1 0 30336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_317
timestamp 1679581782
transform 1 0 31008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_324
timestamp 1679581782
transform 1 0 31680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_331
timestamp 1679581782
transform 1 0 32352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_338
timestamp 1679581782
transform 1 0 33024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_345
timestamp 1679577901
transform 1 0 33696 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_349
timestamp 1677580104
transform 1 0 34080 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_355
timestamp 1677579658
transform 1 0 34656 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_366
timestamp 1679577901
transform 1 0 35712 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_383
timestamp 1679581782
transform 1 0 37344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_390
timestamp 1679581782
transform 1 0 38016 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_397
timestamp 1677579658
transform 1 0 38688 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_411
timestamp 1679581782
transform 1 0 40032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_418
timestamp 1679581782
transform 1 0 40704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_466
timestamp 1679577901
transform 1 0 45312 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_474
timestamp 1679581782
transform 1 0 46080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_481
timestamp 1679581782
transform 1 0 46752 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_488
timestamp 1677580104
transform 1 0 47424 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_490
timestamp 1677579658
transform 1 0 47616 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_505
timestamp 1677579658
transform 1 0 49056 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_511
timestamp 1679581782
transform 1 0 49632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_518
timestamp 1679577901
transform 1 0 50304 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_541
timestamp 1679581782
transform 1 0 52512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_548
timestamp 1679581782
transform 1 0 53184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_555
timestamp 1679581782
transform 1 0 53856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_562
timestamp 1679581782
transform 1 0 54528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_573
timestamp 1679577901
transform 1 0 55584 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_577
timestamp 1677579658
transform 1 0 55968 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_587
timestamp 1677580104
transform 1 0 56928 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_589
timestamp 1677579658
transform 1 0 57120 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_604
timestamp 1677580104
transform 1 0 58560 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_642
timestamp 1679577901
transform 1 0 62208 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_646
timestamp 1677579658
transform 1 0 62592 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_657
timestamp 1677579658
transform 1 0 63648 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_667
timestamp 1679577901
transform 1 0 64608 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_671
timestamp 1677580104
transform 1 0 64992 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_677
timestamp 1679581782
transform 1 0 65568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_684
timestamp 1679581782
transform 1 0 66240 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_691
timestamp 1677580104
transform 1 0 66912 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_693
timestamp 1677579658
transform 1 0 67104 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_698
timestamp 1679581782
transform 1 0 67584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_705
timestamp 1679577901
transform 1 0 68256 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_709
timestamp 1677580104
transform 1 0 68640 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_726
timestamp 1677579658
transform 1 0 70272 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_731
timestamp 1679581782
transform 1 0 70752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_738
timestamp 1679581782
transform 1 0 71424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_745
timestamp 1679577901
transform 1 0 72096 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_776
timestamp 1677579658
transform 1 0 75072 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_787
timestamp 1677580104
transform 1 0 76128 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_789
timestamp 1677579658
transform 1 0 76320 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_803
timestamp 1679581782
transform 1 0 77664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_810
timestamp 1679581782
transform 1 0 78336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_817
timestamp 1679577901
transform 1 0 79008 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_821
timestamp 1677580104
transform 1 0 79392 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_4
timestamp 1677579658
transform 1 0 960 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_27
timestamp 1679581782
transform 1 0 3168 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_34
timestamp 1677579658
transform 1 0 3840 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_39
timestamp 1677580104
transform 1 0 4320 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_58
timestamp 1679581782
transform 1 0 6144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_65
timestamp 1679581782
transform 1 0 6816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_72
timestamp 1679581782
transform 1 0 7488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_79
timestamp 1679581782
transform 1 0 8160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_86
timestamp 1679581782
transform 1 0 8832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_93
timestamp 1679581782
transform 1 0 9504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_100
timestamp 1679581782
transform 1 0 10176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_107
timestamp 1679581782
transform 1 0 10848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_114
timestamp 1679581782
transform 1 0 11520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_121
timestamp 1679581782
transform 1 0 12192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_128
timestamp 1679581782
transform 1 0 12864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_135
timestamp 1679581782
transform 1 0 13536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_142
timestamp 1679581782
transform 1 0 14208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_149
timestamp 1679581782
transform 1 0 14880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_156
timestamp 1679581782
transform 1 0 15552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_163
timestamp 1679581782
transform 1 0 16224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_170
timestamp 1679581782
transform 1 0 16896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_177
timestamp 1679581782
transform 1 0 17568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_184
timestamp 1679581782
transform 1 0 18240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_191
timestamp 1679581782
transform 1 0 18912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_198
timestamp 1679581782
transform 1 0 19584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_205
timestamp 1679581782
transform 1 0 20256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_212
timestamp 1679581782
transform 1 0 20928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_219
timestamp 1679581782
transform 1 0 21600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_226
timestamp 1679581782
transform 1 0 22272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_233
timestamp 1679581782
transform 1 0 22944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_240
timestamp 1679581782
transform 1 0 23616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_247
timestamp 1679581782
transform 1 0 24288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_254
timestamp 1679581782
transform 1 0 24960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_261
timestamp 1679581782
transform 1 0 25632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_268
timestamp 1679581782
transform 1 0 26304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_275
timestamp 1679581782
transform 1 0 26976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_282
timestamp 1679581782
transform 1 0 27648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_289
timestamp 1679581782
transform 1 0 28320 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_296
timestamp 1677580104
transform 1 0 28992 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_323
timestamp 1679581782
transform 1 0 31584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_330
timestamp 1679581782
transform 1 0 32256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_337
timestamp 1679581782
transform 1 0 32928 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_344
timestamp 1677580104
transform 1 0 33600 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_387
timestamp 1679581782
transform 1 0 37728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_394
timestamp 1679581782
transform 1 0 38400 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_428
timestamp 1677580104
transform 1 0 41664 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_439
timestamp 1677579658
transform 1 0 42720 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_444
timestamp 1679581782
transform 1 0 43200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_451
timestamp 1679581782
transform 1 0 43872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_458
timestamp 1679581782
transform 1 0 44544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_519
timestamp 1679577901
transform 1 0 50400 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_523
timestamp 1677579658
transform 1 0 50784 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_528
timestamp 1677580104
transform 1 0 51264 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_530
timestamp 1677579658
transform 1 0 51456 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_562
timestamp 1677580104
transform 1 0 54528 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_591
timestamp 1679577901
transform 1 0 57312 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_603
timestamp 1679581782
transform 1 0 58464 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_610
timestamp 1677579658
transform 1 0 59136 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_615
timestamp 1677579658
transform 1 0 59616 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_620
timestamp 1679581782
transform 1 0 60096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_627
timestamp 1679581782
transform 1 0 60768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_634
timestamp 1679577901
transform 1 0 61440 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_638
timestamp 1677579658
transform 1 0 61824 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_644
timestamp 1679581782
transform 1 0 62400 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_651
timestamp 1677579658
transform 1 0 63072 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_662
timestamp 1677580104
transform 1 0 64128 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_754
timestamp 1679581782
transform 1 0 72960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_761
timestamp 1679577901
transform 1 0 73632 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_765
timestamp 1677580104
transform 1 0 74016 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_777
timestamp 1679581782
transform 1 0 75168 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_784
timestamp 1677579658
transform 1 0 75840 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_789
timestamp 1679577901
transform 1 0 76320 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_793
timestamp 1677579658
transform 1 0 76704 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_821
timestamp 1677580104
transform 1 0 79392 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_35
timestamp 1677580104
transform 1 0 3936 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_55
timestamp 1679581782
transform 1 0 5856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_62
timestamp 1679581782
transform 1 0 6528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_69
timestamp 1679581782
transform 1 0 7200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_76
timestamp 1679581782
transform 1 0 7872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_83
timestamp 1679581782
transform 1 0 8544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_90
timestamp 1679581782
transform 1 0 9216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_97
timestamp 1679581782
transform 1 0 9888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_104
timestamp 1679581782
transform 1 0 10560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_111
timestamp 1679581782
transform 1 0 11232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_118
timestamp 1679581782
transform 1 0 11904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_125
timestamp 1679581782
transform 1 0 12576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_132
timestamp 1679581782
transform 1 0 13248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_139
timestamp 1679581782
transform 1 0 13920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_146
timestamp 1679581782
transform 1 0 14592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_153
timestamp 1679581782
transform 1 0 15264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_160
timestamp 1679581782
transform 1 0 15936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_167
timestamp 1679581782
transform 1 0 16608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_174
timestamp 1679581782
transform 1 0 17280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_181
timestamp 1679581782
transform 1 0 17952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_188
timestamp 1679581782
transform 1 0 18624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_195
timestamp 1679581782
transform 1 0 19296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_202
timestamp 1679581782
transform 1 0 19968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_209
timestamp 1679581782
transform 1 0 20640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_216
timestamp 1679581782
transform 1 0 21312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_223
timestamp 1679581782
transform 1 0 21984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_230
timestamp 1679581782
transform 1 0 22656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_237
timestamp 1679581782
transform 1 0 23328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_244
timestamp 1679581782
transform 1 0 24000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_251
timestamp 1679581782
transform 1 0 24672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_258
timestamp 1679581782
transform 1 0 25344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_265
timestamp 1679581782
transform 1 0 26016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_272
timestamp 1679581782
transform 1 0 26688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_279
timestamp 1679581782
transform 1 0 27360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_286
timestamp 1679581782
transform 1 0 28032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_293
timestamp 1679581782
transform 1 0 28704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_300
timestamp 1679581782
transform 1 0 29376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_307
timestamp 1679581782
transform 1 0 30048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_314
timestamp 1679581782
transform 1 0 30720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_321
timestamp 1679581782
transform 1 0 31392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_328
timestamp 1679581782
transform 1 0 32064 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_340
timestamp 1677580104
transform 1 0 33216 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_342
timestamp 1677579658
transform 1 0 33408 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_347
timestamp 1679581782
transform 1 0 33888 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_354
timestamp 1677580104
transform 1 0 34560 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_356
timestamp 1677579658
transform 1 0 34752 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_362
timestamp 1679581782
transform 1 0 35328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_369
timestamp 1679577901
transform 1 0 36000 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_373
timestamp 1677579658
transform 1 0 36384 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_405
timestamp 1679581782
transform 1 0 39456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_412
timestamp 1679577901
transform 1 0 40128 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_416
timestamp 1677580104
transform 1 0 40512 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_422
timestamp 1677580104
transform 1 0 41088 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_424
timestamp 1677579658
transform 1 0 41280 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_430
timestamp 1679581782
transform 1 0 41856 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_437
timestamp 1677579658
transform 1 0 42528 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_497
timestamp 1677580104
transform 1 0 48288 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_503
timestamp 1677580104
transform 1 0 48864 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_505
timestamp 1677579658
transform 1 0 49056 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_533
timestamp 1677579658
transform 1 0 51744 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_538
timestamp 1677580104
transform 1 0 52224 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_544
timestamp 1679581782
transform 1 0 52800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_551
timestamp 1679581782
transform 1 0 53472 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_558
timestamp 1677580104
transform 1 0 54144 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_565
timestamp 1677580104
transform 1 0 54816 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_572
timestamp 1679577901
transform 1 0 55488 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_576
timestamp 1677579658
transform 1 0 55872 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_587
timestamp 1679581782
transform 1 0 56928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679581782
transform 1 0 59040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679581782
transform 1 0 59712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_623
timestamp 1679577901
transform 1 0 60384 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_645
timestamp 1679581782
transform 1 0 62496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_652
timestamp 1679581782
transform 1 0 63168 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_659
timestamp 1677580104
transform 1 0 63840 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_661
timestamp 1677579658
transform 1 0 64032 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_676
timestamp 1679581782
transform 1 0 65472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_683
timestamp 1679581782
transform 1 0 66144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_690
timestamp 1679581782
transform 1 0 66816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_697
timestamp 1679581782
transform 1 0 67488 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_704
timestamp 1677580104
transform 1 0 68160 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_706
timestamp 1677579658
transform 1 0 68352 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_717
timestamp 1677580104
transform 1 0 69408 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_727
timestamp 1679577901
transform 1 0 70368 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_731
timestamp 1677579658
transform 1 0 70752 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_736
timestamp 1679577901
transform 1 0 71232 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_740
timestamp 1677580104
transform 1 0 71616 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_788
timestamp 1677580104
transform 1 0 76224 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_799
timestamp 1677579658
transform 1 0 77280 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_804
timestamp 1679581782
transform 1 0 77760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679581782
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_818
timestamp 1679577901
transform 1 0 79104 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_822
timestamp 1677579658
transform 1 0 79488 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_20
timestamp 1677579658
transform 1 0 2496 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_36
timestamp 1677580104
transform 1 0 4032 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_38
timestamp 1677579658
transform 1 0 4224 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_71
timestamp 1679581782
transform 1 0 7392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_78
timestamp 1679581782
transform 1 0 8064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_85
timestamp 1679581782
transform 1 0 8736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_92
timestamp 1679581782
transform 1 0 9408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_99
timestamp 1679581782
transform 1 0 10080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_106
timestamp 1679581782
transform 1 0 10752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_113
timestamp 1679581782
transform 1 0 11424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_120
timestamp 1679581782
transform 1 0 12096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_127
timestamp 1679581782
transform 1 0 12768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_134
timestamp 1679581782
transform 1 0 13440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_141
timestamp 1679581782
transform 1 0 14112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_148
timestamp 1679581782
transform 1 0 14784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_155
timestamp 1679581782
transform 1 0 15456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_162
timestamp 1679581782
transform 1 0 16128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_169
timestamp 1679581782
transform 1 0 16800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_176
timestamp 1679581782
transform 1 0 17472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_183
timestamp 1679581782
transform 1 0 18144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_190
timestamp 1679581782
transform 1 0 18816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_197
timestamp 1679581782
transform 1 0 19488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_204
timestamp 1679581782
transform 1 0 20160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_211
timestamp 1679581782
transform 1 0 20832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_218
timestamp 1679581782
transform 1 0 21504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_225
timestamp 1679581782
transform 1 0 22176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_232
timestamp 1679581782
transform 1 0 22848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_239
timestamp 1679581782
transform 1 0 23520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_246
timestamp 1679581782
transform 1 0 24192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_253
timestamp 1679581782
transform 1 0 24864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_260
timestamp 1679581782
transform 1 0 25536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_267
timestamp 1679581782
transform 1 0 26208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_274
timestamp 1679581782
transform 1 0 26880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_281
timestamp 1679581782
transform 1 0 27552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_288
timestamp 1679581782
transform 1 0 28224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_295
timestamp 1679581782
transform 1 0 28896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_302
timestamp 1679581782
transform 1 0 29568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_309
timestamp 1679577901
transform 1 0 30240 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_17_317
timestamp 1679577901
transform 1 0 31008 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_321
timestamp 1677580104
transform 1 0 31392 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_365
timestamp 1679581782
transform 1 0 35616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_372
timestamp 1679581782
transform 1 0 36288 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_379
timestamp 1677580104
transform 1 0 36960 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_399
timestamp 1677580104
transform 1 0 38880 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_406
timestamp 1677580104
transform 1 0 39552 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_454
timestamp 1679577901
transform 1 0 44160 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_494
timestamp 1679581782
transform 1 0 48000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_501
timestamp 1679581782
transform 1 0 48672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_508
timestamp 1679581782
transform 1 0 49344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_515
timestamp 1679581782
transform 1 0 50016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_522
timestamp 1679577901
transform 1 0 50688 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_17_535
timestamp 1679577901
transform 1 0 51936 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_539
timestamp 1677579658
transform 1 0 52320 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_544
timestamp 1679577901
transform 1 0 52800 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_580
timestamp 1677579658
transform 1 0 56256 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_585
timestamp 1679581782
transform 1 0 56736 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_592
timestamp 1677580104
transform 1 0 57408 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_594
timestamp 1677579658
transform 1 0 57600 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_626
timestamp 1677579658
transform 1 0 60672 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_663
timestamp 1677580104
transform 1 0 64224 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_665
timestamp 1677579658
transform 1 0 64416 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_693
timestamp 1677579658
transform 1 0 67104 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_699
timestamp 1677580104
transform 1 0 67680 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_701
timestamp 1677579658
transform 1 0 67872 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_716
timestamp 1677580104
transform 1 0 69312 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_736
timestamp 1679581782
transform 1 0 71232 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_743
timestamp 1677580104
transform 1 0 71904 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_777
timestamp 1679577901
transform 1 0 75168 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_781
timestamp 1677580104
transform 1 0 75552 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_787
timestamp 1679581782
transform 1 0 76128 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_794
timestamp 1677579658
transform 1 0 76800 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_822
timestamp 1677579658
transform 1 0 79488 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_4
timestamp 1677579658
transform 1 0 960 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_13
timestamp 1677579658
transform 1 0 1824 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_33
timestamp 1679581782
transform 1 0 3744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_40
timestamp 1679581782
transform 1 0 4416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_47
timestamp 1679581782
transform 1 0 5088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_54
timestamp 1679581782
transform 1 0 5760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_61
timestamp 1679581782
transform 1 0 6432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_68
timestamp 1679581782
transform 1 0 7104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_75
timestamp 1679581782
transform 1 0 7776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_82
timestamp 1679581782
transform 1 0 8448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_89
timestamp 1679581782
transform 1 0 9120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_96
timestamp 1679581782
transform 1 0 9792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_103
timestamp 1679581782
transform 1 0 10464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_110
timestamp 1679581782
transform 1 0 11136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_117
timestamp 1679581782
transform 1 0 11808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_124
timestamp 1679581782
transform 1 0 12480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_131
timestamp 1679581782
transform 1 0 13152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_138
timestamp 1679581782
transform 1 0 13824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_145
timestamp 1679581782
transform 1 0 14496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_152
timestamp 1679581782
transform 1 0 15168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_159
timestamp 1679581782
transform 1 0 15840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_166
timestamp 1679581782
transform 1 0 16512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_173
timestamp 1679581782
transform 1 0 17184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_180
timestamp 1679581782
transform 1 0 17856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_187
timestamp 1679581782
transform 1 0 18528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_194
timestamp 1679581782
transform 1 0 19200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_201
timestamp 1679581782
transform 1 0 19872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_208
timestamp 1679581782
transform 1 0 20544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_215
timestamp 1679581782
transform 1 0 21216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_222
timestamp 1679581782
transform 1 0 21888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_229
timestamp 1679581782
transform 1 0 22560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_236
timestamp 1679581782
transform 1 0 23232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_243
timestamp 1679581782
transform 1 0 23904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_250
timestamp 1679581782
transform 1 0 24576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_257
timestamp 1679581782
transform 1 0 25248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_264
timestamp 1679581782
transform 1 0 25920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_271
timestamp 1679581782
transform 1 0 26592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_278
timestamp 1679581782
transform 1 0 27264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_285
timestamp 1679581782
transform 1 0 27936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_292
timestamp 1679581782
transform 1 0 28608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_299
timestamp 1679581782
transform 1 0 29280 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_306
timestamp 1677580104
transform 1 0 29952 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_344
timestamp 1679581782
transform 1 0 33600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_351
timestamp 1679577901
transform 1 0 34272 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_355
timestamp 1677579658
transform 1 0 34656 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_415
timestamp 1679581782
transform 1 0 40416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_427
timestamp 1679581782
transform 1 0 41568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_434
timestamp 1679577901
transform 1 0 42240 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_447
timestamp 1679581782
transform 1 0 43488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_454
timestamp 1679581782
transform 1 0 44160 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_461
timestamp 1677580104
transform 1 0 44832 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_467
timestamp 1679577901
transform 1 0 45408 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_471
timestamp 1677580104
transform 1 0 45792 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_478
timestamp 1679577901
transform 1 0 46464 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_492
timestamp 1677579658
transform 1 0 47808 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_520
timestamp 1677580104
transform 1 0 50496 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_574
timestamp 1677580104
transform 1 0 55680 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_595
timestamp 1679581782
transform 1 0 57696 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_602
timestamp 1677580104
transform 1 0 58368 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_608
timestamp 1679581782
transform 1 0 58944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_615
timestamp 1679577901
transform 1 0 59616 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_619
timestamp 1677579658
transform 1 0 60000 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_651
timestamp 1679581782
transform 1 0 63072 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_677
timestamp 1677580104
transform 1 0 65568 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_679
timestamp 1677579658
transform 1 0 65760 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_684
timestamp 1679581782
transform 1 0 66240 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_691
timestamp 1677580104
transform 1 0 66912 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_724
timestamp 1677580104
transform 1 0 70080 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_753
timestamp 1679581782
transform 1 0 72864 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_785
timestamp 1677580104
transform 1 0 75936 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679581782
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_821
timestamp 1677580104
transform 1 0 79392 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_4
timestamp 1677579658
transform 1 0 960 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_36
timestamp 1677580104
transform 1 0 4032 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_43
timestamp 1677580104
transform 1 0 4704 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_45
timestamp 1677579658
transform 1 0 4896 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_50
timestamp 1679581782
transform 1 0 5376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_57
timestamp 1679581782
transform 1 0 6048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_64
timestamp 1679581782
transform 1 0 6720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_71
timestamp 1679581782
transform 1 0 7392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_78
timestamp 1679581782
transform 1 0 8064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_85
timestamp 1679581782
transform 1 0 8736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_92
timestamp 1679581782
transform 1 0 9408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_99
timestamp 1679581782
transform 1 0 10080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_106
timestamp 1679581782
transform 1 0 10752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_113
timestamp 1679581782
transform 1 0 11424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_120
timestamp 1679581782
transform 1 0 12096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_127
timestamp 1679581782
transform 1 0 12768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_134
timestamp 1679581782
transform 1 0 13440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_141
timestamp 1679581782
transform 1 0 14112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_148
timestamp 1679581782
transform 1 0 14784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_155
timestamp 1679581782
transform 1 0 15456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_162
timestamp 1679581782
transform 1 0 16128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_169
timestamp 1679581782
transform 1 0 16800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_176
timestamp 1679581782
transform 1 0 17472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_183
timestamp 1679581782
transform 1 0 18144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_190
timestamp 1679581782
transform 1 0 18816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_197
timestamp 1679581782
transform 1 0 19488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_204
timestamp 1679581782
transform 1 0 20160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_211
timestamp 1679581782
transform 1 0 20832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_218
timestamp 1679581782
transform 1 0 21504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_225
timestamp 1679581782
transform 1 0 22176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_232
timestamp 1679581782
transform 1 0 22848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_239
timestamp 1679581782
transform 1 0 23520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_246
timestamp 1679581782
transform 1 0 24192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_253
timestamp 1679581782
transform 1 0 24864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_260
timestamp 1679581782
transform 1 0 25536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_267
timestamp 1679581782
transform 1 0 26208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_274
timestamp 1679581782
transform 1 0 26880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_281
timestamp 1679581782
transform 1 0 27552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_288
timestamp 1679581782
transform 1 0 28224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_295
timestamp 1679581782
transform 1 0 28896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_302
timestamp 1679581782
transform 1 0 29568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_309
timestamp 1679581782
transform 1 0 30240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_316
timestamp 1679577901
transform 1 0 30912 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_320
timestamp 1677580104
transform 1 0 31296 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_331
timestamp 1679581782
transform 1 0 32352 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_338
timestamp 1677580104
transform 1 0 33024 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_340
timestamp 1677579658
transform 1 0 33216 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_351
timestamp 1679577901
transform 1 0 34272 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_355
timestamp 1677580104
transform 1 0 34656 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_362
timestamp 1677579658
transform 1 0 35328 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_367
timestamp 1679577901
transform 1 0 35808 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_387
timestamp 1677579658
transform 1 0 37728 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_396
timestamp 1679577901
transform 1 0 38592 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_4  FILLER_19_423
timestamp 1679577901
transform 1 0 41184 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_427
timestamp 1677580104
transform 1 0 41568 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_434
timestamp 1679581782
transform 1 0 42240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679581782
transform 1 0 42912 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_448
timestamp 1677580104
transform 1 0 43584 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_454
timestamp 1679581782
transform 1 0 44160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_461
timestamp 1679577901
transform 1 0 44832 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_465
timestamp 1677580104
transform 1 0 45216 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_477
timestamp 1679581782
transform 1 0 46368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_484
timestamp 1679577901
transform 1 0 47040 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_496
timestamp 1677580104
transform 1 0 48192 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_502
timestamp 1677580104
transform 1 0 48768 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_504
timestamp 1677579658
transform 1 0 48960 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_509
timestamp 1679577901
transform 1 0 49440 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_513
timestamp 1677579658
transform 1 0 49824 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_544
timestamp 1677580104
transform 1 0 52800 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_573
timestamp 1679581782
transform 1 0 55584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_580
timestamp 1679581782
transform 1 0 56256 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_587
timestamp 1677579658
transform 1 0 56928 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_615
timestamp 1679577901
transform 1 0 59616 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_619
timestamp 1677579658
transform 1 0 60000 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679581782
transform 1 0 63072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679581782
transform 1 0 63744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_665
timestamp 1679577901
transform 1 0 64416 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_673
timestamp 1677580104
transform 1 0 65184 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_706
timestamp 1677580104
transform 1 0 68352 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_708
timestamp 1677579658
transform 1 0 68544 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_713
timestamp 1679577901
transform 1 0 69024 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_717
timestamp 1677580104
transform 1 0 69408 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_740
timestamp 1679581782
transform 1 0 71616 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_747
timestamp 1677580104
transform 1 0 72288 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_749
timestamp 1677579658
transform 1 0 72480 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_754
timestamp 1679581782
transform 1 0 72960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_761
timestamp 1679581782
transform 1 0 73632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_768
timestamp 1679581782
transform 1 0 74304 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_775
timestamp 1677579658
transform 1 0 74976 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_780
timestamp 1679581782
transform 1 0 75456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_787
timestamp 1679577901
transform 1 0 76128 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_791
timestamp 1677579658
transform 1 0 76512 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_796
timestamp 1679581782
transform 1 0 76992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_803
timestamp 1679581782
transform 1 0 77664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_810
timestamp 1679581782
transform 1 0 78336 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_817
timestamp 1677580104
transform 1 0 79008 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_819
timestamp 1677579658
transform 1 0 79200 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_4
timestamp 1679577901
transform 1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_8
timestamp 1677580104
transform 1 0 1344 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_27
timestamp 1677580104
transform 1 0 3168 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_68
timestamp 1679581782
transform 1 0 7104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_75
timestamp 1679581782
transform 1 0 7776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_82
timestamp 1679581782
transform 1 0 8448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_89
timestamp 1679581782
transform 1 0 9120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_96
timestamp 1679581782
transform 1 0 9792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_103
timestamp 1679581782
transform 1 0 10464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_110
timestamp 1679581782
transform 1 0 11136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_117
timestamp 1679581782
transform 1 0 11808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_124
timestamp 1679581782
transform 1 0 12480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_131
timestamp 1679581782
transform 1 0 13152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_138
timestamp 1679581782
transform 1 0 13824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_145
timestamp 1679581782
transform 1 0 14496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_152
timestamp 1679581782
transform 1 0 15168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_159
timestamp 1679581782
transform 1 0 15840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_166
timestamp 1679581782
transform 1 0 16512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_173
timestamp 1679581782
transform 1 0 17184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_180
timestamp 1679581782
transform 1 0 17856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_187
timestamp 1679581782
transform 1 0 18528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_194
timestamp 1679581782
transform 1 0 19200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_201
timestamp 1679581782
transform 1 0 19872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_208
timestamp 1679581782
transform 1 0 20544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_215
timestamp 1679581782
transform 1 0 21216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_222
timestamp 1679581782
transform 1 0 21888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_229
timestamp 1679581782
transform 1 0 22560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_236
timestamp 1679581782
transform 1 0 23232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_243
timestamp 1679581782
transform 1 0 23904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_250
timestamp 1679581782
transform 1 0 24576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_257
timestamp 1679581782
transform 1 0 25248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_264
timestamp 1679581782
transform 1 0 25920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_271
timestamp 1679581782
transform 1 0 26592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_278
timestamp 1679581782
transform 1 0 27264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_285
timestamp 1679581782
transform 1 0 27936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_292
timestamp 1679581782
transform 1 0 28608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_299
timestamp 1679581782
transform 1 0 29280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_306
timestamp 1679581782
transform 1 0 29952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_313
timestamp 1679577901
transform 1 0 30624 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_358
timestamp 1679581782
transform 1 0 34944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_365
timestamp 1679581782
transform 1 0 35616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_372
timestamp 1679577901
transform 1 0 36288 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_391
timestamp 1679581782
transform 1 0 38112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_398
timestamp 1679581782
transform 1 0 38784 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_405
timestamp 1677580104
transform 1 0 39456 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_407
timestamp 1677579658
transform 1 0 39648 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_439
timestamp 1677580104
transform 1 0 42720 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_477
timestamp 1677580104
transform 1 0 46368 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_479
timestamp 1677579658
transform 1 0 46560 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_488
timestamp 1679581782
transform 1 0 47424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_495
timestamp 1679577901
transform 1 0 48096 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_499
timestamp 1677579658
transform 1 0 48480 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_527
timestamp 1677580104
transform 1 0 51168 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_529
timestamp 1677579658
transform 1 0 51360 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_535
timestamp 1677579658
transform 1 0 51936 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_572
timestamp 1677579658
transform 1 0 55488 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_576
timestamp 1677579658
transform 1 0 55872 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_580
timestamp 1677580104
transform 1 0 56256 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_585
timestamp 1677579658
transform 1 0 56736 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_589
timestamp 1677579658
transform 1 0 57120 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_606
timestamp 1677579658
transform 1 0 58752 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_610
timestamp 1677579658
transform 1 0 59136 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_614
timestamp 1677579658
transform 1 0 59520 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_618
timestamp 1677579658
transform 1 0 59904 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_622
timestamp 1677579658
transform 1 0 60288 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_652
timestamp 1677579658
transform 1 0 63168 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_656
timestamp 1677579658
transform 1 0 63552 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_660
timestamp 1677579658
transform 1 0 63936 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_664
timestamp 1677579658
transform 1 0 64320 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_668
timestamp 1677580104
transform 1 0 64704 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_673
timestamp 1677579658
transform 1 0 65184 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_677
timestamp 1677579658
transform 1 0 65568 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_681
timestamp 1677579658
transform 1 0 65952 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_685
timestamp 1677579658
transform 1 0 66336 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_689
timestamp 1677580104
transform 1 0 66720 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_694
timestamp 1677579658
transform 1 0 67200 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_698
timestamp 1677579658
transform 1 0 67584 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_702
timestamp 1677579658
transform 1 0 67968 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_706
timestamp 1677579658
transform 1 0 68352 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_710
timestamp 1677579658
transform 1 0 68736 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_714
timestamp 1677580104
transform 1 0 69120 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_719
timestamp 1677579658
transform 1 0 69600 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_723
timestamp 1677579658
transform 1 0 69984 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_727
timestamp 1677579658
transform 1 0 70368 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_731
timestamp 1677579658
transform 1 0 70752 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_735
timestamp 1677579658
transform 1 0 71136 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_739
timestamp 1677580104
transform 1 0 71520 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_744
timestamp 1677579658
transform 1 0 72000 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_748
timestamp 1677579658
transform 1 0 72384 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_752
timestamp 1677579658
transform 1 0 72768 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_756
timestamp 1677579658
transform 1 0 73152 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_760
timestamp 1677579658
transform 1 0 73536 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_764
timestamp 1677580104
transform 1 0 73920 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_769
timestamp 1677579658
transform 1 0 74400 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_773
timestamp 1677579658
transform 1 0 74784 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_777
timestamp 1677579658
transform 1 0 75168 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_781
timestamp 1677579658
transform 1 0 75552 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_785
timestamp 1679577901
transform 1 0 75936 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_789
timestamp 1677579658
transform 1 0 76320 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_793
timestamp 1677579658
transform 1 0 76704 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_800
timestamp 1677579658
transform 1 0 77376 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_804
timestamp 1677579658
transform 1 0 77760 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_811
timestamp 1677579658
transform 1 0 78432 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_821
timestamp 1677580104
transform 1 0 79392 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_18
timestamp 1679577901
transform 1 0 2304 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_30
timestamp 1679581782
transform 1 0 3456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_45
timestamp 1679581782
transform 1 0 4896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_52
timestamp 1679581782
transform 1 0 5568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_59
timestamp 1679581782
transform 1 0 6240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_66
timestamp 1679581782
transform 1 0 6912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_73
timestamp 1679581782
transform 1 0 7584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_80
timestamp 1679581782
transform 1 0 8256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_87
timestamp 1679581782
transform 1 0 8928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_94
timestamp 1679581782
transform 1 0 9600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_101
timestamp 1679581782
transform 1 0 10272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_108
timestamp 1679581782
transform 1 0 10944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_115
timestamp 1679581782
transform 1 0 11616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_122
timestamp 1679581782
transform 1 0 12288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_129
timestamp 1679581782
transform 1 0 12960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_136
timestamp 1679581782
transform 1 0 13632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_143
timestamp 1679581782
transform 1 0 14304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_150
timestamp 1679581782
transform 1 0 14976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_157
timestamp 1679581782
transform 1 0 15648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_164
timestamp 1679581782
transform 1 0 16320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_171
timestamp 1679581782
transform 1 0 16992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_178
timestamp 1679581782
transform 1 0 17664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_185
timestamp 1679581782
transform 1 0 18336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_192
timestamp 1679581782
transform 1 0 19008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_199
timestamp 1679581782
transform 1 0 19680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_206
timestamp 1679581782
transform 1 0 20352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_213
timestamp 1679581782
transform 1 0 21024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_220
timestamp 1679581782
transform 1 0 21696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_227
timestamp 1679581782
transform 1 0 22368 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_234
timestamp 1677579658
transform 1 0 23040 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_247
timestamp 1679581782
transform 1 0 24288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_254
timestamp 1679581782
transform 1 0 24960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_261
timestamp 1679581782
transform 1 0 25632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_268
timestamp 1679581782
transform 1 0 26304 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_275
timestamp 1677580104
transform 1 0 26976 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_285
timestamp 1679581782
transform 1 0 27936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_292
timestamp 1679581782
transform 1 0 28608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_299
timestamp 1679581782
transform 1 0 29280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_306
timestamp 1679577901
transform 1 0 29952 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_21_318
timestamp 1679577901
transform 1 0 31104 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_326
timestamp 1679581782
transform 1 0 31872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_333
timestamp 1679581782
transform 1 0 32544 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_340
timestamp 1677579658
transform 1 0 33216 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_377
timestamp 1677579658
transform 1 0 36768 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_409
timestamp 1679581782
transform 1 0 39840 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_416
timestamp 1677580104
transform 1 0 40512 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_418
timestamp 1677579658
transform 1 0 40704 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_446
timestamp 1677579658
transform 1 0 43392 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_455
timestamp 1677580104
transform 1 0 44256 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_502
timestamp 1677580104
transform 1 0 48768 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_504
timestamp 1677579658
transform 1 0 48960 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_510
timestamp 1677579658
transform 1 0 49536 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_516
timestamp 1677579658
transform 1 0 50112 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_535
timestamp 1677580104
transform 1 0 51936 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_537
timestamp 1677579658
transform 1 0 52128 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_158
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_165
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_172
timestamp 1679581782
transform 1 0 17088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_179
timestamp 1679581782
transform 1 0 17760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_186
timestamp 1679581782
transform 1 0 18432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_193
timestamp 1679581782
transform 1 0 19104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_200
timestamp 1679581782
transform 1 0 19776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_207
timestamp 1679581782
transform 1 0 20448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_214
timestamp 1679581782
transform 1 0 21120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_221
timestamp 1679581782
transform 1 0 21792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_264
timestamp 1679581782
transform 1 0 25920 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_303
timestamp 1677579658
transform 1 0 29664 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_336
timestamp 1679577901
transform 1 0 32832 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_22_344
timestamp 1679577901
transform 1 0 33600 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_348
timestamp 1677579658
transform 1 0 33984 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_353
timestamp 1677580104
transform 1 0 34464 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_355
timestamp 1677579658
transform 1 0 34656 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_360
timestamp 1679581782
transform 1 0 35136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_367
timestamp 1679577901
transform 1 0 35808 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_371
timestamp 1677580104
transform 1 0 36192 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_381
timestamp 1679581782
transform 1 0 37152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_392
timestamp 1679581782
transform 1 0 38208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_399
timestamp 1679577901
transform 1 0 38880 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_403
timestamp 1677579658
transform 1 0 39264 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_435
timestamp 1677580104
transform 1 0 42336 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_469
timestamp 1677579658
transform 1 0 45600 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_483
timestamp 1679581782
transform 1 0 46944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_490
timestamp 1679581782
transform 1 0 47616 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_497
timestamp 1677580104
transform 1 0 48288 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_499
timestamp 1677579658
transform 1 0 48480 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_505
timestamp 1677580104
transform 1 0 49056 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_507
timestamp 1677579658
transform 1 0 49248 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_4
timestamp 1679577901
transform 1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_8
timestamp 1677579658
transform 1 0 1344 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_13
timestamp 1679581782
transform 1 0 1824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_20
timestamp 1679581782
transform 1 0 2496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_27
timestamp 1679581782
transform 1 0 3168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_34
timestamp 1679581782
transform 1 0 3840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_41
timestamp 1679581782
transform 1 0 4512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_48
timestamp 1679581782
transform 1 0 5184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_55
timestamp 1679581782
transform 1 0 5856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_62
timestamp 1679581782
transform 1 0 6528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_69
timestamp 1679581782
transform 1 0 7200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_76
timestamp 1679581782
transform 1 0 7872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_83
timestamp 1679581782
transform 1 0 8544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_90
timestamp 1679581782
transform 1 0 9216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_97
timestamp 1679577901
transform 1 0 9888 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_101
timestamp 1677580104
transform 1 0 10272 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_117
timestamp 1677580104
transform 1 0 11808 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679581782
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679581782
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679581782
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679581782
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679581782
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679581782
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679581782
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_172
timestamp 1679581782
transform 1 0 17088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_179
timestamp 1679581782
transform 1 0 17760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_186
timestamp 1679581782
transform 1 0 18432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_193
timestamp 1679581782
transform 1 0 19104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_200
timestamp 1679581782
transform 1 0 19776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_207
timestamp 1679581782
transform 1 0 20448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_214
timestamp 1679581782
transform 1 0 21120 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_221
timestamp 1677579658
transform 1 0 21792 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_256
timestamp 1677580104
transform 1 0 25152 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_258
timestamp 1677579658
transform 1 0 25344 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_263
timestamp 1677580104
transform 1 0 25824 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_265
timestamp 1677579658
transform 1 0 26016 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_271
timestamp 1677579658
transform 1 0 26592 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_286
timestamp 1679577901
transform 1 0 28032 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_290
timestamp 1677580104
transform 1 0 28416 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_297
timestamp 1679577901
transform 1 0 29088 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_301
timestamp 1677579658
transform 1 0 29472 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_329
timestamp 1677580104
transform 1 0 32160 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_363
timestamp 1677580104
transform 1 0 35424 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_424
timestamp 1677580104
transform 1 0 41280 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_444
timestamp 1677580104
transform 1 0 43200 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_446
timestamp 1677579658
transform 1 0 43392 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_460
timestamp 1679581782
transform 1 0 44736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_467
timestamp 1679581782
transform 1 0 45408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_474
timestamp 1679577901
transform 1 0 46080 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_478
timestamp 1677580104
transform 1 0 46464 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_485
timestamp 1677580104
transform 1 0 47136 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_492
timestamp 1679577901
transform 1 0 47808 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_510
timestamp 1677580104
transform 1 0 49536 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_516
timestamp 1677579658
transform 1 0 50112 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_521
timestamp 1677579658
transform 1 0 50592 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_534
timestamp 1679577901
transform 1 0 51840 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_81
timestamp 1679577901
transform 1 0 8352 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_85
timestamp 1677579658
transform 1 0 8736 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_113
timestamp 1677580104
transform 1 0 11424 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_115
timestamp 1677579658
transform 1 0 11616 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_148
timestamp 1679581782
transform 1 0 14784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_155
timestamp 1679581782
transform 1 0 15456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_162
timestamp 1679581782
transform 1 0 16128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_169
timestamp 1679581782
transform 1 0 16800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_176
timestamp 1679581782
transform 1 0 17472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_183
timestamp 1679581782
transform 1 0 18144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_190
timestamp 1679581782
transform 1 0 18816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_197
timestamp 1679581782
transform 1 0 19488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_204
timestamp 1679581782
transform 1 0 20160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_211
timestamp 1679581782
transform 1 0 20832 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_218
timestamp 1677580104
transform 1 0 21504 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_330
timestamp 1679577901
transform 1 0 32256 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_334
timestamp 1677579658
transform 1 0 32640 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_349
timestamp 1679581782
transform 1 0 34080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_356
timestamp 1679581782
transform 1 0 34752 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_363
timestamp 1677580104
transform 1 0 35424 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_383
timestamp 1679581782
transform 1 0 37344 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_390
timestamp 1677579658
transform 1 0 38016 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_410
timestamp 1677580104
transform 1 0 39936 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_425
timestamp 1677579658
transform 1 0 41376 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_435
timestamp 1677580104
transform 1 0 42336 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_437
timestamp 1677579658
transform 1 0 42528 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_502
timestamp 1677579658
transform 1 0 48768 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_508
timestamp 1677580104
transform 1 0 49344 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_537
timestamp 1679581782
transform 1 0 52128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_39
timestamp 1677580104
transform 1 0 4320 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_48
timestamp 1679581782
transform 1 0 5184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_55
timestamp 1679581782
transform 1 0 5856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_62
timestamp 1679581782
transform 1 0 6528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_69
timestamp 1679581782
transform 1 0 7200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_76
timestamp 1679581782
transform 1 0 7872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_83
timestamp 1679581782
transform 1 0 8544 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_90
timestamp 1677579658
transform 1 0 9216 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_95
timestamp 1679581782
transform 1 0 9696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_102
timestamp 1679577901
transform 1 0 10368 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_106
timestamp 1677579658
transform 1 0 10752 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_117
timestamp 1679581782
transform 1 0 11808 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_124
timestamp 1677580104
transform 1 0 12480 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_130
timestamp 1679581782
transform 1 0 13056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_137
timestamp 1679581782
transform 1 0 13728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_144
timestamp 1679581782
transform 1 0 14400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_151
timestamp 1679581782
transform 1 0 15072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_158
timestamp 1679581782
transform 1 0 15744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_165
timestamp 1679581782
transform 1 0 16416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_172
timestamp 1679581782
transform 1 0 17088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_179
timestamp 1679581782
transform 1 0 17760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_186
timestamp 1679581782
transform 1 0 18432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_193
timestamp 1679581782
transform 1 0 19104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_200
timestamp 1679581782
transform 1 0 19776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_207
timestamp 1679581782
transform 1 0 20448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_214
timestamp 1679581782
transform 1 0 21120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_221
timestamp 1679581782
transform 1 0 21792 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_233
timestamp 1677579658
transform 1 0 22944 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_242
timestamp 1679581782
transform 1 0 23808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_249
timestamp 1679581782
transform 1 0 24480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_256
timestamp 1679581782
transform 1 0 25152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_263
timestamp 1679577901
transform 1 0 25824 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_267
timestamp 1677580104
transform 1 0 26208 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_278
timestamp 1679581782
transform 1 0 27264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_285
timestamp 1679581782
transform 1 0 27936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_292
timestamp 1679581782
transform 1 0 28608 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_299
timestamp 1677580104
transform 1 0 29280 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_310
timestamp 1679581782
transform 1 0 30336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_317
timestamp 1679581782
transform 1 0 31008 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_338
timestamp 1677580104
transform 1 0 33024 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_340
timestamp 1677579658
transform 1 0 33216 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_345
timestamp 1679581782
transform 1 0 33696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_352
timestamp 1679577901
transform 1 0 34368 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_361
timestamp 1677580104
transform 1 0 35232 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_373
timestamp 1679581782
transform 1 0 36384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_380
timestamp 1679581782
transform 1 0 37056 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_452
timestamp 1677580104
transform 1 0 43968 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_454
timestamp 1677579658
transform 1 0 44160 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_471
timestamp 1679581782
transform 1 0 45792 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_478
timestamp 1677580104
transform 1 0 46464 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_484
timestamp 1677580104
transform 1 0 47040 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_494
timestamp 1679581782
transform 1 0 48000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_501
timestamp 1679577901
transform 1 0 48672 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_509
timestamp 1679577901
transform 1 0 49440 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_513
timestamp 1677580104
transform 1 0 49824 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_519
timestamp 1679581782
transform 1 0 50400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_526
timestamp 1679581782
transform 1 0 51072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_533
timestamp 1679581782
transform 1 0 51744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_540
timestamp 1679577901
transform 1 0 52416 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_25
timestamp 1679577901
transform 1 0 2976 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_29
timestamp 1677579658
transform 1 0 3360 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_35
timestamp 1679581782
transform 1 0 3936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_42
timestamp 1679577901
transform 1 0 4608 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_50
timestamp 1679581782
transform 1 0 5376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_57
timestamp 1679581782
transform 1 0 6048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_64
timestamp 1679581782
transform 1 0 6720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_71
timestamp 1679581782
transform 1 0 7392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_78
timestamp 1679581782
transform 1 0 8064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_85
timestamp 1679581782
transform 1 0 8736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_92
timestamp 1679581782
transform 1 0 9408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_99
timestamp 1679581782
transform 1 0 10080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_106
timestamp 1679581782
transform 1 0 10752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_113
timestamp 1679581782
transform 1 0 11424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_120
timestamp 1679581782
transform 1 0 12096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_127
timestamp 1679581782
transform 1 0 12768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_134
timestamp 1679581782
transform 1 0 13440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_141
timestamp 1679581782
transform 1 0 14112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_148
timestamp 1679581782
transform 1 0 14784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_155
timestamp 1679581782
transform 1 0 15456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_162
timestamp 1679581782
transform 1 0 16128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_169
timestamp 1679581782
transform 1 0 16800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_176
timestamp 1679581782
transform 1 0 17472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_183
timestamp 1679581782
transform 1 0 18144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_190
timestamp 1679581782
transform 1 0 18816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_197
timestamp 1679581782
transform 1 0 19488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_204
timestamp 1679581782
transform 1 0 20160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_211
timestamp 1679581782
transform 1 0 20832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_218
timestamp 1679581782
transform 1 0 21504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_225
timestamp 1679581782
transform 1 0 22176 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_232
timestamp 1677579658
transform 1 0 22848 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_237
timestamp 1679581782
transform 1 0 23328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_244
timestamp 1679581782
transform 1 0 24000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_251
timestamp 1679581782
transform 1 0 24672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_258
timestamp 1679577901
transform 1 0 25344 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_262
timestamp 1677580104
transform 1 0 25728 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_280
timestamp 1677580104
transform 1 0 27456 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_282
timestamp 1677579658
transform 1 0 27648 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_298
timestamp 1679577901
transform 1 0 29184 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_302
timestamp 1677580104
transform 1 0 29568 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_308
timestamp 1679581782
transform 1 0 30144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_315
timestamp 1679581782
transform 1 0 30816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_322
timestamp 1679581782
transform 1 0 31488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_356
timestamp 1679577901
transform 1 0 34752 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_360
timestamp 1677579658
transform 1 0 35136 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_388
timestamp 1677580104
transform 1 0 37824 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_390
timestamp 1677579658
transform 1 0 38016 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_423
timestamp 1679581782
transform 1 0 41184 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_439
timestamp 1677579658
transform 1 0 42720 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_465
timestamp 1677580104
transform 1 0 45216 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_472
timestamp 1679577901
transform 1 0 45888 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_481
timestamp 1679581782
transform 1 0 46752 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_488
timestamp 1677580104
transform 1 0 47424 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_21
timestamp 1679577901
transform 1 0 2592 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_41
timestamp 1679581782
transform 1 0 4512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_48
timestamp 1679581782
transform 1 0 5184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_55
timestamp 1679581782
transform 1 0 5856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_62
timestamp 1679581782
transform 1 0 6528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_69
timestamp 1679581782
transform 1 0 7200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_76
timestamp 1679581782
transform 1 0 7872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_83
timestamp 1679581782
transform 1 0 8544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_90
timestamp 1679581782
transform 1 0 9216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_97
timestamp 1679581782
transform 1 0 9888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_104
timestamp 1679581782
transform 1 0 10560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_111
timestamp 1679581782
transform 1 0 11232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_118
timestamp 1679581782
transform 1 0 11904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_125
timestamp 1679581782
transform 1 0 12576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_132
timestamp 1679581782
transform 1 0 13248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_139
timestamp 1679581782
transform 1 0 13920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_146
timestamp 1679581782
transform 1 0 14592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_153
timestamp 1679581782
transform 1 0 15264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_160
timestamp 1679581782
transform 1 0 15936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_167
timestamp 1679581782
transform 1 0 16608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_174
timestamp 1679581782
transform 1 0 17280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_181
timestamp 1679581782
transform 1 0 17952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_188
timestamp 1679581782
transform 1 0 18624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_195
timestamp 1679581782
transform 1 0 19296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_202
timestamp 1679581782
transform 1 0 19968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_209
timestamp 1679581782
transform 1 0 20640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_216
timestamp 1679581782
transform 1 0 21312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_223
timestamp 1679581782
transform 1 0 21984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_230
timestamp 1679581782
transform 1 0 22656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_237
timestamp 1679581782
transform 1 0 23328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_244
timestamp 1679581782
transform 1 0 24000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_251
timestamp 1679581782
transform 1 0 24672 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_258
timestamp 1677579658
transform 1 0 25344 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_296
timestamp 1677580104
transform 1 0 28992 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_298
timestamp 1677579658
transform 1 0 29184 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_326
timestamp 1679577901
transform 1 0 31872 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_338
timestamp 1677580104
transform 1 0 33024 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_344
timestamp 1679581782
transform 1 0 33600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_351
timestamp 1679581782
transform 1 0 34272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_358
timestamp 1679581782
transform 1 0 34944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 36864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 37536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 38208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_408
timestamp 1679581782
transform 1 0 39744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_415
timestamp 1679581782
transform 1 0 40416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_426
timestamp 1679581782
transform 1 0 41472 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_433
timestamp 1677580104
transform 1 0 42144 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_499
timestamp 1677580104
transform 1 0 48480 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_501
timestamp 1677579658
transform 1 0 48672 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_507
timestamp 1677580104
transform 1 0 49248 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_532
timestamp 1679577901
transform 1 0 51648 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_536
timestamp 1677580104
transform 1 0 52032 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679581782
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679581782
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679581782
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679581782
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679581782
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679581782
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679581782
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679581782
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_144
timestamp 1679581782
transform 1 0 14400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_151
timestamp 1679581782
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_158
timestamp 1679581782
transform 1 0 15744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_165
timestamp 1679581782
transform 1 0 16416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_172
timestamp 1679581782
transform 1 0 17088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_179
timestamp 1679581782
transform 1 0 17760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_186
timestamp 1679581782
transform 1 0 18432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_193
timestamp 1679581782
transform 1 0 19104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_200
timestamp 1679581782
transform 1 0 19776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_207
timestamp 1679581782
transform 1 0 20448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_214
timestamp 1679581782
transform 1 0 21120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_221
timestamp 1679581782
transform 1 0 21792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_228
timestamp 1679581782
transform 1 0 22464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_235
timestamp 1679581782
transform 1 0 23136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_242
timestamp 1679581782
transform 1 0 23808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_249
timestamp 1679581782
transform 1 0 24480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_256
timestamp 1679581782
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_263
timestamp 1679581782
transform 1 0 25824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_270
timestamp 1679581782
transform 1 0 26496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_277
timestamp 1679577901
transform 1 0 27168 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_281
timestamp 1677579658
transform 1 0 27552 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_298
timestamp 1677580104
transform 1 0 29184 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_300
timestamp 1677579658
transform 1 0 29376 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_306
timestamp 1679577901
transform 1 0 29952 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_310
timestamp 1677580104
transform 1 0 30336 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_327
timestamp 1677579658
transform 1 0 31968 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_333
timestamp 1677580104
transform 1 0 32544 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_362
timestamp 1677580104
transform 1 0 35328 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_364
timestamp 1677579658
transform 1 0 35520 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_392
timestamp 1679577901
transform 1 0 38208 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_405
timestamp 1679581782
transform 1 0 39456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_412
timestamp 1679577901
transform 1 0 40128 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_416
timestamp 1677579658
transform 1 0 40512 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_449
timestamp 1679581782
transform 1 0 43680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_456
timestamp 1679577901
transform 1 0 44352 0 1 21924
box -48 -56 432 834
use sg13g2_decap_4  FILLER_28_473
timestamp 1679577901
transform 1 0 45984 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_481
timestamp 1679581782
transform 1 0 46752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_488
timestamp 1679581782
transform 1 0 47424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_504
timestamp 1679577901
transform 1 0 48960 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_513
timestamp 1677580104
transform 1 0 49824 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_515
timestamp 1677579658
transform 1 0 50016 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_524
timestamp 1679581782
transform 1 0 50880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_4
timestamp 1679577901
transform 1 0 960 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_17
timestamp 1679581782
transform 1 0 2208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_24
timestamp 1679581782
transform 1 0 2880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_31
timestamp 1679581782
transform 1 0 3552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_38
timestamp 1679581782
transform 1 0 4224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_45
timestamp 1679581782
transform 1 0 4896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_52
timestamp 1679581782
transform 1 0 5568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_59
timestamp 1679581782
transform 1 0 6240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_66
timestamp 1679581782
transform 1 0 6912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_73
timestamp 1679581782
transform 1 0 7584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_80
timestamp 1679581782
transform 1 0 8256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_87
timestamp 1679581782
transform 1 0 8928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_94
timestamp 1679581782
transform 1 0 9600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_101
timestamp 1679581782
transform 1 0 10272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_108
timestamp 1679581782
transform 1 0 10944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_115
timestamp 1679581782
transform 1 0 11616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_122
timestamp 1679581782
transform 1 0 12288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_129
timestamp 1679581782
transform 1 0 12960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_136
timestamp 1679581782
transform 1 0 13632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_143
timestamp 1679581782
transform 1 0 14304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_150
timestamp 1679581782
transform 1 0 14976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_157
timestamp 1679581782
transform 1 0 15648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_164
timestamp 1679581782
transform 1 0 16320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_171
timestamp 1679581782
transform 1 0 16992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_178
timestamp 1679581782
transform 1 0 17664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_185
timestamp 1679581782
transform 1 0 18336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_192
timestamp 1679581782
transform 1 0 19008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_199
timestamp 1679581782
transform 1 0 19680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_206
timestamp 1679581782
transform 1 0 20352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_213
timestamp 1679581782
transform 1 0 21024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_220
timestamp 1679581782
transform 1 0 21696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_227
timestamp 1679581782
transform 1 0 22368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_234
timestamp 1679581782
transform 1 0 23040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_241
timestamp 1679581782
transform 1 0 23712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_248
timestamp 1679581782
transform 1 0 24384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_255
timestamp 1679581782
transform 1 0 25056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_262
timestamp 1679581782
transform 1 0 25728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_269
timestamp 1679581782
transform 1 0 26400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_276
timestamp 1679581782
transform 1 0 27072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_283
timestamp 1679577901
transform 1 0 27744 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_287
timestamp 1677580104
transform 1 0 28128 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_321
timestamp 1677580104
transform 1 0 31392 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_323
timestamp 1677579658
transform 1 0 31584 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_337
timestamp 1679577901
transform 1 0 32928 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_345
timestamp 1679581782
transform 1 0 33696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_352
timestamp 1679581782
transform 1 0 34368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_359
timestamp 1679581782
transform 1 0 35040 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_384
timestamp 1677580104
transform 1 0 37440 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_386
timestamp 1677579658
transform 1 0 37632 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_392
timestamp 1677580104
transform 1 0 38208 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_435
timestamp 1679577901
transform 1 0 42336 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_439
timestamp 1677579658
transform 1 0 42720 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_444
timestamp 1679581782
transform 1 0 43200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_451
timestamp 1679581782
transform 1 0 43872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_463
timestamp 1679577901
transform 1 0 45024 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_29_503
timestamp 1679577901
transform 1 0 48864 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_507
timestamp 1677579658
transform 1 0 49248 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_4
timestamp 1679577901
transform 1 0 960 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_8
timestamp 1677580104
transform 1 0 1344 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_18
timestamp 1679581782
transform 1 0 2304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_25
timestamp 1679581782
transform 1 0 2976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_32
timestamp 1679581782
transform 1 0 3648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_39
timestamp 1679581782
transform 1 0 4320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_46
timestamp 1679581782
transform 1 0 4992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_53
timestamp 1679581782
transform 1 0 5664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_60
timestamp 1679581782
transform 1 0 6336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_67
timestamp 1679581782
transform 1 0 7008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_74
timestamp 1679581782
transform 1 0 7680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_81
timestamp 1679581782
transform 1 0 8352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_88
timestamp 1679581782
transform 1 0 9024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_95
timestamp 1679581782
transform 1 0 9696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_102
timestamp 1679581782
transform 1 0 10368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_109
timestamp 1679581782
transform 1 0 11040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_116
timestamp 1679581782
transform 1 0 11712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_123
timestamp 1679581782
transform 1 0 12384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_130
timestamp 1679581782
transform 1 0 13056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_137
timestamp 1679581782
transform 1 0 13728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_144
timestamp 1679581782
transform 1 0 14400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_151
timestamp 1679581782
transform 1 0 15072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_158
timestamp 1679581782
transform 1 0 15744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_165
timestamp 1679581782
transform 1 0 16416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_172
timestamp 1679581782
transform 1 0 17088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_179
timestamp 1679581782
transform 1 0 17760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_186
timestamp 1679581782
transform 1 0 18432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_193
timestamp 1679581782
transform 1 0 19104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_200
timestamp 1679581782
transform 1 0 19776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_207
timestamp 1679581782
transform 1 0 20448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_214
timestamp 1679581782
transform 1 0 21120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_221
timestamp 1679581782
transform 1 0 21792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_228
timestamp 1679581782
transform 1 0 22464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_235
timestamp 1679581782
transform 1 0 23136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_242
timestamp 1679581782
transform 1 0 23808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_249
timestamp 1679581782
transform 1 0 24480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_256
timestamp 1679581782
transform 1 0 25152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_263
timestamp 1679581782
transform 1 0 25824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_270
timestamp 1679581782
transform 1 0 26496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_277
timestamp 1679581782
transform 1 0 27168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_284
timestamp 1679581782
transform 1 0 27840 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_291
timestamp 1677580104
transform 1 0 28512 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_293
timestamp 1677579658
transform 1 0 28704 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_298
timestamp 1679581782
transform 1 0 29184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_305
timestamp 1679581782
transform 1 0 29856 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_312
timestamp 1677580104
transform 1 0 30528 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_314
timestamp 1677579658
transform 1 0 30720 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_334
timestamp 1677580104
transform 1 0 32640 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_367
timestamp 1677580104
transform 1 0 35808 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_379
timestamp 1679581782
transform 1 0 36960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_386
timestamp 1679581782
transform 1 0 37632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_393
timestamp 1679577901
transform 1 0 38304 0 1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_30_407
timestamp 1679577901
transform 1 0 39648 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_427
timestamp 1679581782
transform 1 0 41568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_434
timestamp 1679577901
transform 1 0 42240 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_438
timestamp 1677579658
transform 1 0 42624 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_443
timestamp 1679581782
transform 1 0 43104 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_450
timestamp 1677579658
transform 1 0 43776 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_475
timestamp 1679581782
transform 1 0 46176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_486
timestamp 1679581782
transform 1 0 47232 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_493
timestamp 1677579658
transform 1 0 47904 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_531
timestamp 1677579658
transform 1 0 51552 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_559
timestamp 1679577901
transform 1 0 54240 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_563
timestamp 1677579658
transform 1 0 54624 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_567
timestamp 1677579658
transform 1 0 55008 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_571
timestamp 1677580104
transform 1 0 55392 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_589
timestamp 1677579658
transform 1 0 57120 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_593
timestamp 1677579658
transform 1 0 57504 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_597
timestamp 1677579658
transform 1 0 57888 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_601
timestamp 1677579658
transform 1 0 58272 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_605
timestamp 1677579658
transform 1 0 58656 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_609
timestamp 1677580104
transform 1 0 59040 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_614
timestamp 1677579658
transform 1 0 59520 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_618
timestamp 1677579658
transform 1 0 59904 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_622
timestamp 1677579658
transform 1 0 60288 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_626
timestamp 1677579658
transform 1 0 60672 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_630
timestamp 1677580104
transform 1 0 61056 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_635
timestamp 1677579658
transform 1 0 61536 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_639
timestamp 1677579658
transform 1 0 61920 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_643
timestamp 1677579658
transform 1 0 62304 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_647
timestamp 1677579658
transform 1 0 62688 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_651
timestamp 1677579658
transform 1 0 63072 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_655
timestamp 1677579658
transform 1 0 63456 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_659
timestamp 1677580104
transform 1 0 63840 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_664
timestamp 1677579658
transform 1 0 64320 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_668
timestamp 1677579658
transform 1 0 64704 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_672
timestamp 1677579658
transform 1 0 65088 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_676
timestamp 1677580104
transform 1 0 65472 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_681
timestamp 1677579658
transform 1 0 65952 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_685
timestamp 1677579658
transform 1 0 66336 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_689
timestamp 1677579658
transform 1 0 66720 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_693
timestamp 1677579658
transform 1 0 67104 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_697
timestamp 1677579658
transform 1 0 67488 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_701
timestamp 1677580104
transform 1 0 67872 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_706
timestamp 1677579658
transform 1 0 68352 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_710
timestamp 1677579658
transform 1 0 68736 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_714
timestamp 1677579658
transform 1 0 69120 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_718
timestamp 1677579658
transform 1 0 69504 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_722
timestamp 1677580104
transform 1 0 69888 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_727
timestamp 1677579658
transform 1 0 70368 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_731
timestamp 1677579658
transform 1 0 70752 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_735
timestamp 1677579658
transform 1 0 71136 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_739
timestamp 1677579658
transform 1 0 71520 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_743
timestamp 1677579658
transform 1 0 71904 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_747
timestamp 1677579658
transform 1 0 72288 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_751
timestamp 1677579658
transform 1 0 72672 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_755
timestamp 1677580104
transform 1 0 73056 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_760
timestamp 1677579658
transform 1 0 73536 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_764
timestamp 1677579658
transform 1 0 73920 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_768
timestamp 1677579658
transform 1 0 74304 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_772
timestamp 1677579658
transform 1 0 74688 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_776
timestamp 1677579658
transform 1 0 75072 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_780
timestamp 1677579658
transform 1 0 75456 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_784
timestamp 1677580104
transform 1 0 75840 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_789
timestamp 1679577901
transform 1 0 76320 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_793
timestamp 1677579658
transform 1 0 76704 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_806
timestamp 1677579658
transform 1 0 77952 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_810
timestamp 1677579658
transform 1 0 78336 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_11
timestamp 1679581782
transform 1 0 1632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_18
timestamp 1679581782
transform 1 0 2304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_25
timestamp 1679581782
transform 1 0 2976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_32
timestamp 1679581782
transform 1 0 3648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_39
timestamp 1679581782
transform 1 0 4320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_46
timestamp 1679581782
transform 1 0 4992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_53
timestamp 1679581782
transform 1 0 5664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_60
timestamp 1679581782
transform 1 0 6336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_67
timestamp 1679581782
transform 1 0 7008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_74
timestamp 1679581782
transform 1 0 7680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_81
timestamp 1679581782
transform 1 0 8352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_88
timestamp 1679581782
transform 1 0 9024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_95
timestamp 1679581782
transform 1 0 9696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_102
timestamp 1679581782
transform 1 0 10368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_109
timestamp 1679581782
transform 1 0 11040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_116
timestamp 1679581782
transform 1 0 11712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_123
timestamp 1679581782
transform 1 0 12384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_130
timestamp 1679581782
transform 1 0 13056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_137
timestamp 1679581782
transform 1 0 13728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_144
timestamp 1679581782
transform 1 0 14400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_151
timestamp 1679581782
transform 1 0 15072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_158
timestamp 1679581782
transform 1 0 15744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_165
timestamp 1679581782
transform 1 0 16416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_172
timestamp 1679581782
transform 1 0 17088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_179
timestamp 1679581782
transform 1 0 17760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_186
timestamp 1679581782
transform 1 0 18432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_193
timestamp 1679581782
transform 1 0 19104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_200
timestamp 1679581782
transform 1 0 19776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_207
timestamp 1679581782
transform 1 0 20448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_214
timestamp 1679581782
transform 1 0 21120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_221
timestamp 1679581782
transform 1 0 21792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_228
timestamp 1679581782
transform 1 0 22464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_235
timestamp 1679581782
transform 1 0 23136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_242
timestamp 1679581782
transform 1 0 23808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_249
timestamp 1679581782
transform 1 0 24480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_256
timestamp 1679581782
transform 1 0 25152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_263
timestamp 1679581782
transform 1 0 25824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_270
timestamp 1679581782
transform 1 0 26496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_277
timestamp 1679581782
transform 1 0 27168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_284
timestamp 1679581782
transform 1 0 27840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_291
timestamp 1679581782
transform 1 0 28512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_298
timestamp 1679581782
transform 1 0 29184 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_305
timestamp 1677580104
transform 1 0 29856 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_307
timestamp 1677579658
transform 1 0 30048 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_312
timestamp 1679581782
transform 1 0 30528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_319
timestamp 1679577901
transform 1 0 31200 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_333
timestamp 1677579658
transform 1 0 32544 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_338
timestamp 1677579658
transform 1 0 33024 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_352
timestamp 1679577901
transform 1 0 34368 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_356
timestamp 1677579658
transform 1 0 34752 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_384
timestamp 1677580104
transform 1 0 37440 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_390
timestamp 1679581782
transform 1 0 38016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_397
timestamp 1679577901
transform 1 0 38688 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_31_428
timestamp 1679577901
transform 1 0 41664 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_432
timestamp 1677580104
transform 1 0 42048 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_466
timestamp 1679581782
transform 1 0 45312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_473
timestamp 1679581782
transform 1 0 45984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_485
timestamp 1679581782
transform 1 0 47136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_492
timestamp 1679581782
transform 1 0 47808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_503
timestamp 1679581782
transform 1 0 48864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_510
timestamp 1679577901
transform 1 0 49536 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_31_531
timestamp 1679577901
transform 1 0 51552 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_535
timestamp 1677579658
transform 1 0 51936 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_545
timestamp 1679581782
transform 1 0 52896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_552
timestamp 1679581782
transform 1 0 53568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_559
timestamp 1679577901
transform 1 0 54240 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_563
timestamp 1677580104
transform 1 0 54624 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_592
timestamp 1679577901
transform 1 0 57408 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_596
timestamp 1677580104
transform 1 0 57792 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_603
timestamp 1677580104
transform 1 0 58464 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_605
timestamp 1677579658
transform 1 0 58656 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_632
timestamp 1679581782
transform 1 0 61248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_639
timestamp 1679581782
transform 1 0 61920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_646
timestamp 1679581782
transform 1 0 62592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_653
timestamp 1679577901
transform 1 0 63264 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_657
timestamp 1677580104
transform 1 0 63648 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_676
timestamp 1679581782
transform 1 0 65472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_683
timestamp 1679581782
transform 1 0 66144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_690
timestamp 1679581782
transform 1 0 66816 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_697
timestamp 1677579658
transform 1 0 67488 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_711
timestamp 1679581782
transform 1 0 68832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_718
timestamp 1679581782
transform 1 0 69504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_725
timestamp 1679577901
transform 1 0 70176 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_729
timestamp 1677579658
transform 1 0 70560 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_743
timestamp 1679581782
transform 1 0 71904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_750
timestamp 1679581782
transform 1 0 72576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_757
timestamp 1679581782
transform 1 0 73248 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_764
timestamp 1677580104
transform 1 0 73920 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_766
timestamp 1677579658
transform 1 0 74112 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_772
timestamp 1679577901
transform 1 0 74688 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_776
timestamp 1677580104
transform 1 0 75072 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_788
timestamp 1677579658
transform 1 0 76224 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_793
timestamp 1679577901
transform 1 0 76704 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_801
timestamp 1679581782
transform 1 0 77472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_808
timestamp 1679581782
transform 1 0 78144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_815
timestamp 1679581782
transform 1 0 78816 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_822
timestamp 1677579658
transform 1 0 79488 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1679581782
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_39
timestamp 1679581782
transform 1 0 4320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 4992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 5664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_60
timestamp 1679581782
transform 1 0 6336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679581782
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679581782
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679581782
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679581782
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_109
timestamp 1679581782
transform 1 0 11040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_116
timestamp 1679581782
transform 1 0 11712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_123
timestamp 1679581782
transform 1 0 12384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_130
timestamp 1679581782
transform 1 0 13056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_137
timestamp 1679581782
transform 1 0 13728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_144
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_158
timestamp 1679581782
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679581782
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679581782
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679581782
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679581782
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679581782
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679581782
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679581782
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_221
timestamp 1679581782
transform 1 0 21792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679581782
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679581782
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_249
timestamp 1679581782
transform 1 0 24480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_256
timestamp 1679581782
transform 1 0 25152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_263
timestamp 1679581782
transform 1 0 25824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_270
timestamp 1679581782
transform 1 0 26496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_277
timestamp 1679581782
transform 1 0 27168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_284
timestamp 1679581782
transform 1 0 27840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_291
timestamp 1679581782
transform 1 0 28512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_298
timestamp 1679577901
transform 1 0 29184 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_302
timestamp 1677579658
transform 1 0 29568 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_330
timestamp 1679577901
transform 1 0 32256 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_334
timestamp 1677579658
transform 1 0 32640 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_343
timestamp 1679581782
transform 1 0 33504 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_350
timestamp 1677580104
transform 1 0 34176 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_362
timestamp 1677580104
transform 1 0 35328 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_364
timestamp 1677579658
transform 1 0 35520 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_370
timestamp 1679581782
transform 1 0 36096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_377
timestamp 1679577901
transform 1 0 36768 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_413
timestamp 1677579658
transform 1 0 40224 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_418
timestamp 1677579658
transform 1 0 40704 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_446
timestamp 1679581782
transform 1 0 43392 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_457
timestamp 1677580104
transform 1 0 44448 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_459
timestamp 1677579658
transform 1 0 44640 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_510
timestamp 1679581782
transform 1 0 49536 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_517
timestamp 1677580104
transform 1 0 50208 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_519
timestamp 1677579658
transform 1 0 50400 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_525
timestamp 1677580104
transform 1 0 50976 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_527
timestamp 1677579658
transform 1 0 51168 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_565
timestamp 1679577901
transform 1 0 54816 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_582
timestamp 1679581782
transform 1 0 56448 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_589
timestamp 1677580104
transform 1 0 57120 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_618
timestamp 1677580104
transform 1 0 59904 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_620
timestamp 1677579658
transform 1 0 60096 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_648
timestamp 1677580104
transform 1 0 62784 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_687
timestamp 1679577901
transform 1 0 66528 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_728
timestamp 1677579658
transform 1 0 70464 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_819
timestamp 1679577901
transform 1 0 79200 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_4
timestamp 1679581782
transform 1 0 960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_11
timestamp 1679581782
transform 1 0 1632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_18
timestamp 1679581782
transform 1 0 2304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_25
timestamp 1679581782
transform 1 0 2976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_32
timestamp 1679581782
transform 1 0 3648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_39
timestamp 1679581782
transform 1 0 4320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679581782
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_53
timestamp 1679581782
transform 1 0 5664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_60
timestamp 1679581782
transform 1 0 6336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_67
timestamp 1679581782
transform 1 0 7008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_74
timestamp 1679581782
transform 1 0 7680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_81
timestamp 1679581782
transform 1 0 8352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_88
timestamp 1679581782
transform 1 0 9024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_95
timestamp 1679581782
transform 1 0 9696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_102
timestamp 1679581782
transform 1 0 10368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_109
timestamp 1679581782
transform 1 0 11040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_116
timestamp 1679581782
transform 1 0 11712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_123
timestamp 1679581782
transform 1 0 12384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_130
timestamp 1679581782
transform 1 0 13056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_137
timestamp 1679581782
transform 1 0 13728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_144
timestamp 1679581782
transform 1 0 14400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_151
timestamp 1679581782
transform 1 0 15072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_158
timestamp 1679581782
transform 1 0 15744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_165
timestamp 1679581782
transform 1 0 16416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_172
timestamp 1679581782
transform 1 0 17088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_179
timestamp 1679581782
transform 1 0 17760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_186
timestamp 1679581782
transform 1 0 18432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_193
timestamp 1679581782
transform 1 0 19104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_200
timestamp 1679581782
transform 1 0 19776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_207
timestamp 1679581782
transform 1 0 20448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_214
timestamp 1679581782
transform 1 0 21120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_221
timestamp 1679581782
transform 1 0 21792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_228
timestamp 1679581782
transform 1 0 22464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_235
timestamp 1679581782
transform 1 0 23136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_242
timestamp 1679581782
transform 1 0 23808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_249
timestamp 1679581782
transform 1 0 24480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_256
timestamp 1679581782
transform 1 0 25152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_263
timestamp 1679581782
transform 1 0 25824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_270
timestamp 1679581782
transform 1 0 26496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_277
timestamp 1679581782
transform 1 0 27168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_284
timestamp 1679581782
transform 1 0 27840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_291
timestamp 1679581782
transform 1 0 28512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_298
timestamp 1679581782
transform 1 0 29184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_305
timestamp 1679581782
transform 1 0 29856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_312
timestamp 1679581782
transform 1 0 30528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_319
timestamp 1679581782
transform 1 0 31200 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_326
timestamp 1677580104
transform 1 0 31872 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_328
timestamp 1677579658
transform 1 0 32064 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_375
timestamp 1679581782
transform 1 0 36576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_382
timestamp 1679581782
transform 1 0 37248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_389
timestamp 1679581782
transform 1 0 37920 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_396
timestamp 1677580104
transform 1 0 38592 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_398
timestamp 1677579658
transform 1 0 38784 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_413
timestamp 1677580104
transform 1 0 40224 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_419
timestamp 1677580104
transform 1 0 40800 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_421
timestamp 1677579658
transform 1 0 40992 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_427
timestamp 1679577901
transform 1 0 41568 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_431
timestamp 1677579658
transform 1 0 41952 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_436
timestamp 1679581782
transform 1 0 42432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_443
timestamp 1679577901
transform 1 0 43104 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_447
timestamp 1677579658
transform 1 0 43488 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_475
timestamp 1677579658
transform 1 0 46176 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_528
timestamp 1677580104
transform 1 0 51264 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_534
timestamp 1677579658
transform 1 0 51840 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_547
timestamp 1679581782
transform 1 0 53088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_554
timestamp 1679581782
transform 1 0 53760 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_561
timestamp 1677580104
transform 1 0 54432 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_567
timestamp 1677580104
transform 1 0 55008 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_569
timestamp 1677579658
transform 1 0 55200 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_590
timestamp 1677580104
transform 1 0 57216 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_600
timestamp 1677579658
transform 1 0 58176 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_611
timestamp 1677579658
transform 1 0 59232 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_633
timestamp 1677580104
transform 1 0 61344 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_672
timestamp 1677580104
transform 1 0 65088 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_674
timestamp 1677579658
transform 1 0 65280 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_680
timestamp 1677580104
transform 1 0 65856 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_682
timestamp 1677579658
transform 1 0 66048 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_687
timestamp 1679577901
transform 1 0 66528 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_691
timestamp 1677580104
transform 1 0 66912 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_707
timestamp 1677579658
transform 1 0 68448 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_712
timestamp 1677580104
transform 1 0 68928 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_714
timestamp 1677579658
transform 1 0 69120 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_720
timestamp 1679581782
transform 1 0 69696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_745
timestamp 1679581782
transform 1 0 72096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_752
timestamp 1679577901
transform 1 0 72768 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_760
timestamp 1679577901
transform 1 0 73536 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_764
timestamp 1677580104
transform 1 0 73920 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_781
timestamp 1679581782
transform 1 0 75552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_788
timestamp 1679577901
transform 1 0 76224 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_792
timestamp 1677580104
transform 1 0 76608 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_799
timestamp 1679581782
transform 1 0 77280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_806
timestamp 1679581782
transform 1 0 77952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_813
timestamp 1679581782
transform 1 0 78624 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_820
timestamp 1677580104
transform 1 0 79296 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_822
timestamp 1677579658
transform 1 0 79488 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_35
timestamp 1677580104
transform 1 0 3936 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_40
timestamp 1679581782
transform 1 0 4416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_47
timestamp 1679581782
transform 1 0 5088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_54
timestamp 1679581782
transform 1 0 5760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_61
timestamp 1679581782
transform 1 0 6432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_68
timestamp 1679581782
transform 1 0 7104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_75
timestamp 1679581782
transform 1 0 7776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_82
timestamp 1679581782
transform 1 0 8448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_89
timestamp 1679581782
transform 1 0 9120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_96
timestamp 1679581782
transform 1 0 9792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_103
timestamp 1679581782
transform 1 0 10464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_110
timestamp 1679581782
transform 1 0 11136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_117
timestamp 1679581782
transform 1 0 11808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_124
timestamp 1679581782
transform 1 0 12480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_131
timestamp 1679581782
transform 1 0 13152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_138
timestamp 1679581782
transform 1 0 13824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_145
timestamp 1679581782
transform 1 0 14496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_152
timestamp 1679581782
transform 1 0 15168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_159
timestamp 1679581782
transform 1 0 15840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_166
timestamp 1679581782
transform 1 0 16512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_173
timestamp 1679581782
transform 1 0 17184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_180
timestamp 1679581782
transform 1 0 17856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_187
timestamp 1679581782
transform 1 0 18528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_194
timestamp 1679581782
transform 1 0 19200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_201
timestamp 1679581782
transform 1 0 19872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_208
timestamp 1679581782
transform 1 0 20544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_215
timestamp 1679581782
transform 1 0 21216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_222
timestamp 1679581782
transform 1 0 21888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_229
timestamp 1679581782
transform 1 0 22560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_236
timestamp 1679581782
transform 1 0 23232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_243
timestamp 1679581782
transform 1 0 23904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_250
timestamp 1679581782
transform 1 0 24576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_257
timestamp 1679581782
transform 1 0 25248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_264
timestamp 1679581782
transform 1 0 25920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_271
timestamp 1679581782
transform 1 0 26592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_278
timestamp 1679581782
transform 1 0 27264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_285
timestamp 1679581782
transform 1 0 27936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_292
timestamp 1679581782
transform 1 0 28608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_299
timestamp 1679581782
transform 1 0 29280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_306
timestamp 1679581782
transform 1 0 29952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_313
timestamp 1679581782
transform 1 0 30624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_320
timestamp 1679581782
transform 1 0 31296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_327
timestamp 1679581782
transform 1 0 31968 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_334
timestamp 1677579658
transform 1 0 32640 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_339
timestamp 1679581782
transform 1 0 33120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_346
timestamp 1679581782
transform 1 0 33792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_353
timestamp 1679581782
transform 1 0 34464 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_395
timestamp 1677579658
transform 1 0 38496 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_454
timestamp 1679577901
transform 1 0 44160 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_458
timestamp 1677579658
transform 1 0 44544 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_473
timestamp 1677580104
transform 1 0 45984 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_510
timestamp 1679577901
transform 1 0 49536 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_514
timestamp 1677579658
transform 1 0 49920 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_525
timestamp 1677579658
transform 1 0 50976 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_540
timestamp 1679581782
transform 1 0 52416 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_547
timestamp 1677580104
transform 1 0 53088 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_549
timestamp 1677579658
transform 1 0 53280 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_554
timestamp 1679577901
transform 1 0 53760 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_585
timestamp 1679581782
transform 1 0 56736 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_592
timestamp 1677579658
transform 1 0 57408 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_597
timestamp 1677580104
transform 1 0 57888 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_599
timestamp 1677579658
transform 1 0 58080 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_604
timestamp 1677580104
transform 1 0 58560 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_610
timestamp 1677580104
transform 1 0 59136 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_634
timestamp 1679577901
transform 1 0 61440 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_638
timestamp 1677580104
transform 1 0 61824 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679581782
transform 1 0 62400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679581782
transform 1 0 63072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_663
timestamp 1679581782
transform 1 0 64224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_670
timestamp 1679581782
transform 1 0 64896 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_677
timestamp 1677579658
transform 1 0 65568 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_710
timestamp 1677580104
transform 1 0 68736 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_712
timestamp 1677579658
transform 1 0 68928 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_748
timestamp 1679577901
transform 1 0 72384 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_752
timestamp 1677580104
transform 1 0 72768 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_371
timestamp 1677580104
transform 1 0 36192 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_377
timestamp 1679581782
transform 1 0 36768 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_384
timestamp 1677580104
transform 1 0 37440 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_418
timestamp 1677580104
transform 1 0 40704 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_428
timestamp 1679581782
transform 1 0 41664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_435
timestamp 1679581782
transform 1 0 42336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_442
timestamp 1679577901
transform 1 0 43008 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_446
timestamp 1677579658
transform 1 0 43392 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_493
timestamp 1679581782
transform 1 0 47904 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_500
timestamp 1677580104
transform 1 0 48576 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_529
timestamp 1677580104
transform 1 0 51360 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_578
timestamp 1679581782
transform 1 0 56064 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_585
timestamp 1677580104
transform 1 0 56736 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_587
timestamp 1677579658
transform 1 0 56928 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_620
timestamp 1677580104
transform 1 0 60096 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_622
timestamp 1677579658
transform 1 0 60288 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_650
timestamp 1679581782
transform 1 0 62976 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_657
timestamp 1677579658
transform 1 0 63648 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_663
timestamp 1679581782
transform 1 0 64224 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_670
timestamp 1677580104
transform 1 0 64896 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_681
timestamp 1677580104
transform 1 0 65952 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_687
timestamp 1679581782
transform 1 0 66528 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_694
timestamp 1677579658
transform 1 0 67200 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_699
timestamp 1679581782
transform 1 0 67680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_710
timestamp 1679577901
transform 1 0 68736 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_728
timestamp 1677579658
transform 1 0 70464 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_738
timestamp 1679577901
transform 1 0 71424 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_746
timestamp 1679581782
transform 1 0 72192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_753
timestamp 1679577901
transform 1 0 72864 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_757
timestamp 1677580104
transform 1 0 73248 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_763
timestamp 1679581782
transform 1 0 73824 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_770
timestamp 1677580104
transform 1 0 74496 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_772
timestamp 1677579658
transform 1 0 74688 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_778
timestamp 1677579658
transform 1 0 75264 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_784
timestamp 1679581782
transform 1 0 75840 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_791
timestamp 1677580104
transform 1 0 76512 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_805
timestamp 1679581782
transform 1 0 77856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_812
timestamp 1679581782
transform 1 0 78528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_819
timestamp 1679577901
transform 1 0 79200 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_385
timestamp 1679577901
transform 1 0 37536 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_389
timestamp 1677580104
transform 1 0 37920 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_395
timestamp 1679581782
transform 1 0 38496 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_402
timestamp 1677580104
transform 1 0 39168 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_417
timestamp 1677580104
transform 1 0 40608 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_459
timestamp 1677580104
transform 1 0 44640 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_461
timestamp 1677579658
transform 1 0 44832 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_472
timestamp 1679581782
transform 1 0 45888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_479
timestamp 1679581782
transform 1 0 46560 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_486
timestamp 1677580104
transform 1 0 47232 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_492
timestamp 1679581782
transform 1 0 47808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_499
timestamp 1679577901
transform 1 0 48480 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_503
timestamp 1677579658
transform 1 0 48864 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_523
timestamp 1677580104
transform 1 0 50784 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_529
timestamp 1677580104
transform 1 0 51360 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_531
timestamp 1677579658
transform 1 0 51552 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_583
timestamp 1677580104
transform 1 0 56544 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_589
timestamp 1679581782
transform 1 0 57120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_596
timestamp 1679577901
transform 1 0 57792 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_600
timestamp 1677580104
transform 1 0 58176 0 1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_36_632
timestamp 1679577901
transform 1 0 61248 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_636
timestamp 1677580104
transform 1 0 61632 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_675
timestamp 1677580104
transform 1 0 65376 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_677
timestamp 1677579658
transform 1 0 65568 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_709
timestamp 1679581782
transform 1 0 68640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_716
timestamp 1679577901
transform 1 0 69312 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_720
timestamp 1677579658
transform 1 0 69696 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_735
timestamp 1677580104
transform 1 0 71136 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_764
timestamp 1679581782
transform 1 0 73920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_771
timestamp 1679577901
transform 1 0 74592 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_775
timestamp 1677580104
transform 1 0 74976 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_782
timestamp 1679581782
transform 1 0 75648 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_789
timestamp 1677580104
transform 1 0 76320 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_791
timestamp 1677579658
transform 1 0 76512 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_805
timestamp 1679581782
transform 1 0 77856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_812
timestamp 1679581782
transform 1 0 78528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_819
timestamp 1679577901
transform 1 0 79200 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_392
timestamp 1677579658
transform 1 0 38208 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_439
timestamp 1679581782
transform 1 0 42720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_446
timestamp 1679581782
transform 1 0 43392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_453
timestamp 1679581782
transform 1 0 44064 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_460
timestamp 1677579658
transform 1 0 44736 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_466
timestamp 1679577901
transform 1 0 45312 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_470
timestamp 1677580104
transform 1 0 45696 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_503
timestamp 1679577901
transform 1 0 48864 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_507
timestamp 1677580104
transform 1 0 49248 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_577
timestamp 1677580104
transform 1 0 55968 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_579
timestamp 1677579658
transform 1 0 56160 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_607
timestamp 1677580104
transform 1 0 58848 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_618
timestamp 1677580104
transform 1 0 59904 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_620
timestamp 1677579658
transform 1 0 60096 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_634
timestamp 1679581782
transform 1 0 61440 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_641
timestamp 1677580104
transform 1 0 62112 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_647
timestamp 1679577901
transform 1 0 62688 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_651
timestamp 1677580104
transform 1 0 63072 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_663
timestamp 1679581782
transform 1 0 64224 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_674
timestamp 1677580104
transform 1 0 65280 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_676
timestamp 1677579658
transform 1 0 65472 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_682
timestamp 1679581782
transform 1 0 66048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_689
timestamp 1679581782
transform 1 0 66720 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_696
timestamp 1677580104
transform 1 0 67392 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_698
timestamp 1677579658
transform 1 0 67584 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_735
timestamp 1677579658
transform 1 0 71136 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_744
timestamp 1679581782
transform 1 0 72000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_751
timestamp 1679581782
transform 1 0 72672 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_795
timestamp 1677579658
transform 1 0 76896 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_392
timestamp 1679577901
transform 1 0 38208 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_396
timestamp 1677580104
transform 1 0 38592 0 1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_38_402
timestamp 1679577901
transform 1 0 39168 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_406
timestamp 1677580104
transform 1 0 39552 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_421
timestamp 1677580104
transform 1 0 40992 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_423
timestamp 1677579658
transform 1 0 41184 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_428
timestamp 1679581782
transform 1 0 41664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_435
timestamp 1679581782
transform 1 0 42336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_442
timestamp 1679577901
transform 1 0 43008 0 1 29484
box -48 -56 432 834
use sg13g2_decap_4  FILLER_38_487
timestamp 1679577901
transform 1 0 47328 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_38_554
timestamp 1679581782
transform 1 0 53760 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_570
timestamp 1677579658
transform 1 0 55296 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_580
timestamp 1679581782
transform 1 0 56256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_587
timestamp 1679581782
transform 1 0 56928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_594
timestamp 1679581782
transform 1 0 57600 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_601
timestamp 1677579658
transform 1 0 58272 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_661
timestamp 1679581782
transform 1 0 64032 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_668
timestamp 1677580104
transform 1 0 64704 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_670
timestamp 1677579658
transform 1 0 64896 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_708
timestamp 1679577901
transform 1 0 68544 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_712
timestamp 1677579658
transform 1 0 68928 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_727
timestamp 1677580104
transform 1 0 70368 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_729
timestamp 1677579658
transform 1 0 70560 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_748
timestamp 1679581782
transform 1 0 72384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_755
timestamp 1679581782
transform 1 0 73056 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_762
timestamp 1677579658
transform 1 0 73728 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_767
timestamp 1679577901
transform 1 0 74208 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_771
timestamp 1677580104
transform 1 0 74592 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_787
timestamp 1677580104
transform 1 0 76128 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_789
timestamp 1677579658
transform 1 0 76320 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_794
timestamp 1677580104
transform 1 0 76800 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_801
timestamp 1677579658
transform 1 0 77472 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_806
timestamp 1679581782
transform 1 0 77952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_813
timestamp 1679581782
transform 1 0 78624 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_820
timestamp 1677580104
transform 1 0 79296 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_822
timestamp 1677579658
transform 1 0 79488 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_413
timestamp 1679577901
transform 1 0 40224 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_39_421
timestamp 1679577901
transform 1 0 40992 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_39_430
timestamp 1679577901
transform 1 0 41856 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_447
timestamp 1677580104
transform 1 0 43488 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_463
timestamp 1679581782
transform 1 0 45024 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_470
timestamp 1677580104
transform 1 0 45696 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_472
timestamp 1677579658
transform 1 0 45888 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_478
timestamp 1677580104
transform 1 0 46464 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_480
timestamp 1677579658
transform 1 0 46656 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_485
timestamp 1679581782
transform 1 0 47136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_492
timestamp 1679577901
transform 1 0 47808 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_4  FILLER_39_500
timestamp 1679577901
transform 1 0 48576 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_504
timestamp 1677580104
transform 1 0 48960 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_515
timestamp 1677579658
transform 1 0 50016 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_536
timestamp 1679581782
transform 1 0 52032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_543
timestamp 1679577901
transform 1 0 52704 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_547
timestamp 1677580104
transform 1 0 53088 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679581782
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_560
timestamp 1677580104
transform 1 0 54336 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_581
timestamp 1677580104
transform 1 0 56352 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_587
timestamp 1679581782
transform 1 0 56928 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_594
timestamp 1677580104
transform 1 0 57600 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_596
timestamp 1677579658
transform 1 0 57792 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679581782
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_644
timestamp 1679577901
transform 1 0 62400 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_648
timestamp 1677580104
transform 1 0 62784 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_685
timestamp 1677579658
transform 1 0 66336 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_690
timestamp 1679581782
transform 1 0 66816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_697
timestamp 1679581782
transform 1 0 67488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_767
timestamp 1679577901
transform 1 0 74208 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_771
timestamp 1677580104
transform 1 0 74592 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_783
timestamp 1677580104
transform 1 0 75744 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_785
timestamp 1677579658
transform 1 0 75936 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_406
timestamp 1679577901
transform 1 0 39552 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_410
timestamp 1677580104
transform 1 0 39936 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_454
timestamp 1679581782
transform 1 0 44160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_461
timestamp 1679581782
transform 1 0 44832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_468
timestamp 1679581782
transform 1 0 45504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_475
timestamp 1679577901
transform 1 0 46176 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_497
timestamp 1677580104
transform 1 0 48288 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_508
timestamp 1677580104
transform 1 0 49344 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_510
timestamp 1677579658
transform 1 0 49536 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_535
timestamp 1679581782
transform 1 0 51936 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_542
timestamp 1677580104
transform 1 0 52608 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_571
timestamp 1677580104
transform 1 0 55392 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_605
timestamp 1679581782
transform 1 0 58656 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_612
timestamp 1677580104
transform 1 0 59328 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_623
timestamp 1677580104
transform 1 0 60384 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_629
timestamp 1679581782
transform 1 0 60960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_636
timestamp 1679581782
transform 1 0 61632 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_643
timestamp 1677579658
transform 1 0 62304 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_649
timestamp 1677579658
transform 1 0 62880 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_659
timestamp 1679581782
transform 1 0 63840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_666
timestamp 1679581782
transform 1 0 64512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_673
timestamp 1679581782
transform 1 0 65184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_680
timestamp 1679577901
transform 1 0 65856 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_697
timestamp 1679581782
transform 1 0 67488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_704
timestamp 1679577901
transform 1 0 68160 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_708
timestamp 1677579658
transform 1 0 68544 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_713
timestamp 1679581782
transform 1 0 69024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_720
timestamp 1679581782
transform 1 0 69696 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_727
timestamp 1677579658
transform 1 0 70368 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_750
timestamp 1679581782
transform 1 0 72576 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_757
timestamp 1677580104
transform 1 0 73248 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_759
timestamp 1677579658
transform 1 0 73440 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_787
timestamp 1679581782
transform 1 0 76128 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_794
timestamp 1677579658
transform 1 0 76800 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_799
timestamp 1677579658
transform 1 0 77280 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_808
timestamp 1679581782
transform 1 0 78144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_815
timestamp 1679581782
transform 1 0 78816 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_822
timestamp 1677579658
transform 1 0 79488 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_413
timestamp 1679577901
transform 1 0 40224 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_421
timestamp 1679581782
transform 1 0 40992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_428
timestamp 1679577901
transform 1 0 41664 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_432
timestamp 1677580104
transform 1 0 42048 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_439
timestamp 1677579658
transform 1 0 42720 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_444
timestamp 1677579658
transform 1 0 43200 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_472
timestamp 1677579658
transform 1 0 45888 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_522
timestamp 1679577901
transform 1 0 50688 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_4  FILLER_41_553
timestamp 1679577901
transform 1 0 53664 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_557
timestamp 1677579658
transform 1 0 54048 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_568
timestamp 1679577901
transform 1 0 55104 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_572
timestamp 1677579658
transform 1 0 55488 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_577
timestamp 1679581782
transform 1 0 55968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_584
timestamp 1679581782
transform 1 0 56640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_591
timestamp 1679581782
transform 1 0 57312 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_598
timestamp 1677580104
transform 1 0 57984 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_619
timestamp 1677580104
transform 1 0 60000 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_621
timestamp 1677579658
transform 1 0 60192 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_668
timestamp 1679581782
transform 1 0 64704 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_675
timestamp 1677580104
transform 1 0 65376 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_677
timestamp 1677579658
transform 1 0 65568 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_715
timestamp 1679577901
transform 1 0 69216 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_719
timestamp 1677579658
transform 1 0 69600 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_735
timestamp 1679577901
transform 1 0 71136 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_753
timestamp 1679581782
transform 1 0 72864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_760
timestamp 1679577901
transform 1 0 73536 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_764
timestamp 1677579658
transform 1 0 73920 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_769
timestamp 1679581782
transform 1 0 74400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_776
timestamp 1679581782
transform 1 0 75072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_788
timestamp 1679581782
transform 1 0 76224 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_795
timestamp 1677579658
transform 1 0 76896 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_434
timestamp 1679577901
transform 1 0 42240 0 1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_442
timestamp 1679581782
transform 1 0 43008 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_449
timestamp 1677579658
transform 1 0 43680 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_454
timestamp 1679581782
transform 1 0 44160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_461
timestamp 1679581782
transform 1 0 44832 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_468
timestamp 1677580104
transform 1 0 45504 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_470
timestamp 1677579658
transform 1 0 45696 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_494
timestamp 1679577901
transform 1 0 48000 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_529
timestamp 1677580104
transform 1 0 51360 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_544
timestamp 1679577901
transform 1 0 52800 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_548
timestamp 1677580104
transform 1 0 53184 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_555
timestamp 1679577901
transform 1 0 53856 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_559
timestamp 1677579658
transform 1 0 54240 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_596
timestamp 1677580104
transform 1 0 57792 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_634
timestamp 1679581782
transform 1 0 61440 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_641
timestamp 1677580104
transform 1 0 62112 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_743
timestamp 1677580104
transform 1 0 71904 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_813
timestamp 1679581782
transform 1 0 78624 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_820
timestamp 1677580104
transform 1 0 79296 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_822
timestamp 1677579658
transform 1 0 79488 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_476
timestamp 1679577901
transform 1 0 46272 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_485
timestamp 1679581782
transform 1 0 47136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_492
timestamp 1679581782
transform 1 0 47808 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_499
timestamp 1677580104
transform 1 0 48480 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_501
timestamp 1677579658
transform 1 0 48672 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679581782
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679581782
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_525
timestamp 1679577901
transform 1 0 50976 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_529
timestamp 1677580104
transform 1 0 51360 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_572
timestamp 1677580104
transform 1 0 55488 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_574
timestamp 1677579658
transform 1 0 55680 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_579
timestamp 1679581782
transform 1 0 56160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_586
timestamp 1679581782
transform 1 0 56832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_593
timestamp 1679581782
transform 1 0 57504 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_600
timestamp 1677579658
transform 1 0 58176 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_614
timestamp 1679581782
transform 1 0 59520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_621
timestamp 1679581782
transform 1 0 60192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_628
timestamp 1679581782
transform 1 0 60864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_635
timestamp 1679577901
transform 1 0 61536 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_639
timestamp 1677580104
transform 1 0 61920 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_654
timestamp 1677580104
transform 1 0 63360 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_656
timestamp 1677579658
transform 1 0 63552 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_661
timestamp 1679581782
transform 1 0 64032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_668
timestamp 1679581782
transform 1 0 64704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_675
timestamp 1679581782
transform 1 0 65376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_695
timestamp 1679581782
transform 1 0 67296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_702
timestamp 1679581782
transform 1 0 67968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_709
timestamp 1679581782
transform 1 0 68640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_716
timestamp 1679577901
transform 1 0 69312 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_720
timestamp 1677579658
transform 1 0 69696 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_725
timestamp 1679581782
transform 1 0 70176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_732
timestamp 1679581782
transform 1 0 70848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_756
timestamp 1679581782
transform 1 0 73152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_763
timestamp 1679581782
transform 1 0 73824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_770
timestamp 1679577901
transform 1 0 74496 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_4  FILLER_43_778
timestamp 1679577901
transform 1 0 75264 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_797
timestamp 1677579658
transform 1 0 77088 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_803
timestamp 1677579658
transform 1 0 77664 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_808
timestamp 1679581782
transform 1 0 78144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_815
timestamp 1679581782
transform 1 0 78816 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_822
timestamp 1677579658
transform 1 0 79488 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_469
timestamp 1679577901
transform 1 0 45600 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_473
timestamp 1677579658
transform 1 0 45984 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_518
timestamp 1677579658
transform 1 0 50304 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_529
timestamp 1679577901
transform 1 0 51360 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_542
timestamp 1679581782
transform 1 0 52608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_549
timestamp 1679577901
transform 1 0 53280 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_553
timestamp 1677579658
transform 1 0 53664 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_559
timestamp 1679581782
transform 1 0 54240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_566
timestamp 1679577901
transform 1 0 54912 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_584
timestamp 1679581782
transform 1 0 56640 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_591
timestamp 1677579658
transform 1 0 57312 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_624
timestamp 1679581782
transform 1 0 60480 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_631
timestamp 1677580104
transform 1 0 61152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_633
timestamp 1677579658
transform 1 0 61344 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_644
timestamp 1677580104
transform 1 0 62400 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_678
timestamp 1679577901
transform 1 0 65664 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_687
timestamp 1677580104
transform 1 0 66528 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_689
timestamp 1677579658
transform 1 0 66720 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_703
timestamp 1679581782
transform 1 0 68064 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_737
timestamp 1677580104
transform 1 0 71328 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_775
timestamp 1679577901
transform 1 0 74976 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_779
timestamp 1677579658
transform 1 0 75360 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_809
timestamp 1679581782
transform 1 0 78240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_816
timestamp 1679581782
transform 1 0 78912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_483
timestamp 1677579658
transform 1 0 46944 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_488
timestamp 1679581782
transform 1 0 47424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_495
timestamp 1679577901
transform 1 0 48096 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_545
timestamp 1679581782
transform 1 0 52896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_552
timestamp 1679581782
transform 1 0 53568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_559
timestamp 1679577901
transform 1 0 54240 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_563
timestamp 1677579658
transform 1 0 54624 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_600
timestamp 1677580104
transform 1 0 58176 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_606
timestamp 1679581782
transform 1 0 58752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_613
timestamp 1679577901
transform 1 0 59424 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_654
timestamp 1677580104
transform 1 0 63360 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_660
timestamp 1679581782
transform 1 0 63936 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_667
timestamp 1677580104
transform 1 0 64608 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_673
timestamp 1679581782
transform 1 0 65184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_721
timestamp 1679577901
transform 1 0 69792 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_725
timestamp 1677579658
transform 1 0 70176 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_746
timestamp 1677580104
transform 1 0 72192 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_748
timestamp 1677579658
transform 1 0 72384 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_753
timestamp 1679577901
transform 1 0 72864 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_4  FILLER_45_761
timestamp 1679577901
transform 1 0 73632 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_765
timestamp 1677579658
transform 1 0 74016 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_793
timestamp 1677580104
transform 1 0 76704 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_795
timestamp 1677579658
transform 1 0 76896 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_508
timestamp 1679581782
transform 1 0 49344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_515
timestamp 1679581782
transform 1 0 50016 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_526
timestamp 1677580104
transform 1 0 51072 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_532
timestamp 1677580104
transform 1 0 51648 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_534
timestamp 1677579658
transform 1 0 51840 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_562
timestamp 1679581782
transform 1 0 54528 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_569
timestamp 1677580104
transform 1 0 55200 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_571
timestamp 1677579658
transform 1 0 55392 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_590
timestamp 1679581782
transform 1 0 57216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_597
timestamp 1679577901
transform 1 0 57888 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_601
timestamp 1677580104
transform 1 0 58272 0 1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_46_616
timestamp 1679577901
transform 1 0 59712 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_620
timestamp 1677580104
transform 1 0 60096 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_626
timestamp 1679581782
transform 1 0 60672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_633
timestamp 1679577901
transform 1 0 61344 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_637
timestamp 1677580104
transform 1 0 61728 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_658
timestamp 1679577901
transform 1 0 63744 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_662
timestamp 1677580104
transform 1 0 64128 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_696
timestamp 1679581782
transform 1 0 67392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_703
timestamp 1679581782
transform 1 0 68064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_710
timestamp 1679577901
transform 1 0 68736 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_714
timestamp 1677579658
transform 1 0 69120 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_724
timestamp 1679581782
transform 1 0 70080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_731
timestamp 1679581782
transform 1 0 70752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_747
timestamp 1679577901
transform 1 0 72288 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_769
timestamp 1679581782
transform 1 0 74400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_776
timestamp 1679581782
transform 1 0 75072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_783
timestamp 1679577901
transform 1 0 75744 0 1 35532
box -48 -56 432 834
use sg13g2_decap_4  FILLER_46_792
timestamp 1679577901
transform 1 0 76608 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_808
timestamp 1679581782
transform 1 0 78144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_815
timestamp 1679581782
transform 1 0 78816 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_822
timestamp 1677579658
transform 1 0 79488 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_539
timestamp 1677579658
transform 1 0 52320 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_544
timestamp 1679581782
transform 1 0 52800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_551
timestamp 1679581782
transform 1 0 53472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_558
timestamp 1679577901
transform 1 0 54144 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_562
timestamp 1677579658
transform 1 0 54528 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_595
timestamp 1679577901
transform 1 0 57696 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_646
timestamp 1677580104
transform 1 0 62592 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_666
timestamp 1679581782
transform 1 0 64512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_673
timestamp 1679581782
transform 1 0 65184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_680
timestamp 1679577901
transform 1 0 65856 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_684
timestamp 1677580104
transform 1 0 66240 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_691
timestamp 1677580104
transform 1 0 66912 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_698
timestamp 1677579658
transform 1 0 67584 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_722
timestamp 1679581782
transform 1 0 69888 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_729
timestamp 1677580104
transform 1 0 70560 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_731
timestamp 1677579658
transform 1 0 70752 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_567
timestamp 1677579658
transform 1 0 55008 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_572
timestamp 1677580104
transform 1 0 55488 0 1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_48_625
timestamp 1679577901
transform 1 0 60576 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_629
timestamp 1677579658
transform 1 0 60960 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_711
timestamp 1677580104
transform 1 0 68832 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_713
timestamp 1677579658
transform 1 0 69024 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_741
timestamp 1679581782
transform 1 0 71712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_748
timestamp 1679577901
transform 1 0 72384 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_772
timestamp 1677580104
transform 1 0 74688 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_814
timestamp 1679581782
transform 1 0 78720 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_821
timestamp 1677580104
transform 1 0 79392 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_578
timestamp 1679577901
transform 1 0 56064 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_582
timestamp 1677580104
transform 1 0 56448 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_595
timestamp 1679577901
transform 1 0 57696 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_599
timestamp 1677580104
transform 1 0 58080 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_613
timestamp 1679581782
transform 1 0 59424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679581782
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_627
timestamp 1679581782
transform 1 0 60768 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_634
timestamp 1677579658
transform 1 0 61440 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_639
timestamp 1679581782
transform 1 0 61920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_646
timestamp 1679581782
transform 1 0 62592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_658
timestamp 1679577901
transform 1 0 63744 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_666
timestamp 1679581782
transform 1 0 64512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_673
timestamp 1679581782
transform 1 0 65184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_680
timestamp 1679577901
transform 1 0 65856 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_4  FILLER_49_688
timestamp 1679577901
transform 1 0 66624 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_719
timestamp 1677579658
transform 1 0 69600 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_745
timestamp 1679581782
transform 1 0 72096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_752
timestamp 1679581782
transform 1 0 72768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_759
timestamp 1679581782
transform 1 0 73440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_779
timestamp 1679577901
transform 1 0 75360 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_783
timestamp 1677579658
transform 1 0 75744 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_788
timestamp 1679577901
transform 1 0 76224 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_792
timestamp 1677580104
transform 1 0 76608 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_804
timestamp 1679581782
transform 1 0 77760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_811
timestamp 1679581782
transform 1 0 78432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_818
timestamp 1679577901
transform 1 0 79104 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_822
timestamp 1677579658
transform 1 0 79488 0 -1 38556
box -48 -56 144 834
use sg13g2_tiehi  heichips25_pudding_458
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_459
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_460
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_461
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_462
timestamp 1680000651
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_463
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_464
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 1344 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 1344 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use analog_wires  wires
timestamp 0
transform 1 0 80000 0 1 800
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 99920 21586 100000 21726 0 FreeSans 640 0 0 0 i_in
port 4 nsew signal bidirectional
flabel metal3 s 99920 19949 100000 20089 0 FreeSans 640 0 0 0 i_out
port 5 nsew signal bidirectional
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 6 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 7 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 8 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 9 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 10 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 11 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 12 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 13 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 14 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 15 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 16 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 17 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 18 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 19 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 20 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 21 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 22 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 23 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 24 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 25 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 26 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 27 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 28 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 29 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 30 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 31 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 32 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 33 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 34 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 35 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 36 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 37 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 38 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 39 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 40 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 41 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 42 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 43 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 44 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 45 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 46 nsew signal output
rlabel via5 65100 22479 65100 22479 0 VGND
rlabel via5 78980 19603 78980 19603 0 VPWR
rlabel metal2 54048 16926 54048 16926 0 _0000_
rlabel metal2 64734 22764 64734 22764 0 _0001_
rlabel metal2 64342 22764 64342 22764 0 _0002_
rlabel metal2 63950 22764 63950 22764 0 _0003_
rlabel metal2 63565 22828 63565 22828 0 _0004_
rlabel metal2 63165 22828 63165 22828 0 _0005_
rlabel metal2 62726 22764 62726 22764 0 _0006_
rlabel metal2 62334 22764 62334 22764 0 _0007_
rlabel metal2 61942 22764 61942 22764 0 _0008_
rlabel metal2 61550 22764 61550 22764 0 _0009_
rlabel metal2 61165 22828 61165 22828 0 _0010_
rlabel metal2 58080 16758 58080 16758 0 _0011_
rlabel metal2 60670 22764 60670 22764 0 _0012_
rlabel metal2 60365 22828 60365 22828 0 _0013_
rlabel metal2 59934 22764 59934 22764 0 _0014_
rlabel metal2 59542 22764 59542 22764 0 _0015_
rlabel metal2 59150 22764 59150 22764 0 _0016_
rlabel metal2 58765 22828 58765 22828 0 _0017_
rlabel metal2 58270 22764 58270 22764 0 _0018_
rlabel metal2 57965 22828 57965 22828 0 _0019_
rlabel metal2 57565 22828 57565 22828 0 _0020_
rlabel metal2 57142 22764 57142 22764 0 _0021_
rlabel metal2 58368 16758 58368 16758 0 _0022_
rlabel metal2 56750 22764 56750 22764 0 _0023_
rlabel metal2 56365 22828 56365 22828 0 _0024_
rlabel metal2 55965 22828 55965 22828 0 _0025_
rlabel metal2 55526 22764 55526 22764 0 _0026_
rlabel metal2 55165 22828 55165 22828 0 _0027_
rlabel metal2 54765 22828 54765 22828 0 _0028_
rlabel metal2 54365 22828 54365 22828 0 _0029_
rlabel metal2 53965 22690 53965 22690 0 _0030_
rlabel metal2 58656 16758 58656 16758 0 _0031_
rlabel metal2 59040 16590 59040 16590 0 _0032_
rlabel metal2 59520 16044 59520 16044 0 _0033_
rlabel metal2 59904 16044 59904 16044 0 _0034_
rlabel metal2 60192 16590 60192 16590 0 _0035_
rlabel metal2 60576 16590 60576 16590 0 _0036_
rlabel metal3 61056 16464 61056 16464 0 _0037_
rlabel metal2 61536 16758 61536 16758 0 _0038_
rlabel metal3 54528 17094 54528 17094 0 _0039_
rlabel metal2 62208 16758 62208 16758 0 _0040_
rlabel metal2 62496 16758 62496 16758 0 _0041_
rlabel metal2 62784 16758 62784 16758 0 _0042_
rlabel metal2 63072 16758 63072 16758 0 _0043_
rlabel metal2 63456 16758 63456 16758 0 _0044_
rlabel metal2 63840 16170 63840 16170 0 _0045_
rlabel metal2 64320 16044 64320 16044 0 _0046_
rlabel metal2 64608 16800 64608 16800 0 _0047_
rlabel metal2 65088 16758 65088 16758 0 _0048_
rlabel metal2 65472 16758 65472 16758 0 _0049_
rlabel metal2 54816 16758 54816 16758 0 _0050_
rlabel metal2 65856 16758 65856 16758 0 _0051_
rlabel metal2 66336 16044 66336 16044 0 _0052_
rlabel metal2 66624 16800 66624 16800 0 _0053_
rlabel metal2 67104 16758 67104 16758 0 _0054_
rlabel metal2 67584 16464 67584 16464 0 _0055_
rlabel metal2 67872 16758 67872 16758 0 _0056_
rlabel metal2 68256 16758 68256 16758 0 _0057_
rlabel metal2 68736 16044 68736 16044 0 _0058_
rlabel metal2 69024 16590 69024 16590 0 _0059_
rlabel metal2 69504 16758 69504 16758 0 _0060_
rlabel metal2 55104 16758 55104 16758 0 _0061_
rlabel metal2 69888 16758 69888 16758 0 _0062_
rlabel metal2 70272 16758 70272 16758 0 _0063_
rlabel metal2 70656 16758 70656 16758 0 _0064_
rlabel metal2 71040 16758 71040 16758 0 _0065_
rlabel metal2 71424 16800 71424 16800 0 _0066_
rlabel metal2 71904 16758 71904 16758 0 _0067_
rlabel metal2 72288 16758 72288 16758 0 _0068_
rlabel metal2 72672 16758 72672 16758 0 _0069_
rlabel metal2 73056 16758 73056 16758 0 _0070_
rlabel metal2 73536 16758 73536 16758 0 _0071_
rlabel metal2 55392 16758 55392 16758 0 _0072_
rlabel metal2 73920 16044 73920 16044 0 _0073_
rlabel metal2 74304 16758 74304 16758 0 _0074_
rlabel metal2 74784 16464 74784 16464 0 _0075_
rlabel metal2 75072 16758 75072 16758 0 _0076_
rlabel metal2 75456 16758 75456 16758 0 _0077_
rlabel metal2 75936 16044 75936 16044 0 _0078_
rlabel metal2 76512 16758 76512 16758 0 _0079_
rlabel metal2 76896 16758 76896 16758 0 _0080_
rlabel metal2 77280 16758 77280 16758 0 _0081_
rlabel metal2 77664 16758 77664 16758 0 _0082_
rlabel metal2 55776 16758 55776 16758 0 _0083_
rlabel metal2 78048 16758 78048 16758 0 _0084_
rlabel metal2 78336 16758 78336 16758 0 _0085_
rlabel metal2 78720 16758 78720 16758 0 _0086_
rlabel metal2 79296 16800 79296 16800 0 _0087_
rlabel metal2 79165 22828 79165 22828 0 _0088_
rlabel metal2 78765 22828 78765 22828 0 _0089_
rlabel metal2 78350 22764 78350 22764 0 _0090_
rlabel metal2 77965 22828 77965 22828 0 _0091_
rlabel metal2 77565 22828 77565 22828 0 _0092_
rlabel metal2 77165 22828 77165 22828 0 _0093_
rlabel metal2 56304 16044 56304 16044 0 _0094_
rlabel metal2 76765 22828 76765 22828 0 _0095_
rlabel metal2 76365 22828 76365 22828 0 _0096_
rlabel metal2 75950 22764 75950 22764 0 _0097_
rlabel metal2 75565 22828 75565 22828 0 _0098_
rlabel metal2 75165 22828 75165 22828 0 _0099_
rlabel metal2 74765 22828 74765 22828 0 _0100_
rlabel metal2 74334 22764 74334 22764 0 _0101_
rlabel metal2 73942 22764 73942 22764 0 _0102_
rlabel metal2 73550 22764 73550 22764 0 _0103_
rlabel metal2 73165 22828 73165 22828 0 _0104_
rlabel metal2 56640 16590 56640 16590 0 _0105_
rlabel metal2 72670 22764 72670 22764 0 _0106_
rlabel metal2 72326 22764 72326 22764 0 _0107_
rlabel metal2 71934 22764 71934 22764 0 _0108_
rlabel metal2 71542 22764 71542 22764 0 _0109_
rlabel metal2 71150 22764 71150 22764 0 _0110_
rlabel metal2 70765 22828 70765 22828 0 _0111_
rlabel metal2 70365 22828 70365 22828 0 _0112_
rlabel metal2 69926 22764 69926 22764 0 _0113_
rlabel metal2 69534 22764 69534 22764 0 _0114_
rlabel metal2 69142 22764 69142 22764 0 _0115_
rlabel metal2 57120 16044 57120 16044 0 _0116_
rlabel metal2 68750 22764 68750 22764 0 _0117_
rlabel metal2 68365 22828 68365 22828 0 _0118_
rlabel metal2 67965 22828 67965 22828 0 _0119_
rlabel metal2 67526 22764 67526 22764 0 _0120_
rlabel metal2 67134 22764 67134 22764 0 _0121_
rlabel metal2 66742 22764 66742 22764 0 _0122_
rlabel metal2 66350 22764 66350 22764 0 _0123_
rlabel metal2 65965 22828 65965 22828 0 _0124_
rlabel metal2 65565 22828 65565 22828 0 _0125_
rlabel metal2 65126 22764 65126 22764 0 _0126_
rlabel metal2 57408 16590 57408 16590 0 _0127_
rlabel metal2 22608 19236 22608 19236 0 _0128_
rlabel metal2 26304 18942 26304 18942 0 _0129_
rlabel metal2 29280 19320 29280 19320 0 _0130_
rlabel metal2 32304 20244 32304 20244 0 _0131_
rlabel metal2 35520 20244 35520 20244 0 _0132_
rlabel metal2 38688 20832 38688 20832 0 _0133_
rlabel metal3 41808 19152 41808 19152 0 _0134_
rlabel metal3 40896 17724 40896 17724 0 _0135_
rlabel metal3 40944 13104 40944 13104 0 _0136_
rlabel metal2 39840 14784 39840 14784 0 _0137_
rlabel metal3 37008 14700 37008 14700 0 _0138_
rlabel metal2 33984 15792 33984 15792 0 _0139_
rlabel metal2 32832 13482 32832 13482 0 _0140_
rlabel metal3 34368 11928 34368 11928 0 _0141_
rlabel metal3 36864 10164 36864 10164 0 _0142_
rlabel metal2 40224 9702 40224 9702 0 _0143_
rlabel metal2 41568 8652 41568 8652 0 _0144_
rlabel metal3 44544 8148 44544 8148 0 _0145_
rlabel metal2 45408 7434 45408 7434 0 _0146_
rlabel metal3 46608 5040 46608 5040 0 _0147_
rlabel metal2 50304 3780 50304 3780 0 _0148_
rlabel metal2 52512 6006 52512 6006 0 _0149_
rlabel metal2 52896 7266 52896 7266 0 _0150_
rlabel metal3 51168 10164 51168 10164 0 _0151_
rlabel metal2 50592 10920 50592 10920 0 _0152_
rlabel metal3 46800 11928 46800 11928 0 _0153_
rlabel metal2 46176 13734 46176 13734 0 _0154_
rlabel metal2 46080 15792 46080 15792 0 _0155_
rlabel metal3 46656 18396 46656 18396 0 _0156_
rlabel metal2 48672 16254 48672 16254 0 _0157_
rlabel metal2 51456 13734 51456 13734 0 _0158_
rlabel metal2 54624 13482 54624 13482 0 _0159_
rlabel metal3 55728 12600 55728 12600 0 _0160_
rlabel metal3 57312 10416 57312 10416 0 _0161_
rlabel metal2 55968 8316 55968 8316 0 _0162_
rlabel metal3 57504 6300 57504 6300 0 _0163_
rlabel metal2 58944 5250 58944 5250 0 _0164_
rlabel metal3 56784 3528 56784 3528 0 _0165_
rlabel metal3 54480 1344 54480 1344 0 _0166_
rlabel metal2 59088 1344 59088 1344 0 _0167_
rlabel metal3 62160 1344 62160 1344 0 _0168_
rlabel metal2 62880 3822 62880 3822 0 _0169_
rlabel metal2 64704 5250 64704 5250 0 _0170_
rlabel metal2 62208 7434 62208 7434 0 _0171_
rlabel metal3 63552 9576 63552 9576 0 _0172_
rlabel metal2 63360 11298 63360 11298 0 _0173_
rlabel metal2 61200 13440 61200 13440 0 _0174_
rlabel metal2 64560 13440 64560 13440 0 _0175_
rlabel metal4 68352 14112 68352 14112 0 _0176_
rlabel metal3 68160 11928 68160 11928 0 _0177_
rlabel metal2 66912 9828 66912 9828 0 _0178_
rlabel metal3 68880 8064 68880 8064 0 _0179_
rlabel metal3 69552 5880 69552 5880 0 _0180_
rlabel metal3 66720 1092 66720 1092 0 _0181_
rlabel metal3 69216 3612 69216 3612 0 _0182_
rlabel metal3 71952 1344 71952 1344 0 _0183_
rlabel metal2 75648 1848 75648 1848 0 _0184_
rlabel metal3 74544 3528 74544 3528 0 _0185_
rlabel metal3 74976 5544 74976 5544 0 _0186_
rlabel metal3 74976 8064 74976 8064 0 _0187_
rlabel metal2 76032 9198 76032 9198 0 _0188_
rlabel metal2 72576 11382 72576 11382 0 _0189_
rlabel metal2 74400 12894 74400 12894 0 _0190_
rlabel metal2 72192 14322 72192 14322 0 _0191_
rlabel metal2 73248 25620 73248 25620 0 _0192_
rlabel metal2 74880 27132 74880 27132 0 _0193_
rlabel metal2 75360 28476 75360 28476 0 _0194_
rlabel metal3 74544 30828 74544 30828 0 _0195_
rlabel metal3 75408 33432 75408 33432 0 _0196_
rlabel metal2 76032 34860 76032 34860 0 _0197_
rlabel metal2 76080 36540 76080 36540 0 _0198_
rlabel metal2 73344 37002 73344 37002 0 _0199_
rlabel metal2 71232 34440 71232 34440 0 _0200_
rlabel metal2 66336 37674 66336 37674 0 _0201_
rlabel metal3 65472 35868 65472 35868 0 _0202_
rlabel metal2 66288 32844 66288 32844 0 _0203_
rlabel metal3 69744 32004 69744 32004 0 _0204_
rlabel metal3 69456 30744 69456 30744 0 _0205_
rlabel metal3 68976 29232 68976 29232 0 _0206_
rlabel metal2 69120 27090 69120 27090 0 _0207_
rlabel metal2 67824 26292 67824 26292 0 _0208_
rlabel metal3 63216 26208 63216 26208 0 _0209_
rlabel metal2 61920 28014 61920 28014 0 _0210_
rlabel metal2 63072 30450 63072 30450 0 _0211_
rlabel metal3 61488 31248 61488 31248 0 _0212_
rlabel metal3 60912 34524 60912 34524 0 _0213_
rlabel metal2 62304 37086 62304 37086 0 _0214_
rlabel metal3 59040 37296 59040 37296 0 _0215_
rlabel metal3 55296 36792 55296 36792 0 _0216_
rlabel metal2 57984 34440 57984 34440 0 _0217_
rlabel metal2 60384 30576 60384 30576 0 _0218_
rlabel metal2 57120 27930 57120 27930 0 _0219_
rlabel metal2 57408 25620 57408 25620 0 _0220_
rlabel metal2 56544 26292 56544 26292 0 _0221_
rlabel metal2 54816 28140 54816 28140 0 _0222_
rlabel metal2 52896 30870 52896 30870 0 _0223_
rlabel metal2 53952 33978 53952 33978 0 _0224_
rlabel metal2 50976 34902 50976 34902 0 _0225_
rlabel metal2 46656 34440 46656 34440 0 _0226_
rlabel metal3 48816 33432 48816 33432 0 _0227_
rlabel metal3 48672 28980 48672 28980 0 _0228_
rlabel metal2 48864 27930 48864 27930 0 _0229_
rlabel metal2 48768 26418 48768 26418 0 _0230_
rlabel metal3 49440 23688 49440 23688 0 _0231_
rlabel metal2 47712 21042 47712 21042 0 _0232_
rlabel metal3 42816 21672 42816 21672 0 _0233_
rlabel metal2 44448 24318 44448 24318 0 _0234_
rlabel metal2 45120 25830 45120 25830 0 _0235_
rlabel metal3 44592 27720 44592 27720 0 _0236_
rlabel metal3 44256 29316 44256 29316 0 _0237_
rlabel metal3 41520 30828 41520 30828 0 _0238_
rlabel metal3 39696 28224 39696 28224 0 _0239_
rlabel metal3 39072 27720 39072 27720 0 _0240_
rlabel metal3 38304 25284 38304 25284 0 _0241_
rlabel metal2 39120 22512 39120 22512 0 _0242_
rlabel metal2 36576 24444 36576 24444 0 _0243_
rlabel metal2 34896 25536 34896 25536 0 _0244_
rlabel metal3 31008 24780 31008 24780 0 _0245_
rlabel metal3 29712 23100 29712 23100 0 _0246_
rlabel metal2 28224 21000 28224 21000 0 _0247_
rlabel metal2 11376 19236 11376 19236 0 _0248_
rlabel metal3 1968 2520 1968 2520 0 _0249_
rlabel metal3 1776 5124 1776 5124 0 _0250_
rlabel metal3 1776 6300 1776 6300 0 _0251_
rlabel metal3 1680 8568 1680 8568 0 _0252_
rlabel metal3 2304 10920 2304 10920 0 _0253_
rlabel metal3 1920 12684 1920 12684 0 _0254_
rlabel metal3 3216 15624 3216 15624 0 _0255_
rlabel metal2 23424 17808 23424 17808 0 _0256_
rlabel metal2 27168 17598 27168 17598 0 _0257_
rlabel metal3 30144 17640 30144 17640 0 _0258_
rlabel metal2 32544 18774 32544 18774 0 _0259_
rlabel metal3 36000 18648 36000 18648 0 _0260_
rlabel metal2 38784 18858 38784 18858 0 _0261_
rlabel metal2 44016 18732 44016 18732 0 _0262_
rlabel metal3 42912 17640 42912 17640 0 _0263_
rlabel metal2 43104 13545 43104 13545 0 _0264_
rlabel metal2 40512 15834 40512 15834 0 _0265_
rlabel metal3 37680 16464 37680 16464 0 _0266_
rlabel metal2 34272 16968 34272 16968 0 _0267_
rlabel metal2 30240 15036 30240 15036 0 _0268_
rlabel metal2 36912 11928 36912 11928 0 _0269_
rlabel metal2 38880 11970 38880 11970 0 _0270_
rlabel metal2 42432 11970 42432 11970 0 _0271_
rlabel metal2 44736 10416 44736 10416 0 _0272_
rlabel metal2 46848 10248 46848 10248 0 _0273_
rlabel metal2 48768 7182 48768 7182 0 _0274_
rlabel metal2 49056 6174 49056 6174 0 _0275_
rlabel metal2 52416 4410 52416 4410 0 _0276_
rlabel metal3 54432 6552 54432 6552 0 _0277_
rlabel metal2 54048 7938 54048 7938 0 _0278_
rlabel metal2 53952 10920 53952 10920 0 _0279_
rlabel metal2 51888 11928 51888 11928 0 _0280_
rlabel metal2 49104 12684 49104 12684 0 _0281_
rlabel metal2 47712 14007 47712 14007 0 _0282_
rlabel metal2 46272 16758 46272 16758 0 _0283_
rlabel metal2 49632 19446 49632 19446 0 _0284_
rlabel metal2 50304 17850 50304 17850 0 _0285_
rlabel metal2 53136 15624 53136 15624 0 _0286_
rlabel metal2 56928 15246 56928 15246 0 _0287_
rlabel metal2 58944 13650 58944 13650 0 _0288_
rlabel metal3 59136 11592 59136 11592 0 _0289_
rlabel metal2 59280 8484 59280 8484 0 _0290_
rlabel metal2 60624 6972 60624 6972 0 _0291_
rlabel metal2 61344 5502 61344 5502 0 _0292_
rlabel metal2 55968 5124 55968 5124 0 _0293_
rlabel metal2 56544 2226 56544 2226 0 _0294_
rlabel metal3 59424 2856 59424 2856 0 _0295_
rlabel metal2 64464 1932 64464 1932 0 _0296_
rlabel metal2 66240 3822 66240 3822 0 _0297_
rlabel metal2 66480 5880 66480 5880 0 _0298_
rlabel metal2 65664 8358 65664 8358 0 _0299_
rlabel metal2 65280 10458 65280 10458 0 _0300_
rlabel metal3 64512 11928 64512 11928 0 _0301_
rlabel metal2 60576 15246 60576 15246 0 _0302_
rlabel metal2 65472 15246 65472 15246 0 _0303_
rlabel metal2 70368 14994 70368 14994 0 _0304_
rlabel metal2 70464 12474 70464 12474 0 _0305_
rlabel metal3 70272 9324 70272 9324 0 _0306_
rlabel metal2 71520 8358 71520 8358 0 _0307_
rlabel metal2 71808 6552 71808 6552 0 _0308_
rlabel metal2 68880 1344 68880 1344 0 _0309_
rlabel metal2 72000 4620 72000 4620 0 _0310_
rlabel metal3 74832 1092 74832 1092 0 _0311_
rlabel metal2 79488 1176 79488 1176 0 _0312_
rlabel metal2 77184 3612 77184 3612 0 _0313_
rlabel metal2 77088 6174 77088 6174 0 _0314_
rlabel metal2 77088 8358 77088 8358 0 _0315_
rlabel metal2 77136 9660 77136 9660 0 _0316_
rlabel metal2 76512 12222 76512 12222 0 _0317_
rlabel metal2 76512 13734 76512 13734 0 _0318_
rlabel metal2 76224 14784 76224 14784 0 _0319_
rlabel metal2 76704 25368 76704 25368 0 _0320_
rlabel metal2 76992 26502 76992 26502 0 _0321_
rlabel metal2 76704 28602 76704 28602 0 _0322_
rlabel metal2 77088 30366 77088 30366 0 _0323_
rlabel metal2 77088 32298 77088 32298 0 _0324_
rlabel metal2 77424 34524 77424 34524 0 _0325_
rlabel metal3 76848 36540 76848 36540 0 _0326_
rlabel metal2 73536 36834 73536 36834 0 _0327_
rlabel metal2 72096 34440 72096 34440 0 _0328_
rlabel metal2 69072 36456 69072 36456 0 _0329_
rlabel metal2 66912 34650 66912 34650 0 _0330_
rlabel metal2 66336 31878 66336 31878 0 _0331_
rlabel metal2 72000 33276 72000 33276 0 _0332_
rlabel metal2 71712 30912 71712 30912 0 _0333_
rlabel metal2 71136 27594 71136 27594 0 _0334_
rlabel metal2 70704 24444 70704 24444 0 _0335_
rlabel metal2 67776 24990 67776 24990 0 _0336_
rlabel metal2 64032 24990 64032 24990 0 _0337_
rlabel metal3 65520 27720 65520 27720 0 _0338_
rlabel metal2 65760 29106 65760 29106 0 _0339_
rlabel metal2 63264 32550 63264 32550 0 _0340_
rlabel metal3 62976 34272 62976 34272 0 _0341_
rlabel metal2 63600 37380 63600 37380 0 _0342_
rlabel metal2 59040 35910 59040 35910 0 _0343_
rlabel metal2 55200 35490 55200 35490 0 _0344_
rlabel metal3 58368 32760 58368 32760 0 _0345_
rlabel metal2 60528 29316 60528 29316 0 _0346_
rlabel metal2 60336 27720 60336 27720 0 _0347_
rlabel metal2 60288 25578 60288 25578 0 _0348_
rlabel metal2 54912 24780 54912 24780 0 _0349_
rlabel metal3 56160 29232 56160 29232 0 _0350_
rlabel metal2 56160 31206 56160 31206 0 _0351_
rlabel metal2 55296 32928 55296 32928 0 _0352_
rlabel metal2 52128 35364 52128 35364 0 _0353_
rlabel metal2 46032 32256 46032 32256 0 _0354_
rlabel metal2 51312 31584 51312 31584 0 _0355_
rlabel metal2 51264 29610 51264 29610 0 _0356_
rlabel metal3 51936 27720 51936 27720 0 _0357_
rlabel metal2 52272 24780 52272 24780 0 _0358_
rlabel metal2 51744 23856 51744 23856 0 _0359_
rlabel metal2 50352 20748 50352 20748 0 _0360_
rlabel metal2 45792 20580 45792 20580 0 _0361_
rlabel metal2 46272 22932 46272 22932 0 _0362_
rlabel metal2 46848 24822 46848 24822 0 _0363_
rlabel metal2 47088 26796 47088 26796 0 _0364_
rlabel metal2 46320 29232 46320 29232 0 _0365_
rlabel metal2 44064 31626 44064 31626 0 _0366_
rlabel metal2 41760 28560 41760 28560 0 _0367_
rlabel metal2 41568 25956 41568 25956 0 _0368_
rlabel metal2 40608 24822 40608 24822 0 _0369_
rlabel metal2 41184 22344 41184 22344 0 _0370_
rlabel metal2 36240 21756 36240 21756 0 _0371_
rlabel metal2 35952 26292 35952 26292 0 _0372_
rlabel metal3 32784 23268 32784 23268 0 _0373_
rlabel metal3 32544 22176 32544 22176 0 _0374_
rlabel metal2 29088 21294 29088 21294 0 _0375_
rlabel metal3 12096 19152 12096 19152 0 _0376_
rlabel metal2 4848 3612 4848 3612 0 _0377_
rlabel metal2 4848 3948 4848 3948 0 _0378_
rlabel metal2 4608 8148 4608 8148 0 _0379_
rlabel metal2 4656 9660 4656 9660 0 _0380_
rlabel metal2 4992 11760 4992 11760 0 _0381_
rlabel metal2 4896 13944 4896 13944 0 _0382_
rlabel metal2 4656 15708 4656 15708 0 _0383_
rlabel metal2 64416 8610 64416 8610 0 _0384_
rlabel metal2 64128 9156 64128 9156 0 _0385_
rlabel metal2 64032 11970 64032 11970 0 _0386_
rlabel metal3 64176 11676 64176 11676 0 _0387_
rlabel metal2 63456 10626 63456 10626 0 _0388_
rlabel metal2 63168 11676 63168 11676 0 _0389_
rlabel metal2 61824 14028 61824 14028 0 _0390_
rlabel via2 60960 13440 60960 13440 0 _0391_
rlabel metal3 61488 12684 61488 12684 0 _0392_
rlabel metal2 61248 13188 61248 13188 0 _0393_
rlabel metal2 64032 14784 64032 14784 0 _0394_
rlabel metal2 65280 14742 65280 14742 0 _0395_
rlabel metal2 64176 13188 64176 13188 0 _0396_
rlabel metal2 64608 13188 64608 13188 0 _0397_
rlabel metal2 70320 13188 70320 13188 0 _0398_
rlabel metal2 70224 13440 70224 13440 0 _0399_
rlabel metal2 68064 14070 68064 14070 0 _0400_
rlabel metal2 68448 14028 68448 14028 0 _0401_
rlabel metal2 70032 11928 70032 11928 0 _0402_
rlabel metal2 70080 12432 70080 12432 0 _0403_
rlabel metal2 69216 12348 69216 12348 0 _0404_
rlabel metal2 68736 11676 68736 11676 0 _0405_
rlabel metal2 70032 8652 70032 8652 0 _0406_
rlabel metal2 70176 9786 70176 9786 0 _0407_
rlabel metal2 69024 10458 69024 10458 0 _0408_
rlabel metal2 68256 10038 68256 10038 0 _0409_
rlabel metal2 71520 9198 71520 9198 0 _0410_
rlabel metal2 69504 8694 69504 8694 0 _0411_
rlabel metal2 69600 8946 69600 8946 0 _0412_
rlabel metal2 69552 6972 69552 6972 0 _0413_
rlabel metal2 71232 6510 71232 6510 0 _0414_
rlabel metal3 70656 7056 70656 7056 0 _0415_
rlabel metal2 70128 5628 70128 5628 0 _0416_
rlabel metal2 69696 5628 69696 5628 0 _0417_
rlabel metal2 68640 2184 68640 2184 0 _0418_
rlabel metal2 68736 1008 68736 1008 0 _0419_
rlabel metal2 67680 2406 67680 2406 0 _0420_
rlabel metal2 67392 2184 67392 2184 0 _0421_
rlabel metal2 71808 3696 71808 3696 0 _0422_
rlabel metal3 70512 4032 70512 4032 0 _0423_
rlabel metal2 69216 3360 69216 3360 0 _0424_
rlabel metal2 69648 3444 69648 3444 0 _0425_
rlabel metal2 75168 2688 75168 2688 0 _0426_
rlabel metal2 74160 1932 74160 1932 0 _0427_
rlabel metal2 72768 1986 72768 1986 0 _0428_
rlabel metal3 72192 1092 72192 1092 0 _0429_
rlabel metal2 77568 2604 77568 2604 0 _0430_
rlabel metal2 78432 2142 78432 2142 0 _0431_
rlabel metal2 75168 1848 75168 1848 0 _0432_
rlabel metal2 75936 1512 75936 1512 0 _0433_
rlabel via1 76983 4962 76983 4962 0 _0434_
rlabel metal2 77376 3738 77376 3738 0 _0435_
rlabel metal3 75984 3612 75984 3612 0 _0436_
rlabel metal2 75648 4200 75648 4200 0 _0437_
rlabel metal2 76896 6720 76896 6720 0 _0438_
rlabel metal2 77280 6132 77280 6132 0 _0439_
rlabel metal3 76320 5124 76320 5124 0 _0440_
rlabel metal3 75936 5628 75936 5628 0 _0441_
rlabel metal2 77664 8400 77664 8400 0 _0442_
rlabel metal3 76800 7980 76800 7980 0 _0443_
rlabel metal2 76032 7140 76032 7140 0 _0444_
rlabel metal2 75744 7518 75744 7518 0 _0445_
rlabel metal2 76992 11004 76992 11004 0 _0446_
rlabel metal2 77232 10752 77232 10752 0 _0447_
rlabel metal3 76128 8904 76128 8904 0 _0448_
rlabel metal2 76032 9744 76032 9744 0 _0449_
rlabel metal2 76128 11424 76128 11424 0 _0450_
rlabel metal2 76224 11382 76224 11382 0 _0451_
rlabel metal2 75456 10920 75456 10920 0 _0452_
rlabel metal3 74928 11004 74928 11004 0 _0453_
rlabel metal2 76128 13158 76128 13158 0 _0454_
rlabel metal2 76128 12642 76128 12642 0 _0455_
rlabel metal2 74592 12432 74592 12432 0 _0456_
rlabel metal3 74592 13020 74592 13020 0 _0457_
rlabel metal2 75360 15246 75360 15246 0 _0458_
rlabel metal3 74784 14700 74784 14700 0 _0459_
rlabel metal2 74736 13860 74736 13860 0 _0460_
rlabel metal2 74112 14784 74112 14784 0 _0461_
rlabel metal2 75980 25299 75980 25299 0 _0462_
rlabel metal3 75120 25536 75120 25536 0 _0463_
rlabel metal2 74304 24780 74304 24780 0 _0464_
rlabel metal3 74592 26124 74592 26124 0 _0465_
rlabel metal2 76992 27342 76992 27342 0 _0466_
rlabel metal3 75984 27636 75984 27636 0 _0467_
rlabel metal2 75264 26334 75264 26334 0 _0468_
rlabel metal3 75216 26796 75216 26796 0 _0469_
rlabel metal2 76704 29400 76704 29400 0 _0470_
rlabel metal3 76752 28308 76752 28308 0 _0471_
rlabel metal2 75552 28056 75552 28056 0 _0472_
rlabel metal2 75264 28980 75264 28980 0 _0473_
rlabel metal2 76944 31332 76944 31332 0 _0474_
rlabel metal2 77280 30366 77280 30366 0 _0475_
rlabel metal2 75696 30072 75696 30072 0 _0476_
rlabel metal2 75360 30786 75360 30786 0 _0477_
rlabel metal2 78528 32928 78528 32928 0 _0478_
rlabel metal3 77952 33684 77952 33684 0 _0479_
rlabel metal2 75840 32340 75840 32340 0 _0480_
rlabel metal2 76128 33684 76128 33684 0 _0481_
rlabel metal2 77280 35238 77280 35238 0 _0482_
rlabel metal2 77664 34440 77664 34440 0 _0483_
rlabel metal2 76704 33390 76704 33390 0 _0484_
rlabel metal3 75792 34188 75792 34188 0 _0485_
rlabel metal2 77664 36918 77664 36918 0 _0486_
rlabel metal2 76800 36750 76800 36750 0 _0487_
rlabel metal2 76320 35910 76320 35910 0 _0488_
rlabel metal2 76128 36960 76128 36960 0 _0489_
rlabel metal2 73536 35616 73536 35616 0 _0490_
rlabel metal3 73776 37380 73776 37380 0 _0491_
rlabel metal2 74160 37380 74160 37380 0 _0492_
rlabel metal2 73776 37464 73776 37464 0 _0493_
rlabel metal2 71520 35448 71520 35448 0 _0494_
rlabel metal2 72000 35280 72000 35280 0 _0495_
rlabel metal2 72096 35448 72096 35448 0 _0496_
rlabel metal3 71232 35196 71232 35196 0 _0497_
rlabel metal2 71040 38178 71040 38178 0 _0498_
rlabel metal2 69312 36876 69312 36876 0 _0499_
rlabel metal3 68832 35784 68832 35784 0 _0500_
rlabel metal3 67728 38220 67728 38220 0 _0501_
rlabel metal2 66144 35112 66144 35112 0 _0502_
rlabel metal2 66048 35406 66048 35406 0 _0503_
rlabel metal2 66816 36624 66816 36624 0 _0504_
rlabel metal2 67296 35994 67296 35994 0 _0505_
rlabel metal2 66672 33012 66672 33012 0 _0506_
rlabel metal2 66336 33402 66336 33402 0 _0507_
rlabel metal2 66432 33810 66432 33810 0 _0508_
rlabel metal3 65952 33348 65952 33348 0 _0509_
rlabel metal2 72480 33402 72480 33402 0 _0510_
rlabel metal3 71088 33684 71088 33684 0 _0511_
rlabel metal2 69792 32424 69792 32424 0 _0512_
rlabel metal2 70176 32172 70176 32172 0 _0513_
rlabel metal2 71040 31206 71040 31206 0 _0514_
rlabel metal3 71376 31500 71376 31500 0 _0515_
rlabel metal2 70848 31626 70848 31626 0 _0516_
rlabel metal3 70704 30828 70704 30828 0 _0517_
rlabel metal2 70848 28056 70848 28056 0 _0518_
rlabel metal2 71232 28224 71232 28224 0 _0519_
rlabel metal2 69984 29778 69984 29778 0 _0520_
rlabel metal2 70320 29316 70320 29316 0 _0521_
rlabel metal2 71808 26040 71808 26040 0 _0522_
rlabel metal2 71904 26250 71904 26250 0 _0523_
rlabel metal2 69888 27552 69888 27552 0 _0524_
rlabel metal2 69648 26292 69648 26292 0 _0525_
rlabel metal2 68352 25830 68352 25830 0 _0526_
rlabel metal2 67872 25914 67872 25914 0 _0527_
rlabel metal2 67968 26250 67968 26250 0 _0528_
rlabel metal2 67584 26124 67584 26124 0 _0529_
rlabel metal3 64320 24612 64320 24612 0 _0530_
rlabel metal3 65088 24696 65088 24696 0 _0531_
rlabel metal2 64992 26040 64992 26040 0 _0532_
rlabel metal2 64704 26076 64704 26076 0 _0533_
rlabel metal2 65232 29148 65232 29148 0 _0534_
rlabel metal2 65376 27888 65376 27888 0 _0535_
rlabel metal2 63936 27048 63936 27048 0 _0536_
rlabel metal2 64128 28392 64128 28392 0 _0537_
rlabel metal2 65856 30366 65856 30366 0 _0538_
rlabel metal2 65856 29484 65856 29484 0 _0539_
rlabel metal2 63696 29316 63696 29316 0 _0540_
rlabel metal3 63168 29778 63168 29778 0 _0541_
rlabel metal2 62880 32424 62880 32424 0 _0542_
rlabel metal2 62976 32508 62976 32508 0 _0543_
rlabel metal2 62784 31416 62784 31416 0 _0544_
rlabel metal2 62496 32004 62496 32004 0 _0545_
rlabel metal2 62640 33684 62640 33684 0 _0546_
rlabel metal2 62880 34188 62880 34188 0 _0547_
rlabel metal2 62304 34104 62304 34104 0 _0548_
rlabel metal3 61776 34356 61776 34356 0 _0549_
rlabel metal2 63840 36624 63840 36624 0 _0550_
rlabel metal2 63936 36960 63936 36960 0 _0551_
rlabel metal2 62400 36120 62400 36120 0 _0552_
rlabel metal2 62112 36708 62112 36708 0 _0553_
rlabel metal2 58560 36162 58560 36162 0 _0554_
rlabel metal3 59232 35868 59232 35868 0 _0555_
rlabel metal2 59616 37338 59616 37338 0 _0556_
rlabel metal2 59232 37380 59232 37380 0 _0557_
rlabel metal2 56736 35532 56736 35532 0 _0558_
rlabel metal2 55680 36624 55680 36624 0 _0559_
rlabel metal3 56688 36540 56688 36540 0 _0560_
rlabel metal2 56016 35868 56016 35868 0 _0561_
rlabel metal2 59232 32256 59232 32256 0 _0562_
rlabel metal2 58272 32424 58272 32424 0 _0563_
rlabel metal2 57504 34482 57504 34482 0 _0564_
rlabel metal2 58368 33936 58368 33936 0 _0565_
rlabel metal2 60768 29568 60768 29568 0 _0566_
rlabel metal2 60864 29694 60864 29694 0 _0567_
rlabel metal2 60864 30828 60864 30828 0 _0568_
rlabel metal2 60576 30912 60576 30912 0 _0569_
rlabel metal2 59712 28140 59712 28140 0 _0570_
rlabel metal2 60048 28476 60048 28476 0 _0571_
rlabel metal2 59520 28602 59520 28602 0 _0572_
rlabel metal3 59472 27804 59472 27804 0 _0573_
rlabel metal2 59616 25662 59616 25662 0 _0574_
rlabel metal3 59040 26124 59040 26124 0 _0575_
rlabel metal2 58656 26040 58656 26040 0 _0576_
rlabel metal2 58320 24780 58320 24780 0 _0577_
rlabel metal2 56160 25578 56160 25578 0 _0578_
rlabel metal2 56400 25536 56400 25536 0 _0579_
rlabel metal2 56640 26040 56640 26040 0 _0580_
rlabel metal2 56352 26880 56352 26880 0 _0581_
rlabel metal2 55488 29190 55488 29190 0 _0582_
rlabel metal2 55296 29988 55296 29988 0 _0583_
rlabel metal2 55008 27552 55008 27552 0 _0584_
rlabel metal2 54720 28224 54720 28224 0 _0585_
rlabel metal2 55872 31836 55872 31836 0 _0586_
rlabel metal2 55872 30996 55872 30996 0 _0587_
rlabel metal2 54912 30366 54912 30366 0 _0588_
rlabel metal2 54672 30660 54672 30660 0 _0589_
rlabel metal2 55392 33768 55392 33768 0 _0590_
rlabel metal3 55296 33726 55296 33726 0 _0591_
rlabel metal2 54192 32004 54192 32004 0 _0592_
rlabel metal2 53808 32844 53808 32844 0 _0593_
rlabel metal2 51360 35448 51360 35448 0 _0594_
rlabel metal3 51264 35784 51264 35784 0 _0595_
rlabel metal2 51264 34440 51264 34440 0 _0596_
rlabel metal2 50880 34356 50880 34356 0 _0597_
rlabel metal3 47520 32844 47520 32844 0 _0598_
rlabel metal2 46080 32886 46080 32886 0 _0599_
rlabel metal2 46176 34440 46176 34440 0 _0600_
rlabel metal2 46656 33852 46656 33852 0 _0601_
rlabel metal2 50400 31878 50400 31878 0 _0602_
rlabel metal2 50496 32298 50496 32298 0 _0603_
rlabel metal2 49248 31710 49248 31710 0 _0604_
rlabel metal3 49152 33684 49152 33684 0 _0605_
rlabel metal2 50784 30324 50784 30324 0 _0606_
rlabel metal2 50880 29463 50880 29463 0 _0607_
rlabel metal2 49824 29232 49824 29232 0 _0608_
rlabel metal2 49584 29148 49584 29148 0 _0609_
rlabel metal2 51984 28308 51984 28308 0 _0610_
rlabel metal3 50928 28308 50928 28308 0 _0611_
rlabel metal2 49920 28224 49920 28224 0 _0612_
rlabel metal2 50400 28098 50400 28098 0 _0613_
rlabel metal2 52224 25830 52224 25830 0 _0614_
rlabel metal2 52128 26250 52128 26250 0 _0615_
rlabel metal2 50592 26754 50592 26754 0 _0616_
rlabel metal2 50880 26040 50880 26040 0 _0617_
rlabel metal2 51072 23961 51072 23961 0 _0618_
rlabel metal2 50880 24066 50880 24066 0 _0619_
rlabel metal2 50976 23814 50976 23814 0 _0620_
rlabel via2 50116 23268 50116 23268 0 _0621_
rlabel metal2 49728 21504 49728 21504 0 _0622_
rlabel metal3 50304 21588 50304 21588 0 _0623_
rlabel metal2 49152 21840 49152 21840 0 _0624_
rlabel metal2 48864 21840 48864 21840 0 _0625_
rlabel metal2 45024 21840 45024 21840 0 _0626_
rlabel metal2 45408 22008 45408 22008 0 _0627_
rlabel metal2 46320 21000 46320 21000 0 _0628_
rlabel metal2 45168 20748 45168 20748 0 _0629_
rlabel metal2 45888 23856 45888 23856 0 _0630_
rlabel metal3 45312 23772 45312 23772 0 _0631_
rlabel metal2 44736 23520 44736 23520 0 _0632_
rlabel metal3 44208 23604 44208 23604 0 _0633_
rlabel metal2 46848 26166 46848 26166 0 _0634_
rlabel metal2 46944 24990 46944 24990 0 _0635_
rlabel metal2 44928 24780 44928 24780 0 _0636_
rlabel metal2 45216 25284 45216 25284 0 _0637_
rlabel via1 46263 26789 46263 26789 0 _0638_
rlabel metal2 46368 27678 46368 27678 0 _0639_
rlabel metal2 45840 27048 45840 27048 0 _0640_
rlabel metal2 45456 26796 45456 26796 0 _0641_
rlabel metal2 45984 29568 45984 29568 0 _0642_
rlabel metal2 46080 29400 46080 29400 0 _0643_
rlabel metal2 45264 28560 45264 28560 0 _0644_
rlabel metal2 44928 29904 44928 29904 0 _0645_
rlabel metal2 42864 32172 42864 32172 0 _0646_
rlabel metal2 42912 31290 42912 31290 0 _0647_
rlabel metal2 43008 30576 43008 30576 0 _0648_
rlabel metal2 42720 31416 42720 31416 0 _0649_
rlabel metal2 41568 29736 41568 29736 0 _0650_
rlabel metal2 42048 29064 42048 29064 0 _0651_
rlabel metal2 41184 29358 41184 29358 0 _0652_
rlabel metal2 40896 28980 40896 28980 0 _0653_
rlabel metal2 41184 27342 41184 27342 0 _0654_
rlabel metal3 41184 27384 41184 27384 0 _0655_
rlabel metal2 40608 27888 40608 27888 0 _0656_
rlabel metal2 39840 27216 39840 27216 0 _0657_
rlabel metal2 40320 24066 40320 24066 0 _0658_
rlabel metal2 40704 25158 40704 25158 0 _0659_
rlabel metal2 39648 26082 39648 26082 0 _0660_
rlabel metal2 40128 25326 40128 25326 0 _0661_
rlabel metal2 41088 23541 41088 23541 0 _0662_
rlabel metal3 40032 22260 40032 22260 0 _0663_
rlabel metal2 39360 22932 39360 22932 0 _0664_
rlabel metal2 39024 22260 39024 22260 0 _0665_
rlabel metal2 37008 22932 37008 22932 0 _0666_
rlabel metal3 36624 22596 36624 22596 0 _0667_
rlabel metal3 37392 23268 37392 23268 0 _0668_
rlabel metal2 36480 23772 36480 23772 0 _0669_
rlabel metal2 35424 26376 35424 26376 0 _0670_
rlabel metal2 35136 26124 35136 26124 0 _0671_
rlabel metal2 35232 25368 35232 25368 0 _0672_
rlabel metal2 34848 25284 34848 25284 0 _0673_
rlabel metal2 32352 23520 32352 23520 0 _0674_
rlabel metal2 32256 23352 32256 23352 0 _0675_
rlabel metal2 33216 24864 33216 24864 0 _0676_
rlabel metal2 32064 24612 32064 24612 0 _0677_
rlabel metal2 31920 22512 31920 22512 0 _0678_
rlabel metal3 31536 23100 31536 23100 0 _0679_
rlabel metal2 31296 23352 31296 23352 0 _0680_
rlabel metal2 30960 23100 30960 23100 0 _0681_
rlabel metal2 28752 22260 28752 22260 0 _0682_
rlabel metal2 28464 20748 28464 20748 0 _0683_
rlabel metal2 28656 20748 28656 20748 0 _0684_
rlabel metal2 28224 20748 28224 20748 0 _0685_
rlabel metal2 11520 18480 11520 18480 0 _0686_
rlabel metal2 12000 19320 12000 19320 0 _0687_
rlabel metal3 17280 20034 17280 20034 0 _0688_
rlabel metal2 11328 20076 11328 20076 0 _0689_
rlabel metal2 4224 3864 4224 3864 0 _0690_
rlabel metal3 3456 2604 3456 2604 0 _0691_
rlabel metal2 2688 2520 2688 2520 0 _0692_
rlabel metal2 2400 3276 2400 3276 0 _0693_
rlabel metal2 3744 5586 3744 5586 0 _0694_
rlabel metal2 2400 4872 2400 4872 0 _0695_
rlabel metal2 2592 4620 2592 4620 0 _0696_
rlabel metal2 2208 5061 2208 5061 0 _0697_
rlabel metal2 4032 7434 4032 7434 0 _0698_
rlabel metal2 2400 6762 2400 6762 0 _0699_
rlabel metal2 2496 6384 2496 6384 0 _0700_
rlabel metal2 2256 6468 2256 6468 0 _0701_
rlabel metal2 3648 9198 3648 9198 0 _0702_
rlabel metal2 3744 8946 3744 8946 0 _0703_
rlabel metal2 2544 7728 2544 7728 0 _0704_
rlabel metal2 2016 8610 2016 8610 0 _0705_
rlabel metal2 3936 11256 3936 11256 0 _0706_
rlabel metal2 4032 11298 4032 11298 0 _0707_
rlabel metal2 2592 10710 2592 10710 0 _0708_
rlabel metal2 2208 11004 2208 11004 0 _0709_
rlabel metal2 3984 13776 3984 13776 0 _0710_
rlabel metal3 4368 13020 4368 13020 0 _0711_
rlabel metal2 2592 12432 2592 12432 0 _0712_
rlabel metal2 2400 13494 2400 13494 0 _0713_
rlabel metal2 3696 15540 3696 15540 0 _0714_
rlabel metal2 3840 15666 3840 15666 0 _0715_
rlabel metal2 2880 14784 2880 14784 0 _0716_
rlabel metal2 2736 14700 2736 14700 0 _0717_
rlabel metal2 23712 17430 23712 17430 0 _0718_
rlabel metal2 27360 17472 27360 17472 0 _0719_
rlabel metal3 30336 17136 30336 17136 0 _0720_
rlabel metal2 32736 18270 32736 18270 0 _0721_
rlabel metal2 36576 18018 36576 18018 0 _0722_
rlabel metal2 38880 19530 38880 19530 0 _0723_
rlabel metal2 44256 18480 44256 18480 0 _0724_
rlabel metal3 42960 16380 42960 16380 0 _0725_
rlabel metal3 43152 14700 43152 14700 0 _0726_
rlabel metal2 40704 15456 40704 15456 0 _0727_
rlabel metal3 37392 16212 37392 16212 0 _0728_
rlabel metal2 33792 16968 33792 16968 0 _0729_
rlabel metal2 31872 15582 31872 15582 0 _0730_
rlabel metal2 36624 12348 36624 12348 0 _0731_
rlabel metal2 39168 11760 39168 11760 0 _0732_
rlabel metal3 42240 12516 42240 12516 0 _0733_
rlabel metal2 44544 10458 44544 10458 0 _0734_
rlabel metal2 46704 10164 46704 10164 0 _0735_
rlabel metal2 48960 7770 48960 7770 0 _0736_
rlabel metal2 49344 5544 49344 5544 0 _0737_
rlabel metal2 52704 3948 52704 3948 0 _0738_
rlabel metal2 54816 5754 54816 5754 0 _0739_
rlabel metal2 54240 8610 54240 8610 0 _0740_
rlabel metal3 53328 11004 53328 11004 0 _0741_
rlabel metal2 52032 13032 52032 13032 0 _0742_
rlabel metal2 49152 12474 49152 12474 0 _0743_
rlabel metal2 47904 14658 47904 14658 0 _0744_
rlabel metal2 45936 16212 45936 16212 0 _0745_
rlabel metal2 49248 19530 49248 19530 0 _0746_
rlabel metal2 49824 17766 49824 17766 0 _0747_
rlabel metal2 53376 16296 53376 16296 0 _0748_
rlabel metal2 57216 14784 57216 14784 0 _0749_
rlabel metal2 58656 13314 58656 13314 0 _0750_
rlabel metal2 59136 11970 59136 11970 0 _0751_
rlabel metal2 59328 9156 59328 9156 0 _0752_
rlabel metal2 60576 7854 60576 7854 0 _0753_
rlabel metal2 61152 5922 61152 5922 0 _0754_
rlabel metal3 56160 4956 56160 4956 0 _0755_
rlabel metal2 56544 2688 56544 2688 0 _0756_
rlabel metal3 59136 3192 59136 3192 0 _0757_
rlabel metal2 64512 2646 64512 2646 0 _0758_
rlabel metal2 66432 3360 66432 3360 0 _0759_
rlabel metal2 66768 5628 66768 5628 0 _0760_
rlabel metal2 65856 7896 65856 7896 0 _0761_
rlabel metal2 65376 10290 65376 10290 0 _0762_
rlabel metal2 64512 11970 64512 11970 0 _0763_
rlabel metal3 61680 14700 61680 14700 0 _0764_
rlabel metal2 65184 14994 65184 14994 0 _0765_
rlabel metal3 70560 15540 70560 15540 0 _0766_
rlabel metal2 70560 12222 70560 12222 0 _0767_
rlabel metal3 70608 9492 70608 9492 0 _0768_
rlabel metal2 71760 7980 71760 7980 0 _0769_
rlabel metal2 72192 6426 72192 6426 0 _0770_
rlabel metal2 68640 1344 68640 1344 0 _0771_
rlabel metal3 72048 4956 72048 4956 0 _0772_
rlabel metal2 74304 2058 74304 2058 0 _0773_
rlabel metal2 78528 1848 78528 1848 0 _0774_
rlabel metal2 77520 3444 77520 3444 0 _0775_
rlabel metal2 77376 5544 77376 5544 0 _0776_
rlabel metal3 77376 7392 77376 7392 0 _0777_
rlabel metal2 77424 9492 77424 9492 0 _0778_
rlabel metal2 76848 11676 76848 11676 0 _0779_
rlabel metal2 76800 13272 76800 13272 0 _0780_
rlabel metal2 75936 14154 75936 14154 0 _0781_
rlabel metal2 76512 24738 76512 24738 0 _0782_
rlabel metal2 77232 26124 77232 26124 0 _0783_
rlabel metal2 76992 28266 76992 28266 0 _0784_
rlabel metal2 77376 30324 77376 30324 0 _0785_
rlabel metal2 77760 33684 77760 33684 0 _0786_
rlabel metal2 77760 34272 77760 34272 0 _0787_
rlabel metal2 76896 37002 76896 37002 0 _0788_
rlabel metal2 73728 36120 73728 36120 0 _0789_
rlabel metal2 71712 33810 71712 33810 0 _0790_
rlabel metal2 69408 36624 69408 36624 0 _0791_
rlabel metal2 67200 34440 67200 34440 0 _0792_
rlabel metal2 66624 31416 66624 31416 0 _0793_
rlabel metal2 72672 31878 72672 31878 0 _0794_
rlabel metal2 72192 30156 72192 30156 0 _0795_
rlabel metal2 71328 28266 71328 28266 0 _0796_
rlabel metal3 71184 24612 71184 24612 0 _0797_
rlabel metal2 67968 24696 67968 24696 0 _0798_
rlabel metal2 64224 24696 64224 24696 0 _0799_
rlabel metal2 65472 27594 65472 27594 0 _0800_
rlabel metal2 65952 29778 65952 29778 0 _0801_
rlabel metal2 64224 32088 64224 32088 0 _0802_
rlabel metal2 63168 33810 63168 33810 0 _0803_
rlabel metal2 64320 37506 64320 37506 0 _0804_
rlabel metal2 59232 35826 59232 35826 0 _0805_
rlabel metal2 54912 35574 54912 35574 0 _0806_
rlabel metal3 58656 33432 58656 33432 0 _0807_
rlabel metal2 60288 29778 60288 29778 0 _0808_
rlabel metal3 60528 28308 60528 28308 0 _0809_
rlabel metal2 60288 24822 60288 24822 0 _0810_
rlabel metal3 55680 24024 55680 24024 0 _0811_
rlabel metal2 56352 28182 56352 28182 0 _0812_
rlabel metal2 56160 30870 56160 30870 0 _0813_
rlabel metal3 54672 32844 54672 32844 0 _0814_
rlabel metal2 52416 35280 52416 35280 0 _0815_
rlabel metal3 46464 31584 46464 31584 0 _0816_
rlabel metal2 51120 31332 51120 31332 0 _0817_
rlabel metal2 50784 29862 50784 29862 0 _0818_
rlabel metal3 52080 27636 52080 27636 0 _0819_
rlabel metal2 52416 25242 52416 25242 0 _0820_
rlabel metal3 51264 23184 51264 23184 0 _0821_
rlabel metal2 50880 21546 50880 21546 0 _0822_
rlabel metal2 45792 21462 45792 21462 0 _0823_
rlabel metal2 45888 23184 45888 23184 0 _0824_
rlabel metal2 47088 24612 47088 24612 0 _0825_
rlabel metal3 47568 27636 47568 27636 0 _0826_
rlabel metal2 47136 30198 47136 30198 0 _0827_
rlabel metal2 43296 30828 43296 30828 0 _0828_
rlabel metal3 41712 28560 41712 28560 0 _0829_
rlabel metal2 41184 26250 41184 26250 0 _0830_
rlabel metal2 40800 24570 40800 24570 0 _0831_
rlabel metal3 40992 21672 40992 21672 0 _0832_
rlabel metal2 36384 21504 36384 21504 0 _0833_
rlabel metal2 36096 26208 36096 26208 0 _0834_
rlabel metal2 32832 23730 32832 23730 0 _0835_
rlabel metal2 32448 21966 32448 21966 0 _0836_
rlabel metal2 28800 21000 28800 21000 0 _0837_
rlabel metal2 12192 18942 12192 18942 0 _0838_
rlabel metal2 4896 3360 4896 3360 0 _0839_
rlabel metal2 4896 5166 4896 5166 0 _0840_
rlabel metal2 4752 7392 4752 7392 0 _0841_
rlabel metal2 4704 9408 4704 9408 0 _0842_
rlabel metal2 4992 11130 4992 11130 0 _0843_
rlabel metal2 4368 13440 4368 13440 0 _0844_
rlabel metal2 4224 15540 4224 15540 0 _0845_
rlabel metal2 4224 24066 4224 24066 0 _0846_
rlabel metal2 4704 19824 4704 19824 0 _0847_
rlabel metal2 22560 17850 22560 17850 0 _0848_
rlabel metal2 22656 17850 22656 17850 0 _0849_
rlabel metal3 2496 21504 2496 21504 0 _0850_
rlabel metal3 2256 22848 2256 22848 0 _0851_
rlabel metal2 22848 20328 22848 20328 0 _0852_
rlabel metal2 22176 19656 22176 19656 0 _0853_
rlabel metal2 27744 18480 27744 18480 0 _0854_
rlabel metal3 27120 18564 27120 18564 0 _0855_
rlabel metal2 26496 18816 26496 18816 0 _0856_
rlabel metal2 26208 18648 26208 18648 0 _0857_
rlabel metal2 29856 18480 29856 18480 0 _0858_
rlabel metal2 29760 18690 29760 18690 0 _0859_
rlabel metal2 28896 18690 28896 18690 0 _0860_
rlabel metal2 29088 19194 29088 19194 0 _0861_
rlabel metal2 33792 19320 33792 19320 0 _0862_
rlabel metal2 33888 18942 33888 18942 0 _0863_
rlabel metal2 32160 19782 32160 19782 0 _0864_
rlabel metal2 32544 20076 32544 20076 0 _0865_
rlabel metal2 36000 19236 36000 19236 0 _0866_
rlabel metal2 35712 19488 35712 19488 0 _0867_
rlabel metal2 35520 19992 35520 19992 0 _0868_
rlabel metal2 35904 20076 35904 20076 0 _0869_
rlabel metal2 38496 19950 38496 19950 0 _0870_
rlabel metal2 38400 19740 38400 19740 0 _0871_
rlabel metal2 38112 20244 38112 20244 0 _0872_
rlabel metal3 38736 20748 38736 20748 0 _0873_
rlabel metal2 43584 18984 43584 18984 0 _0874_
rlabel metal2 42048 18984 42048 18984 0 _0875_
rlabel metal2 41952 19320 41952 19320 0 _0876_
rlabel metal2 42240 19908 42240 19908 0 _0877_
rlabel metal2 42912 16968 42912 16968 0 _0878_
rlabel metal2 42816 18144 42816 18144 0 _0879_
rlabel metal2 42240 18438 42240 18438 0 _0880_
rlabel metal2 41664 17514 41664 17514 0 _0881_
rlabel metal2 42912 13482 42912 13482 0 _0882_
rlabel metal2 42816 13608 42816 13608 0 _0883_
rlabel metal2 41760 14238 41760 14238 0 _0884_
rlabel metal2 41472 13860 41472 13860 0 _0885_
rlabel metal2 39072 15414 39072 15414 0 _0886_
rlabel metal2 40560 15540 40560 15540 0 _0887_
rlabel metal2 40176 14196 40176 14196 0 _0888_
rlabel metal2 39456 14322 39456 14322 0 _0889_
rlabel metal2 38496 15960 38496 15960 0 _0890_
rlabel metal2 37824 15918 37824 15918 0 _0891_
rlabel metal2 38592 14322 38592 14322 0 _0892_
rlabel metal2 36672 15540 36672 15540 0 _0893_
rlabel metal2 34656 16296 34656 16296 0 _0894_
rlabel metal3 34320 16464 34320 16464 0 _0895_
rlabel metal2 34176 15456 34176 15456 0 _0896_
rlabel metal2 33792 15540 33792 15540 0 _0897_
rlabel metal2 33024 14280 33024 14280 0 _0898_
rlabel metal3 32352 14952 32352 14952 0 _0899_
rlabel metal2 33138 13235 33138 13235 0 _0900_
rlabel metal3 32256 13188 32256 13188 0 _0901_
rlabel metal2 36432 11676 36432 11676 0 _0902_
rlabel metal3 35664 11844 35664 11844 0 _0903_
rlabel metal2 35136 12990 35136 12990 0 _0904_
rlabel metal3 35088 11676 35088 11676 0 _0905_
rlabel metal2 39648 10836 39648 10836 0 _0906_
rlabel metal3 38304 10920 38304 10920 0 _0907_
rlabel metal2 36960 10920 36960 10920 0 _0908_
rlabel metal2 37344 11004 37344 11004 0 _0909_
rlabel metal2 42912 11214 42912 11214 0 _0910_
rlabel metal2 43008 10248 43008 10248 0 _0911_
rlabel metal2 40032 9408 40032 9408 0 _0912_
rlabel metal2 40512 9492 40512 9492 0 _0913_
rlabel metal2 43872 9492 43872 9492 0 _0914_
rlabel metal2 42336 9366 42336 9366 0 _0915_
rlabel metal2 42240 9408 42240 9408 0 _0916_
rlabel metal2 42528 9660 42528 9660 0 _0917_
rlabel metal2 46752 8946 46752 8946 0 _0918_
rlabel metal3 45840 8568 45840 8568 0 _0919_
rlabel metal2 44736 7896 44736 7896 0 _0920_
rlabel metal2 45216 7980 45216 7980 0 _0921_
rlabel metal2 48672 8232 48672 8232 0 _0922_
rlabel metal2 48576 8274 48576 8274 0 _0923_
rlabel metal2 47232 7896 47232 7896 0 _0924_
rlabel metal2 47328 6636 47328 6636 0 _0925_
rlabel metal2 48672 5166 48672 5166 0 _0926_
rlabel metal3 48000 4788 48000 4788 0 _0927_
rlabel metal2 47520 5922 47520 5922 0 _0928_
rlabel metal2 47328 4116 47328 4116 0 _0929_
rlabel metal2 52512 4116 52512 4116 0 _0930_
rlabel metal2 51648 4368 51648 4368 0 _0931_
rlabel metal2 49824 3444 49824 3444 0 _0932_
rlabel metal2 50544 3444 50544 3444 0 _0933_
rlabel metal2 54480 7140 54480 7140 0 _0934_
rlabel metal2 54336 6762 54336 6762 0 _0935_
rlabel metal2 52272 5124 52272 5124 0 _0936_
rlabel metal2 52704 5628 52704 5628 0 _0937_
rlabel metal2 53856 9198 53856 9198 0 _0938_
rlabel metal2 54144 8022 54144 8022 0 _0939_
rlabel via2 53087 7056 53087 7056 0 _0940_
rlabel metal2 52800 7560 52800 7560 0 _0941_
rlabel metal2 53664 10248 53664 10248 0 _0942_
rlabel metal2 53568 10710 53568 10710 0 _0943_
rlabel metal2 52848 9660 52848 9660 0 _0944_
rlabel metal2 52464 9660 52464 9660 0 _0945_
rlabel metal3 51888 11676 51888 11676 0 _0946_
rlabel metal2 51936 11634 51936 11634 0 _0947_
rlabel metal2 51552 10332 51552 10332 0 _0948_
rlabel metal2 51168 11004 51168 11004 0 _0949_
rlabel metal2 48720 12348 48720 12348 0 _0950_
rlabel metal2 49056 12096 49056 12096 0 _0951_
rlabel metal2 48576 11760 48576 11760 0 _0952_
rlabel metal2 48192 11676 48192 11676 0 _0953_
rlabel metal2 47712 15246 47712 15246 0 _0954_
rlabel metal3 47088 14028 47088 14028 0 _0955_
rlabel metal2 46464 13146 46464 13146 0 _0956_
rlabel metal3 45936 13188 45936 13188 0 _0957_
rlabel metal2 47136 16506 47136 16506 0 _0958_
rlabel metal3 46656 16212 46656 16212 0 _0959_
rlabel metal2 46320 14952 46320 14952 0 _0960_
rlabel metal2 45888 15540 45888 15540 0 _0961_
rlabel metal2 49440 18522 49440 18522 0 _0962_
rlabel metal3 48096 18648 48096 18648 0 _0963_
rlabel metal2 46464 18270 46464 18270 0 _0964_
rlabel metal2 47232 18564 47232 18564 0 _0965_
rlabel metal3 51360 17052 51360 17052 0 _0966_
rlabel metal2 49920 17640 49920 17640 0 _0967_
rlabel metal2 49056 17052 49056 17052 0 _0968_
rlabel metal2 49584 17052 49584 17052 0 _0969_
rlabel metal2 52416 14028 52416 14028 0 _0970_
rlabel metal2 52608 14154 52608 14154 0 _0971_
rlabel metal2 51120 14028 51120 14028 0 _0972_
rlabel metal2 51456 15036 51456 15036 0 _0973_
rlabel metal2 56640 14448 56640 14448 0 _0974_
rlabel metal3 56304 13776 56304 13776 0 _0975_
rlabel metal3 54000 13188 54000 13188 0 _0976_
rlabel metal3 54912 13188 54912 13188 0 _0977_
rlabel metal2 58416 13356 58416 13356 0 _0978_
rlabel metal3 57696 13188 57696 13188 0 _0979_
rlabel metal2 56832 13230 56832 13230 0 _0980_
rlabel metal2 56544 12432 56544 12432 0 _0981_
rlabel metal2 59136 10458 59136 10458 0 _0982_
rlabel metal2 59232 10500 59232 10500 0 _0983_
rlabel metal2 57744 10164 57744 10164 0 _0984_
rlabel metal2 58128 10164 58128 10164 0 _0985_
rlabel metal2 58848 8946 58848 8946 0 _0986_
rlabel metal3 58752 8778 58752 8778 0 _0987_
rlabel metal2 58080 9576 58080 9576 0 _0988_
rlabel metal2 57744 8652 57744 8652 0 _0989_
rlabel metal2 60384 6699 60384 6699 0 _0990_
rlabel metal3 59280 6300 59280 6300 0 _0991_
rlabel metal2 58368 7098 58368 7098 0 _0992_
rlabel metal2 58080 6510 58080 6510 0 _0993_
rlabel metal2 62208 4662 62208 4662 0 _0994_
rlabel metal3 61056 5586 61056 5586 0 _0995_
rlabel metal2 59520 5922 59520 5922 0 _0996_
rlabel metal2 59328 4452 59328 4452 0 _0997_
rlabel metal2 56928 3864 56928 3864 0 _0998_
rlabel metal2 57312 4242 57312 4242 0 _0999_
rlabel metal2 57408 4200 57408 4200 0 _1000_
rlabel metal3 56400 4116 56400 4116 0 _1001_
rlabel metal2 56160 1638 56160 1638 0 _1002_
rlabel metal2 56256 1554 56256 1554 0 _1003_
rlabel metal2 55728 1092 55728 1092 0 _1004_
rlabel metal2 55344 1092 55344 1092 0 _1005_
rlabel metal2 60192 2604 60192 2604 0 _1006_
rlabel metal3 59664 2604 59664 2604 0 _1007_
rlabel metal2 59328 1176 59328 1176 0 _1008_
rlabel metal2 58752 924 58752 924 0 _1009_
rlabel metal2 64608 1176 64608 1176 0 _1010_
rlabel metal2 62400 1176 62400 1176 0 _1011_
rlabel metal2 62304 1176 62304 1176 0 _1012_
rlabel metal2 62688 1092 62688 1092 0 _1013_
rlabel metal2 66432 4662 66432 4662 0 _1014_
rlabel metal2 66336 3486 66336 3486 0 _1015_
rlabel metal2 63936 3192 63936 3192 0 _1016_
rlabel metal3 64224 3444 64224 3444 0 _1017_
rlabel metal2 66432 6720 66432 6720 0 _1018_
rlabel metal3 66480 5628 66480 5628 0 _1019_
rlabel metal2 65856 5292 65856 5292 0 _1020_
rlabel metal2 65088 5712 65088 5712 0 _1021_
rlabel metal2 65472 7434 65472 7434 0 _1022_
rlabel metal2 65760 8022 65760 8022 0 _1023_
rlabel metal3 64464 7056 64464 7056 0 _1024_
rlabel metal2 63648 8064 63648 8064 0 _1025_
rlabel metal2 64512 10710 64512 10710 0 _1026_
rlabel metal2 65088 10500 65088 10500 0 _1027_
rlabel metal3 16974 36708 16974 36708 0 clk
rlabel metal2 53136 22764 53136 22764 0 clknet_0_clk
rlabel metal2 59616 4536 59616 4536 0 clknet_2_0__leaf_clk
rlabel metal2 30096 12516 30096 12516 0 clknet_2_1__leaf_clk
rlabel metal2 54768 13020 54768 13020 0 clknet_2_2__leaf_clk
rlabel metal3 58464 33852 58464 33852 0 clknet_2_3__leaf_clk
rlabel metal2 6192 14028 6192 14028 0 clknet_leaf_0_clk
rlabel metal2 43008 18522 43008 18522 0 clknet_leaf_10_clk
rlabel metal2 77424 13860 77424 13860 0 clknet_leaf_11_clk
rlabel metal2 62112 10248 62112 10248 0 clknet_leaf_12_clk
rlabel metal2 78288 1092 78288 1092 0 clknet_leaf_13_clk
rlabel metal2 60432 1932 60432 1932 0 clknet_leaf_14_clk
rlabel metal3 56304 1932 56304 1932 0 clknet_leaf_15_clk
rlabel metal3 40992 14028 40992 14028 0 clknet_leaf_16_clk
rlabel metal3 40560 18564 40560 18564 0 clknet_leaf_17_clk
rlabel metal2 2496 5376 2496 5376 0 clknet_leaf_18_clk
rlabel metal2 29808 23100 29808 23100 0 clknet_leaf_1_clk
rlabel metal3 11808 19236 11808 19236 0 clknet_leaf_2_clk
rlabel metal2 42960 26796 42960 26796 0 clknet_leaf_3_clk
rlabel metal2 47952 34356 47952 34356 0 clknet_leaf_4_clk
rlabel metal3 56208 36708 56208 36708 0 clknet_leaf_5_clk
rlabel metal2 60384 36792 60384 36792 0 clknet_leaf_6_clk
rlabel metal2 75408 35196 75408 35196 0 clknet_leaf_7_clk
rlabel metal3 62448 28308 62448 28308 0 clknet_leaf_8_clk
rlabel metal2 53568 24948 53568 24948 0 clknet_leaf_9_clk
rlabel metal2 22464 18984 22464 18984 0 daisychain\[0\]
rlabel metal2 50208 29316 50208 29316 0 daisychain\[100\]
rlabel metal2 51264 27846 51264 27846 0 daisychain\[101\]
rlabel metal2 50592 25200 50592 25200 0 daisychain\[102\]
rlabel metal3 50640 23184 50640 23184 0 daisychain\[103\]
rlabel metal3 47664 22260 47664 22260 0 daisychain\[104\]
rlabel metal2 44784 21756 44784 21756 0 daisychain\[105\]
rlabel metal2 44736 24318 44736 24318 0 daisychain\[106\]
rlabel metal3 45840 25872 45840 25872 0 daisychain\[107\]
rlabel metal3 45504 27804 45504 27804 0 daisychain\[108\]
rlabel metal2 44352 30660 44352 30660 0 daisychain\[109\]
rlabel metal2 36288 15624 36288 15624 0 daisychain\[10\]
rlabel metal2 42624 30912 42624 30912 0 daisychain\[110\]
rlabel metal2 40800 28602 40800 28602 0 daisychain\[111\]
rlabel metal2 40128 27090 40128 27090 0 daisychain\[112\]
rlabel metal2 39600 25116 39600 25116 0 daisychain\[113\]
rlabel metal3 38448 23772 38448 23772 0 daisychain\[114\]
rlabel metal2 36048 23772 36048 23772 0 daisychain\[115\]
rlabel metal2 34464 25704 34464 25704 0 daisychain\[116\]
rlabel metal2 31680 24864 31680 24864 0 daisychain\[117\]
rlabel metal3 31104 22260 31104 22260 0 daisychain\[118\]
rlabel metal2 26784 20118 26784 20118 0 daisychain\[119\]
rlabel metal2 33504 16002 33504 16002 0 daisychain\[11\]
rlabel metal2 3168 2646 3168 2646 0 daisychain\[120\]
rlabel metal2 2112 3738 2112 3738 0 daisychain\[121\]
rlabel metal2 1728 5250 1728 5250 0 daisychain\[122\]
rlabel metal2 2016 7812 2016 7812 0 daisychain\[123\]
rlabel metal2 1728 8694 1728 8694 0 daisychain\[124\]
rlabel metal2 1824 11046 1824 11046 0 daisychain\[125\]
rlabel metal3 1920 14028 1920 14028 0 daisychain\[126\]
rlabel metal2 1344 15036 1344 15036 0 daisychain\[127\]
rlabel metal2 34944 13230 34944 13230 0 daisychain\[12\]
rlabel metal3 36528 12348 36528 12348 0 daisychain\[13\]
rlabel metal3 38352 11004 38352 11004 0 daisychain\[14\]
rlabel metal2 41904 10416 41904 10416 0 daisychain\[15\]
rlabel metal2 43104 9576 43104 9576 0 daisychain\[16\]
rlabel metal2 46608 8904 46608 8904 0 daisychain\[17\]
rlabel metal3 48096 7392 48096 7392 0 daisychain\[18\]
rlabel metal2 48288 4410 48288 4410 0 daisychain\[19\]
rlabel metal2 27264 18732 27264 18732 0 daisychain\[1\]
rlabel metal3 51552 3528 51552 3528 0 daisychain\[20\]
rlabel metal2 53808 6216 53808 6216 0 daisychain\[21\]
rlabel metal2 53376 8274 53376 8274 0 daisychain\[22\]
rlabel metal2 52224 10038 52224 10038 0 daisychain\[23\]
rlabel metal2 49536 11634 49536 11634 0 daisychain\[24\]
rlabel metal2 48192 13074 48192 13074 0 daisychain\[25\]
rlabel metal2 46032 14700 46032 14700 0 daisychain\[26\]
rlabel metal3 45984 17136 45984 17136 0 daisychain\[27\]
rlabel metal2 48816 18564 48816 18564 0 daisychain\[28\]
rlabel metal3 50400 17052 50400 17052 0 daisychain\[29\]
rlabel metal2 30288 18648 30288 18648 0 daisychain\[2\]
rlabel metal3 52128 16212 52128 16212 0 daisychain\[30\]
rlabel metal2 56160 14238 56160 14238 0 daisychain\[31\]
rlabel via2 57696 12684 57696 12684 0 daisychain\[32\]
rlabel metal3 58704 11172 58704 11172 0 daisychain\[33\]
rlabel metal2 58080 8778 58080 8778 0 daisychain\[34\]
rlabel metal3 59328 7014 59328 7014 0 daisychain\[35\]
rlabel metal2 61296 4116 61296 4116 0 daisychain\[36\]
rlabel metal2 55968 3864 55968 3864 0 daisychain\[37\]
rlabel metal3 55776 2100 55776 2100 0 daisychain\[38\]
rlabel metal2 59808 2478 59808 2478 0 daisychain\[39\]
rlabel metal2 33312 19320 33312 19320 0 daisychain\[3\]
rlabel metal2 64128 1386 64128 1386 0 daisychain\[40\]
rlabel metal2 65280 3696 65280 3696 0 daisychain\[41\]
rlabel metal2 66144 6846 66144 6846 0 daisychain\[42\]
rlabel metal2 64416 7686 64416 7686 0 daisychain\[43\]
rlabel metal2 64608 9072 64608 9072 0 daisychain\[44\]
rlabel metal3 61872 11676 61872 11676 0 daisychain\[45\]
rlabel metal2 61632 13482 61632 13482 0 daisychain\[46\]
rlabel metal2 65136 13188 65136 13188 0 daisychain\[47\]
rlabel metal2 70080 14322 70080 14322 0 daisychain\[48\]
rlabel metal3 69216 13188 69216 13188 0 daisychain\[49\]
rlabel metal2 37776 20076 37776 20076 0 daisychain\[4\]
rlabel metal3 69120 10164 69120 10164 0 daisychain\[50\]
rlabel metal2 70752 8358 70752 8358 0 daisychain\[51\]
rlabel metal2 71424 5670 71424 5670 0 daisychain\[52\]
rlabel metal2 68400 1932 68400 1932 0 daisychain\[53\]
rlabel metal3 70848 3444 70848 3444 0 daisychain\[54\]
rlabel metal2 73824 2352 73824 2352 0 daisychain\[55\]
rlabel metal2 78048 2310 78048 2310 0 daisychain\[56\]
rlabel metal2 75936 4536 75936 4536 0 daisychain\[57\]
rlabel metal2 76608 6174 76608 6174 0 daisychain\[58\]
rlabel metal3 75744 7728 75744 7728 0 daisychain\[59\]
rlabel metal2 39360 20412 39360 20412 0 daisychain\[5\]
rlabel metal2 75936 10710 75936 10710 0 daisychain\[60\]
rlabel metal2 75024 11928 75024 11928 0 daisychain\[61\]
rlabel metal3 75504 13188 75504 13188 0 daisychain\[62\]
rlabel metal3 74592 13818 74592 13818 0 daisychain\[63\]
rlabel metal2 75744 25116 75744 25116 0 daisychain\[64\]
rlabel metal3 76272 26796 76272 26796 0 daisychain\[65\]
rlabel metal3 75792 29820 75792 29820 0 daisychain\[66\]
rlabel metal2 76032 30912 76032 30912 0 daisychain\[67\]
rlabel metal2 76992 33558 76992 33558 0 daisychain\[68\]
rlabel metal3 76416 34356 76416 34356 0 daisychain\[69\]
rlabel metal2 42624 20370 42624 20370 0 daisychain\[6\]
rlabel metal2 77376 37716 77376 37716 0 daisychain\[70\]
rlabel metal2 72192 36162 72192 36162 0 daisychain\[71\]
rlabel metal2 70368 34902 70368 34902 0 daisychain\[72\]
rlabel metal3 68064 36708 68064 36708 0 daisychain\[73\]
rlabel metal2 66624 34776 66624 34776 0 daisychain\[74\]
rlabel metal2 66144 32760 66144 32760 0 daisychain\[75\]
rlabel metal2 72096 32340 72096 32340 0 daisychain\[76\]
rlabel metal3 70416 29820 70416 29820 0 daisychain\[77\]
rlabel metal2 70656 29106 70656 29106 0 daisychain\[78\]
rlabel metal2 69312 26460 69312 26460 0 daisychain\[79\]
rlabel metal2 41952 16464 41952 16464 0 daisychain\[7\]
rlabel metal2 65760 26376 65760 26376 0 daisychain\[80\]
rlabel metal2 64032 25704 64032 25704 0 daisychain\[81\]
rlabel metal2 64320 28182 64320 28182 0 daisychain\[82\]
rlabel metal2 63264 30450 63264 30450 0 daisychain\[83\]
rlabel metal2 62496 33402 62496 33402 0 daisychain\[84\]
rlabel metal3 62064 34944 62064 34944 0 daisychain\[85\]
rlabel metal3 61152 36708 61152 36708 0 daisychain\[86\]
rlabel metal2 57600 36960 57600 36960 0 daisychain\[87\]
rlabel metal2 56352 35238 56352 35238 0 daisychain\[88\]
rlabel metal2 58656 33936 58656 33936 0 daisychain\[89\]
rlabel metal2 41184 14448 41184 14448 0 daisychain\[8\]
rlabel metal2 59616 31080 59616 31080 0 daisychain\[90\]
rlabel metal2 59712 26670 59712 26670 0 daisychain\[91\]
rlabel metal2 58080 24864 58080 24864 0 daisychain\[92\]
rlabel metal2 55680 27342 55680 27342 0 daisychain\[93\]
rlabel metal2 55392 29568 55392 29568 0 daisychain\[94\]
rlabel metal3 55440 31164 55440 31164 0 daisychain\[95\]
rlabel metal2 52512 33936 52512 33936 0 daisychain\[96\]
rlabel metal3 49248 34356 49248 34356 0 daisychain\[97\]
rlabel metal2 47040 33936 47040 33936 0 daisychain\[98\]
rlabel metal2 50496 31542 50496 31542 0 daisychain\[99\]
rlabel metal2 39168 14196 39168 14196 0 daisychain\[9\]
rlabel metal2 53675 17336 53675 17336 0 digitalen.g\[0\].u.OUTN
rlabel metal2 53565 17378 53565 17378 0 digitalen.g\[0\].u.OUTP
rlabel metal2 79008 16800 79008 16800 0 digitalen.g\[1\].u.OUTN
rlabel metal2 79488 16380 79488 16380 0 digitalen.g\[1\].u.OUTP
rlabel metal2 79565 22828 79565 22828 0 digitalen.g\[2\].u.OUTN
rlabel metal2 79675 22828 79675 22828 0 digitalen.g\[2\].u.OUTP
rlabel metal2 53565 22732 53565 22732 0 digitalen.g\[3\].u.OUTN
rlabel metal2 53675 22828 53675 22828 0 digitalen.g\[3\].u.OUTP
rlabel metal3 99924 21672 99924 21672 0 i_in
rlabel metal3 99924 19992 99924 19992 0 i_out
rlabel metal2 58608 14868 58608 14868 0 net
rlabel metal3 3024 20832 3024 20832 0 net1
rlabel metal2 912 10920 912 10920 0 net10
rlabel metal3 48096 13146 48096 13146 0 net100
rlabel metal2 40032 15834 40032 15834 0 net101
rlabel metal2 42912 18228 42912 18228 0 net102
rlabel metal3 57024 2604 57024 2604 0 net103
rlabel metal2 53472 6468 53472 6468 0 net104
rlabel metal2 53376 15036 53376 15036 0 net105
rlabel metal3 43008 18480 43008 18480 0 net106
rlabel metal2 45888 21882 45888 21882 0 net107
rlabel metal2 41184 20412 41184 20412 0 net108
rlabel metal2 49392 34356 49392 34356 0 net109
rlabel metal2 864 12390 864 12390 0 net11
rlabel metal2 57024 26208 57024 26208 0 net110
rlabel metal2 57984 35154 57984 35154 0 net111
rlabel metal2 52416 33768 52416 33768 0 net112
rlabel metal2 55392 27300 55392 27300 0 net113
rlabel metal2 42816 20832 42816 20832 0 net114
rlabel metal3 64272 2604 64272 2604 0 net115
rlabel metal2 59520 10122 59520 10122 0 net116
rlabel metal2 59328 12474 59328 12474 0 net117
rlabel metal2 70848 10080 70848 10080 0 net118
rlabel metal2 78672 1932 78672 1932 0 net119
rlabel metal2 864 13314 864 13314 0 net12
rlabel metal2 77376 6720 77376 6720 0 net120
rlabel metal2 76512 9534 76512 9534 0 net121
rlabel via2 74980 13020 74980 13020 0 net122
rlabel metal2 62208 14868 62208 14868 0 net123
rlabel metal3 61056 33684 61056 33684 0 net124
rlabel metal3 59760 34104 59760 34104 0 net125
rlabel metal2 60576 28434 60576 28434 0 net126
rlabel metal2 74496 24780 74496 24780 0 net127
rlabel metal3 72096 35826 72096 35826 0 net128
rlabel metal3 76416 35910 76416 35910 0 net129
rlabel metal2 1296 14196 1296 14196 0 net13
rlabel metal2 77952 35868 77952 35868 0 net130
rlabel metal2 60960 27090 60960 27090 0 net131
rlabel metal2 4416 21000 4416 21000 0 net132
rlabel metal2 22176 18480 22176 18480 0 net133
rlabel metal2 21984 17934 21984 17934 0 net134
rlabel metal2 2592 16506 2592 16506 0 net135
rlabel metal2 31776 23268 31776 23268 0 net136
rlabel metal2 42288 17052 42288 17052 0 net137
rlabel metal3 46896 17052 46896 17052 0 net138
rlabel metal3 56832 2520 56832 2520 0 net139
rlabel metal3 1200 14952 1200 14952 0 net14
rlabel metal2 56064 15288 56064 15288 0 net140
rlabel metal2 51264 16884 51264 16884 0 net141
rlabel metal2 41760 23394 41760 23394 0 net142
rlabel metal2 55920 34356 55920 34356 0 net143
rlabel metal2 51840 35154 51840 35154 0 net144
rlabel metal2 41088 30114 41088 30114 0 net145
rlabel metal2 60864 4158 60864 4158 0 net146
rlabel metal2 61152 14658 61152 14658 0 net147
rlabel metal2 76800 2730 76800 2730 0 net148
rlabel metal2 75360 11592 75360 11592 0 net149
rlabel metal2 864 2730 864 2730 0 net15
rlabel metal2 60912 13944 60912 13944 0 net150
rlabel metal3 59472 24612 59472 24612 0 net151
rlabel metal2 62976 36666 62976 36666 0 net152
rlabel metal2 76224 30534 76224 30534 0 net153
rlabel metal2 76608 34524 76608 34524 0 net154
rlabel metal2 58896 24528 58896 24528 0 net155
rlabel metal2 3360 17010 3360 17010 0 net156
rlabel metal2 3936 15792 3936 15792 0 net157
rlabel metal3 22752 17766 22752 17766 0 net158
rlabel metal2 32160 23142 32160 23142 0 net159
rlabel metal2 864 3318 864 3318 0 net16
rlabel metal3 3120 23100 3120 23100 0 net160
rlabel metal2 39264 16002 39264 16002 0 net161
rlabel metal2 44352 19362 44352 19362 0 net162
rlabel metal2 56208 2436 56208 2436 0 net163
rlabel metal2 56448 14070 56448 14070 0 net164
rlabel metal2 40128 23604 40128 23604 0 net165
rlabel metal2 56688 36036 56688 36036 0 net166
rlabel metal2 51648 35868 51648 35868 0 net167
rlabel metal2 43104 30282 43104 30282 0 net168
rlabel metal3 58896 8652 58896 8652 0 net169
rlabel metal2 1248 4452 1248 4452 0 net17
rlabel metal3 62784 14490 62784 14490 0 net170
rlabel metal3 76608 3108 76608 3108 0 net171
rlabel via1 76331 11003 76331 11003 0 net172
rlabel metal3 59088 34608 59088 34608 0 net173
rlabel metal3 59904 28350 59904 28350 0 net174
rlabel metal2 77184 31668 77184 31668 0 net175
rlabel metal2 75840 25704 75840 25704 0 net176
rlabel metal2 62976 14826 62976 14826 0 net177
rlabel metal2 1824 23730 1824 23730 0 net178
rlabel metal2 2592 14784 2592 14784 0 net179
rlabel metal2 816 4200 816 4200 0 net18
rlabel metal2 22272 19110 22272 19110 0 net180
rlabel metal2 28032 20958 28032 20958 0 net181
rlabel metal2 4800 20076 4800 20076 0 net182
rlabel metal2 41376 14490 41376 14490 0 net183
rlabel metal2 47520 18522 47520 18522 0 net184
rlabel metal2 55776 4158 55776 4158 0 net185
rlabel metal3 43104 16926 43104 16926 0 net186
rlabel metal2 42432 20832 42432 20832 0 net187
rlabel metal2 46752 33684 46752 33684 0 net188
rlabel metal2 56160 35700 56160 35700 0 net189
rlabel metal2 912 4872 912 4872 0 net19
rlabel metal2 50688 33768 50688 33768 0 net190
rlabel metal3 50688 35952 50688 35952 0 net191
rlabel metal2 62880 1986 62880 1986 0 net192
rlabel metal2 57888 13116 57888 13116 0 net193
rlabel metal2 75888 924 75888 924 0 net194
rlabel metal2 74880 13272 74880 13272 0 net195
rlabel metal2 59040 37464 59040 37464 0 net196
rlabel metal3 60864 37968 60864 37968 0 net197
rlabel metal3 74976 30702 74976 30702 0 net198
rlabel metal2 75168 37212 75168 37212 0 net199
rlabel metal3 2208 20748 2208 20748 0 net2
rlabel metal2 816 6384 816 6384 0 net20
rlabel metal2 58560 38094 58560 38094 0 net200
rlabel metal2 5088 19866 5088 19866 0 net201
rlabel metal2 72672 14700 72672 14700 0 net202
rlabel metal2 68544 24864 68544 24864 0 net203
rlabel metal2 72384 13356 72384 13356 0 net204
rlabel metal2 57552 16380 57552 16380 0 net205
rlabel metal2 73008 10836 73008 10836 0 net206
rlabel metal2 51360 21084 51360 21084 0 net207
rlabel metal2 74016 9744 74016 9744 0 net208
rlabel metal2 53952 16170 53952 16170 0 net209
rlabel metal3 720 7224 720 7224 0 net21
rlabel metal2 74304 8400 74304 8400 0 net210
rlabel metal2 71616 24612 71616 24612 0 net211
rlabel metal2 74496 5964 74496 5964 0 net212
rlabel metal2 50784 18060 50784 18060 0 net213
rlabel metal2 74256 4788 74256 4788 0 net214
rlabel metal2 36480 27132 36480 27132 0 net215
rlabel metal2 76128 2352 76128 2352 0 net216
rlabel metal2 50112 19572 50112 19572 0 net217
rlabel metal2 71520 2352 71520 2352 0 net218
rlabel metal2 71904 27888 71904 27888 0 net219
rlabel metal2 1152 13746 1152 13746 0 net22
rlabel metal2 69408 4452 69408 4452 0 net220
rlabel metal2 46704 16380 46704 16380 0 net221
rlabel metal2 66528 1932 66528 1932 0 net222
rlabel metal2 52608 24108 52608 24108 0 net223
rlabel metal2 69408 6888 69408 6888 0 net224
rlabel metal2 48432 15372 48432 15372 0 net225
rlabel metal3 69456 8820 69456 8820 0 net226
rlabel metal2 72288 31080 72288 31080 0 net227
rlabel metal3 67584 10332 67584 10332 0 net228
rlabel metal2 49584 13188 49584 13188 0 net229
rlabel metal2 22368 19194 22368 19194 0 net23
rlabel metal2 67488 12180 67488 12180 0 net230
rlabel metal2 5424 6300 5424 6300 0 net231
rlabel metal2 68064 15036 68064 15036 0 net232
rlabel metal2 52512 13158 52512 13158 0 net233
rlabel metal2 65088 13356 65088 13356 0 net234
rlabel metal2 72720 32844 72720 32844 0 net235
rlabel metal2 62208 13713 62208 13713 0 net236
rlabel metal2 54384 10332 54384 10332 0 net237
rlabel metal2 62160 11844 62160 11844 0 net238
rlabel metal2 52800 25620 52800 25620 0 net239
rlabel metal2 31776 23982 31776 23982 0 net24
rlabel metal2 62400 9912 62400 9912 0 net240
rlabel metal2 54816 8988 54816 8988 0 net241
rlabel metal2 63072 7476 63072 7476 0 net242
rlabel metal2 67200 31836 67200 31836 0 net243
rlabel metal2 63264 5628 63264 5628 0 net244
rlabel metal2 55296 7056 55296 7056 0 net245
rlabel metal2 63264 3906 63264 3906 0 net246
rlabel metal2 36048 22932 36048 22932 0 net247
rlabel metal2 62160 2772 62160 2772 0 net248
rlabel metal2 52896 4452 52896 4452 0 net249
rlabel metal2 2496 15372 2496 15372 0 net25
rlabel metal3 60144 1260 60144 1260 0 net250
rlabel metal2 67824 34524 67824 34524 0 net251
rlabel metal2 54000 2772 54000 2772 0 net252
rlabel metal2 49536 6132 49536 6132 0 net253
rlabel metal2 55200 3864 55200 3864 0 net254
rlabel metal2 52512 28056 52512 28056 0 net255
rlabel metal2 59712 5502 59712 5502 0 net256
rlabel metal2 49344 7980 49344 7980 0 net257
rlabel metal2 57408 6720 57408 6720 0 net258
rlabel metal2 71424 37632 71424 37632 0 net259
rlabel metal2 41088 16968 41088 16968 0 net26
rlabel metal2 56448 8652 56448 8652 0 net260
rlabel metal2 47328 9744 47328 9744 0 net261
rlabel metal2 56352 11634 56352 11634 0 net262
rlabel metal3 5616 12348 5616 12348 0 net263
rlabel metal2 55296 12180 55296 12180 0 net264
rlabel metal2 45024 11424 45024 11424 0 net265
rlabel metal2 54288 16380 54288 16380 0 net266
rlabel metal2 72576 34692 72576 34692 0 net267
rlabel metal2 51648 13881 51648 13881 0 net268
rlabel metal2 42912 12012 42912 12012 0 net269
rlabel metal2 45600 15456 45600 15456 0 net27
rlabel metal2 49104 15372 49104 15372 0 net270
rlabel metal2 51696 30492 51696 30492 0 net271
rlabel metal2 46704 19908 46704 19908 0 net272
rlabel metal2 39744 12180 39744 12180 0 net273
rlabel metal2 43872 15792 43872 15792 0 net274
rlabel metal2 74112 36372 74112 36372 0 net275
rlabel metal2 45072 14868 45072 14868 0 net276
rlabel metal2 37344 13074 37344 13074 0 net277
rlabel metal2 45744 11844 45744 11844 0 net278
rlabel metal3 41808 22932 41808 22932 0 net279
rlabel metal2 55872 4032 55872 4032 0 net28
rlabel metal2 48960 11424 48960 11424 0 net280
rlabel metal2 30672 13860 30672 13860 0 net281
rlabel metal2 50304 9324 50304 9324 0 net282
rlabel metal2 78432 37464 78432 37464 0 net283
rlabel metal2 50976 8400 50976 8400 0 net284
rlabel metal2 34944 17892 34944 17892 0 net285
rlabel metal2 51888 7308 51888 7308 0 net286
rlabel metal2 51648 31836 51648 31836 0 net287
rlabel metal2 50112 4788 50112 4788 0 net288
rlabel metal2 37920 17472 37920 17472 0 net289
rlabel metal2 40416 19362 40416 19362 0 net29
rlabel metal2 46368 5376 46368 5376 0 net290
rlabel metal2 77808 36036 77808 36036 0 net291
rlabel metal2 45984 7476 45984 7476 0 net292
rlabel metal2 40896 15456 40896 15456 0 net293
rlabel metal2 44640 8988 44640 8988 0 net294
rlabel metal2 5520 4788 5520 4788 0 net295
rlabel metal3 41760 9324 41760 9324 0 net296
rlabel metal3 43680 13860 43680 13860 0 net297
rlabel metal2 40032 10500 40032 10500 0 net298
rlabel metal2 77856 33318 77856 33318 0 net299
rlabel metal2 1488 22932 1488 22932 0 net3
rlabel metal2 42528 21168 42528 21168 0 net30
rlabel metal2 37104 11844 37104 11844 0 net300
rlabel metal2 43584 17304 43584 17304 0 net301
rlabel metal2 34320 11844 34320 11844 0 net302
rlabel metal2 47328 32802 47328 32802 0 net303
rlabel metal2 33600 13398 33600 13398 0 net304
rlabel metal3 44400 19908 44400 19908 0 net305
rlabel metal2 31584 16548 31584 16548 0 net306
rlabel metal2 77664 30324 77664 30324 0 net307
rlabel metal2 35712 15246 35712 15246 0 net308
rlabel metal2 39456 18228 39456 18228 0 net309
rlabel metal2 42432 32340 42432 32340 0 net31
rlabel metal2 38112 15036 38112 15036 0 net310
rlabel metal2 41328 24444 41328 24444 0 net311
rlabel metal2 40800 13692 40800 13692 0 net312
rlabel metal2 36864 19404 36864 19404 0 net313
rlabel metal2 38400 19026 38400 19026 0 net314
rlabel metal2 77520 28476 77520 28476 0 net315
rlabel metal2 41952 20496 41952 20496 0 net316
rlabel metal2 33312 19908 33312 19908 0 net317
rlabel metal2 39456 21084 39456 21084 0 net318
rlabel metal2 52512 36204 52512 36204 0 net319
rlabel metal2 56304 34440 56304 34440 0 net32
rlabel metal2 35712 21084 35712 21084 0 net320
rlabel metal2 30816 17304 30816 17304 0 net321
rlabel metal2 32736 21084 32736 21084 0 net322
rlabel metal2 77520 27468 77520 27468 0 net323
rlabel metal2 29760 19572 29760 19572 0 net324
rlabel metal2 27600 16884 27600 16884 0 net325
rlabel metal3 26784 19908 26784 19908 0 net326
rlabel metal2 23040 19422 23040 19422 0 net327
rlabel metal2 24000 17304 24000 17304 0 net328
rlabel metal2 77136 24444 77136 24444 0 net329
rlabel metal2 48864 32382 48864 32382 0 net33
rlabel metal2 1824 15960 1824 15960 0 net330
rlabel metal2 55776 32844 55776 32844 0 net331
rlabel metal2 1872 13860 1872 13860 0 net332
rlabel metal2 76704 15036 76704 15036 0 net333
rlabel metal2 1920 12012 1920 12012 0 net334
rlabel metal2 42144 26376 42144 26376 0 net335
rlabel metal2 1488 8820 1488 8820 0 net336
rlabel metal3 77376 13356 77376 13356 0 net337
rlabel metal2 1392 7812 1392 7812 0 net338
rlabel metal2 56592 30492 56592 30492 0 net339
rlabel metal2 39168 26712 39168 26712 0 net34
rlabel metal2 1728 5964 1728 5964 0 net340
rlabel metal2 77376 12180 77376 12180 0 net341
rlabel metal2 1872 4284 1872 4284 0 net342
rlabel metal2 12720 19908 12720 19908 0 net343
rlabel metal2 9600 19740 9600 19740 0 net344
rlabel metal2 77664 10500 77664 10500 0 net345
rlabel metal3 26880 20916 26880 20916 0 net346
rlabel metal2 56784 28476 56784 28476 0 net347
rlabel metal2 28896 23520 28896 23520 0 net348
rlabel metal2 77856 8232 77856 8232 0 net349
rlabel metal2 62976 1428 62976 1428 0 net35
rlabel metal2 30240 24864 30240 24864 0 net350
rlabel metal2 42432 28644 42432 28644 0 net351
rlabel metal2 34272 26544 34272 26544 0 net352
rlabel metal2 77856 7266 77856 7266 0 net353
rlabel metal2 35424 23940 35424 23940 0 net354
rlabel metal2 55776 25284 55776 25284 0 net355
rlabel metal2 38880 22764 38880 22764 0 net356
rlabel metal3 77664 4788 77664 4788 0 net357
rlabel metal2 37680 24444 37680 24444 0 net358
rlabel metal2 5280 9744 5280 9744 0 net359
rlabel metal2 61536 13164 61536 13164 0 net36
rlabel metal2 38208 28056 38208 28056 0 net360
rlabel metal3 78720 2772 78720 2772 0 net361
rlabel metal2 38880 29568 38880 29568 0 net362
rlabel metal2 60960 24780 60960 24780 0 net363
rlabel metal2 40704 31668 40704 31668 0 net364
rlabel metal2 74976 2436 74976 2436 0 net365
rlabel metal2 44256 30156 44256 30156 0 net366
rlabel metal2 43872 32592 43872 32592 0 net367
rlabel metal2 44352 28056 44352 28056 0 net368
rlabel metal2 72432 4788 72432 4788 0 net369
rlabel metal3 75984 1092 75984 1092 0 net37
rlabel metal2 44112 25452 44112 25452 0 net370
rlabel metal2 61152 27300 61152 27300 0 net371
rlabel metal2 42816 24276 42816 24276 0 net372
rlabel metal2 69312 1596 69312 1596 0 net373
rlabel metal2 42912 22260 42912 22260 0 net374
rlabel metal2 29808 20916 29808 20916 0 net375
rlabel metal2 48144 22428 48144 22428 0 net376
rlabel metal2 72384 6888 72384 6888 0 net377
rlabel metal2 48576 24402 48576 24402 0 net378
rlabel metal2 61440 30366 61440 30366 0 net379
rlabel metal3 75696 7140 75696 7140 0 net38
rlabel metal3 48864 25956 48864 25956 0 net380
rlabel metal2 72192 8988 72192 8988 0 net381
rlabel metal2 49248 28056 49248 28056 0 net382
rlabel metal2 46848 29820 46848 29820 0 net383
rlabel metal2 48288 30156 48288 30156 0 net384
rlabel metal2 71328 10500 71328 10500 0 net385
rlabel metal2 48912 33516 48912 33516 0 net386
rlabel metal3 59088 33264 59088 33264 0 net387
rlabel metal2 47136 34692 47136 34692 0 net388
rlabel metal2 70944 13158 70944 13158 0 net389
rlabel metal2 61824 36834 61824 36834 0 net39
rlabel metal3 49920 36036 49920 36036 0 net390
rlabel metal2 5568 13692 5568 13692 0 net391
rlabel metal2 52032 34104 52032 34104 0 net392
rlabel metal2 71328 15288 71328 15288 0 net393
rlabel metal2 53376 30744 53376 30744 0 net394
rlabel metal2 55584 34860 55584 34860 0 net395
rlabel metal2 53472 28056 53472 28056 0 net396
rlabel metal2 65904 14868 65904 14868 0 net397
rlabel metal3 55584 25956 55584 25956 0 net398
rlabel metal2 47520 27636 47520 27636 0 net399
rlabel metal3 1440 23856 1440 23856 0 net4
rlabel metal2 60096 31458 60096 31458 0 net40
rlabel metal2 57840 25956 57840 25956 0 net400
rlabel metal2 61008 16380 61008 16380 0 net401
rlabel metal2 57552 26964 57552 26964 0 net402
rlabel metal2 59808 37338 59808 37338 0 net403
rlabel metal2 58656 30324 58656 30324 0 net404
rlabel metal2 65232 11844 65232 11844 0 net405
rlabel metal2 58464 34692 58464 34692 0 net406
rlabel metal2 33312 21840 33312 21840 0 net407
rlabel metal2 55200 37128 55200 37128 0 net408
rlabel metal2 65712 10836 65712 10836 0 net409
rlabel metal2 75072 30576 75072 30576 0 net41
rlabel metal3 57600 38052 57600 38052 0 net410
rlabel metal2 64224 37716 64224 37716 0 net411
rlabel metal2 61584 38052 61584 38052 0 net412
rlabel metal2 66480 7812 66480 7812 0 net413
rlabel metal2 60384 35616 60384 35616 0 net414
rlabel metal2 47568 25956 47568 25956 0 net415
rlabel metal2 61152 32592 61152 32592 0 net416
rlabel metal2 67152 5796 67152 5796 0 net417
rlabel metal2 63552 31080 63552 31080 0 net418
rlabel metal2 63552 35028 63552 35028 0 net419
rlabel metal2 75072 37254 75072 37254 0 net42
rlabel metal2 62400 28644 62400 28644 0 net420
rlabel metal2 66864 4788 66864 4788 0 net421
rlabel metal2 62112 26544 62112 26544 0 net422
rlabel metal2 5280 8400 5280 8400 0 net423
rlabel metal2 66432 26376 66432 26376 0 net424
rlabel metal2 64992 1596 64992 1596 0 net425
rlabel metal2 69456 27468 69456 27468 0 net426
rlabel metal2 63600 33516 63600 33516 0 net427
rlabel metal2 68256 28476 68256 28476 0 net428
rlabel metal2 60192 3864 60192 3864 0 net429
rlabel metal2 74304 15036 74304 15036 0 net43
rlabel metal2 68688 31500 68688 31500 0 net430
rlabel metal2 46848 23940 46848 23940 0 net431
rlabel metal2 69888 33318 69888 33318 0 net432
rlabel metal2 57120 2352 57120 2352 0 net433
rlabel metal3 66864 32844 66864 32844 0 net434
rlabel metal2 66528 30156 66528 30156 0 net435
rlabel metal2 64896 35196 64896 35196 0 net436
rlabel metal2 56640 5376 56640 5376 0 net437
rlabel metal2 66624 38052 66624 38052 0 net438
rlabel metal2 33408 22986 33408 22986 0 net439
rlabel metal4 22368 18522 22368 18522 0 net44
rlabel metal3 70176 36036 70176 36036 0 net440
rlabel metal2 61824 5208 61824 5208 0 net441
rlabel metal2 72192 38052 72192 38052 0 net442
rlabel metal2 66192 27468 66192 27468 0 net443
rlabel metal2 75888 38052 75888 38052 0 net444
rlabel metal2 60960 7308 60960 7308 0 net445
rlabel metal2 74688 34860 74688 34860 0 net446
rlabel metal2 46464 22008 46464 22008 0 net447
rlabel metal2 75168 33180 75168 33180 0 net448
rlabel metal2 60096 9156 60096 9156 0 net449
rlabel metal2 33216 14784 33216 14784 0 net45
rlabel metal2 74064 32004 74064 32004 0 net450
rlabel metal3 64944 24444 64944 24444 0 net451
rlabel metal2 73920 29568 73920 29568 0 net452
rlabel metal2 59808 12012 59808 12012 0 net453
rlabel metal2 73536 27300 73536 27300 0 net454
rlabel metal2 5040 15372 5040 15372 0 net455
rlabel metal2 73536 25452 73536 25452 0 net456
rlabel metal3 366 15708 366 15708 0 net457
rlabel metal3 366 16548 366 16548 0 net458
rlabel metal3 366 17388 366 17388 0 net459
rlabel metal2 35088 20076 35088 20076 0 net46
rlabel metal3 366 18228 366 18228 0 net460
rlabel metal3 366 19068 366 19068 0 net461
rlabel metal3 366 19908 366 19908 0 net462
rlabel metal3 366 20748 366 20748 0 net463
rlabel metal3 366 21588 366 21588 0 net464
rlabel metal2 31248 23772 31248 23772 0 net47
rlabel metal2 2832 2604 2832 2604 0 net48
rlabel via2 42048 18396 42048 18396 0 net49
rlabel metal3 2400 25116 2400 25116 0 net5
rlabel metal2 55776 2646 55776 2646 0 net50
rlabel metal2 56352 13146 56352 13146 0 net51
rlabel metal2 41760 18228 41760 18228 0 net52
rlabel metal2 41520 21168 41520 21168 0 net53
rlabel metal2 49248 34314 49248 34314 0 net54
rlabel metal2 55200 27678 55200 27678 0 net55
rlabel metal2 41472 30618 41472 30618 0 net56
rlabel metal2 62016 1050 62016 1050 0 net57
rlabel metal2 58752 10290 58752 10290 0 net58
rlabel metal3 75648 3444 75648 3444 0 net59
rlabel metal3 4032 25956 4032 25956 0 net6
rlabel metal2 74784 12558 74784 12558 0 net60
rlabel metal2 58848 26376 58848 26376 0 net61
rlabel metal2 75744 29862 75744 29862 0 net62
rlabel metal2 74304 36666 74304 36666 0 net63
rlabel metal2 60048 35028 60048 35028 0 net64
rlabel metal2 74784 14406 74784 14406 0 net65
rlabel metal2 3648 21462 3648 21462 0 net66
rlabel metal2 38592 18858 38592 18858 0 net67
rlabel metal2 34080 17094 34080 17094 0 net68
rlabel metal2 35808 22314 35808 22314 0 net69
rlabel metal2 1536 17796 1536 17796 0 net7
rlabel metal2 4032 16548 4032 16548 0 net70
rlabel metal3 42480 14700 42480 14700 0 net71
rlabel metal2 46272 16254 46272 16254 0 net72
rlabel metal2 53760 11382 53760 11382 0 net73
rlabel metal2 58896 13188 58896 13188 0 net74
rlabel metal2 50496 18396 50496 18396 0 net75
rlabel metal2 41136 22092 41136 22092 0 net76
rlabel metal2 52128 35112 52128 35112 0 net77
rlabel metal2 51552 29610 51552 29610 0 net78
rlabel metal2 42192 29148 42192 29148 0 net79
rlabel metal2 720 9660 720 9660 0 net8
rlabel metal2 59088 2604 59088 2604 0 net80
rlabel metal2 78144 2394 78144 2394 0 net81
rlabel metal2 76560 13188 76560 13188 0 net82
rlabel metal2 60576 14742 60576 14742 0 net83
rlabel metal2 60480 25494 60480 25494 0 net84
rlabel metal2 62688 36246 62688 36246 0 net85
rlabel metal2 77040 29820 77040 29820 0 net86
rlabel metal3 74496 37338 74496 37338 0 net87
rlabel metal2 60384 14994 60384 14994 0 net88
rlabel metal2 4224 16338 4224 16338 0 net89
rlabel metal2 1248 10878 1248 10878 0 net9
rlabel metal2 3024 2604 3024 2604 0 net90
rlabel metal3 4416 17052 4416 17052 0 net91
rlabel metal3 36864 13188 36864 13188 0 net92
rlabel metal3 37680 17976 37680 17976 0 net93
rlabel metal3 37920 17808 37920 17808 0 net94
rlabel metal2 32976 24612 32976 24612 0 net95
rlabel metal3 37584 22932 37584 22932 0 net96
rlabel metal2 30912 23898 30912 23898 0 net97
rlabel metal2 3648 20622 3648 20622 0 net98
rlabel metal2 42336 10668 42336 10668 0 net99
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal2 23616 17304 23616 17304 0 state\[0\]
rlabel metal2 54048 26754 54048 26754 0 state\[100\]
rlabel metal2 54528 27888 54528 27888 0 state\[101\]
rlabel metal2 54720 25620 54720 25620 0 state\[102\]
rlabel metal2 63264 23688 63264 23688 0 state\[103\]
rlabel metal2 63275 22828 63275 22828 0 state\[104\]
rlabel metal2 62875 22828 62875 22828 0 state\[105\]
rlabel metal2 62475 22828 62475 22828 0 state\[106\]
rlabel metal2 62075 22828 62075 22828 0 state\[107\]
rlabel metal2 61675 22828 61675 22828 0 state\[108\]
rlabel metal2 61275 22828 61275 22828 0 state\[109\]
rlabel metal2 37152 16968 37152 16968 0 state\[10\]
rlabel metal2 43199 30880 43199 30880 0 state\[110\]
rlabel metal2 41376 28056 41376 28056 0 state\[111\]
rlabel metal2 41472 26586 41472 26586 0 state\[112\]
rlabel metal2 41184 24738 41184 24738 0 state\[113\]
rlabel metal2 41376 21756 41376 21756 0 state\[114\]
rlabel metal2 38112 22134 38112 22134 0 state\[115\]
rlabel metal2 38400 25872 38400 25872 0 state\[116\]
rlabel metal2 32736 24444 32736 24444 0 state\[117\]
rlabel metal2 35232 21882 35232 21882 0 state\[118\]
rlabel metal2 57275 22828 57275 22828 0 state\[119\]
rlabel metal2 34080 16464 34080 16464 0 state\[11\]
rlabel metal2 10944 18522 10944 18522 0 state\[120\]
rlabel metal2 56475 22828 56475 22828 0 state\[121\]
rlabel metal2 56062 23016 56062 23016 0 state\[122\]
rlabel metal2 55675 22828 55675 22828 0 state\[123\]
rlabel metal2 55275 22828 55275 22828 0 state\[124\]
rlabel metal3 2400 13272 2400 13272 0 state\[125\]
rlabel metal2 3552 14112 3552 14112 0 state\[126\]
rlabel metal2 3264 14658 3264 14658 0 state\[127\]
rlabel metal4 58560 15372 58560 15372 0 state\[12\]
rlabel metal2 36768 13272 36768 13272 0 state\[13\]
rlabel metal2 59280 16212 59280 16212 0 state\[14\]
rlabel metal2 59965 17294 59965 17294 0 state\[15\]
rlabel metal2 60365 17252 60365 17252 0 state\[16\]
rlabel metal2 60765 17294 60765 17294 0 state\[17\]
rlabel metal2 60768 15876 60768 15876 0 state\[18\]
rlabel metal2 61440 15876 61440 15876 0 state\[19\]
rlabel metal2 54365 17294 54365 17294 0 state\[1\]
rlabel metal2 62112 15204 62112 15204 0 state\[20\]
rlabel metal2 62352 16212 62352 16212 0 state\[21\]
rlabel metal3 62880 16212 62880 16212 0 state\[22\]
rlabel metal2 62928 16212 62928 16212 0 state\[23\]
rlabel metal2 63347 16038 63347 16038 0 state\[24\]
rlabel metal2 55776 14742 55776 14742 0 state\[25\]
rlabel metal2 50400 14994 50400 14994 0 state\[26\]
rlabel metal3 49728 16968 49728 16968 0 state\[27\]
rlabel metal3 51888 19068 51888 19068 0 state\[28\]
rlabel metal2 50688 17178 50688 17178 0 state\[29\]
rlabel metal4 54720 16422 54720 16422 0 state\[2\]
rlabel metal2 55488 16044 55488 16044 0 state\[30\]
rlabel metal2 59520 15792 59520 15792 0 state\[31\]
rlabel metal2 60576 14238 60576 14238 0 state\[32\]
rlabel metal2 61728 11970 61728 11970 0 state\[33\]
rlabel metal2 62016 9954 62016 9954 0 state\[34\]
rlabel via2 62880 8652 62880 8652 0 state\[35\]
rlabel metal2 61632 6174 61632 6174 0 state\[36\]
rlabel metal2 56544 4452 56544 4452 0 state\[37\]
rlabel metal2 56880 2604 56880 2604 0 state\[38\]
rlabel metal2 59712 2646 59712 2646 0 state\[39\]
rlabel metal2 35328 18564 35328 18564 0 state\[3\]
rlabel metal3 65088 2604 65088 2604 0 state\[40\]
rlabel metal2 70365 17294 70365 17294 0 state\[41\]
rlabel metal2 70560 16128 70560 16128 0 state\[42\]
rlabel metal2 70944 16044 70944 16044 0 state\[43\]
rlabel metal2 71376 16212 71376 16212 0 state\[44\]
rlabel metal2 71965 17294 71965 17294 0 state\[45\]
rlabel metal3 62976 15666 62976 15666 0 state\[46\]
rlabel metal2 72576 16674 72576 16674 0 state\[47\]
rlabel metal2 72960 16674 72960 16674 0 state\[48\]
rlabel metal2 73565 17336 73565 17336 0 state\[49\]
rlabel metal2 38592 18270 38592 18270 0 state\[4\]
rlabel metal2 73632 16212 73632 16212 0 state\[50\]
rlabel metal2 74352 16212 74352 16212 0 state\[51\]
rlabel metal2 74592 15078 74592 15078 0 state\[52\]
rlabel metal2 74976 16674 74976 16674 0 state\[53\]
rlabel metal2 75408 16212 75408 16212 0 state\[54\]
rlabel metal2 74400 2646 74400 2646 0 state\[55\]
rlabel metal3 78912 1974 78912 1974 0 state\[56\]
rlabel metal3 77376 16212 77376 16212 0 state\[57\]
rlabel metal2 77184 15876 77184 15876 0 state\[58\]
rlabel metal2 77565 17252 77565 17252 0 state\[59\]
rlabel metal2 41184 17808 41184 17808 0 state\[5\]
rlabel metal2 77965 17252 77965 17252 0 state\[60\]
rlabel metal2 78288 16212 78288 16212 0 state\[61\]
rlabel metal2 78624 16674 78624 16674 0 state\[62\]
rlabel metal2 79200 16632 79200 16632 0 state\[63\]
rlabel metal2 79275 22828 79275 22828 0 state\[64\]
rlabel metal3 78749 22764 78749 22764 0 state\[65\]
rlabel metal2 78453 22848 78453 22848 0 state\[66\]
rlabel metal2 78075 22828 78075 22828 0 state\[67\]
rlabel metal2 77675 22828 77675 22828 0 state\[68\]
rlabel metal3 78816 34356 78816 34356 0 state\[69\]
rlabel metal2 43104 19068 43104 19068 0 state\[6\]
rlabel metal2 76875 22690 76875 22690 0 state\[70\]
rlabel metal2 76475 22828 76475 22828 0 state\[71\]
rlabel metal2 74496 33852 74496 33852 0 state\[72\]
rlabel metal2 75675 22828 75675 22828 0 state\[73\]
rlabel metal2 75275 22828 75275 22828 0 state\[74\]
rlabel metal2 74875 22732 74875 22732 0 state\[75\]
rlabel metal2 74475 22828 74475 22828 0 state\[76\]
rlabel metal2 74075 22828 74075 22828 0 state\[77\]
rlabel metal2 73675 22828 73675 22828 0 state\[78\]
rlabel metal2 73275 22828 73275 22828 0 state\[79\]
rlabel metal2 43193 16261 43193 16261 0 state\[7\]
rlabel metal2 72875 22828 72875 22828 0 state\[80\]
rlabel metal2 72475 22828 72475 22828 0 state\[81\]
rlabel metal2 72075 22828 72075 22828 0 state\[82\]
rlabel metal2 71675 22828 71675 22828 0 state\[83\]
rlabel metal2 71275 22828 71275 22828 0 state\[84\]
rlabel metal2 70875 22828 70875 22828 0 state\[85\]
rlabel metal2 63264 36582 63264 36582 0 state\[86\]
rlabel metal2 61536 36078 61536 36078 0 state\[87\]
rlabel metal2 57600 34902 57600 34902 0 state\[88\]
rlabel metal2 60960 32550 60960 32550 0 state\[89\]
rlabel metal2 56880 16212 56880 16212 0 state\[8\]
rlabel metal2 62976 29316 62976 29316 0 state\[90\]
rlabel metal2 62880 26964 62880 26964 0 state\[91\]
rlabel metal2 62688 24948 62688 24948 0 state\[92\]
rlabel metal2 57312 24234 57312 24234 0 state\[93\]
rlabel metal2 58752 28770 58752 28770 0 state\[94\]
rlabel metal2 58560 30744 58560 30744 0 state\[95\]
rlabel metal2 57696 31710 57696 31710 0 state\[96\]
rlabel metal2 52800 35238 52800 35238 0 state\[97\]
rlabel metal2 57216 28014 57216 28014 0 state\[98\]
rlabel metal2 53568 31878 53568 31878 0 state\[99\]
rlabel metal2 39840 16128 39840 16128 0 state\[9\]
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 25788 366 25788 0 ui_in[4]
rlabel metal2 672 8946 672 8946 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 558 10668 558 10668 0 uio_out[2]
rlabel metal2 672 11340 672 11340 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 558 3948 558 3948 0 uo_out[2]
rlabel metal2 672 4536 672 4536 0 uo_out[3]
rlabel metal2 672 5376 672 5376 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
