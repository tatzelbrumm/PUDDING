magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771901320
<< metal1 >>
rect 576 38576 79584 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 79584 38576
rect 576 38512 79584 38536
rect 57667 38240 57725 38241
rect 57667 38200 57676 38240
rect 57716 38200 57725 38240
rect 57667 38199 57725 38200
rect 59875 38240 59933 38241
rect 59875 38200 59884 38240
rect 59924 38200 59933 38240
rect 59875 38199 59933 38200
rect 61227 38240 61269 38249
rect 61227 38200 61228 38240
rect 61268 38200 61269 38240
rect 61227 38191 61269 38200
rect 61419 38240 61461 38249
rect 61419 38200 61420 38240
rect 61460 38200 61461 38240
rect 61419 38191 61461 38200
rect 61507 38240 61565 38241
rect 61507 38200 61516 38240
rect 61556 38200 61565 38240
rect 61507 38199 61565 38200
rect 64675 38240 64733 38241
rect 64675 38200 64684 38240
rect 64724 38200 64733 38240
rect 64675 38199 64733 38200
rect 65259 38240 65301 38249
rect 65259 38200 65260 38240
rect 65300 38200 65301 38240
rect 65259 38191 65301 38200
rect 65451 38240 65493 38249
rect 65451 38200 65452 38240
rect 65492 38200 65493 38240
rect 65451 38191 65493 38200
rect 65539 38240 65597 38241
rect 65539 38200 65548 38240
rect 65588 38200 65597 38240
rect 65539 38199 65597 38200
rect 65731 38240 65789 38241
rect 65731 38200 65740 38240
rect 65780 38200 65789 38240
rect 65731 38199 65789 38200
rect 66891 38240 66933 38249
rect 66891 38200 66892 38240
rect 66932 38200 66933 38240
rect 66891 38191 66933 38200
rect 68331 38240 68373 38249
rect 68331 38200 68332 38240
rect 68372 38200 68373 38240
rect 68331 38191 68373 38200
rect 68707 38240 68765 38241
rect 68707 38200 68716 38240
rect 68756 38200 68765 38240
rect 68707 38199 68765 38200
rect 69579 38240 69621 38249
rect 69579 38200 69580 38240
rect 69620 38200 69621 38240
rect 69579 38191 69621 38200
rect 69963 38240 70005 38249
rect 69963 38200 69964 38240
rect 70004 38200 70005 38240
rect 69963 38191 70005 38200
rect 70059 38240 70101 38249
rect 70059 38200 70060 38240
rect 70100 38200 70101 38240
rect 70059 38191 70101 38200
rect 70155 38240 70197 38249
rect 70155 38200 70156 38240
rect 70196 38200 70197 38240
rect 70155 38191 70197 38200
rect 70251 38240 70293 38249
rect 70251 38200 70252 38240
rect 70292 38200 70293 38240
rect 70251 38191 70293 38200
rect 73995 38240 74037 38249
rect 73995 38200 73996 38240
rect 74036 38200 74037 38240
rect 73995 38191 74037 38200
rect 74187 38240 74229 38249
rect 74187 38200 74188 38240
rect 74228 38200 74229 38240
rect 74187 38191 74229 38200
rect 74275 38240 74333 38241
rect 74275 38200 74284 38240
rect 74324 38200 74333 38240
rect 74275 38199 74333 38200
rect 74475 38240 74517 38249
rect 74475 38200 74476 38240
rect 74516 38200 74517 38240
rect 74475 38191 74517 38200
rect 74571 38240 74613 38249
rect 74571 38200 74572 38240
rect 74612 38200 74613 38240
rect 74571 38191 74613 38200
rect 74667 38240 74709 38249
rect 74667 38200 74668 38240
rect 74708 38200 74709 38240
rect 74667 38191 74709 38200
rect 74763 38240 74805 38249
rect 74763 38200 74764 38240
rect 74804 38200 74805 38240
rect 74763 38191 74805 38200
rect 75619 38240 75677 38241
rect 75619 38200 75628 38240
rect 75668 38200 75677 38240
rect 75619 38199 75677 38200
rect 75907 38240 75965 38241
rect 75907 38200 75916 38240
rect 75956 38200 75965 38240
rect 75907 38199 75965 38200
rect 643 38156 701 38157
rect 643 38116 652 38156
rect 692 38116 701 38156
rect 643 38115 701 38116
rect 64867 38156 64925 38157
rect 64867 38116 64876 38156
rect 64916 38116 64925 38156
rect 64867 38115 64925 38116
rect 70435 38156 70493 38157
rect 70435 38116 70444 38156
rect 70484 38116 70493 38156
rect 70435 38115 70493 38116
rect 71011 38156 71069 38157
rect 71011 38116 71020 38156
rect 71060 38116 71069 38156
rect 71011 38115 71069 38116
rect 77251 38156 77309 38157
rect 77251 38116 77260 38156
rect 77300 38116 77309 38156
rect 77251 38115 77309 38116
rect 67755 38072 67797 38081
rect 67755 38032 67756 38072
rect 67796 38032 67797 38072
rect 67755 38023 67797 38032
rect 843 37988 885 37997
rect 843 37948 844 37988
rect 884 37948 885 37988
rect 843 37939 885 37948
rect 57579 37988 57621 37997
rect 57579 37948 57580 37988
rect 57620 37948 57621 37988
rect 57579 37939 57621 37948
rect 59979 37988 60021 37997
rect 59979 37948 59980 37988
rect 60020 37948 60021 37988
rect 59979 37939 60021 37948
rect 61227 37988 61269 37997
rect 61227 37948 61228 37988
rect 61268 37948 61269 37988
rect 61227 37939 61269 37948
rect 65067 37988 65109 37997
rect 65067 37948 65068 37988
rect 65108 37948 65109 37988
rect 65067 37939 65109 37948
rect 65259 37988 65301 37997
rect 65259 37948 65260 37988
rect 65300 37948 65301 37988
rect 65259 37939 65301 37948
rect 65835 37988 65877 37997
rect 65835 37948 65836 37988
rect 65876 37948 65877 37988
rect 65835 37939 65877 37948
rect 66699 37988 66741 37997
rect 66699 37948 66700 37988
rect 66740 37948 66741 37988
rect 66699 37939 66741 37948
rect 70635 37988 70677 37997
rect 70635 37948 70636 37988
rect 70676 37948 70677 37988
rect 70635 37939 70677 37948
rect 70827 37988 70869 37997
rect 70827 37948 70828 37988
rect 70868 37948 70869 37988
rect 70827 37939 70869 37948
rect 73995 37988 74037 37997
rect 73995 37948 73996 37988
rect 74036 37948 74037 37988
rect 73995 37939 74037 37948
rect 76203 37988 76245 37997
rect 76203 37948 76204 37988
rect 76244 37948 76245 37988
rect 76203 37939 76245 37948
rect 77451 37988 77493 37997
rect 77451 37948 77452 37988
rect 77492 37948 77493 37988
rect 77451 37939 77493 37948
rect 576 37820 79584 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 79584 37820
rect 576 37756 79584 37780
rect 73131 37568 73173 37577
rect 73131 37528 73132 37568
rect 73172 37528 73173 37568
rect 73131 37519 73173 37528
rect 56619 37484 56661 37493
rect 56619 37444 56620 37484
rect 56660 37444 56661 37484
rect 56619 37435 56661 37444
rect 56811 37484 56853 37493
rect 56811 37444 56812 37484
rect 56852 37444 56853 37484
rect 56811 37435 56853 37444
rect 57091 37484 57149 37485
rect 57091 37444 57100 37484
rect 57140 37444 57149 37484
rect 57091 37443 57149 37444
rect 60259 37484 60317 37485
rect 60259 37444 60268 37484
rect 60308 37444 60317 37484
rect 60259 37443 60317 37444
rect 64203 37484 64245 37493
rect 64203 37444 64204 37484
rect 64244 37444 64245 37484
rect 64099 37442 64157 37443
rect 56515 37400 56573 37401
rect 56515 37360 56524 37400
rect 56564 37360 56573 37400
rect 56515 37359 56573 37360
rect 56907 37400 56949 37409
rect 64099 37402 64108 37442
rect 64148 37402 64157 37442
rect 64203 37435 64245 37444
rect 64395 37484 64437 37493
rect 64395 37444 64396 37484
rect 64436 37444 64437 37484
rect 64395 37435 64437 37444
rect 67363 37484 67421 37485
rect 67363 37444 67372 37484
rect 67412 37444 67421 37484
rect 67363 37443 67421 37444
rect 64099 37401 64157 37402
rect 56907 37360 56908 37400
rect 56948 37360 56949 37400
rect 56907 37351 56949 37360
rect 58627 37400 58685 37401
rect 58627 37360 58636 37400
rect 58676 37360 58685 37400
rect 58627 37359 58685 37360
rect 59491 37400 59549 37401
rect 59491 37360 59500 37400
rect 59540 37360 59549 37400
rect 59491 37359 59549 37360
rect 60931 37400 60989 37401
rect 60931 37360 60940 37400
rect 60980 37360 60989 37400
rect 60931 37359 60989 37360
rect 61795 37400 61853 37401
rect 61795 37360 61804 37400
rect 61844 37360 61853 37400
rect 61795 37359 61853 37360
rect 64491 37400 64533 37409
rect 64491 37360 64492 37400
rect 64532 37360 64533 37400
rect 64491 37351 64533 37360
rect 65923 37400 65981 37401
rect 65923 37360 65932 37400
rect 65972 37360 65981 37400
rect 65923 37359 65981 37360
rect 66787 37400 66845 37401
rect 66787 37360 66796 37400
rect 66836 37360 66845 37400
rect 66787 37359 66845 37360
rect 68899 37400 68957 37401
rect 68899 37360 68908 37400
rect 68948 37360 68957 37400
rect 68899 37359 68957 37360
rect 69763 37400 69821 37401
rect 69763 37360 69772 37400
rect 69812 37360 69821 37400
rect 69763 37359 69821 37360
rect 70155 37400 70197 37409
rect 70155 37360 70156 37400
rect 70196 37360 70197 37400
rect 70155 37351 70197 37360
rect 71491 37400 71549 37401
rect 71491 37360 71500 37400
rect 71540 37360 71549 37400
rect 71491 37359 71549 37360
rect 72355 37400 72413 37401
rect 72355 37360 72364 37400
rect 72404 37360 72413 37400
rect 72355 37359 72413 37360
rect 73419 37400 73461 37409
rect 73419 37360 73420 37400
rect 73460 37360 73461 37400
rect 73419 37351 73461 37360
rect 73507 37400 73565 37401
rect 73507 37360 73516 37400
rect 73556 37360 73565 37400
rect 73507 37359 73565 37360
rect 74179 37400 74237 37401
rect 74179 37360 74188 37400
rect 74228 37360 74237 37400
rect 74179 37359 74237 37360
rect 75043 37400 75101 37401
rect 75043 37360 75052 37400
rect 75092 37360 75101 37400
rect 75043 37359 75101 37360
rect 76579 37400 76637 37401
rect 76579 37360 76588 37400
rect 76628 37360 76637 37400
rect 76579 37359 76637 37360
rect 77155 37400 77213 37401
rect 77155 37360 77164 37400
rect 77204 37360 77213 37400
rect 77155 37359 77213 37360
rect 78019 37400 78077 37401
rect 78019 37360 78028 37400
rect 78068 37360 78077 37400
rect 78019 37359 78077 37360
rect 59883 37316 59925 37325
rect 56715 37274 56757 37283
rect 56715 37234 56716 37274
rect 56756 37234 56757 37274
rect 59883 37276 59884 37316
rect 59924 37276 59925 37316
rect 59883 37267 59925 37276
rect 60555 37316 60597 37325
rect 60555 37276 60556 37316
rect 60596 37276 60597 37316
rect 67179 37316 67221 37325
rect 60555 37267 60597 37276
rect 64299 37274 64341 37283
rect 56715 37225 56757 37234
rect 57291 37232 57333 37241
rect 57291 37192 57292 37232
rect 57332 37192 57333 37232
rect 57291 37183 57333 37192
rect 57475 37232 57533 37233
rect 57475 37192 57484 37232
rect 57524 37192 57533 37232
rect 57475 37191 57533 37192
rect 60075 37232 60117 37241
rect 64299 37234 64300 37274
rect 64340 37234 64341 37274
rect 67179 37276 67180 37316
rect 67220 37276 67221 37316
rect 67179 37267 67221 37276
rect 72747 37316 72789 37325
rect 72747 37276 72748 37316
rect 72788 37276 72789 37316
rect 72747 37267 72789 37276
rect 73803 37316 73845 37325
rect 73803 37276 73804 37316
rect 73844 37276 73845 37316
rect 73803 37267 73845 37276
rect 76779 37316 76821 37325
rect 76779 37276 76780 37316
rect 76820 37276 76821 37316
rect 76779 37267 76821 37276
rect 60075 37192 60076 37232
rect 60116 37192 60117 37232
rect 60075 37183 60117 37192
rect 62947 37232 63005 37233
rect 62947 37192 62956 37232
rect 62996 37192 63005 37232
rect 64299 37225 64341 37234
rect 64771 37232 64829 37233
rect 62947 37191 63005 37192
rect 64771 37192 64780 37232
rect 64820 37192 64829 37232
rect 64771 37191 64829 37192
rect 67563 37232 67605 37241
rect 67563 37192 67564 37232
rect 67604 37192 67605 37232
rect 67563 37183 67605 37192
rect 67747 37232 67805 37233
rect 67747 37192 67756 37232
rect 67796 37192 67805 37232
rect 67747 37191 67805 37192
rect 70339 37232 70397 37233
rect 70339 37192 70348 37232
rect 70388 37192 70397 37232
rect 70339 37191 70397 37192
rect 76195 37232 76253 37233
rect 76195 37192 76204 37232
rect 76244 37192 76253 37232
rect 76195 37191 76253 37192
rect 76491 37232 76533 37241
rect 76491 37192 76492 37232
rect 76532 37192 76533 37232
rect 76491 37183 76533 37192
rect 79171 37232 79229 37233
rect 79171 37192 79180 37232
rect 79220 37192 79229 37232
rect 79171 37191 79229 37192
rect 73611 37174 73653 37183
rect 73611 37134 73612 37174
rect 73652 37134 73653 37174
rect 73611 37125 73653 37134
rect 576 37064 79584 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 79584 37064
rect 576 37000 79584 37024
rect 67659 36954 67701 36963
rect 67659 36914 67660 36954
rect 67700 36914 67701 36954
rect 59403 36896 59445 36905
rect 59403 36856 59404 36896
rect 59444 36856 59445 36896
rect 59403 36847 59445 36856
rect 60171 36900 60213 36909
rect 67659 36905 67701 36914
rect 60171 36860 60172 36900
rect 60212 36860 60213 36900
rect 60171 36851 60213 36860
rect 60835 36896 60893 36897
rect 60835 36856 60844 36896
rect 60884 36856 60893 36896
rect 60835 36855 60893 36856
rect 69387 36896 69429 36905
rect 69387 36856 69388 36896
rect 69428 36856 69429 36896
rect 69387 36847 69429 36856
rect 74083 36896 74141 36897
rect 74083 36856 74092 36896
rect 74132 36856 74141 36896
rect 74083 36855 74141 36856
rect 56235 36812 56277 36821
rect 56235 36772 56236 36812
rect 56276 36772 56277 36812
rect 56235 36763 56277 36772
rect 64107 36812 64149 36821
rect 64107 36772 64108 36812
rect 64148 36772 64149 36812
rect 64107 36763 64149 36772
rect 73323 36812 73365 36821
rect 73323 36772 73324 36812
rect 73364 36772 73365 36812
rect 73323 36763 73365 36772
rect 56611 36728 56669 36729
rect 56611 36688 56620 36728
rect 56660 36688 56669 36728
rect 56611 36687 56669 36688
rect 57475 36728 57533 36729
rect 57475 36688 57484 36728
rect 57524 36688 57533 36728
rect 57475 36687 57533 36688
rect 59595 36728 59637 36737
rect 59595 36688 59596 36728
rect 59636 36688 59637 36728
rect 59595 36679 59637 36688
rect 59971 36728 60029 36729
rect 59971 36688 59980 36728
rect 60020 36688 60029 36728
rect 59971 36687 60029 36688
rect 60259 36728 60317 36729
rect 60259 36688 60268 36728
rect 60308 36688 60317 36728
rect 60259 36687 60317 36688
rect 60363 36728 60405 36737
rect 60363 36688 60364 36728
rect 60404 36688 60405 36728
rect 60363 36679 60405 36688
rect 60939 36728 60981 36737
rect 60939 36688 60940 36728
rect 60980 36688 60981 36728
rect 60939 36679 60981 36688
rect 61035 36728 61077 36737
rect 61035 36688 61036 36728
rect 61076 36688 61077 36728
rect 61035 36679 61077 36688
rect 61131 36728 61173 36737
rect 61131 36688 61132 36728
rect 61172 36688 61173 36728
rect 61131 36679 61173 36688
rect 62851 36728 62909 36729
rect 62851 36688 62860 36728
rect 62900 36688 62909 36728
rect 62851 36687 62909 36688
rect 63715 36728 63773 36729
rect 63715 36688 63724 36728
rect 63764 36688 63773 36728
rect 63715 36687 63773 36688
rect 64299 36728 64341 36737
rect 64299 36688 64300 36728
rect 64340 36688 64341 36728
rect 64299 36679 64341 36688
rect 64675 36728 64733 36729
rect 64675 36688 64684 36728
rect 64724 36688 64733 36728
rect 64675 36687 64733 36688
rect 65539 36728 65597 36729
rect 65539 36688 65548 36728
rect 65588 36688 65597 36728
rect 65539 36687 65597 36688
rect 67083 36728 67125 36737
rect 67083 36688 67084 36728
rect 67124 36688 67125 36728
rect 67083 36679 67125 36688
rect 67459 36728 67517 36729
rect 67459 36688 67468 36728
rect 67508 36688 67517 36728
rect 67459 36687 67517 36688
rect 67747 36728 67805 36729
rect 67747 36688 67756 36728
rect 67796 36688 67805 36728
rect 67747 36687 67805 36688
rect 67851 36728 67893 36737
rect 67851 36688 67852 36728
rect 67892 36688 67893 36728
rect 67851 36679 67893 36688
rect 68331 36728 68373 36737
rect 68331 36688 68332 36728
rect 68372 36688 68373 36728
rect 68331 36679 68373 36688
rect 68523 36728 68565 36737
rect 68523 36688 68524 36728
rect 68564 36688 68565 36728
rect 68523 36679 68565 36688
rect 68611 36728 68669 36729
rect 68611 36688 68620 36728
rect 68660 36688 68669 36728
rect 68611 36687 68669 36688
rect 68811 36728 68853 36737
rect 68811 36688 68812 36728
rect 68852 36688 68853 36728
rect 68811 36679 68853 36688
rect 68907 36728 68949 36737
rect 68907 36688 68908 36728
rect 68948 36688 68949 36728
rect 68907 36679 68949 36688
rect 69003 36728 69045 36737
rect 69003 36688 69004 36728
rect 69044 36688 69045 36728
rect 69003 36679 69045 36688
rect 69099 36728 69141 36737
rect 69099 36688 69100 36728
rect 69140 36688 69141 36728
rect 69099 36679 69141 36688
rect 69283 36728 69341 36729
rect 69283 36688 69292 36728
rect 69332 36688 69341 36728
rect 69283 36687 69341 36688
rect 70723 36728 70781 36729
rect 70723 36688 70732 36728
rect 70772 36688 70781 36728
rect 70723 36687 70781 36688
rect 71587 36728 71645 36729
rect 71587 36688 71596 36728
rect 71636 36688 71645 36728
rect 71587 36687 71645 36688
rect 71979 36728 72021 36737
rect 71979 36688 71980 36728
rect 72020 36688 72021 36728
rect 71979 36679 72021 36688
rect 72171 36728 72213 36737
rect 72171 36688 72172 36728
rect 72212 36688 72213 36728
rect 72171 36679 72213 36688
rect 72547 36728 72605 36729
rect 72547 36688 72556 36728
rect 72596 36688 72605 36728
rect 72547 36687 72605 36688
rect 72747 36728 72789 36737
rect 72747 36688 72748 36728
rect 72788 36688 72789 36728
rect 72747 36679 72789 36688
rect 72939 36728 72981 36737
rect 72939 36688 72940 36728
rect 72980 36688 72981 36728
rect 72939 36679 72981 36688
rect 73027 36728 73085 36729
rect 73027 36688 73036 36728
rect 73076 36688 73085 36728
rect 73027 36687 73085 36688
rect 73219 36728 73277 36729
rect 73219 36688 73228 36728
rect 73268 36688 73277 36728
rect 73219 36687 73277 36688
rect 73507 36728 73565 36729
rect 73507 36688 73516 36728
rect 73556 36688 73565 36728
rect 73507 36687 73565 36688
rect 73899 36728 73941 36737
rect 73899 36688 73900 36728
rect 73940 36688 73941 36728
rect 73899 36679 73941 36688
rect 74187 36728 74229 36737
rect 74187 36688 74188 36728
rect 74228 36688 74229 36728
rect 74187 36679 74229 36688
rect 74283 36728 74325 36737
rect 74283 36688 74284 36728
rect 74324 36688 74325 36728
rect 74283 36679 74325 36688
rect 74379 36728 74421 36737
rect 74379 36688 74380 36728
rect 74420 36688 74421 36728
rect 74379 36679 74421 36688
rect 75331 36728 75389 36729
rect 75331 36688 75340 36728
rect 75380 36688 75389 36728
rect 75331 36687 75389 36688
rect 75627 36728 75669 36737
rect 75627 36688 75628 36728
rect 75668 36688 75669 36728
rect 75627 36679 75669 36688
rect 75723 36728 75765 36737
rect 75723 36688 75724 36728
rect 75764 36688 75765 36728
rect 75723 36679 75765 36688
rect 75819 36728 75861 36737
rect 75819 36688 75820 36728
rect 75860 36688 75861 36728
rect 75819 36679 75861 36688
rect 75915 36728 75957 36737
rect 75915 36688 75916 36728
rect 75956 36688 75957 36728
rect 75915 36679 75957 36688
rect 76099 36728 76157 36729
rect 76099 36688 76108 36728
rect 76148 36688 76157 36728
rect 76099 36687 76157 36688
rect 76491 36728 76533 36737
rect 76491 36688 76492 36728
rect 76532 36688 76533 36728
rect 76491 36679 76533 36688
rect 76683 36728 76725 36737
rect 76683 36688 76684 36728
rect 76724 36688 76725 36728
rect 76683 36679 76725 36688
rect 77059 36728 77117 36729
rect 77059 36688 77068 36728
rect 77108 36688 77117 36728
rect 77059 36687 77117 36688
rect 77923 36728 77981 36729
rect 77923 36688 77932 36728
rect 77972 36688 77981 36728
rect 77923 36687 77981 36688
rect 58819 36644 58877 36645
rect 58819 36604 58828 36644
rect 58868 36604 58877 36644
rect 58819 36603 58877 36604
rect 59203 36644 59261 36645
rect 59203 36604 59212 36644
rect 59252 36604 59261 36644
rect 59203 36603 59261 36604
rect 59691 36644 59733 36653
rect 59691 36604 59692 36644
rect 59732 36604 59733 36644
rect 59691 36595 59733 36604
rect 59883 36644 59925 36653
rect 59883 36604 59884 36644
rect 59924 36604 59925 36644
rect 59883 36595 59925 36604
rect 67179 36644 67221 36653
rect 67179 36604 67180 36644
rect 67220 36604 67221 36644
rect 67179 36595 67221 36604
rect 67371 36644 67413 36653
rect 67371 36604 67372 36644
rect 67412 36604 67413 36644
rect 67371 36595 67413 36604
rect 72267 36644 72309 36653
rect 72267 36604 72268 36644
rect 72308 36604 72309 36644
rect 72267 36595 72309 36604
rect 72459 36644 72501 36653
rect 72459 36604 72460 36644
rect 72500 36604 72501 36644
rect 72459 36595 72501 36604
rect 73611 36644 73653 36653
rect 73611 36604 73612 36644
rect 73652 36604 73653 36644
rect 73611 36595 73653 36604
rect 73803 36644 73845 36653
rect 73803 36604 73804 36644
rect 73844 36604 73845 36644
rect 73803 36595 73845 36604
rect 74563 36644 74621 36645
rect 74563 36604 74572 36644
rect 74612 36604 74621 36644
rect 74563 36603 74621 36604
rect 76203 36644 76245 36653
rect 76203 36604 76204 36644
rect 76244 36604 76245 36644
rect 76203 36595 76245 36604
rect 76395 36644 76437 36653
rect 76395 36604 76396 36644
rect 76436 36604 76437 36644
rect 76395 36595 76437 36604
rect 58627 36560 58685 36561
rect 58627 36520 58636 36560
rect 58676 36520 58685 36560
rect 58627 36519 58685 36520
rect 59787 36560 59829 36569
rect 59787 36520 59788 36560
rect 59828 36520 59829 36560
rect 59787 36511 59829 36520
rect 60651 36560 60693 36569
rect 60651 36520 60652 36560
rect 60692 36520 60693 36560
rect 60651 36511 60693 36520
rect 67275 36560 67317 36569
rect 67275 36520 67276 36560
rect 67316 36520 67317 36560
rect 67275 36511 67317 36520
rect 68139 36560 68181 36569
rect 68139 36520 68140 36560
rect 68180 36520 68181 36560
rect 68139 36511 68181 36520
rect 68331 36560 68373 36569
rect 68331 36520 68332 36560
rect 68372 36520 68373 36560
rect 68331 36511 68373 36520
rect 72363 36560 72405 36569
rect 72363 36520 72364 36560
rect 72404 36520 72405 36560
rect 72363 36511 72405 36520
rect 72747 36560 72789 36569
rect 72747 36520 72748 36560
rect 72788 36520 72789 36560
rect 72747 36511 72789 36520
rect 73707 36560 73749 36569
rect 73707 36520 73708 36560
rect 73748 36520 73749 36560
rect 73707 36511 73749 36520
rect 74763 36560 74805 36569
rect 74763 36520 74764 36560
rect 74804 36520 74805 36560
rect 74763 36511 74805 36520
rect 76299 36560 76341 36569
rect 76299 36520 76300 36560
rect 76340 36520 76341 36560
rect 76299 36511 76341 36520
rect 59019 36476 59061 36485
rect 59019 36436 59020 36476
rect 59060 36436 59061 36476
rect 59019 36427 59061 36436
rect 59403 36476 59445 36485
rect 59403 36436 59404 36476
rect 59444 36436 59445 36476
rect 59403 36427 59445 36436
rect 61699 36476 61757 36477
rect 61699 36436 61708 36476
rect 61748 36436 61757 36476
rect 61699 36435 61757 36436
rect 66691 36476 66749 36477
rect 66691 36436 66700 36476
rect 66740 36436 66749 36476
rect 66691 36435 66749 36436
rect 69571 36476 69629 36477
rect 69571 36436 69580 36476
rect 69620 36436 69629 36476
rect 69571 36435 69629 36436
rect 75435 36476 75477 36485
rect 75435 36436 75436 36476
rect 75476 36436 75477 36476
rect 75435 36427 75477 36436
rect 79075 36476 79133 36477
rect 79075 36436 79084 36476
rect 79124 36436 79133 36476
rect 79075 36435 79133 36436
rect 576 36308 79584 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 79584 36308
rect 576 36244 79584 36268
rect 56427 36140 56469 36149
rect 56427 36100 56428 36140
rect 56468 36100 56469 36140
rect 56427 36091 56469 36100
rect 63915 36140 63957 36149
rect 63915 36100 63916 36140
rect 63956 36100 63957 36140
rect 63915 36091 63957 36100
rect 72171 36140 72213 36149
rect 72171 36100 72172 36140
rect 72212 36100 72213 36140
rect 72171 36091 72213 36100
rect 72939 36140 72981 36149
rect 72939 36100 72940 36140
rect 72980 36100 72981 36140
rect 72939 36091 72981 36100
rect 77259 36140 77301 36149
rect 77259 36100 77260 36140
rect 77300 36100 77301 36140
rect 77259 36091 77301 36100
rect 77451 36140 77493 36149
rect 77451 36100 77452 36140
rect 77492 36100 77493 36140
rect 77451 36091 77493 36100
rect 64587 36056 64629 36065
rect 64587 36016 64588 36056
rect 64628 36016 64629 36056
rect 64587 36007 64629 36016
rect 74275 35972 74333 35973
rect 74275 35932 74284 35972
rect 74324 35932 74333 35972
rect 74275 35931 74333 35932
rect 74659 35972 74717 35973
rect 74659 35932 74668 35972
rect 74708 35932 74717 35972
rect 74659 35931 74717 35932
rect 56043 35888 56085 35897
rect 56043 35848 56044 35888
rect 56084 35848 56085 35888
rect 56043 35839 56085 35848
rect 56139 35888 56181 35897
rect 56139 35848 56140 35888
rect 56180 35848 56181 35888
rect 56139 35839 56181 35848
rect 56235 35888 56277 35897
rect 56235 35848 56236 35888
rect 56276 35848 56277 35888
rect 56235 35839 56277 35848
rect 56715 35888 56757 35897
rect 56715 35848 56716 35888
rect 56756 35848 56757 35888
rect 56715 35839 56757 35848
rect 56803 35888 56861 35889
rect 56803 35848 56812 35888
rect 56852 35848 56861 35888
rect 56803 35847 56861 35848
rect 57099 35888 57141 35897
rect 57099 35848 57100 35888
rect 57140 35848 57141 35888
rect 57099 35839 57141 35848
rect 57195 35888 57237 35897
rect 57195 35848 57196 35888
rect 57236 35848 57237 35888
rect 57195 35839 57237 35848
rect 57291 35888 57333 35897
rect 57291 35848 57292 35888
rect 57332 35848 57333 35888
rect 57675 35888 57717 35897
rect 57291 35839 57333 35848
rect 57387 35867 57429 35876
rect 57387 35827 57388 35867
rect 57428 35827 57429 35867
rect 57675 35848 57676 35888
rect 57716 35848 57717 35888
rect 57675 35839 57717 35848
rect 57867 35888 57909 35897
rect 57867 35848 57868 35888
rect 57908 35848 57909 35888
rect 57867 35839 57909 35848
rect 57955 35888 58013 35889
rect 57955 35848 57964 35888
rect 58004 35848 58013 35888
rect 57955 35847 58013 35848
rect 58147 35888 58205 35889
rect 58147 35848 58156 35888
rect 58196 35848 58205 35888
rect 58147 35847 58205 35848
rect 58251 35888 58293 35897
rect 58251 35848 58252 35888
rect 58292 35848 58293 35888
rect 58251 35839 58293 35848
rect 58443 35888 58485 35897
rect 58443 35848 58444 35888
rect 58484 35848 58485 35888
rect 58443 35839 58485 35848
rect 59011 35888 59069 35889
rect 59011 35848 59020 35888
rect 59060 35848 59069 35888
rect 59011 35847 59069 35848
rect 59875 35888 59933 35889
rect 59875 35848 59884 35888
rect 59924 35848 59933 35888
rect 59875 35847 59933 35848
rect 61227 35888 61269 35897
rect 61227 35848 61228 35888
rect 61268 35848 61269 35888
rect 61227 35839 61269 35848
rect 61323 35888 61365 35897
rect 61323 35848 61324 35888
rect 61364 35848 61365 35888
rect 61323 35839 61365 35848
rect 61419 35888 61461 35897
rect 61419 35848 61420 35888
rect 61460 35848 61461 35888
rect 61419 35839 61461 35848
rect 61515 35888 61557 35897
rect 61515 35848 61516 35888
rect 61556 35848 61557 35888
rect 63811 35888 63869 35889
rect 61515 35839 61557 35848
rect 61699 35877 61757 35878
rect 61699 35837 61708 35877
rect 61748 35837 61757 35877
rect 63811 35848 63820 35888
rect 63860 35848 63869 35888
rect 63811 35847 63869 35848
rect 64195 35888 64253 35889
rect 64195 35848 64204 35888
rect 64244 35848 64253 35888
rect 64195 35847 64253 35848
rect 64299 35888 64341 35897
rect 64299 35848 64300 35888
rect 64340 35848 64341 35888
rect 64299 35839 64341 35848
rect 64779 35888 64821 35897
rect 64779 35848 64780 35888
rect 64820 35848 64821 35888
rect 64779 35839 64821 35848
rect 64875 35888 64917 35897
rect 64875 35848 64876 35888
rect 64916 35848 64917 35888
rect 64875 35839 64917 35848
rect 64971 35888 65013 35897
rect 64971 35848 64972 35888
rect 65012 35848 65013 35888
rect 64971 35839 65013 35848
rect 65067 35888 65109 35897
rect 65067 35848 65068 35888
rect 65108 35848 65109 35888
rect 65067 35839 65109 35848
rect 65259 35888 65301 35897
rect 65259 35848 65260 35888
rect 65300 35848 65301 35888
rect 65259 35839 65301 35848
rect 65355 35888 65397 35897
rect 65355 35848 65356 35888
rect 65396 35848 65397 35888
rect 65355 35839 65397 35848
rect 65451 35888 65493 35897
rect 65451 35848 65452 35888
rect 65492 35848 65493 35888
rect 65451 35839 65493 35848
rect 65547 35888 65589 35897
rect 65547 35848 65548 35888
rect 65588 35848 65589 35888
rect 65547 35839 65589 35848
rect 65827 35888 65885 35889
rect 65827 35848 65836 35888
rect 65876 35848 65885 35888
rect 65827 35847 65885 35848
rect 66787 35888 66845 35889
rect 66787 35848 66796 35888
rect 66836 35848 66845 35888
rect 66787 35847 66845 35848
rect 67651 35888 67709 35889
rect 67651 35848 67660 35888
rect 67700 35848 67709 35888
rect 67651 35847 67709 35848
rect 71299 35888 71357 35889
rect 71299 35848 71308 35888
rect 71348 35848 71357 35888
rect 71299 35847 71357 35848
rect 71403 35888 71445 35897
rect 71403 35848 71404 35888
rect 71444 35848 71445 35888
rect 71403 35839 71445 35848
rect 71595 35888 71637 35897
rect 71595 35848 71596 35888
rect 71636 35848 71637 35888
rect 71595 35839 71637 35848
rect 72067 35888 72125 35889
rect 72067 35848 72076 35888
rect 72116 35848 72125 35888
rect 72067 35847 72125 35848
rect 72547 35888 72605 35889
rect 72547 35848 72556 35888
rect 72596 35848 72605 35888
rect 72547 35847 72605 35848
rect 72651 35888 72693 35897
rect 72651 35848 72652 35888
rect 72692 35848 72693 35888
rect 72651 35839 72693 35848
rect 73803 35888 73845 35897
rect 73803 35848 73804 35888
rect 73844 35848 73845 35888
rect 73803 35839 73845 35848
rect 73899 35888 73941 35897
rect 73899 35848 73900 35888
rect 73940 35848 73941 35888
rect 73899 35839 73941 35848
rect 73995 35888 74037 35897
rect 73995 35848 73996 35888
rect 74036 35848 74037 35888
rect 73995 35839 74037 35848
rect 74091 35888 74133 35897
rect 74091 35848 74092 35888
rect 74132 35848 74133 35888
rect 74091 35839 74133 35848
rect 76299 35888 76341 35897
rect 76299 35848 76300 35888
rect 76340 35848 76341 35888
rect 76299 35839 76341 35848
rect 76395 35888 76437 35897
rect 76395 35848 76396 35888
rect 76436 35848 76437 35888
rect 76395 35839 76437 35848
rect 76491 35888 76533 35897
rect 76491 35848 76492 35888
rect 76532 35848 76533 35888
rect 76491 35839 76533 35848
rect 76587 35888 76629 35897
rect 76587 35848 76588 35888
rect 76628 35848 76629 35888
rect 76587 35839 76629 35848
rect 76867 35888 76925 35889
rect 76867 35848 76876 35888
rect 76916 35848 76925 35888
rect 76867 35847 76925 35848
rect 76971 35888 77013 35897
rect 76971 35848 76972 35888
rect 77012 35848 77013 35888
rect 76971 35839 77013 35848
rect 77451 35888 77493 35897
rect 77451 35848 77452 35888
rect 77492 35848 77493 35888
rect 77451 35839 77493 35848
rect 77643 35888 77685 35897
rect 77643 35848 77644 35888
rect 77684 35848 77685 35888
rect 77643 35839 77685 35848
rect 77731 35888 77789 35889
rect 77731 35848 77740 35888
rect 77780 35848 77789 35888
rect 77731 35847 77789 35848
rect 78019 35888 78077 35889
rect 78019 35848 78028 35888
rect 78068 35848 78077 35888
rect 78019 35847 78077 35848
rect 61699 35836 61757 35837
rect 57387 35818 57429 35827
rect 57771 35804 57813 35813
rect 57771 35764 57772 35804
rect 57812 35764 57813 35804
rect 57771 35755 57813 35764
rect 58635 35804 58677 35813
rect 58635 35764 58636 35804
rect 58676 35764 58677 35804
rect 58635 35755 58677 35764
rect 66411 35804 66453 35813
rect 66411 35764 66412 35804
rect 66452 35764 66453 35804
rect 66411 35755 66453 35764
rect 55939 35720 55997 35721
rect 55939 35680 55948 35720
rect 55988 35680 55997 35720
rect 55939 35679 55997 35680
rect 56907 35716 56949 35725
rect 56907 35676 56908 35716
rect 56948 35676 56949 35716
rect 58339 35720 58397 35721
rect 58339 35680 58348 35720
rect 58388 35680 58397 35720
rect 58339 35679 58397 35680
rect 61027 35720 61085 35721
rect 61027 35680 61036 35720
rect 61076 35680 61085 35720
rect 61027 35679 61085 35680
rect 61803 35720 61845 35729
rect 61803 35680 61804 35720
rect 61844 35680 61845 35720
rect 56907 35667 56949 35676
rect 61803 35671 61845 35680
rect 63915 35720 63957 35729
rect 63915 35680 63916 35720
rect 63956 35680 63957 35720
rect 63915 35671 63957 35680
rect 64107 35716 64149 35725
rect 64107 35676 64108 35716
rect 64148 35676 64149 35716
rect 64107 35667 64149 35676
rect 65739 35720 65781 35729
rect 65739 35680 65740 35720
rect 65780 35680 65781 35720
rect 65739 35671 65781 35680
rect 68803 35720 68861 35721
rect 68803 35680 68812 35720
rect 68852 35680 68861 35720
rect 68803 35679 68861 35680
rect 71491 35720 71549 35721
rect 71491 35680 71500 35720
rect 71540 35680 71549 35720
rect 71491 35679 71549 35680
rect 72459 35716 72501 35725
rect 72459 35676 72460 35716
rect 72500 35676 72501 35716
rect 72459 35667 72501 35676
rect 74475 35720 74517 35729
rect 74475 35680 74476 35720
rect 74516 35680 74517 35720
rect 74475 35671 74517 35680
rect 74859 35720 74901 35729
rect 74859 35680 74860 35720
rect 74900 35680 74901 35720
rect 74859 35671 74901 35680
rect 76779 35716 76821 35725
rect 76779 35676 76780 35716
rect 76820 35676 76821 35716
rect 76779 35667 76821 35676
rect 77931 35720 77973 35729
rect 77931 35680 77932 35720
rect 77972 35680 77973 35720
rect 77931 35671 77973 35680
rect 576 35552 79584 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 79584 35552
rect 576 35488 79584 35512
rect 59403 35388 59445 35397
rect 57475 35384 57533 35385
rect 57475 35344 57484 35384
rect 57524 35344 57533 35384
rect 57475 35343 57533 35344
rect 59403 35348 59404 35388
rect 59444 35348 59445 35388
rect 59403 35339 59445 35348
rect 60171 35384 60213 35393
rect 60171 35344 60172 35384
rect 60212 35344 60213 35384
rect 60171 35335 60213 35344
rect 75715 35384 75773 35385
rect 75715 35344 75724 35384
rect 75764 35344 75773 35384
rect 75715 35343 75773 35344
rect 79459 35384 79517 35385
rect 79459 35344 79468 35384
rect 79508 35344 79517 35384
rect 79459 35343 79517 35344
rect 55083 35300 55125 35309
rect 55083 35260 55084 35300
rect 55124 35260 55125 35300
rect 55083 35251 55125 35260
rect 72843 35300 72885 35309
rect 72843 35260 72844 35300
rect 72884 35260 72885 35300
rect 72843 35251 72885 35260
rect 73323 35300 73365 35309
rect 73323 35260 73324 35300
rect 73364 35260 73365 35300
rect 73323 35251 73365 35260
rect 55459 35216 55517 35217
rect 55459 35176 55468 35216
rect 55508 35176 55517 35216
rect 55459 35175 55517 35176
rect 56323 35216 56381 35217
rect 56323 35176 56332 35216
rect 56372 35176 56381 35216
rect 56323 35175 56381 35176
rect 58347 35216 58389 35225
rect 58347 35176 58348 35216
rect 58388 35176 58389 35216
rect 58347 35167 58389 35176
rect 58723 35216 58781 35217
rect 58723 35176 58732 35216
rect 58772 35176 58781 35216
rect 58723 35175 58781 35176
rect 59211 35216 59253 35225
rect 59211 35176 59212 35216
rect 59252 35176 59253 35216
rect 59211 35167 59253 35176
rect 59299 35216 59357 35217
rect 59299 35176 59308 35216
rect 59348 35176 59357 35216
rect 59299 35175 59357 35176
rect 60259 35216 60317 35217
rect 60259 35176 60268 35216
rect 60308 35176 60317 35216
rect 60259 35175 60317 35176
rect 61123 35216 61181 35217
rect 61123 35176 61132 35216
rect 61172 35176 61181 35216
rect 61123 35175 61181 35176
rect 61227 35216 61269 35225
rect 61227 35176 61228 35216
rect 61268 35176 61269 35216
rect 61227 35167 61269 35176
rect 61419 35216 61461 35225
rect 61419 35176 61420 35216
rect 61460 35176 61461 35216
rect 61419 35167 61461 35176
rect 61611 35216 61653 35225
rect 61611 35176 61612 35216
rect 61652 35176 61653 35216
rect 61611 35167 61653 35176
rect 61987 35216 62045 35217
rect 61987 35176 61996 35216
rect 62036 35176 62045 35216
rect 61987 35175 62045 35176
rect 62851 35216 62909 35217
rect 62851 35176 62860 35216
rect 62900 35176 62909 35216
rect 62851 35175 62909 35176
rect 68227 35216 68285 35217
rect 68227 35176 68236 35216
rect 68276 35176 68285 35216
rect 68227 35175 68285 35176
rect 70243 35216 70301 35217
rect 70243 35176 70252 35216
rect 70292 35176 70301 35216
rect 70243 35175 70301 35176
rect 71107 35216 71165 35217
rect 71107 35176 71116 35216
rect 71156 35176 71165 35216
rect 71107 35175 71165 35176
rect 71499 35216 71541 35225
rect 71499 35176 71500 35216
rect 71540 35176 71541 35216
rect 71499 35167 71541 35176
rect 71691 35216 71733 35225
rect 71691 35176 71692 35216
rect 71732 35176 71733 35216
rect 71691 35167 71733 35176
rect 72067 35216 72125 35217
rect 72067 35176 72076 35216
rect 72116 35176 72125 35216
rect 72067 35175 72125 35176
rect 72939 35216 72981 35225
rect 72939 35176 72940 35216
rect 72980 35176 72981 35216
rect 72939 35167 72981 35176
rect 73035 35216 73077 35225
rect 73035 35176 73036 35216
rect 73076 35176 73077 35216
rect 73035 35167 73077 35176
rect 73131 35216 73173 35225
rect 73131 35176 73132 35216
rect 73172 35176 73173 35216
rect 73131 35167 73173 35176
rect 73699 35216 73757 35217
rect 73699 35176 73708 35216
rect 73748 35176 73757 35216
rect 73699 35175 73757 35176
rect 74563 35216 74621 35217
rect 74563 35176 74572 35216
rect 74612 35176 74621 35216
rect 74563 35175 74621 35176
rect 76867 35216 76925 35217
rect 76867 35176 76876 35216
rect 76916 35176 76925 35216
rect 76867 35175 76925 35176
rect 77067 35216 77109 35225
rect 77067 35176 77068 35216
rect 77108 35176 77109 35216
rect 77067 35167 77109 35176
rect 77443 35216 77501 35217
rect 77443 35176 77452 35216
rect 77492 35176 77501 35216
rect 77443 35175 77501 35176
rect 78307 35216 78365 35217
rect 78307 35176 78316 35216
rect 78356 35176 78365 35216
rect 78307 35175 78365 35176
rect 58443 35132 58485 35141
rect 58443 35092 58444 35132
rect 58484 35092 58485 35132
rect 58443 35083 58485 35092
rect 58635 35132 58677 35141
rect 58635 35092 58636 35132
rect 58676 35092 58677 35132
rect 58635 35083 58677 35092
rect 71787 35132 71829 35141
rect 71787 35092 71788 35132
rect 71828 35092 71829 35132
rect 71787 35083 71829 35092
rect 71979 35132 72021 35141
rect 71979 35092 71980 35132
rect 72020 35092 72021 35132
rect 71979 35083 72021 35092
rect 58539 35048 58581 35057
rect 58539 35008 58540 35048
rect 58580 35008 58581 35048
rect 58539 34999 58581 35008
rect 58923 35048 58965 35057
rect 58923 35008 58924 35048
rect 58964 35008 58965 35048
rect 58923 34999 58965 35008
rect 71883 35048 71925 35057
rect 71883 35008 71884 35048
rect 71924 35008 71925 35048
rect 71883 34999 71925 35008
rect 57475 34964 57533 34965
rect 57475 34924 57484 34964
rect 57524 34924 57533 34964
rect 57475 34923 57533 34924
rect 61419 34964 61461 34973
rect 61419 34924 61420 34964
rect 61460 34924 61461 34964
rect 61419 34915 61461 34924
rect 64003 34964 64061 34965
rect 64003 34924 64012 34964
rect 64052 34924 64061 34964
rect 64003 34923 64061 34924
rect 68139 34964 68181 34973
rect 68139 34924 68140 34964
rect 68180 34924 68181 34964
rect 68139 34915 68181 34924
rect 69091 34964 69149 34965
rect 69091 34924 69100 34964
rect 69140 34924 69149 34964
rect 69091 34923 69149 34924
rect 76779 34964 76821 34973
rect 76779 34924 76780 34964
rect 76820 34924 76821 34964
rect 76779 34915 76821 34924
rect 576 34796 79584 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 79584 34796
rect 576 34732 79584 34756
rect 57291 34628 57333 34637
rect 57291 34588 57292 34628
rect 57332 34588 57333 34628
rect 57291 34579 57333 34588
rect 71019 34628 71061 34637
rect 71019 34588 71020 34628
rect 71060 34588 71061 34628
rect 71019 34579 71061 34588
rect 52107 34544 52149 34553
rect 52107 34504 52108 34544
rect 52148 34504 52149 34544
rect 52107 34495 52149 34504
rect 62475 34544 62517 34553
rect 62475 34504 62476 34544
rect 62516 34504 62517 34544
rect 62475 34495 62517 34504
rect 64011 34544 64053 34553
rect 64011 34504 64012 34544
rect 64052 34504 64053 34544
rect 67275 34544 67317 34553
rect 64011 34495 64053 34504
rect 67179 34502 67221 34511
rect 52011 34460 52053 34469
rect 52011 34420 52012 34460
rect 52052 34420 52053 34460
rect 52011 34411 52053 34420
rect 52203 34460 52245 34469
rect 52203 34420 52204 34460
rect 52244 34420 52245 34460
rect 52203 34411 52245 34420
rect 62379 34460 62421 34469
rect 62379 34420 62380 34460
rect 62420 34420 62421 34460
rect 62379 34411 62421 34420
rect 62571 34460 62613 34469
rect 62571 34420 62572 34460
rect 62612 34420 62613 34460
rect 67179 34462 67180 34502
rect 67220 34462 67221 34502
rect 67275 34504 67276 34544
rect 67316 34504 67317 34544
rect 67275 34495 67317 34504
rect 67659 34544 67701 34553
rect 67659 34504 67660 34544
rect 67700 34504 67701 34544
rect 67659 34495 67701 34504
rect 71691 34544 71733 34553
rect 71691 34504 71692 34544
rect 71732 34504 71733 34544
rect 71691 34495 71733 34504
rect 77547 34544 77589 34553
rect 77547 34504 77548 34544
rect 77588 34504 77589 34544
rect 77547 34495 77589 34504
rect 67179 34453 67221 34462
rect 67371 34460 67413 34469
rect 62571 34411 62613 34420
rect 67371 34420 67372 34460
rect 67412 34420 67413 34460
rect 67371 34411 67413 34420
rect 63341 34395 63399 34396
rect 51907 34376 51965 34377
rect 51907 34336 51916 34376
rect 51956 34336 51965 34376
rect 51907 34335 51965 34336
rect 52299 34376 52341 34385
rect 52299 34336 52300 34376
rect 52340 34336 52341 34376
rect 52299 34327 52341 34336
rect 52963 34376 53021 34377
rect 52963 34336 52972 34376
rect 53012 34336 53021 34376
rect 52963 34335 53021 34336
rect 53827 34376 53885 34377
rect 53827 34336 53836 34376
rect 53876 34336 53885 34376
rect 53827 34335 53885 34336
rect 55171 34376 55229 34377
rect 55171 34336 55180 34376
rect 55220 34336 55229 34376
rect 55171 34335 55229 34336
rect 55947 34376 55989 34385
rect 55947 34336 55948 34376
rect 55988 34336 55989 34376
rect 55947 34327 55989 34336
rect 56043 34376 56085 34385
rect 56043 34336 56044 34376
rect 56084 34336 56085 34376
rect 56043 34327 56085 34336
rect 56139 34376 56181 34385
rect 56139 34336 56140 34376
rect 56180 34336 56181 34376
rect 56139 34327 56181 34336
rect 57187 34376 57245 34377
rect 57187 34336 57196 34376
rect 57236 34336 57245 34376
rect 57187 34335 57245 34336
rect 58539 34376 58581 34385
rect 58539 34336 58540 34376
rect 58580 34336 58581 34376
rect 58539 34327 58581 34336
rect 58635 34376 58677 34385
rect 58635 34336 58636 34376
rect 58676 34336 58677 34376
rect 58635 34327 58677 34336
rect 58731 34376 58773 34385
rect 58731 34336 58732 34376
rect 58772 34336 58773 34376
rect 58731 34327 58773 34336
rect 59299 34376 59357 34377
rect 59299 34336 59308 34376
rect 59348 34336 59357 34376
rect 59299 34335 59357 34336
rect 60163 34376 60221 34377
rect 60163 34336 60172 34376
rect 60212 34336 60221 34376
rect 60163 34335 60221 34336
rect 62283 34376 62325 34385
rect 62283 34336 62284 34376
rect 62324 34336 62325 34376
rect 62283 34327 62325 34336
rect 62659 34376 62717 34377
rect 62659 34336 62668 34376
rect 62708 34336 62717 34376
rect 62659 34335 62717 34336
rect 63051 34376 63093 34385
rect 63051 34336 63052 34376
rect 63092 34336 63093 34376
rect 63051 34327 63093 34336
rect 63243 34376 63285 34385
rect 63243 34336 63244 34376
rect 63284 34336 63285 34376
rect 63341 34355 63350 34395
rect 63390 34355 63399 34395
rect 63341 34354 63399 34355
rect 63619 34376 63677 34377
rect 63243 34327 63285 34336
rect 63619 34336 63628 34376
rect 63668 34336 63677 34376
rect 63619 34335 63677 34336
rect 63723 34376 63765 34385
rect 63723 34336 63724 34376
rect 63764 34336 63765 34376
rect 63723 34327 63765 34336
rect 64675 34376 64733 34377
rect 64675 34336 64684 34376
rect 64724 34336 64733 34376
rect 64675 34335 64733 34336
rect 65539 34376 65597 34377
rect 65539 34336 65548 34376
rect 65588 34336 65597 34376
rect 65539 34335 65597 34336
rect 67083 34376 67125 34385
rect 67083 34336 67084 34376
rect 67124 34336 67125 34376
rect 67083 34327 67125 34336
rect 67459 34376 67517 34377
rect 67459 34336 67468 34376
rect 67508 34336 67517 34376
rect 67459 34335 67517 34336
rect 67947 34376 67989 34385
rect 67947 34336 67948 34376
rect 67988 34336 67989 34376
rect 67947 34327 67989 34336
rect 68035 34376 68093 34377
rect 68035 34336 68044 34376
rect 68084 34336 68093 34376
rect 68035 34335 68093 34336
rect 68619 34376 68661 34385
rect 68619 34336 68620 34376
rect 68660 34336 68661 34376
rect 68619 34327 68661 34336
rect 68715 34376 68757 34385
rect 68715 34336 68716 34376
rect 68756 34336 68757 34376
rect 68715 34327 68757 34336
rect 68811 34376 68853 34385
rect 68811 34336 68812 34376
rect 68852 34336 68853 34376
rect 68811 34327 68853 34336
rect 68907 34376 68949 34385
rect 68907 34336 68908 34376
rect 68948 34336 68949 34376
rect 68907 34327 68949 34336
rect 69667 34376 69725 34377
rect 69667 34336 69676 34376
rect 69716 34336 69725 34376
rect 69667 34335 69725 34336
rect 70915 34376 70973 34377
rect 70915 34336 70924 34376
rect 70964 34336 70973 34376
rect 70915 34335 70973 34336
rect 71299 34376 71357 34377
rect 71299 34336 71308 34376
rect 71348 34336 71357 34376
rect 71299 34335 71357 34336
rect 71403 34376 71445 34385
rect 71403 34336 71404 34376
rect 71444 34336 71445 34376
rect 71403 34327 71445 34336
rect 71979 34376 72021 34385
rect 71979 34336 71980 34376
rect 72020 34336 72021 34376
rect 71979 34327 72021 34336
rect 72075 34376 72117 34385
rect 72075 34336 72076 34376
rect 72116 34336 72117 34376
rect 72075 34327 72117 34336
rect 72171 34376 72213 34385
rect 72171 34336 72172 34376
rect 72212 34336 72213 34376
rect 72171 34327 72213 34336
rect 72739 34376 72797 34377
rect 72739 34336 72748 34376
rect 72788 34336 72797 34376
rect 72739 34335 72797 34336
rect 73603 34376 73661 34377
rect 73603 34336 73612 34376
rect 73652 34336 73661 34376
rect 73603 34335 73661 34336
rect 76099 34376 76157 34377
rect 76099 34336 76108 34376
rect 76148 34336 76157 34376
rect 76099 34335 76157 34336
rect 76963 34376 77021 34377
rect 76963 34336 76972 34376
rect 77012 34336 77021 34376
rect 76963 34335 77021 34336
rect 77835 34376 77877 34385
rect 77835 34336 77836 34376
rect 77876 34336 77877 34376
rect 77835 34327 77877 34336
rect 77923 34376 77981 34377
rect 77923 34336 77932 34376
rect 77972 34336 77981 34376
rect 77923 34335 77981 34336
rect 78219 34376 78261 34385
rect 78219 34336 78220 34376
rect 78260 34336 78261 34376
rect 78219 34327 78261 34336
rect 78315 34376 78357 34385
rect 78315 34336 78316 34376
rect 78356 34336 78357 34376
rect 78315 34327 78357 34336
rect 78411 34376 78453 34385
rect 78411 34336 78412 34376
rect 78452 34336 78453 34376
rect 78411 34327 78453 34336
rect 78507 34376 78549 34385
rect 78507 34336 78508 34376
rect 78548 34336 78549 34376
rect 78507 34327 78549 34336
rect 52587 34292 52629 34301
rect 52587 34252 52588 34292
rect 52628 34252 52629 34292
rect 52587 34243 52629 34252
rect 58923 34292 58965 34301
rect 58923 34252 58924 34292
rect 58964 34252 58965 34292
rect 58923 34243 58965 34252
rect 64299 34292 64341 34301
rect 64299 34252 64300 34292
rect 64340 34252 64341 34292
rect 64299 34243 64341 34252
rect 71883 34292 71925 34301
rect 71883 34252 71884 34292
rect 71924 34252 71925 34292
rect 71883 34243 71925 34252
rect 72363 34292 72405 34301
rect 72363 34252 72364 34292
rect 72404 34252 72405 34292
rect 72363 34243 72405 34252
rect 77355 34292 77397 34301
rect 77355 34252 77356 34292
rect 77396 34252 77397 34292
rect 77355 34243 77397 34252
rect 54979 34208 55037 34209
rect 54979 34168 54988 34208
rect 55028 34168 55037 34208
rect 54979 34167 55037 34168
rect 55275 34208 55317 34217
rect 55275 34168 55276 34208
rect 55316 34168 55317 34208
rect 55275 34159 55317 34168
rect 55843 34208 55901 34209
rect 55843 34168 55852 34208
rect 55892 34168 55901 34208
rect 55843 34167 55901 34168
rect 57291 34208 57333 34217
rect 57291 34168 57292 34208
rect 57332 34168 57333 34208
rect 57291 34159 57333 34168
rect 58435 34208 58493 34209
rect 58435 34168 58444 34208
rect 58484 34168 58493 34208
rect 58435 34167 58493 34168
rect 61315 34208 61373 34209
rect 61315 34168 61324 34208
rect 61364 34168 61373 34208
rect 61315 34167 61373 34168
rect 63139 34208 63197 34209
rect 63139 34168 63148 34208
rect 63188 34168 63197 34208
rect 63139 34167 63197 34168
rect 66691 34208 66749 34209
rect 66691 34168 66700 34208
rect 66740 34168 66749 34208
rect 66691 34167 66749 34168
rect 68139 34204 68181 34213
rect 68139 34164 68140 34204
rect 68180 34164 68181 34204
rect 63531 34150 63573 34159
rect 68139 34155 68181 34164
rect 69579 34208 69621 34217
rect 69579 34168 69580 34208
rect 69620 34168 69621 34208
rect 69579 34159 69621 34168
rect 71211 34204 71253 34213
rect 71211 34164 71212 34204
rect 71252 34164 71253 34204
rect 74755 34208 74813 34209
rect 74755 34168 74764 34208
rect 74804 34168 74813 34208
rect 74755 34167 74813 34168
rect 74947 34208 75005 34209
rect 74947 34168 74956 34208
rect 74996 34168 75005 34208
rect 74947 34167 75005 34168
rect 78027 34204 78069 34213
rect 71211 34155 71253 34164
rect 78027 34164 78028 34204
rect 78068 34164 78069 34204
rect 78027 34155 78069 34164
rect 63531 34110 63532 34150
rect 63572 34110 63573 34150
rect 63531 34101 63573 34110
rect 576 34040 79584 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 79584 34040
rect 576 33976 79584 34000
rect 52011 33872 52053 33881
rect 52011 33832 52012 33872
rect 52052 33832 52053 33872
rect 52011 33823 52053 33832
rect 55467 33876 55509 33885
rect 55467 33836 55468 33876
rect 55508 33836 55509 33876
rect 55467 33827 55509 33836
rect 58051 33872 58109 33873
rect 58051 33832 58060 33872
rect 58100 33832 58109 33872
rect 58051 33831 58109 33832
rect 59299 33872 59357 33873
rect 59299 33832 59308 33872
rect 59348 33832 59357 33872
rect 59299 33831 59357 33832
rect 59979 33872 60021 33881
rect 59979 33832 59980 33872
rect 60020 33832 60021 33872
rect 59979 33823 60021 33832
rect 61995 33872 62037 33881
rect 61995 33832 61996 33872
rect 62036 33832 62037 33872
rect 61995 33823 62037 33832
rect 63531 33872 63573 33881
rect 63531 33832 63532 33872
rect 63572 33832 63573 33872
rect 63531 33823 63573 33832
rect 64003 33872 64061 33873
rect 64003 33832 64012 33872
rect 64052 33832 64061 33872
rect 64003 33831 64061 33832
rect 64483 33872 64541 33873
rect 64483 33832 64492 33872
rect 64532 33832 64541 33872
rect 64483 33831 64541 33832
rect 67363 33872 67421 33873
rect 67363 33832 67372 33872
rect 67412 33832 67421 33872
rect 67363 33831 67421 33832
rect 70147 33872 70205 33873
rect 70147 33832 70156 33872
rect 70196 33832 70205 33872
rect 70147 33831 70205 33832
rect 71779 33872 71837 33873
rect 71779 33832 71788 33872
rect 71828 33832 71837 33872
rect 71779 33831 71837 33832
rect 72651 33872 72693 33881
rect 72651 33832 72652 33872
rect 72692 33832 72693 33872
rect 72651 33823 72693 33832
rect 76867 33872 76925 33873
rect 76867 33832 76876 33872
rect 76916 33832 76925 33872
rect 76867 33831 76925 33832
rect 51723 33788 51765 33797
rect 51723 33748 51724 33788
rect 51764 33748 51765 33788
rect 51723 33739 51765 33748
rect 50467 33704 50525 33705
rect 50467 33664 50476 33704
rect 50516 33664 50525 33704
rect 50467 33663 50525 33664
rect 51331 33704 51389 33705
rect 51331 33664 51340 33704
rect 51380 33664 51389 33704
rect 51331 33663 51389 33664
rect 51907 33704 51965 33705
rect 51907 33664 51916 33704
rect 51956 33664 51965 33704
rect 51907 33663 51965 33664
rect 53443 33704 53501 33705
rect 53443 33664 53452 33704
rect 53492 33664 53501 33704
rect 53443 33663 53501 33664
rect 54307 33704 54365 33705
rect 54307 33664 54316 33704
rect 54356 33664 54365 33704
rect 54307 33663 54365 33664
rect 54699 33704 54741 33713
rect 54699 33664 54700 33704
rect 54740 33664 54741 33704
rect 54699 33655 54741 33664
rect 55275 33704 55317 33713
rect 55275 33664 55276 33704
rect 55316 33664 55317 33704
rect 55275 33655 55317 33664
rect 55363 33704 55421 33705
rect 55363 33664 55372 33704
rect 55412 33664 55421 33704
rect 55363 33663 55421 33664
rect 55659 33704 55701 33713
rect 55659 33664 55660 33704
rect 55700 33664 55701 33704
rect 55659 33655 55701 33664
rect 56035 33704 56093 33705
rect 56035 33664 56044 33704
rect 56084 33664 56093 33704
rect 56035 33663 56093 33664
rect 56899 33704 56957 33705
rect 56899 33664 56908 33704
rect 56948 33664 56957 33704
rect 56899 33663 56957 33664
rect 59403 33704 59445 33713
rect 59403 33664 59404 33704
rect 59444 33664 59445 33704
rect 59403 33655 59445 33664
rect 59499 33704 59541 33713
rect 59499 33664 59500 33704
rect 59540 33664 59541 33704
rect 59499 33655 59541 33664
rect 59595 33704 59637 33713
rect 59595 33664 59596 33704
rect 59636 33664 59637 33704
rect 59595 33655 59637 33664
rect 59875 33704 59933 33705
rect 59875 33664 59884 33704
rect 59924 33664 59933 33704
rect 59875 33663 59933 33664
rect 63619 33704 63677 33705
rect 63619 33664 63628 33704
rect 63668 33664 63677 33704
rect 63619 33663 63677 33664
rect 64107 33704 64149 33713
rect 64107 33664 64108 33704
rect 64148 33664 64149 33704
rect 64107 33655 64149 33664
rect 64203 33704 64245 33713
rect 64203 33664 64204 33704
rect 64244 33664 64245 33704
rect 64203 33655 64245 33664
rect 64299 33704 64341 33713
rect 64299 33664 64300 33704
rect 64340 33664 64341 33704
rect 64299 33655 64341 33664
rect 64587 33704 64629 33713
rect 64587 33664 64588 33704
rect 64628 33664 64629 33704
rect 64587 33655 64629 33664
rect 64683 33704 64725 33713
rect 64683 33664 64684 33704
rect 64724 33664 64725 33704
rect 64683 33655 64725 33664
rect 64779 33704 64821 33713
rect 64779 33664 64780 33704
rect 64820 33664 64821 33704
rect 64779 33655 64821 33664
rect 66795 33704 66837 33713
rect 66795 33664 66796 33704
rect 66836 33664 66837 33704
rect 66795 33655 66837 33664
rect 66891 33704 66933 33713
rect 66891 33664 66892 33704
rect 66932 33664 66933 33704
rect 66891 33655 66933 33664
rect 66987 33704 67029 33713
rect 66987 33664 66988 33704
rect 67028 33664 67029 33704
rect 66987 33655 67029 33664
rect 67083 33704 67125 33713
rect 67083 33664 67084 33704
rect 67124 33664 67125 33704
rect 67083 33655 67125 33664
rect 67275 33704 67317 33713
rect 67275 33664 67276 33704
rect 67316 33664 67317 33704
rect 67275 33655 67317 33664
rect 67467 33704 67509 33713
rect 67467 33664 67468 33704
rect 67508 33664 67509 33704
rect 67467 33655 67509 33664
rect 67555 33704 67613 33705
rect 67555 33664 67564 33704
rect 67604 33664 67613 33704
rect 67555 33663 67613 33664
rect 67755 33704 67797 33713
rect 67755 33664 67756 33704
rect 67796 33664 67797 33704
rect 67755 33655 67797 33664
rect 68131 33704 68189 33705
rect 68131 33664 68140 33704
rect 68180 33664 68189 33704
rect 68131 33663 68189 33664
rect 68995 33704 69053 33705
rect 68995 33664 69004 33704
rect 69044 33664 69053 33704
rect 68995 33663 69053 33664
rect 71299 33704 71357 33705
rect 71299 33664 71308 33704
rect 71348 33664 71357 33704
rect 71299 33663 71357 33664
rect 71403 33704 71445 33713
rect 71403 33664 71404 33704
rect 71444 33664 71445 33704
rect 71403 33655 71445 33664
rect 71595 33704 71637 33713
rect 71595 33664 71596 33704
rect 71636 33664 71637 33704
rect 71595 33655 71637 33664
rect 71883 33704 71925 33713
rect 71883 33664 71884 33704
rect 71924 33664 71925 33704
rect 71883 33655 71925 33664
rect 71979 33704 72021 33713
rect 71979 33664 71980 33704
rect 72020 33664 72021 33704
rect 71979 33655 72021 33664
rect 72075 33704 72117 33713
rect 72075 33664 72076 33704
rect 72116 33664 72117 33704
rect 72075 33655 72117 33664
rect 72547 33704 72605 33705
rect 72547 33664 72556 33704
rect 72596 33664 72605 33704
rect 72547 33663 72605 33664
rect 74755 33704 74813 33705
rect 74755 33664 74764 33704
rect 74804 33664 74813 33704
rect 74755 33663 74813 33664
rect 76291 33704 76349 33705
rect 76291 33664 76300 33704
rect 76340 33664 76349 33704
rect 76291 33663 76349 33664
rect 76395 33704 76437 33713
rect 76395 33664 76396 33704
rect 76436 33664 76437 33704
rect 76395 33655 76437 33664
rect 76587 33704 76629 33713
rect 76587 33664 76588 33704
rect 76628 33664 76629 33704
rect 76587 33655 76629 33664
rect 76683 33704 76725 33713
rect 76683 33664 76684 33704
rect 76724 33664 76725 33704
rect 76683 33655 76725 33664
rect 76779 33704 76821 33713
rect 76779 33664 76780 33704
rect 76820 33664 76821 33704
rect 76779 33655 76821 33664
rect 77059 33704 77117 33705
rect 77059 33664 77068 33704
rect 77108 33664 77117 33704
rect 77059 33663 77117 33664
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77451 33655 77493 33664
rect 77643 33704 77685 33713
rect 77643 33664 77644 33704
rect 77684 33664 77685 33704
rect 77643 33655 77685 33664
rect 77835 33704 77877 33713
rect 77835 33664 77836 33704
rect 77876 33664 77877 33704
rect 77835 33655 77877 33664
rect 77923 33704 77981 33705
rect 77923 33664 77932 33704
rect 77972 33664 77981 33704
rect 77923 33663 77981 33664
rect 78211 33704 78269 33705
rect 78211 33664 78220 33704
rect 78260 33664 78269 33704
rect 78211 33663 78269 33664
rect 61795 33620 61853 33621
rect 61795 33580 61804 33620
rect 61844 33580 61853 33620
rect 61795 33579 61853 33580
rect 77163 33620 77205 33629
rect 77163 33580 77164 33620
rect 77204 33580 77205 33620
rect 77163 33571 77205 33580
rect 77355 33620 77397 33629
rect 77355 33580 77356 33620
rect 77396 33580 77397 33620
rect 77355 33571 77397 33580
rect 77259 33536 77301 33545
rect 77259 33496 77260 33536
rect 77300 33496 77301 33536
rect 77259 33487 77301 33496
rect 77643 33536 77685 33545
rect 77643 33496 77644 33536
rect 77684 33496 77685 33536
rect 77643 33487 77685 33496
rect 49315 33452 49373 33453
rect 49315 33412 49324 33452
rect 49364 33412 49373 33452
rect 49315 33411 49373 33412
rect 52011 33452 52053 33461
rect 52011 33412 52012 33452
rect 52052 33412 52053 33452
rect 52011 33403 52053 33412
rect 52291 33452 52349 33453
rect 52291 33412 52300 33452
rect 52340 33412 52349 33452
rect 52291 33411 52349 33412
rect 54987 33452 55029 33461
rect 54987 33412 54988 33452
rect 55028 33412 55029 33452
rect 54987 33403 55029 33412
rect 58051 33452 58109 33453
rect 58051 33412 58060 33452
rect 58100 33412 58109 33452
rect 58051 33411 58109 33412
rect 59979 33452 60021 33461
rect 59979 33412 59980 33452
rect 60020 33412 60021 33452
rect 59979 33403 60021 33412
rect 61995 33452 62037 33461
rect 61995 33412 61996 33452
rect 62036 33412 62037 33452
rect 61995 33403 62037 33412
rect 71595 33452 71637 33461
rect 71595 33412 71596 33452
rect 71636 33412 71637 33452
rect 71595 33403 71637 33412
rect 72651 33452 72693 33461
rect 72651 33412 72652 33452
rect 72692 33412 72693 33452
rect 72651 33403 72693 33412
rect 74859 33452 74901 33461
rect 74859 33412 74860 33452
rect 74900 33412 74901 33452
rect 74859 33403 74901 33412
rect 78123 33452 78165 33461
rect 78123 33412 78124 33452
rect 78164 33412 78165 33452
rect 78123 33403 78165 33412
rect 576 33284 79584 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 75112 33284
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75480 33244 79584 33284
rect 576 33220 79584 33244
rect 50955 33116 50997 33125
rect 50955 33076 50956 33116
rect 50996 33076 50997 33116
rect 50955 33067 50997 33076
rect 52107 33116 52149 33125
rect 52107 33076 52108 33116
rect 52148 33076 52149 33116
rect 52107 33067 52149 33076
rect 53835 33116 53877 33125
rect 53835 33076 53836 33116
rect 53876 33076 53877 33116
rect 53835 33067 53877 33076
rect 67843 33116 67901 33117
rect 67843 33076 67852 33116
rect 67892 33076 67901 33116
rect 67843 33075 67901 33076
rect 78787 33116 78845 33117
rect 78787 33076 78796 33116
rect 78836 33076 78845 33116
rect 78787 33075 78845 33076
rect 51915 33032 51957 33041
rect 51915 32992 51916 33032
rect 51956 32992 51957 33032
rect 51915 32983 51957 32992
rect 55275 33032 55317 33041
rect 55275 32992 55276 33032
rect 55316 32992 55317 33032
rect 55275 32983 55317 32992
rect 55851 33032 55893 33041
rect 55851 32992 55852 33032
rect 55892 32992 55893 33032
rect 55851 32983 55893 32992
rect 63531 33032 63573 33041
rect 63531 32992 63532 33032
rect 63572 32992 63573 33032
rect 63531 32983 63573 32992
rect 72843 33032 72885 33041
rect 72843 32992 72844 33032
rect 72884 32992 72885 33032
rect 72843 32983 72885 32992
rect 49987 32948 50045 32949
rect 49987 32908 49996 32948
rect 50036 32908 50045 32948
rect 49987 32907 50045 32908
rect 55179 32948 55221 32957
rect 55179 32908 55180 32948
rect 55220 32908 55221 32948
rect 55179 32899 55221 32908
rect 55371 32948 55413 32957
rect 55371 32908 55372 32948
rect 55412 32908 55413 32948
rect 55371 32899 55413 32908
rect 63811 32948 63869 32949
rect 63811 32908 63820 32948
rect 63860 32908 63869 32948
rect 63811 32907 63869 32908
rect 50467 32864 50525 32865
rect 50467 32824 50476 32864
rect 50516 32824 50525 32864
rect 50467 32823 50525 32824
rect 50571 32864 50613 32873
rect 50571 32824 50572 32864
rect 50612 32824 50613 32864
rect 50571 32815 50613 32824
rect 50763 32864 50805 32873
rect 50763 32824 50764 32864
rect 50804 32824 50805 32864
rect 50763 32815 50805 32824
rect 51243 32864 51285 32873
rect 51243 32824 51244 32864
rect 51284 32824 51285 32864
rect 51243 32815 51285 32824
rect 51331 32864 51389 32865
rect 51331 32824 51340 32864
rect 51380 32824 51389 32864
rect 51331 32823 51389 32824
rect 52579 32864 52637 32865
rect 52579 32824 52588 32864
rect 52628 32824 52637 32864
rect 52579 32823 52637 32824
rect 52875 32864 52917 32873
rect 52875 32824 52876 32864
rect 52916 32824 52917 32864
rect 52875 32815 52917 32824
rect 52971 32864 53013 32873
rect 52971 32824 52972 32864
rect 53012 32824 53013 32864
rect 52971 32815 53013 32824
rect 53067 32864 53109 32873
rect 53067 32824 53068 32864
rect 53108 32824 53109 32864
rect 53067 32815 53109 32824
rect 53163 32864 53205 32873
rect 53163 32824 53164 32864
rect 53204 32824 53205 32864
rect 53163 32815 53205 32824
rect 53355 32864 53397 32873
rect 53355 32824 53356 32864
rect 53396 32824 53397 32864
rect 53355 32815 53397 32824
rect 53451 32864 53493 32873
rect 53451 32824 53452 32864
rect 53492 32824 53493 32864
rect 53451 32815 53493 32824
rect 53547 32864 53589 32873
rect 53547 32824 53548 32864
rect 53588 32824 53589 32864
rect 53547 32815 53589 32824
rect 53643 32864 53685 32873
rect 53643 32824 53644 32864
rect 53684 32824 53685 32864
rect 53643 32815 53685 32824
rect 53835 32864 53877 32873
rect 53835 32824 53836 32864
rect 53876 32824 53877 32864
rect 53835 32815 53877 32824
rect 54027 32864 54069 32873
rect 54027 32824 54028 32864
rect 54068 32824 54069 32864
rect 54027 32815 54069 32824
rect 54115 32864 54173 32865
rect 54115 32824 54124 32864
rect 54164 32824 54173 32864
rect 54115 32823 54173 32824
rect 54603 32864 54645 32873
rect 54603 32824 54604 32864
rect 54644 32824 54645 32864
rect 54603 32815 54645 32824
rect 54699 32864 54741 32873
rect 54699 32824 54700 32864
rect 54740 32824 54741 32864
rect 54699 32815 54741 32824
rect 54795 32864 54837 32873
rect 54795 32824 54796 32864
rect 54836 32824 54837 32864
rect 54795 32815 54837 32824
rect 54891 32864 54933 32873
rect 54891 32824 54892 32864
rect 54932 32824 54933 32864
rect 54891 32815 54933 32824
rect 55075 32864 55133 32865
rect 55075 32824 55084 32864
rect 55124 32824 55133 32864
rect 55075 32823 55133 32824
rect 55467 32864 55509 32873
rect 55467 32824 55468 32864
rect 55508 32824 55509 32864
rect 56043 32864 56085 32873
rect 55467 32815 55509 32824
rect 55851 32822 55893 32831
rect 55851 32782 55852 32822
rect 55892 32782 55893 32822
rect 56043 32824 56044 32864
rect 56084 32824 56085 32864
rect 56043 32815 56085 32824
rect 56131 32864 56189 32865
rect 56131 32824 56140 32864
rect 56180 32824 56189 32864
rect 56131 32823 56189 32824
rect 61315 32864 61373 32865
rect 61315 32824 61324 32864
rect 61364 32824 61373 32864
rect 61315 32823 61373 32824
rect 62179 32864 62237 32865
rect 62179 32824 62188 32864
rect 62228 32824 62237 32864
rect 62179 32823 62237 32824
rect 62755 32864 62813 32865
rect 62755 32824 62764 32864
rect 62804 32824 62813 32864
rect 62755 32823 62813 32824
rect 63139 32864 63197 32865
rect 63139 32824 63148 32864
rect 63188 32824 63197 32864
rect 63139 32823 63197 32824
rect 63243 32864 63285 32873
rect 63243 32824 63244 32864
rect 63284 32824 63285 32864
rect 63243 32815 63285 32824
rect 65827 32864 65885 32865
rect 65827 32824 65836 32864
rect 65876 32824 65885 32864
rect 65827 32823 65885 32824
rect 66691 32864 66749 32865
rect 66691 32824 66700 32864
rect 66740 32824 66749 32864
rect 66691 32823 66749 32824
rect 68035 32864 68093 32865
rect 68035 32824 68044 32864
rect 68084 32824 68093 32864
rect 68035 32823 68093 32824
rect 70147 32864 70205 32865
rect 70147 32824 70156 32864
rect 70196 32824 70205 32864
rect 70147 32823 70205 32824
rect 71011 32864 71069 32865
rect 71011 32824 71020 32864
rect 71060 32824 71069 32864
rect 71011 32823 71069 32824
rect 72451 32864 72509 32865
rect 72451 32824 72460 32864
rect 72500 32824 72509 32864
rect 72451 32823 72509 32824
rect 72555 32864 72597 32873
rect 72555 32824 72556 32864
rect 72596 32824 72597 32864
rect 72555 32815 72597 32824
rect 76771 32864 76829 32865
rect 76771 32824 76780 32864
rect 76820 32824 76829 32864
rect 76771 32823 76829 32824
rect 77635 32864 77693 32865
rect 77635 32824 77644 32864
rect 77684 32824 77693 32864
rect 77635 32823 77693 32824
rect 55851 32773 55893 32782
rect 62571 32780 62613 32789
rect 62571 32740 62572 32780
rect 62612 32740 62613 32780
rect 62571 32731 62613 32740
rect 65451 32780 65493 32789
rect 65451 32740 65452 32780
rect 65492 32740 65493 32780
rect 65451 32731 65493 32740
rect 69771 32780 69813 32789
rect 69771 32740 69772 32780
rect 69812 32740 69813 32780
rect 69771 32731 69813 32740
rect 76395 32780 76437 32789
rect 76395 32740 76396 32780
rect 76436 32740 76437 32780
rect 76395 32731 76437 32740
rect 49803 32696 49845 32705
rect 49803 32656 49804 32696
rect 49844 32656 49845 32696
rect 49803 32647 49845 32656
rect 50659 32696 50717 32697
rect 50659 32656 50668 32696
rect 50708 32656 50717 32696
rect 50659 32655 50717 32656
rect 51435 32692 51477 32701
rect 51435 32652 51436 32692
rect 51476 32652 51477 32692
rect 60163 32696 60221 32697
rect 60163 32656 60172 32696
rect 60212 32656 60221 32696
rect 60163 32655 60221 32656
rect 62859 32696 62901 32705
rect 62859 32656 62860 32696
rect 62900 32656 62901 32696
rect 51435 32643 51477 32652
rect 62859 32647 62901 32656
rect 63051 32692 63093 32701
rect 63051 32652 63052 32692
rect 63092 32652 63093 32692
rect 63051 32643 63093 32652
rect 64011 32696 64053 32705
rect 64011 32656 64012 32696
rect 64052 32656 64053 32696
rect 64011 32647 64053 32656
rect 68139 32696 68181 32705
rect 68139 32656 68140 32696
rect 68180 32656 68181 32696
rect 68139 32647 68181 32656
rect 72163 32696 72221 32697
rect 72163 32656 72172 32696
rect 72212 32656 72221 32696
rect 72163 32655 72221 32656
rect 72363 32638 72405 32647
rect 72363 32598 72364 32638
rect 72404 32598 72405 32638
rect 72363 32589 72405 32598
rect 576 32528 79584 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 76352 32528
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76720 32488 79584 32528
rect 576 32464 79584 32488
rect 67659 32418 67701 32427
rect 67659 32378 67660 32418
rect 67700 32378 67701 32418
rect 67659 32369 67701 32378
rect 76779 32418 76821 32427
rect 76779 32378 76780 32418
rect 76820 32378 76821 32418
rect 76779 32369 76821 32378
rect 68427 32360 68469 32369
rect 68427 32320 68428 32360
rect 68468 32320 68469 32360
rect 68427 32311 68469 32320
rect 68811 32360 68853 32369
rect 68811 32320 68812 32360
rect 68852 32320 68853 32360
rect 68811 32311 68853 32320
rect 72651 32360 72693 32369
rect 72651 32320 72652 32360
rect 72692 32320 72693 32360
rect 72651 32311 72693 32320
rect 56907 32276 56949 32285
rect 56907 32236 56908 32276
rect 56948 32236 56949 32276
rect 56907 32227 56949 32236
rect 50571 32192 50613 32201
rect 50571 32152 50572 32192
rect 50612 32152 50613 32192
rect 50571 32143 50613 32152
rect 50947 32192 51005 32193
rect 50947 32152 50956 32192
rect 50996 32152 51005 32192
rect 50947 32151 51005 32152
rect 51811 32192 51869 32193
rect 51811 32152 51820 32192
rect 51860 32152 51869 32192
rect 51811 32151 51869 32152
rect 53355 32192 53397 32201
rect 53355 32152 53356 32192
rect 53396 32152 53397 32192
rect 53355 32143 53397 32152
rect 55651 32192 55709 32193
rect 55651 32152 55660 32192
rect 55700 32152 55709 32192
rect 55651 32151 55709 32152
rect 56515 32192 56573 32193
rect 56515 32152 56524 32192
rect 56564 32152 56573 32192
rect 56515 32151 56573 32152
rect 57187 32192 57245 32193
rect 57187 32152 57196 32192
rect 57236 32152 57245 32192
rect 57187 32151 57245 32152
rect 57579 32192 57621 32201
rect 57579 32152 57580 32192
rect 57620 32152 57621 32192
rect 57579 32143 57621 32152
rect 58915 32192 58973 32193
rect 58915 32152 58924 32192
rect 58964 32152 58973 32192
rect 58915 32151 58973 32152
rect 59779 32192 59837 32193
rect 59779 32152 59788 32192
rect 59828 32152 59837 32192
rect 59779 32151 59837 32152
rect 60171 32192 60213 32201
rect 60171 32152 60172 32192
rect 60212 32152 60213 32192
rect 60171 32143 60213 32152
rect 60355 32192 60413 32193
rect 60355 32152 60364 32192
rect 60404 32152 60413 32192
rect 60355 32151 60413 32152
rect 60739 32192 60797 32193
rect 60739 32152 60748 32192
rect 60788 32152 60797 32192
rect 60739 32151 60797 32152
rect 61131 32192 61173 32201
rect 61131 32152 61132 32192
rect 61172 32152 61173 32192
rect 61131 32143 61173 32152
rect 61515 32192 61557 32201
rect 61515 32152 61516 32192
rect 61556 32152 61557 32192
rect 61515 32143 61557 32152
rect 61707 32192 61749 32201
rect 61707 32152 61708 32192
rect 61748 32152 61749 32192
rect 61707 32143 61749 32152
rect 61795 32192 61853 32193
rect 61795 32152 61804 32192
rect 61844 32152 61853 32192
rect 61795 32151 61853 32152
rect 62763 32192 62805 32201
rect 62763 32152 62764 32192
rect 62804 32152 62805 32192
rect 62763 32143 62805 32152
rect 63139 32192 63197 32193
rect 63139 32152 63148 32192
rect 63188 32152 63197 32192
rect 63139 32151 63197 32152
rect 63339 32192 63381 32201
rect 63339 32152 63340 32192
rect 63380 32152 63381 32192
rect 63339 32143 63381 32152
rect 63715 32192 63773 32193
rect 63715 32152 63724 32192
rect 63764 32152 63773 32192
rect 63715 32151 63773 32152
rect 64579 32192 64637 32193
rect 64579 32152 64588 32192
rect 64628 32152 64637 32192
rect 64579 32151 64637 32152
rect 66411 32192 66453 32201
rect 66411 32152 66412 32192
rect 66452 32152 66453 32192
rect 66411 32143 66453 32152
rect 66787 32192 66845 32193
rect 66787 32152 66796 32192
rect 66836 32152 66845 32192
rect 66787 32151 66845 32152
rect 67467 32192 67509 32201
rect 67467 32152 67468 32192
rect 67508 32152 67509 32192
rect 67467 32143 67509 32152
rect 67555 32192 67613 32193
rect 67555 32152 67564 32192
rect 67604 32152 67613 32192
rect 67555 32151 67613 32152
rect 71499 32192 71541 32201
rect 71499 32152 71500 32192
rect 71540 32152 71541 32192
rect 71499 32143 71541 32152
rect 71875 32192 71933 32193
rect 71875 32152 71884 32192
rect 71924 32152 71933 32192
rect 71875 32151 71933 32152
rect 72075 32192 72117 32201
rect 72075 32152 72076 32192
rect 72116 32152 72117 32192
rect 72075 32143 72117 32152
rect 72267 32192 72309 32201
rect 72267 32152 72268 32192
rect 72308 32152 72309 32192
rect 72267 32143 72309 32152
rect 72355 32192 72413 32193
rect 72355 32152 72364 32192
rect 72404 32152 72413 32192
rect 72355 32151 72413 32152
rect 72547 32192 72605 32193
rect 72547 32152 72556 32192
rect 72596 32152 72605 32192
rect 72547 32151 72605 32152
rect 72843 32192 72885 32201
rect 72843 32152 72844 32192
rect 72884 32152 72885 32192
rect 72843 32143 72885 32152
rect 73219 32192 73277 32193
rect 73219 32152 73228 32192
rect 73268 32152 73277 32192
rect 73219 32151 73277 32152
rect 74083 32192 74141 32193
rect 74083 32152 74092 32192
rect 74132 32152 74141 32192
rect 74083 32151 74141 32152
rect 76587 32192 76629 32201
rect 76587 32152 76588 32192
rect 76628 32152 76629 32192
rect 76587 32143 76629 32152
rect 76675 32192 76733 32193
rect 76675 32152 76684 32192
rect 76724 32152 76733 32192
rect 76675 32151 76733 32152
rect 76971 32192 77013 32201
rect 76971 32152 76972 32192
rect 77012 32152 77013 32192
rect 76971 32143 77013 32152
rect 77347 32192 77405 32193
rect 77347 32152 77356 32192
rect 77396 32152 77405 32192
rect 77347 32151 77405 32152
rect 78211 32192 78269 32193
rect 78211 32152 78220 32192
rect 78260 32152 78269 32192
rect 78211 32151 78269 32152
rect 57291 32108 57333 32117
rect 57291 32068 57292 32108
rect 57332 32068 57333 32108
rect 57291 32059 57333 32068
rect 57483 32108 57525 32117
rect 57483 32068 57484 32108
rect 57524 32068 57525 32108
rect 57483 32059 57525 32068
rect 60843 32108 60885 32117
rect 60843 32068 60844 32108
rect 60884 32068 60885 32108
rect 60843 32059 60885 32068
rect 61035 32108 61077 32117
rect 61035 32068 61036 32108
rect 61076 32068 61077 32108
rect 61035 32059 61077 32068
rect 62859 32108 62901 32117
rect 62859 32068 62860 32108
rect 62900 32068 62901 32108
rect 62859 32059 62901 32068
rect 63051 32108 63093 32117
rect 63051 32068 63052 32108
rect 63092 32068 63093 32108
rect 63051 32059 63093 32068
rect 66507 32108 66549 32117
rect 66507 32068 66508 32108
rect 66548 32068 66549 32108
rect 66507 32059 66549 32068
rect 66699 32108 66741 32117
rect 66699 32068 66700 32108
rect 66740 32068 66741 32108
rect 66699 32059 66741 32068
rect 68611 32108 68669 32109
rect 68611 32068 68620 32108
rect 68660 32068 68669 32108
rect 68611 32067 68669 32068
rect 68995 32108 69053 32109
rect 68995 32068 69004 32108
rect 69044 32068 69053 32108
rect 68995 32067 69053 32068
rect 71595 32108 71637 32117
rect 71595 32068 71596 32108
rect 71636 32068 71637 32108
rect 71595 32059 71637 32068
rect 71787 32108 71829 32117
rect 71787 32068 71788 32108
rect 71828 32068 71829 32108
rect 71787 32059 71829 32068
rect 57387 32024 57429 32033
rect 57387 31984 57388 32024
rect 57428 31984 57429 32024
rect 57387 31975 57429 31984
rect 60939 32024 60981 32033
rect 60939 31984 60940 32024
rect 60980 31984 60981 32024
rect 60939 31975 60981 31984
rect 61515 32024 61557 32033
rect 61515 31984 61516 32024
rect 61556 31984 61557 32024
rect 61515 31975 61557 31984
rect 62955 32024 62997 32033
rect 62955 31984 62956 32024
rect 62996 31984 62997 32024
rect 62955 31975 62997 31984
rect 66603 32024 66645 32033
rect 66603 31984 66604 32024
rect 66644 31984 66645 32024
rect 66603 31975 66645 31984
rect 71691 32024 71733 32033
rect 71691 31984 71692 32024
rect 71732 31984 71733 32024
rect 71691 31975 71733 31984
rect 52963 31940 53021 31941
rect 52963 31900 52972 31940
rect 53012 31900 53021 31940
rect 52963 31899 53021 31900
rect 54499 31940 54557 31941
rect 54499 31900 54508 31940
rect 54548 31900 54557 31940
rect 54499 31899 54557 31900
rect 57763 31940 57821 31941
rect 57763 31900 57772 31940
rect 57812 31900 57821 31940
rect 57763 31899 57821 31900
rect 60459 31940 60501 31949
rect 60459 31900 60460 31940
rect 60500 31900 60501 31940
rect 60459 31891 60501 31900
rect 65731 31940 65789 31941
rect 65731 31900 65740 31940
rect 65780 31900 65789 31940
rect 65731 31899 65789 31900
rect 67179 31940 67221 31949
rect 67179 31900 67180 31940
rect 67220 31900 67221 31940
rect 67179 31891 67221 31900
rect 68427 31940 68469 31949
rect 68427 31900 68428 31940
rect 68468 31900 68469 31940
rect 68427 31891 68469 31900
rect 72075 31940 72117 31949
rect 72075 31900 72076 31940
rect 72116 31900 72117 31940
rect 72075 31891 72117 31900
rect 75235 31940 75293 31941
rect 75235 31900 75244 31940
rect 75284 31900 75293 31940
rect 75235 31899 75293 31900
rect 76299 31940 76341 31949
rect 76299 31900 76300 31940
rect 76340 31900 76341 31940
rect 76299 31891 76341 31900
rect 79363 31940 79421 31941
rect 79363 31900 79372 31940
rect 79412 31900 79421 31940
rect 79363 31899 79421 31900
rect 576 31772 79584 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 75112 31772
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75480 31732 79584 31772
rect 576 31708 79584 31732
rect 50187 31604 50229 31613
rect 50187 31564 50188 31604
rect 50228 31564 50229 31604
rect 50187 31555 50229 31564
rect 51819 31604 51861 31613
rect 51819 31564 51820 31604
rect 51860 31564 51861 31604
rect 51819 31555 51861 31564
rect 54603 31604 54645 31613
rect 54603 31564 54604 31604
rect 54644 31564 54645 31604
rect 54603 31555 54645 31564
rect 57195 31604 57237 31613
rect 57195 31564 57196 31604
rect 57236 31564 57237 31604
rect 57195 31555 57237 31564
rect 57867 31604 57909 31613
rect 57867 31564 57868 31604
rect 57908 31564 57909 31604
rect 57867 31555 57909 31564
rect 58635 31604 58677 31613
rect 58635 31564 58636 31604
rect 58676 31564 58677 31604
rect 58635 31555 58677 31564
rect 66219 31604 66261 31613
rect 66219 31564 66220 31604
rect 66260 31564 66261 31604
rect 66219 31555 66261 31564
rect 71595 31604 71637 31613
rect 71595 31564 71596 31604
rect 71636 31564 71637 31604
rect 71595 31555 71637 31564
rect 50571 31520 50613 31529
rect 50571 31480 50572 31520
rect 50612 31480 50613 31520
rect 50571 31471 50613 31480
rect 50955 31520 50997 31529
rect 50955 31480 50956 31520
rect 50996 31480 50997 31520
rect 50955 31471 50997 31480
rect 52491 31520 52533 31529
rect 52491 31480 52492 31520
rect 52532 31480 52533 31520
rect 52491 31471 52533 31480
rect 60843 31520 60885 31529
rect 60843 31480 60844 31520
rect 60884 31480 60885 31520
rect 60843 31471 60885 31480
rect 70443 31520 70485 31529
rect 70443 31480 70444 31520
rect 70484 31480 70485 31520
rect 70443 31471 70485 31480
rect 76683 31520 76725 31529
rect 76683 31480 76684 31520
rect 76724 31480 76725 31520
rect 76683 31471 76725 31480
rect 77067 31520 77109 31529
rect 77067 31480 77068 31520
rect 77108 31480 77109 31520
rect 77067 31471 77109 31480
rect 49987 31436 50045 31437
rect 49987 31396 49996 31436
rect 50036 31396 50045 31436
rect 49987 31395 50045 31396
rect 50475 31436 50517 31445
rect 50475 31396 50476 31436
rect 50516 31396 50517 31436
rect 50475 31387 50517 31396
rect 50667 31436 50709 31445
rect 50667 31396 50668 31436
rect 50708 31396 50709 31436
rect 50667 31387 50709 31396
rect 52395 31436 52437 31445
rect 52395 31396 52396 31436
rect 52436 31396 52437 31436
rect 52395 31387 52437 31396
rect 52587 31436 52629 31445
rect 52587 31396 52588 31436
rect 52628 31396 52629 31436
rect 52587 31387 52629 31396
rect 71395 31436 71453 31437
rect 71395 31396 71404 31436
rect 71444 31396 71453 31436
rect 71395 31395 71453 31396
rect 73219 31436 73277 31437
rect 73219 31396 73228 31436
rect 73268 31396 73277 31436
rect 73219 31395 73277 31396
rect 76587 31436 76629 31445
rect 76587 31396 76588 31436
rect 76628 31396 76629 31436
rect 63331 31394 63389 31395
rect 51819 31363 51861 31372
rect 50371 31352 50429 31353
rect 50371 31312 50380 31352
rect 50420 31312 50429 31352
rect 50371 31311 50429 31312
rect 50763 31352 50805 31361
rect 50763 31312 50764 31352
rect 50804 31312 50805 31352
rect 50763 31303 50805 31312
rect 51243 31352 51285 31361
rect 51243 31312 51244 31352
rect 51284 31312 51285 31352
rect 51243 31303 51285 31312
rect 51331 31352 51389 31353
rect 51331 31312 51340 31352
rect 51380 31312 51389 31352
rect 51819 31323 51820 31363
rect 51860 31323 51861 31363
rect 51819 31314 51861 31323
rect 52011 31352 52053 31361
rect 51331 31311 51389 31312
rect 52011 31312 52012 31352
rect 52052 31312 52053 31352
rect 52011 31303 52053 31312
rect 52099 31352 52157 31353
rect 52099 31312 52108 31352
rect 52148 31312 52157 31352
rect 52099 31311 52157 31312
rect 52299 31352 52341 31361
rect 52299 31312 52300 31352
rect 52340 31312 52341 31352
rect 52299 31303 52341 31312
rect 52675 31352 52733 31353
rect 52675 31312 52684 31352
rect 52724 31312 52733 31352
rect 52675 31311 52733 31312
rect 52963 31352 53021 31353
rect 52963 31312 52972 31352
rect 53012 31312 53021 31352
rect 52963 31311 53021 31312
rect 55275 31352 55317 31361
rect 55275 31312 55276 31352
rect 55316 31312 55317 31352
rect 55275 31303 55317 31312
rect 55363 31352 55421 31353
rect 55363 31312 55372 31352
rect 55412 31312 55421 31352
rect 55363 31311 55421 31312
rect 57091 31352 57149 31353
rect 57091 31312 57100 31352
rect 57140 31312 57149 31352
rect 57091 31311 57149 31312
rect 57475 31352 57533 31353
rect 57475 31312 57484 31352
rect 57524 31312 57533 31352
rect 57475 31311 57533 31312
rect 57579 31352 57621 31361
rect 57579 31312 57580 31352
rect 57620 31312 57621 31352
rect 57579 31303 57621 31312
rect 58059 31352 58101 31361
rect 58059 31312 58060 31352
rect 58100 31312 58101 31352
rect 58059 31303 58101 31312
rect 58155 31352 58197 31361
rect 58155 31312 58156 31352
rect 58196 31312 58197 31352
rect 58155 31303 58197 31312
rect 58251 31352 58293 31361
rect 58251 31312 58252 31352
rect 58292 31312 58293 31352
rect 58251 31303 58293 31312
rect 58347 31352 58389 31361
rect 58347 31312 58348 31352
rect 58388 31312 58389 31352
rect 58347 31303 58389 31312
rect 58635 31352 58677 31361
rect 58635 31312 58636 31352
rect 58676 31312 58677 31352
rect 58635 31303 58677 31312
rect 58827 31352 58869 31361
rect 58827 31312 58828 31352
rect 58868 31312 58869 31352
rect 58827 31303 58869 31312
rect 58915 31352 58973 31353
rect 58915 31312 58924 31352
rect 58964 31312 58973 31352
rect 58915 31311 58973 31312
rect 59203 31352 59261 31353
rect 59203 31312 59212 31352
rect 59252 31312 59261 31352
rect 59203 31311 59261 31312
rect 61131 31352 61173 31361
rect 61131 31312 61132 31352
rect 61172 31312 61173 31352
rect 61131 31303 61173 31312
rect 61219 31352 61277 31353
rect 61219 31312 61228 31352
rect 61268 31312 61277 31352
rect 61219 31311 61277 31312
rect 61515 31352 61557 31361
rect 61515 31312 61516 31352
rect 61556 31312 61557 31352
rect 61515 31303 61557 31312
rect 61611 31352 61653 31361
rect 61611 31312 61612 31352
rect 61652 31312 61653 31352
rect 61611 31303 61653 31312
rect 61707 31352 61749 31361
rect 61707 31312 61708 31352
rect 61748 31312 61749 31352
rect 61707 31303 61749 31312
rect 61803 31352 61845 31361
rect 61803 31312 61804 31352
rect 61844 31312 61845 31352
rect 61803 31303 61845 31312
rect 63243 31352 63285 31361
rect 63331 31354 63340 31394
rect 63380 31354 63389 31394
rect 76587 31387 76629 31396
rect 76779 31436 76821 31445
rect 76779 31396 76780 31436
rect 76820 31396 76821 31436
rect 76779 31387 76821 31396
rect 63331 31353 63389 31354
rect 63243 31312 63244 31352
rect 63284 31312 63285 31352
rect 63243 31303 63285 31312
rect 63435 31352 63477 31361
rect 63435 31312 63436 31352
rect 63476 31312 63477 31352
rect 63435 31303 63477 31312
rect 63531 31352 63573 31361
rect 63531 31312 63532 31352
rect 63572 31312 63573 31352
rect 63531 31303 63573 31312
rect 63723 31352 63765 31361
rect 63723 31312 63724 31352
rect 63764 31312 63765 31352
rect 63723 31303 63765 31312
rect 63819 31352 63861 31361
rect 63819 31312 63820 31352
rect 63860 31312 63861 31352
rect 63819 31303 63861 31312
rect 63915 31352 63957 31361
rect 63915 31312 63916 31352
rect 63956 31312 63957 31352
rect 63915 31303 63957 31312
rect 64011 31352 64053 31361
rect 64011 31312 64012 31352
rect 64052 31312 64053 31352
rect 64011 31303 64053 31312
rect 66219 31352 66261 31361
rect 66219 31312 66220 31352
rect 66260 31312 66261 31352
rect 66219 31303 66261 31312
rect 66411 31352 66453 31361
rect 66411 31312 66412 31352
rect 66452 31312 66453 31352
rect 66411 31303 66453 31312
rect 66499 31352 66557 31353
rect 66499 31312 66508 31352
rect 66548 31312 66557 31352
rect 66499 31311 66557 31312
rect 67179 31352 67221 31361
rect 67179 31312 67180 31352
rect 67220 31312 67221 31352
rect 67179 31303 67221 31312
rect 67275 31352 67317 31361
rect 67275 31312 67276 31352
rect 67316 31312 67317 31352
rect 67275 31303 67317 31312
rect 67371 31352 67413 31361
rect 67371 31312 67372 31352
rect 67412 31312 67413 31352
rect 67371 31303 67413 31312
rect 67939 31352 67997 31353
rect 67939 31312 67948 31352
rect 67988 31312 67997 31352
rect 67939 31311 67997 31312
rect 68803 31352 68861 31353
rect 68803 31312 68812 31352
rect 68852 31312 68861 31352
rect 68803 31311 68861 31312
rect 71779 31352 71837 31353
rect 71779 31312 71788 31352
rect 71828 31312 71837 31352
rect 71779 31311 71837 31312
rect 72363 31352 72405 31361
rect 72363 31312 72364 31352
rect 72404 31312 72405 31352
rect 72363 31303 72405 31312
rect 72459 31352 72501 31361
rect 72459 31312 72460 31352
rect 72500 31312 72501 31352
rect 72459 31303 72501 31312
rect 72555 31352 72597 31361
rect 72555 31312 72556 31352
rect 72596 31312 72597 31352
rect 72555 31303 72597 31312
rect 72747 31352 72789 31361
rect 72747 31312 72748 31352
rect 72788 31312 72789 31352
rect 72747 31303 72789 31312
rect 72843 31352 72885 31361
rect 72843 31312 72844 31352
rect 72884 31312 72885 31352
rect 72843 31303 72885 31312
rect 72939 31352 72981 31361
rect 72939 31312 72940 31352
rect 72980 31312 72981 31352
rect 72939 31303 72981 31312
rect 73035 31352 73077 31361
rect 73035 31312 73036 31352
rect 73076 31312 73077 31352
rect 73035 31303 73077 31312
rect 73611 31352 73653 31361
rect 73611 31312 73612 31352
rect 73652 31312 73653 31352
rect 73611 31303 73653 31312
rect 73707 31352 73749 31361
rect 73707 31312 73708 31352
rect 73748 31312 73749 31352
rect 73899 31352 73941 31361
rect 73707 31303 73749 31312
rect 73803 31331 73845 31340
rect 73803 31291 73804 31331
rect 73844 31291 73845 31331
rect 73899 31312 73900 31352
rect 73940 31312 73941 31352
rect 73899 31303 73941 31312
rect 74467 31352 74525 31353
rect 74467 31312 74476 31352
rect 74516 31312 74525 31352
rect 74467 31311 74525 31312
rect 76011 31352 76053 31361
rect 76011 31312 76012 31352
rect 76052 31312 76053 31352
rect 76011 31303 76053 31312
rect 76107 31352 76149 31361
rect 76107 31312 76108 31352
rect 76148 31312 76149 31352
rect 76107 31303 76149 31312
rect 76203 31352 76245 31361
rect 76203 31312 76204 31352
rect 76244 31312 76245 31352
rect 76203 31303 76245 31312
rect 76483 31352 76541 31353
rect 76483 31312 76492 31352
rect 76532 31312 76541 31352
rect 76483 31311 76541 31312
rect 76875 31352 76917 31361
rect 76875 31312 76876 31352
rect 76916 31312 76917 31352
rect 76875 31303 76917 31312
rect 77067 31352 77109 31361
rect 77067 31312 77068 31352
rect 77108 31312 77109 31352
rect 77067 31303 77109 31312
rect 77259 31352 77301 31361
rect 77259 31312 77260 31352
rect 77300 31312 77301 31352
rect 77259 31303 77301 31312
rect 77347 31352 77405 31353
rect 77347 31312 77356 31352
rect 77396 31312 77405 31352
rect 77347 31311 77405 31312
rect 77547 31352 77589 31361
rect 77547 31312 77548 31352
rect 77588 31312 77589 31352
rect 77547 31303 77589 31312
rect 77643 31352 77685 31361
rect 77643 31312 77644 31352
rect 77684 31312 77685 31352
rect 77643 31303 77685 31312
rect 77739 31352 77781 31361
rect 77739 31312 77740 31352
rect 77780 31312 77781 31352
rect 77739 31303 77781 31312
rect 77835 31352 77877 31361
rect 77835 31312 77836 31352
rect 77876 31312 77877 31352
rect 77835 31303 77877 31312
rect 78115 31352 78173 31353
rect 78115 31312 78124 31352
rect 78164 31312 78173 31352
rect 78115 31311 78173 31312
rect 73803 31282 73845 31291
rect 67563 31268 67605 31277
rect 67563 31228 67564 31268
rect 67604 31228 67605 31268
rect 57763 31226 57821 31227
rect 57195 31184 57237 31193
rect 57195 31144 57196 31184
rect 57236 31144 57237 31184
rect 57195 31135 57237 31144
rect 57387 31180 57429 31189
rect 57763 31186 57772 31226
rect 57812 31186 57821 31226
rect 67563 31219 67605 31228
rect 57763 31185 57821 31186
rect 57387 31140 57388 31180
rect 57428 31140 57429 31180
rect 51435 31126 51477 31135
rect 57387 31131 57429 31140
rect 59115 31184 59157 31193
rect 59115 31144 59116 31184
rect 59156 31144 59157 31184
rect 59115 31135 59157 31144
rect 61323 31180 61365 31189
rect 61323 31140 61324 31180
rect 61364 31140 61365 31180
rect 67075 31184 67133 31185
rect 67075 31144 67084 31184
rect 67124 31144 67133 31184
rect 67075 31143 67133 31144
rect 69955 31184 70013 31185
rect 69955 31144 69964 31184
rect 70004 31144 70013 31184
rect 69955 31143 70013 31144
rect 71595 31184 71637 31193
rect 71595 31144 71596 31184
rect 71636 31144 71637 31184
rect 61323 31131 61365 31140
rect 71595 31135 71637 31144
rect 71883 31184 71925 31193
rect 71883 31144 71884 31184
rect 71924 31144 71925 31184
rect 71883 31135 71925 31144
rect 72259 31184 72317 31185
rect 72259 31144 72268 31184
rect 72308 31144 72317 31184
rect 72259 31143 72317 31144
rect 73419 31184 73461 31193
rect 73419 31144 73420 31184
rect 73460 31144 73461 31184
rect 73419 31135 73461 31144
rect 74379 31184 74421 31193
rect 74379 31144 74380 31184
rect 74420 31144 74421 31184
rect 74379 31135 74421 31144
rect 76291 31184 76349 31185
rect 76291 31144 76300 31184
rect 76340 31144 76349 31184
rect 76291 31143 76349 31144
rect 78027 31184 78069 31193
rect 78027 31144 78028 31184
rect 78068 31144 78069 31184
rect 78027 31135 78069 31144
rect 51435 31086 51436 31126
rect 51476 31086 51477 31126
rect 51435 31077 51477 31086
rect 576 31016 79584 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 76352 31016
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76720 30976 79584 31016
rect 576 30952 79584 30976
rect 56035 30848 56093 30849
rect 56035 30808 56044 30848
rect 56084 30808 56093 30848
rect 56035 30807 56093 30808
rect 56427 30848 56469 30857
rect 56427 30808 56428 30848
rect 56468 30808 56469 30848
rect 56427 30799 56469 30808
rect 57667 30848 57725 30849
rect 57667 30808 57676 30848
rect 57716 30808 57725 30848
rect 57667 30807 57725 30808
rect 60835 30848 60893 30849
rect 60835 30808 60844 30848
rect 60884 30808 60893 30848
rect 60835 30807 60893 30808
rect 66403 30848 66461 30849
rect 66403 30808 66412 30848
rect 66452 30808 66461 30848
rect 66403 30807 66461 30808
rect 68419 30848 68477 30849
rect 68419 30808 68428 30848
rect 68468 30808 68477 30848
rect 68419 30807 68477 30808
rect 69099 30848 69141 30857
rect 69099 30808 69100 30848
rect 69140 30808 69141 30848
rect 69099 30799 69141 30808
rect 74851 30848 74909 30849
rect 74851 30808 74860 30848
rect 74900 30808 74909 30848
rect 74851 30807 74909 30808
rect 77443 30848 77501 30849
rect 77443 30808 77452 30848
rect 77492 30808 77501 30848
rect 77443 30807 77501 30808
rect 53643 30764 53685 30773
rect 53643 30724 53644 30764
rect 53684 30724 53685 30764
rect 53643 30715 53685 30724
rect 57867 30764 57909 30773
rect 57867 30724 57868 30764
rect 57908 30724 57909 30764
rect 57867 30715 57909 30724
rect 61323 30764 61365 30773
rect 61323 30724 61324 30764
rect 61364 30724 61365 30764
rect 61323 30715 61365 30724
rect 72459 30764 72501 30773
rect 72459 30724 72460 30764
rect 72500 30724 72501 30764
rect 72459 30715 72501 30724
rect 48075 30680 48117 30689
rect 48075 30640 48076 30680
rect 48116 30640 48117 30680
rect 48075 30631 48117 30640
rect 48451 30680 48509 30681
rect 48451 30640 48460 30680
rect 48500 30640 48509 30680
rect 48451 30639 48509 30640
rect 50187 30680 50229 30689
rect 50187 30640 50188 30680
rect 50228 30640 50229 30680
rect 50187 30631 50229 30640
rect 50283 30680 50325 30689
rect 50283 30640 50284 30680
rect 50324 30640 50325 30680
rect 50283 30631 50325 30640
rect 50379 30680 50421 30689
rect 50379 30640 50380 30680
rect 50420 30640 50421 30680
rect 50379 30631 50421 30640
rect 50475 30680 50517 30689
rect 50475 30640 50476 30680
rect 50516 30640 50517 30680
rect 50475 30631 50517 30640
rect 50667 30680 50709 30689
rect 50667 30640 50668 30680
rect 50708 30640 50709 30680
rect 50667 30631 50709 30640
rect 51043 30680 51101 30681
rect 51043 30640 51052 30680
rect 51092 30640 51101 30680
rect 51043 30639 51101 30640
rect 51907 30680 51965 30681
rect 51907 30640 51916 30680
rect 51956 30640 51965 30680
rect 51907 30639 51965 30640
rect 54019 30680 54077 30681
rect 54019 30640 54028 30680
rect 54068 30640 54077 30680
rect 54019 30639 54077 30640
rect 54883 30680 54941 30681
rect 54883 30640 54892 30680
rect 54932 30640 54941 30680
rect 54883 30639 54941 30640
rect 57387 30680 57429 30689
rect 57387 30640 57388 30680
rect 57428 30640 57429 30680
rect 57387 30631 57429 30640
rect 57483 30680 57525 30689
rect 57483 30640 57484 30680
rect 57524 30640 57525 30680
rect 57483 30631 57525 30640
rect 57579 30680 57621 30689
rect 57579 30640 57580 30680
rect 57620 30640 57621 30680
rect 57579 30631 57621 30640
rect 58243 30680 58301 30681
rect 58243 30640 58252 30680
rect 58292 30640 58301 30680
rect 58243 30639 58301 30640
rect 59107 30680 59165 30681
rect 59107 30640 59116 30680
rect 59156 30640 59165 30680
rect 59107 30639 59165 30640
rect 60939 30680 60981 30689
rect 60939 30640 60940 30680
rect 60980 30640 60981 30680
rect 60939 30631 60981 30640
rect 61035 30680 61077 30689
rect 61035 30640 61036 30680
rect 61076 30640 61077 30680
rect 61035 30631 61077 30640
rect 61131 30680 61173 30689
rect 61131 30640 61132 30680
rect 61172 30640 61173 30680
rect 61131 30631 61173 30640
rect 61699 30680 61757 30681
rect 61699 30640 61708 30680
rect 61748 30640 61757 30680
rect 61699 30639 61757 30640
rect 62563 30680 62621 30681
rect 62563 30640 62572 30680
rect 62612 30640 62621 30680
rect 62563 30639 62621 30640
rect 64011 30680 64053 30689
rect 64011 30640 64012 30680
rect 64052 30640 64053 30680
rect 64011 30631 64053 30640
rect 64387 30680 64445 30681
rect 64387 30640 64396 30680
rect 64436 30640 64445 30680
rect 64387 30639 64445 30640
rect 65251 30680 65309 30681
rect 65251 30640 65260 30680
rect 65300 30640 65309 30680
rect 65251 30639 65309 30640
rect 66603 30680 66645 30689
rect 66603 30640 66604 30680
rect 66644 30640 66645 30680
rect 66603 30631 66645 30640
rect 66699 30680 66741 30689
rect 66699 30640 66700 30680
rect 66740 30640 66741 30680
rect 66699 30631 66741 30640
rect 66795 30680 66837 30689
rect 66795 30640 66796 30680
rect 66836 30640 66837 30680
rect 66795 30631 66837 30640
rect 66891 30680 66933 30689
rect 66891 30640 66892 30680
rect 66932 30640 66933 30680
rect 66891 30631 66933 30640
rect 67075 30680 67133 30681
rect 67075 30640 67084 30680
rect 67124 30640 67133 30680
rect 67075 30639 67133 30640
rect 68139 30680 68181 30689
rect 68139 30640 68140 30680
rect 68180 30640 68181 30680
rect 68139 30631 68181 30640
rect 68235 30680 68277 30689
rect 68235 30640 68236 30680
rect 68276 30640 68277 30680
rect 68235 30631 68277 30640
rect 68331 30680 68373 30689
rect 68331 30640 68332 30680
rect 68372 30640 68373 30680
rect 68331 30631 68373 30640
rect 68995 30680 69053 30681
rect 68995 30640 69004 30680
rect 69044 30640 69053 30680
rect 68995 30639 69053 30640
rect 70435 30680 70493 30681
rect 70435 30640 70444 30680
rect 70484 30640 70493 30680
rect 70435 30639 70493 30640
rect 71299 30680 71357 30681
rect 71299 30640 71308 30680
rect 71348 30640 71357 30680
rect 71299 30639 71357 30640
rect 71691 30680 71733 30689
rect 71691 30640 71692 30680
rect 71732 30640 71733 30680
rect 71691 30631 71733 30640
rect 71875 30680 71933 30681
rect 71875 30640 71884 30680
rect 71924 30640 71933 30680
rect 71875 30639 71933 30640
rect 72267 30680 72309 30689
rect 72267 30640 72268 30680
rect 72308 30640 72309 30680
rect 72267 30631 72309 30640
rect 72835 30680 72893 30681
rect 72835 30640 72844 30680
rect 72884 30640 72893 30680
rect 72835 30639 72893 30640
rect 73699 30680 73757 30681
rect 73699 30640 73708 30680
rect 73748 30640 73757 30680
rect 73699 30639 73757 30640
rect 75051 30680 75093 30689
rect 75051 30640 75052 30680
rect 75092 30640 75093 30680
rect 75051 30631 75093 30640
rect 75427 30680 75485 30681
rect 75427 30640 75436 30680
rect 75476 30640 75485 30680
rect 75427 30639 75485 30640
rect 76291 30680 76349 30681
rect 76291 30640 76300 30680
rect 76340 30640 76349 30680
rect 76291 30639 76349 30640
rect 77635 30680 77693 30681
rect 77635 30640 77644 30680
rect 77684 30640 77693 30680
rect 77635 30639 77693 30640
rect 48171 30596 48213 30605
rect 48171 30556 48172 30596
rect 48212 30556 48213 30596
rect 48171 30547 48213 30556
rect 48363 30596 48405 30605
rect 48363 30556 48364 30596
rect 48404 30556 48405 30596
rect 48363 30547 48405 30556
rect 56227 30596 56285 30597
rect 56227 30556 56236 30596
rect 56276 30556 56285 30596
rect 56227 30555 56285 30556
rect 71979 30596 72021 30605
rect 71979 30556 71980 30596
rect 72020 30556 72021 30596
rect 71979 30547 72021 30556
rect 72171 30596 72213 30605
rect 72171 30556 72172 30596
rect 72212 30556 72213 30596
rect 72171 30547 72213 30556
rect 48267 30512 48309 30521
rect 48267 30472 48268 30512
rect 48308 30472 48309 30512
rect 48267 30463 48309 30472
rect 72075 30512 72117 30521
rect 72075 30472 72076 30512
rect 72116 30472 72117 30512
rect 72075 30463 72117 30472
rect 53059 30428 53117 30429
rect 53059 30388 53068 30428
rect 53108 30388 53117 30428
rect 53059 30387 53117 30388
rect 56035 30428 56093 30429
rect 56035 30388 56044 30428
rect 56084 30388 56093 30428
rect 56035 30387 56093 30388
rect 56427 30428 56469 30437
rect 56427 30388 56428 30428
rect 56468 30388 56469 30428
rect 56427 30379 56469 30388
rect 60259 30428 60317 30429
rect 60259 30388 60268 30428
rect 60308 30388 60317 30428
rect 60259 30387 60317 30388
rect 63715 30428 63773 30429
rect 63715 30388 63724 30428
rect 63764 30388 63773 30428
rect 63715 30387 63773 30388
rect 67179 30428 67221 30437
rect 67179 30388 67180 30428
rect 67220 30388 67221 30428
rect 67179 30379 67221 30388
rect 69099 30428 69141 30437
rect 69099 30388 69100 30428
rect 69140 30388 69141 30428
rect 69099 30379 69141 30388
rect 69283 30428 69341 30429
rect 69283 30388 69292 30428
rect 69332 30388 69341 30428
rect 69283 30387 69341 30388
rect 77739 30428 77781 30437
rect 77739 30388 77740 30428
rect 77780 30388 77781 30428
rect 77739 30379 77781 30388
rect 576 30260 79584 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 75112 30260
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75480 30220 79584 30260
rect 576 30196 79584 30220
rect 53931 30092 53973 30101
rect 53931 30052 53932 30092
rect 53972 30052 53973 30092
rect 53931 30043 53973 30052
rect 55467 30092 55509 30101
rect 55467 30052 55468 30092
rect 55508 30052 55509 30092
rect 55467 30043 55509 30052
rect 59211 30092 59253 30101
rect 59211 30052 59212 30092
rect 59252 30052 59253 30092
rect 59211 30043 59253 30052
rect 59595 30092 59637 30101
rect 59595 30052 59596 30092
rect 59636 30052 59637 30092
rect 59595 30043 59637 30052
rect 60939 30092 60981 30101
rect 60939 30052 60940 30092
rect 60980 30052 60981 30092
rect 60939 30043 60981 30052
rect 61323 30092 61365 30101
rect 61323 30052 61324 30092
rect 61364 30052 61365 30092
rect 61323 30043 61365 30052
rect 70923 30092 70965 30101
rect 70923 30052 70924 30092
rect 70964 30052 70965 30092
rect 70923 30043 70965 30052
rect 71787 30092 71829 30101
rect 71787 30052 71788 30092
rect 71828 30052 71829 30092
rect 71787 30043 71829 30052
rect 72459 30092 72501 30101
rect 72459 30052 72460 30092
rect 72500 30052 72501 30092
rect 72459 30043 72501 30052
rect 72651 30092 72693 30101
rect 72651 30052 72652 30092
rect 72692 30052 72693 30092
rect 72651 30043 72693 30052
rect 73611 30092 73653 30101
rect 73611 30052 73612 30092
rect 73652 30052 73653 30092
rect 73611 30043 73653 30052
rect 74091 30092 74133 30101
rect 74091 30052 74092 30092
rect 74132 30052 74133 30092
rect 74091 30043 74133 30052
rect 61899 30008 61941 30017
rect 61899 29968 61900 30008
rect 61940 29968 61941 30008
rect 61899 29959 61941 29968
rect 65067 30008 65109 30017
rect 65067 29968 65068 30008
rect 65108 29968 65109 30008
rect 65067 29959 65109 29968
rect 65451 30008 65493 30017
rect 65451 29968 65452 30008
rect 65492 29968 65493 30008
rect 65451 29959 65493 29968
rect 65931 30008 65973 30017
rect 65931 29968 65932 30008
rect 65972 29968 65973 30008
rect 65931 29959 65973 29968
rect 75627 30008 75669 30017
rect 75627 29968 75628 30008
rect 75668 29968 75669 30008
rect 75627 29959 75669 29968
rect 76011 30008 76053 30017
rect 76011 29968 76012 30008
rect 76052 29968 76053 30008
rect 76011 29959 76053 29968
rect 76395 30008 76437 30017
rect 76395 29968 76396 30008
rect 76436 29968 76437 30008
rect 76395 29959 76437 29968
rect 40387 29924 40445 29925
rect 40387 29884 40396 29924
rect 40436 29884 40445 29924
rect 40387 29883 40445 29884
rect 48075 29924 48117 29933
rect 48075 29884 48076 29924
rect 48116 29884 48117 29924
rect 48075 29875 48117 29884
rect 51139 29924 51197 29925
rect 51139 29884 51148 29924
rect 51188 29884 51197 29924
rect 51139 29883 51197 29884
rect 55075 29924 55133 29925
rect 55075 29884 55084 29924
rect 55124 29884 55133 29924
rect 55075 29883 55133 29884
rect 55651 29924 55709 29925
rect 55651 29884 55660 29924
rect 55700 29884 55709 29924
rect 55651 29883 55709 29884
rect 59395 29924 59453 29925
rect 59395 29884 59404 29924
rect 59444 29884 59453 29924
rect 59395 29883 59453 29884
rect 59779 29924 59837 29925
rect 59779 29884 59788 29924
rect 59828 29884 59837 29924
rect 59779 29883 59837 29884
rect 60739 29924 60797 29925
rect 60739 29884 60748 29924
rect 60788 29884 60797 29924
rect 60739 29883 60797 29884
rect 61123 29924 61181 29925
rect 61123 29884 61132 29924
rect 61172 29884 61181 29924
rect 61123 29883 61181 29884
rect 61699 29924 61757 29925
rect 61699 29884 61708 29924
rect 61748 29884 61757 29924
rect 61699 29883 61757 29884
rect 62083 29924 62141 29925
rect 62083 29884 62092 29924
rect 62132 29884 62141 29924
rect 65355 29924 65397 29933
rect 62083 29883 62141 29884
rect 65259 29882 65301 29891
rect 46531 29840 46589 29841
rect 46531 29800 46540 29840
rect 46580 29800 46589 29840
rect 46531 29799 46589 29800
rect 47395 29840 47453 29841
rect 47395 29800 47404 29840
rect 47444 29800 47453 29840
rect 47395 29799 47453 29800
rect 47787 29840 47829 29849
rect 47787 29800 47788 29840
rect 47828 29800 47829 29840
rect 47787 29791 47829 29800
rect 47971 29840 48029 29841
rect 47971 29800 47980 29840
rect 48020 29800 48029 29840
rect 47971 29799 48029 29800
rect 48739 29840 48797 29841
rect 48739 29800 48748 29840
rect 48788 29800 48797 29840
rect 48739 29799 48797 29800
rect 49603 29840 49661 29841
rect 49603 29800 49612 29840
rect 49652 29800 49661 29840
rect 49603 29799 49661 29800
rect 51435 29840 51477 29849
rect 51435 29800 51436 29840
rect 51476 29800 51477 29840
rect 51435 29791 51477 29800
rect 51531 29840 51573 29849
rect 51531 29800 51532 29840
rect 51572 29800 51573 29840
rect 51531 29791 51573 29800
rect 51627 29840 51669 29849
rect 51627 29800 51628 29840
rect 51668 29800 51669 29840
rect 51627 29791 51669 29800
rect 51723 29840 51765 29849
rect 51723 29800 51724 29840
rect 51764 29800 51765 29840
rect 51723 29791 51765 29800
rect 52195 29840 52253 29841
rect 52195 29800 52204 29840
rect 52244 29800 52253 29840
rect 52195 29799 52253 29800
rect 54219 29840 54261 29849
rect 54219 29800 54220 29840
rect 54260 29800 54261 29840
rect 54219 29791 54261 29800
rect 54307 29840 54365 29841
rect 54307 29800 54316 29840
rect 54356 29800 54365 29840
rect 54307 29799 54365 29800
rect 54603 29840 54645 29849
rect 54603 29800 54604 29840
rect 54644 29800 54645 29840
rect 54603 29791 54645 29800
rect 54699 29840 54741 29849
rect 54699 29800 54700 29840
rect 54740 29800 54741 29840
rect 54699 29791 54741 29800
rect 54795 29840 54837 29849
rect 54795 29800 54796 29840
rect 54836 29800 54837 29840
rect 54795 29791 54837 29800
rect 54891 29840 54933 29849
rect 54891 29800 54892 29840
rect 54932 29800 54933 29840
rect 54891 29791 54933 29800
rect 56035 29840 56093 29841
rect 56035 29800 56044 29840
rect 56084 29800 56093 29840
rect 56035 29799 56093 29800
rect 56139 29840 56181 29849
rect 56139 29800 56140 29840
rect 56180 29800 56181 29840
rect 56139 29791 56181 29800
rect 56331 29840 56373 29849
rect 56331 29800 56332 29840
rect 56372 29800 56373 29840
rect 56331 29791 56373 29800
rect 56995 29840 57053 29841
rect 56995 29800 57004 29840
rect 57044 29800 57053 29840
rect 56995 29799 57053 29800
rect 57859 29840 57917 29841
rect 57859 29800 57868 29840
rect 57908 29800 57917 29840
rect 57859 29799 57917 29800
rect 64771 29840 64829 29841
rect 64771 29800 64780 29840
rect 64820 29800 64829 29840
rect 64771 29799 64829 29800
rect 64875 29840 64917 29849
rect 64875 29800 64876 29840
rect 64916 29800 64917 29840
rect 64875 29791 64917 29800
rect 65067 29840 65109 29849
rect 65067 29800 65068 29840
rect 65108 29800 65109 29840
rect 65259 29842 65260 29882
rect 65300 29842 65301 29882
rect 65355 29884 65356 29924
rect 65396 29884 65397 29924
rect 65355 29875 65397 29884
rect 65547 29924 65589 29933
rect 65547 29884 65548 29924
rect 65588 29884 65589 29924
rect 65547 29875 65589 29884
rect 70723 29924 70781 29925
rect 70723 29884 70732 29924
rect 70772 29884 70781 29924
rect 70723 29883 70781 29884
rect 71587 29924 71645 29925
rect 71587 29884 71596 29924
rect 71636 29884 71645 29924
rect 71587 29883 71645 29884
rect 72835 29924 72893 29925
rect 72835 29884 72844 29924
rect 72884 29884 72893 29924
rect 73795 29924 73853 29925
rect 72835 29883 72893 29884
rect 73419 29885 73461 29894
rect 65259 29833 65301 29842
rect 65635 29840 65693 29841
rect 65067 29791 65109 29800
rect 65635 29800 65644 29840
rect 65684 29800 65693 29840
rect 65635 29799 65693 29800
rect 66219 29840 66261 29849
rect 66219 29800 66220 29840
rect 66260 29800 66261 29840
rect 66219 29791 66261 29800
rect 66307 29840 66365 29841
rect 66307 29800 66316 29840
rect 66356 29800 66365 29840
rect 66307 29799 66365 29800
rect 67075 29840 67133 29841
rect 67075 29800 67084 29840
rect 67124 29800 67133 29840
rect 67075 29799 67133 29800
rect 67939 29840 67997 29841
rect 67939 29800 67948 29840
rect 67988 29800 67997 29840
rect 67939 29799 67997 29800
rect 71115 29840 71157 29849
rect 71115 29800 71116 29840
rect 71156 29800 71157 29840
rect 71115 29791 71157 29800
rect 71307 29840 71349 29849
rect 71307 29800 71308 29840
rect 71348 29800 71349 29840
rect 71307 29791 71349 29800
rect 71395 29840 71453 29841
rect 71395 29800 71404 29840
rect 71444 29800 71453 29840
rect 71395 29799 71453 29800
rect 72067 29840 72125 29841
rect 72067 29800 72076 29840
rect 72116 29800 72125 29840
rect 72067 29799 72125 29800
rect 72171 29840 72213 29849
rect 72171 29800 72172 29840
rect 72212 29800 72213 29840
rect 72171 29791 72213 29800
rect 73131 29840 73173 29849
rect 73131 29800 73132 29840
rect 73172 29800 73173 29840
rect 73131 29791 73173 29800
rect 73227 29840 73269 29849
rect 73227 29800 73228 29840
rect 73268 29800 73269 29840
rect 73227 29791 73269 29800
rect 73323 29840 73365 29849
rect 73323 29800 73324 29840
rect 73364 29800 73365 29840
rect 73419 29845 73420 29885
rect 73460 29845 73461 29885
rect 73795 29884 73804 29924
rect 73844 29884 73853 29924
rect 73795 29883 73853 29884
rect 75427 29924 75485 29925
rect 75427 29884 75436 29924
rect 75476 29884 75485 29924
rect 75427 29883 75485 29884
rect 75915 29924 75957 29933
rect 75915 29884 75916 29924
rect 75956 29884 75957 29924
rect 75915 29875 75957 29884
rect 76107 29924 76149 29933
rect 76107 29884 76108 29924
rect 76148 29884 76149 29924
rect 76107 29875 76149 29884
rect 73419 29836 73461 29845
rect 73987 29840 74045 29841
rect 73323 29791 73365 29800
rect 73987 29800 73996 29840
rect 74036 29800 74045 29840
rect 73987 29799 74045 29800
rect 75819 29840 75861 29849
rect 75819 29800 75820 29840
rect 75860 29800 75861 29840
rect 75819 29791 75861 29800
rect 76195 29840 76253 29841
rect 76195 29800 76204 29840
rect 76244 29800 76253 29840
rect 76195 29799 76253 29800
rect 76683 29840 76725 29849
rect 76683 29800 76684 29840
rect 76724 29800 76725 29840
rect 76683 29791 76725 29800
rect 76771 29840 76829 29841
rect 76771 29800 76780 29840
rect 76820 29800 76829 29840
rect 76771 29799 76829 29800
rect 77443 29840 77501 29841
rect 77443 29800 77452 29840
rect 77492 29800 77501 29840
rect 77443 29799 77501 29800
rect 78307 29840 78365 29841
rect 78307 29800 78316 29840
rect 78356 29800 78365 29840
rect 78307 29799 78365 29800
rect 48363 29756 48405 29765
rect 48363 29716 48364 29756
rect 48404 29716 48405 29756
rect 48363 29707 48405 29716
rect 56619 29756 56661 29765
rect 56619 29716 56620 29756
rect 56660 29716 56661 29756
rect 56619 29707 56661 29716
rect 66699 29756 66741 29765
rect 66699 29716 66700 29756
rect 66740 29716 66741 29756
rect 66699 29707 66741 29716
rect 77067 29756 77109 29765
rect 77067 29716 77068 29756
rect 77108 29716 77109 29756
rect 77067 29707 77109 29716
rect 40587 29672 40629 29681
rect 40587 29632 40588 29672
rect 40628 29632 40629 29672
rect 40587 29623 40629 29632
rect 45379 29672 45437 29673
rect 45379 29632 45388 29672
rect 45428 29632 45437 29672
rect 45379 29631 45437 29632
rect 50755 29672 50813 29673
rect 50755 29632 50764 29672
rect 50804 29632 50813 29672
rect 50755 29631 50813 29632
rect 50955 29672 50997 29681
rect 50955 29632 50956 29672
rect 50996 29632 50997 29672
rect 50955 29623 50997 29632
rect 52107 29672 52149 29681
rect 52107 29632 52108 29672
rect 52148 29632 52149 29672
rect 52107 29623 52149 29632
rect 54411 29668 54453 29677
rect 54411 29628 54412 29668
rect 54452 29628 54453 29668
rect 54411 29619 54453 29628
rect 55275 29672 55317 29681
rect 55275 29632 55276 29672
rect 55316 29632 55317 29672
rect 55275 29623 55317 29632
rect 56227 29672 56285 29673
rect 56227 29632 56236 29672
rect 56276 29632 56285 29672
rect 56227 29631 56285 29632
rect 59011 29672 59069 29673
rect 59011 29632 59020 29672
rect 59060 29632 59069 29672
rect 59011 29631 59069 29632
rect 59211 29672 59253 29681
rect 59211 29632 59212 29672
rect 59252 29632 59253 29672
rect 59211 29623 59253 29632
rect 60939 29672 60981 29681
rect 60939 29632 60940 29672
rect 60980 29632 60981 29672
rect 60939 29623 60981 29632
rect 61323 29672 61365 29681
rect 61323 29632 61324 29672
rect 61364 29632 61365 29672
rect 61323 29623 61365 29632
rect 61515 29672 61557 29681
rect 61515 29632 61516 29672
rect 61556 29632 61557 29672
rect 61515 29623 61557 29632
rect 66411 29668 66453 29677
rect 66411 29628 66412 29668
rect 66452 29628 66453 29668
rect 69091 29672 69149 29673
rect 69091 29632 69100 29672
rect 69140 29632 69149 29672
rect 69091 29631 69149 29632
rect 71203 29672 71261 29673
rect 71203 29632 71212 29672
rect 71252 29632 71261 29672
rect 71203 29631 71261 29632
rect 71787 29672 71829 29681
rect 71787 29632 71788 29672
rect 71828 29632 71829 29672
rect 66411 29619 66453 29628
rect 71787 29623 71829 29632
rect 71979 29668 72021 29677
rect 71979 29628 71980 29668
rect 72020 29628 72021 29668
rect 71979 29619 72021 29628
rect 72651 29672 72693 29681
rect 72651 29632 72652 29672
rect 72692 29632 72693 29672
rect 72651 29623 72693 29632
rect 74091 29672 74133 29681
rect 74091 29632 74092 29672
rect 74132 29632 74133 29672
rect 74091 29623 74133 29632
rect 76875 29668 76917 29677
rect 76875 29628 76876 29668
rect 76916 29628 76917 29668
rect 79459 29672 79517 29673
rect 79459 29632 79468 29672
rect 79508 29632 79517 29672
rect 79459 29631 79517 29632
rect 76875 29619 76917 29628
rect 576 29504 79584 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 76352 29504
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76720 29464 79584 29504
rect 576 29440 79584 29464
rect 47979 29394 48021 29403
rect 47979 29354 47980 29394
rect 48020 29354 48021 29394
rect 47979 29345 48021 29354
rect 39915 29336 39957 29345
rect 39915 29296 39916 29336
rect 39956 29296 39957 29336
rect 39915 29287 39957 29296
rect 46723 29336 46781 29337
rect 46723 29296 46732 29336
rect 46772 29296 46781 29336
rect 46723 29295 46781 29296
rect 51043 29336 51101 29337
rect 51043 29296 51052 29336
rect 51092 29296 51101 29336
rect 51043 29295 51101 29296
rect 51819 29336 51861 29345
rect 51819 29296 51820 29336
rect 51860 29296 51861 29336
rect 51819 29287 51861 29296
rect 57483 29340 57525 29349
rect 57483 29300 57484 29340
rect 57524 29300 57525 29340
rect 57483 29291 57525 29300
rect 58155 29336 58197 29345
rect 58155 29296 58156 29336
rect 58196 29296 58197 29336
rect 58155 29287 58197 29296
rect 65451 29336 65493 29345
rect 65451 29296 65452 29336
rect 65492 29296 65493 29336
rect 65451 29287 65493 29296
rect 66307 29336 66365 29337
rect 66307 29296 66316 29336
rect 66356 29296 66365 29336
rect 66307 29295 66365 29296
rect 66987 29336 67029 29345
rect 66987 29296 66988 29336
rect 67028 29296 67029 29336
rect 66987 29287 67029 29296
rect 71115 29336 71157 29345
rect 71115 29296 71116 29336
rect 71156 29296 71157 29336
rect 71115 29287 71157 29296
rect 71307 29340 71349 29349
rect 71307 29300 71308 29340
rect 71348 29300 71349 29340
rect 71307 29291 71349 29300
rect 76579 29336 76637 29337
rect 76579 29296 76588 29336
rect 76628 29296 76637 29336
rect 76579 29295 76637 29296
rect 77443 29336 77501 29337
rect 77443 29296 77452 29336
rect 77492 29296 77501 29336
rect 77443 29295 77501 29296
rect 48651 29252 48693 29261
rect 48651 29212 48652 29252
rect 48692 29212 48693 29252
rect 48651 29203 48693 29212
rect 76971 29252 77013 29261
rect 76971 29212 76972 29252
rect 77012 29212 77013 29252
rect 76971 29203 77013 29212
rect 42603 29168 42645 29177
rect 42603 29128 42604 29168
rect 42644 29128 42645 29168
rect 42603 29119 42645 29128
rect 42699 29168 42741 29177
rect 42699 29128 42700 29168
rect 42740 29128 42741 29168
rect 42699 29119 42741 29128
rect 42795 29168 42837 29177
rect 42795 29128 42796 29168
rect 42836 29128 42837 29168
rect 42795 29119 42837 29128
rect 42891 29168 42933 29177
rect 42891 29128 42892 29168
rect 42932 29128 42933 29168
rect 42891 29119 42933 29128
rect 43083 29168 43125 29177
rect 43083 29128 43084 29168
rect 43124 29128 43125 29168
rect 43083 29119 43125 29128
rect 43275 29168 43317 29177
rect 43275 29128 43276 29168
rect 43316 29128 43317 29168
rect 43171 29126 43229 29127
rect 43171 29086 43180 29126
rect 43220 29086 43229 29126
rect 43275 29119 43317 29128
rect 43371 29168 43413 29177
rect 43371 29128 43372 29168
rect 43412 29128 43413 29168
rect 43371 29119 43413 29128
rect 46635 29168 46677 29177
rect 46635 29128 46636 29168
rect 46676 29128 46677 29168
rect 46635 29119 46677 29128
rect 46827 29168 46869 29177
rect 46827 29128 46828 29168
rect 46868 29128 46869 29168
rect 46827 29119 46869 29128
rect 46915 29168 46973 29169
rect 46915 29128 46924 29168
rect 46964 29128 46973 29168
rect 46915 29127 46973 29128
rect 47115 29168 47157 29177
rect 47115 29128 47116 29168
rect 47156 29128 47157 29168
rect 47115 29119 47157 29128
rect 47491 29168 47549 29169
rect 47491 29128 47500 29168
rect 47540 29128 47549 29168
rect 47491 29127 47549 29128
rect 48067 29168 48125 29169
rect 48067 29128 48076 29168
rect 48116 29128 48125 29168
rect 48067 29127 48125 29128
rect 48171 29168 48213 29177
rect 48171 29128 48172 29168
rect 48212 29128 48213 29168
rect 48171 29119 48213 29128
rect 48747 29168 48789 29177
rect 48747 29128 48748 29168
rect 48788 29128 48789 29168
rect 48747 29119 48789 29128
rect 48843 29168 48885 29177
rect 48843 29128 48844 29168
rect 48884 29128 48885 29168
rect 48843 29119 48885 29128
rect 48939 29168 48981 29177
rect 48939 29128 48940 29168
rect 48980 29128 48981 29168
rect 48939 29119 48981 29128
rect 49699 29168 49757 29169
rect 49699 29128 49708 29168
rect 49748 29128 49757 29168
rect 49699 29127 49757 29128
rect 50571 29168 50613 29177
rect 50571 29128 50572 29168
rect 50612 29128 50613 29168
rect 50571 29119 50613 29128
rect 50955 29168 50997 29177
rect 50955 29128 50956 29168
rect 50996 29128 50997 29168
rect 50955 29119 50997 29128
rect 51147 29168 51189 29177
rect 51147 29128 51148 29168
rect 51188 29128 51189 29168
rect 51147 29119 51189 29128
rect 51235 29168 51293 29169
rect 51235 29128 51244 29168
rect 51284 29128 51293 29168
rect 51235 29127 51293 29128
rect 52195 29168 52253 29169
rect 52195 29128 52204 29168
rect 52244 29128 52253 29168
rect 52195 29127 52253 29128
rect 53163 29168 53205 29177
rect 53163 29128 53164 29168
rect 53204 29128 53205 29168
rect 53163 29119 53205 29128
rect 53355 29168 53397 29177
rect 53355 29128 53356 29168
rect 53396 29128 53397 29168
rect 53251 29126 53309 29127
rect 43171 29085 43229 29086
rect 39715 29084 39773 29085
rect 39715 29044 39724 29084
rect 39764 29044 39773 29084
rect 39715 29043 39773 29044
rect 40099 29084 40157 29085
rect 40099 29044 40108 29084
rect 40148 29044 40157 29084
rect 40099 29043 40157 29044
rect 40675 29084 40733 29085
rect 40675 29044 40684 29084
rect 40724 29044 40733 29084
rect 40675 29043 40733 29044
rect 47211 29084 47253 29093
rect 47211 29044 47212 29084
rect 47252 29044 47253 29084
rect 47211 29035 47253 29044
rect 47403 29084 47445 29093
rect 53251 29086 53260 29126
rect 53300 29086 53309 29126
rect 53355 29119 53397 29128
rect 53451 29168 53493 29177
rect 53451 29128 53452 29168
rect 53492 29128 53493 29168
rect 53451 29119 53493 29128
rect 53643 29168 53685 29177
rect 53643 29128 53644 29168
rect 53684 29128 53685 29168
rect 53643 29119 53685 29128
rect 54019 29168 54077 29169
rect 54019 29128 54028 29168
rect 54068 29128 54077 29168
rect 54019 29127 54077 29128
rect 54883 29168 54941 29169
rect 54883 29128 54892 29168
rect 54932 29128 54941 29168
rect 54883 29127 54941 29128
rect 56427 29168 56469 29177
rect 56427 29128 56428 29168
rect 56468 29128 56469 29168
rect 56427 29119 56469 29128
rect 56803 29168 56861 29169
rect 56803 29128 56812 29168
rect 56852 29128 56861 29168
rect 56803 29127 56861 29128
rect 57291 29168 57333 29177
rect 57291 29128 57292 29168
rect 57332 29128 57333 29168
rect 57291 29119 57333 29128
rect 57379 29168 57437 29169
rect 57379 29128 57388 29168
rect 57428 29128 57437 29168
rect 57379 29127 57437 29128
rect 58243 29168 58301 29169
rect 58243 29128 58252 29168
rect 58292 29128 58301 29168
rect 58243 29127 58301 29128
rect 58819 29168 58877 29169
rect 58819 29128 58828 29168
rect 58868 29128 58877 29168
rect 58819 29127 58877 29128
rect 58923 29168 58965 29177
rect 58923 29128 58924 29168
rect 58964 29128 58965 29168
rect 58923 29119 58965 29128
rect 59115 29168 59157 29177
rect 59115 29128 59116 29168
rect 59156 29128 59157 29168
rect 59115 29119 59157 29128
rect 59307 29168 59349 29177
rect 59307 29128 59308 29168
rect 59348 29128 59349 29168
rect 59307 29119 59349 29128
rect 59683 29168 59741 29169
rect 59683 29128 59692 29168
rect 59732 29128 59741 29168
rect 59683 29127 59741 29128
rect 60547 29168 60605 29169
rect 60547 29128 60556 29168
rect 60596 29128 60605 29168
rect 60547 29127 60605 29128
rect 61899 29168 61941 29177
rect 61899 29128 61900 29168
rect 61940 29128 61941 29168
rect 61899 29119 61941 29128
rect 62275 29168 62333 29169
rect 62275 29128 62284 29168
rect 62324 29128 62333 29168
rect 62275 29127 62333 29128
rect 63139 29168 63197 29169
rect 63139 29128 63148 29168
rect 63188 29128 63197 29168
rect 63139 29127 63197 29128
rect 64491 29168 64533 29177
rect 64491 29128 64492 29168
rect 64532 29128 64533 29168
rect 64491 29119 64533 29128
rect 64867 29168 64925 29169
rect 64867 29128 64876 29168
rect 64916 29128 64925 29168
rect 64867 29127 64925 29128
rect 65835 29168 65877 29177
rect 65835 29128 65836 29168
rect 65876 29128 65877 29168
rect 65835 29119 65877 29128
rect 65931 29168 65973 29177
rect 65931 29128 65932 29168
rect 65972 29128 65973 29168
rect 65931 29119 65973 29128
rect 66027 29168 66069 29177
rect 66027 29128 66028 29168
rect 66068 29128 66069 29168
rect 66027 29119 66069 29128
rect 66123 29168 66165 29177
rect 66123 29128 66124 29168
rect 66164 29128 66165 29168
rect 66123 29119 66165 29128
rect 66411 29168 66453 29177
rect 66411 29128 66412 29168
rect 66452 29128 66453 29168
rect 66411 29119 66453 29128
rect 66507 29168 66549 29177
rect 66507 29128 66508 29168
rect 66548 29128 66549 29168
rect 66507 29119 66549 29128
rect 66603 29168 66645 29177
rect 66603 29128 66604 29168
rect 66644 29128 66645 29168
rect 66603 29119 66645 29128
rect 67363 29168 67421 29169
rect 67363 29128 67372 29168
rect 67412 29128 67421 29168
rect 67363 29127 67421 29128
rect 69571 29168 69629 29169
rect 69571 29128 69580 29168
rect 69620 29128 69629 29168
rect 69571 29127 69629 29128
rect 70435 29168 70493 29169
rect 70435 29128 70444 29168
rect 70484 29128 70493 29168
rect 70435 29127 70493 29128
rect 70827 29168 70869 29177
rect 70827 29128 70828 29168
rect 70868 29128 70869 29168
rect 70827 29119 70869 29128
rect 71011 29168 71069 29169
rect 71011 29128 71020 29168
rect 71060 29128 71069 29168
rect 71011 29127 71069 29128
rect 71395 29168 71453 29169
rect 71395 29128 71404 29168
rect 71444 29128 71453 29168
rect 71395 29127 71453 29128
rect 71499 29168 71541 29177
rect 71499 29128 71500 29168
rect 71540 29128 71541 29168
rect 71499 29119 71541 29128
rect 72171 29168 72213 29177
rect 72171 29128 72172 29168
rect 72212 29128 72213 29168
rect 72171 29119 72213 29128
rect 72547 29168 72605 29169
rect 72547 29128 72556 29168
rect 72596 29128 72605 29168
rect 72547 29127 72605 29128
rect 73452 29168 73494 29177
rect 73452 29128 73453 29168
rect 73493 29128 73494 29168
rect 73452 29119 73494 29128
rect 76491 29168 76533 29177
rect 76491 29128 76492 29168
rect 76532 29128 76533 29168
rect 76491 29119 76533 29128
rect 76683 29168 76725 29177
rect 76683 29128 76684 29168
rect 76724 29128 76725 29168
rect 76683 29119 76725 29128
rect 76771 29168 76829 29169
rect 76771 29128 76780 29168
rect 76820 29128 76829 29168
rect 76771 29127 76829 29128
rect 77067 29160 77109 29169
rect 77067 29120 77068 29160
rect 77108 29120 77109 29160
rect 77259 29168 77301 29177
rect 77259 29128 77260 29168
rect 77300 29128 77301 29168
rect 77067 29111 77109 29120
rect 77155 29126 77213 29127
rect 53251 29085 53309 29086
rect 47403 29044 47404 29084
rect 47444 29044 47445 29084
rect 47403 29035 47445 29044
rect 49507 29084 49565 29085
rect 49507 29044 49516 29084
rect 49556 29044 49565 29084
rect 49507 29043 49565 29044
rect 51619 29084 51677 29085
rect 51619 29044 51628 29084
rect 51668 29044 51677 29084
rect 51619 29043 51677 29044
rect 52003 29084 52061 29085
rect 52003 29044 52012 29084
rect 52052 29044 52061 29084
rect 52003 29043 52061 29044
rect 56523 29084 56565 29093
rect 56523 29044 56524 29084
rect 56564 29044 56565 29084
rect 56523 29035 56565 29044
rect 56715 29084 56757 29093
rect 56715 29044 56716 29084
rect 56756 29044 56757 29084
rect 56715 29035 56757 29044
rect 64587 29084 64629 29093
rect 64587 29044 64588 29084
rect 64628 29044 64629 29084
rect 64587 29035 64629 29044
rect 64779 29084 64821 29093
rect 77155 29086 77164 29126
rect 77204 29086 77213 29126
rect 77259 29119 77301 29128
rect 77547 29168 77589 29177
rect 77547 29128 77548 29168
rect 77588 29128 77589 29168
rect 77547 29119 77589 29128
rect 77643 29168 77685 29177
rect 77643 29128 77644 29168
rect 77684 29128 77685 29168
rect 77643 29119 77685 29128
rect 77739 29168 77781 29177
rect 77739 29128 77740 29168
rect 77780 29128 77781 29168
rect 77739 29119 77781 29128
rect 78019 29168 78077 29169
rect 78019 29128 78028 29168
rect 78068 29128 78077 29168
rect 78019 29127 78077 29128
rect 77155 29085 77213 29086
rect 64779 29044 64780 29084
rect 64820 29044 64821 29084
rect 64779 29035 64821 29044
rect 65251 29084 65309 29085
rect 65251 29044 65260 29084
rect 65300 29044 65309 29084
rect 65251 29043 65309 29044
rect 66787 29084 66845 29085
rect 66787 29044 66796 29084
rect 66836 29044 66845 29084
rect 66787 29043 66845 29044
rect 47307 29000 47349 29009
rect 47307 28960 47308 29000
rect 47348 28960 47349 29000
rect 47307 28951 47349 28960
rect 48459 29000 48501 29009
rect 48459 28960 48460 29000
rect 48500 28960 48501 29000
rect 48459 28951 48501 28960
rect 51435 29000 51477 29009
rect 51435 28960 51436 29000
rect 51476 28960 51477 29000
rect 51435 28951 51477 28960
rect 56619 29000 56661 29009
rect 56619 28960 56620 29000
rect 56660 28960 56661 29000
rect 56619 28951 56661 28960
rect 57003 29000 57045 29009
rect 57003 28960 57004 29000
rect 57044 28960 57045 29000
rect 57003 28951 57045 28960
rect 64683 29000 64725 29009
rect 64683 28960 64684 29000
rect 64724 28960 64725 29000
rect 64683 28951 64725 28960
rect 40299 28916 40341 28925
rect 40299 28876 40300 28916
rect 40340 28876 40341 28916
rect 40299 28867 40341 28876
rect 40491 28916 40533 28925
rect 40491 28876 40492 28916
rect 40532 28876 40533 28916
rect 40491 28867 40533 28876
rect 49323 28916 49365 28925
rect 49323 28876 49324 28916
rect 49364 28876 49365 28916
rect 49323 28867 49365 28876
rect 49995 28916 50037 28925
rect 49995 28876 49996 28916
rect 50036 28876 50037 28916
rect 49995 28867 50037 28876
rect 50379 28916 50421 28925
rect 50379 28876 50380 28916
rect 50420 28876 50421 28916
rect 50379 28867 50421 28876
rect 52299 28916 52341 28925
rect 52299 28876 52300 28916
rect 52340 28876 52341 28916
rect 52299 28867 52341 28876
rect 56035 28916 56093 28917
rect 56035 28876 56044 28916
rect 56084 28876 56093 28916
rect 56035 28875 56093 28876
rect 59115 28916 59157 28925
rect 59115 28876 59116 28916
rect 59156 28876 59157 28916
rect 59115 28867 59157 28876
rect 61699 28916 61757 28917
rect 61699 28876 61708 28916
rect 61748 28876 61757 28916
rect 61699 28875 61757 28876
rect 64291 28916 64349 28917
rect 64291 28876 64300 28916
rect 64340 28876 64349 28916
rect 64291 28875 64349 28876
rect 67467 28916 67509 28925
rect 67467 28876 67468 28916
rect 67508 28876 67509 28916
rect 67467 28867 67509 28876
rect 68419 28916 68477 28917
rect 68419 28876 68428 28916
rect 68468 28876 68477 28916
rect 68419 28875 68477 28876
rect 71115 28916 71157 28925
rect 71115 28876 71116 28916
rect 71156 28876 71157 28916
rect 71115 28867 71157 28876
rect 71787 28916 71829 28925
rect 71787 28876 71788 28916
rect 71828 28876 71829 28916
rect 71787 28867 71829 28876
rect 74563 28916 74621 28917
rect 74563 28876 74572 28916
rect 74612 28876 74621 28916
rect 74563 28875 74621 28876
rect 77931 28916 77973 28925
rect 77931 28876 77932 28916
rect 77972 28876 77973 28916
rect 77931 28867 77973 28876
rect 576 28748 79584 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 75112 28748
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75480 28708 79584 28748
rect 576 28684 79584 28708
rect 45187 28580 45245 28581
rect 45187 28540 45196 28580
rect 45236 28540 45245 28580
rect 45187 28539 45245 28540
rect 49699 28580 49757 28581
rect 49699 28540 49708 28580
rect 49748 28540 49757 28580
rect 49699 28539 49757 28540
rect 55179 28580 55221 28589
rect 55179 28540 55180 28580
rect 55220 28540 55221 28580
rect 55179 28531 55221 28540
rect 65443 28580 65501 28581
rect 65443 28540 65452 28580
rect 65492 28540 65501 28580
rect 65443 28539 65501 28540
rect 65739 28580 65781 28589
rect 65739 28540 65740 28580
rect 65780 28540 65781 28580
rect 65739 28531 65781 28540
rect 72267 28580 72309 28589
rect 72267 28540 72268 28580
rect 72308 28540 72309 28580
rect 72267 28531 72309 28540
rect 76867 28580 76925 28581
rect 76867 28540 76876 28580
rect 76916 28540 76925 28580
rect 76867 28539 76925 28540
rect 42411 28496 42453 28505
rect 42411 28456 42412 28496
rect 42452 28456 42453 28496
rect 42411 28447 42453 28456
rect 52779 28496 52821 28505
rect 52779 28456 52780 28496
rect 52820 28456 52821 28496
rect 52779 28447 52821 28456
rect 59979 28496 60021 28505
rect 59979 28456 59980 28496
rect 60020 28456 60021 28496
rect 59979 28447 60021 28456
rect 61323 28496 61365 28505
rect 61323 28456 61324 28496
rect 61364 28456 61365 28496
rect 61323 28447 61365 28456
rect 70731 28496 70773 28505
rect 70731 28456 70732 28496
rect 70772 28456 70773 28496
rect 70731 28447 70773 28456
rect 71115 28496 71157 28505
rect 71115 28456 71116 28496
rect 71156 28456 71157 28496
rect 71115 28447 71157 28456
rect 77067 28496 77109 28505
rect 77067 28456 77068 28496
rect 77108 28456 77109 28496
rect 77067 28447 77109 28456
rect 42315 28412 42357 28421
rect 42315 28372 42316 28412
rect 42356 28372 42357 28412
rect 42315 28363 42357 28372
rect 42507 28412 42549 28421
rect 42507 28372 42508 28412
rect 42548 28372 42549 28412
rect 42507 28363 42549 28372
rect 59883 28412 59925 28421
rect 59883 28372 59884 28412
rect 59924 28372 59925 28412
rect 52483 28370 52541 28371
rect 43171 28364 43229 28365
rect 40771 28328 40829 28329
rect 40771 28288 40780 28328
rect 40820 28288 40829 28328
rect 40771 28287 40829 28288
rect 41635 28328 41693 28329
rect 41635 28288 41644 28328
rect 41684 28288 41693 28328
rect 41635 28287 41693 28288
rect 42027 28328 42069 28337
rect 42027 28288 42028 28328
rect 42068 28288 42069 28328
rect 42027 28279 42069 28288
rect 42219 28328 42261 28337
rect 42219 28288 42220 28328
rect 42260 28288 42261 28328
rect 42219 28279 42261 28288
rect 42595 28328 42653 28329
rect 42595 28288 42604 28328
rect 42644 28288 42653 28328
rect 42595 28287 42653 28288
rect 42795 28328 42837 28337
rect 42795 28288 42796 28328
rect 42836 28288 42837 28328
rect 43171 28324 43180 28364
rect 43220 28324 43229 28364
rect 43171 28323 43229 28324
rect 44035 28328 44093 28329
rect 42795 28279 42837 28288
rect 44035 28288 44044 28328
rect 44084 28288 44093 28328
rect 44035 28287 44093 28288
rect 45387 28328 45429 28337
rect 45387 28288 45388 28328
rect 45428 28288 45429 28328
rect 45387 28279 45429 28288
rect 45763 28328 45821 28329
rect 45763 28288 45772 28328
rect 45812 28288 45821 28328
rect 45763 28287 45821 28288
rect 46627 28328 46685 28329
rect 46627 28288 46636 28328
rect 46676 28288 46685 28328
rect 46627 28287 46685 28288
rect 48171 28328 48213 28337
rect 48171 28288 48172 28328
rect 48212 28288 48213 28328
rect 48171 28279 48213 28288
rect 48267 28328 48309 28337
rect 48267 28288 48268 28328
rect 48308 28288 48309 28328
rect 48267 28279 48309 28288
rect 48363 28328 48405 28337
rect 48363 28288 48364 28328
rect 48404 28288 48405 28328
rect 48363 28279 48405 28288
rect 48459 28328 48501 28337
rect 52483 28330 52492 28370
rect 52532 28330 52541 28370
rect 59883 28363 59925 28372
rect 60075 28412 60117 28421
rect 60075 28372 60076 28412
rect 60116 28372 60117 28412
rect 60075 28363 60117 28372
rect 69091 28412 69149 28413
rect 69091 28372 69100 28412
rect 69140 28372 69149 28412
rect 69091 28371 69149 28372
rect 71019 28412 71061 28421
rect 71019 28372 71020 28412
rect 71060 28372 71061 28412
rect 71019 28363 71061 28372
rect 71211 28412 71253 28421
rect 71211 28372 71212 28412
rect 71252 28372 71253 28412
rect 71211 28363 71253 28372
rect 72451 28412 72509 28413
rect 72451 28372 72460 28412
rect 72500 28372 72509 28412
rect 72451 28371 72509 28372
rect 70531 28342 70589 28343
rect 52483 28329 52541 28330
rect 48459 28288 48460 28328
rect 48500 28288 48501 28328
rect 48459 28279 48501 28288
rect 50851 28328 50909 28329
rect 50851 28288 50860 28328
rect 50900 28288 50909 28328
rect 50851 28287 50909 28288
rect 51715 28328 51773 28329
rect 51715 28288 51724 28328
rect 51764 28288 51773 28328
rect 51715 28287 51773 28288
rect 52387 28328 52445 28329
rect 52387 28288 52396 28328
rect 52436 28288 52445 28328
rect 52387 28287 52445 28288
rect 53067 28328 53109 28337
rect 53067 28288 53068 28328
rect 53108 28288 53109 28328
rect 53067 28279 53109 28288
rect 53163 28328 53205 28337
rect 53163 28288 53164 28328
rect 53204 28288 53205 28328
rect 53163 28279 53205 28288
rect 53259 28328 53301 28337
rect 53259 28288 53260 28328
rect 53300 28288 53301 28328
rect 53259 28279 53301 28288
rect 55075 28328 55133 28329
rect 55075 28288 55084 28328
rect 55124 28288 55133 28328
rect 55075 28287 55133 28288
rect 56139 28328 56181 28337
rect 56139 28288 56140 28328
rect 56180 28288 56181 28328
rect 56139 28279 56181 28288
rect 56235 28328 56277 28337
rect 56235 28288 56236 28328
rect 56276 28288 56277 28328
rect 56235 28279 56277 28288
rect 56331 28328 56373 28337
rect 56331 28288 56332 28328
rect 56372 28288 56373 28328
rect 56331 28279 56373 28288
rect 56995 28328 57053 28329
rect 56995 28288 57004 28328
rect 57044 28288 57053 28328
rect 56995 28287 57053 28288
rect 57859 28328 57917 28329
rect 57859 28288 57868 28328
rect 57908 28288 57917 28328
rect 57859 28287 57917 28288
rect 59787 28328 59829 28337
rect 59787 28288 59788 28328
rect 59828 28288 59829 28328
rect 59787 28279 59829 28288
rect 60163 28328 60221 28329
rect 60163 28288 60172 28328
rect 60212 28288 60221 28328
rect 60163 28287 60221 28288
rect 60555 28328 60597 28337
rect 60555 28288 60556 28328
rect 60596 28288 60597 28328
rect 60555 28279 60597 28288
rect 60643 28328 60701 28329
rect 60643 28288 60652 28328
rect 60692 28288 60701 28328
rect 60643 28287 60701 28288
rect 60931 28328 60989 28329
rect 60931 28288 60940 28328
rect 60980 28288 60989 28328
rect 60931 28287 60989 28288
rect 61035 28328 61077 28337
rect 61035 28288 61036 28328
rect 61076 28288 61077 28328
rect 61035 28279 61077 28288
rect 61515 28328 61557 28337
rect 61515 28288 61516 28328
rect 61556 28288 61557 28328
rect 61515 28279 61557 28288
rect 61611 28328 61653 28337
rect 61611 28288 61612 28328
rect 61652 28288 61653 28328
rect 61611 28279 61653 28288
rect 61707 28328 61749 28337
rect 61707 28288 61708 28328
rect 61748 28288 61749 28328
rect 61707 28279 61749 28288
rect 61803 28328 61845 28337
rect 61803 28288 61804 28328
rect 61844 28288 61845 28328
rect 61803 28279 61845 28288
rect 61995 28328 62037 28337
rect 61995 28288 61996 28328
rect 62036 28288 62037 28328
rect 61995 28279 62037 28288
rect 62091 28328 62133 28337
rect 62091 28288 62092 28328
rect 62132 28288 62133 28328
rect 62091 28279 62133 28288
rect 62187 28328 62229 28337
rect 62187 28288 62188 28328
rect 62228 28288 62229 28328
rect 62187 28279 62229 28288
rect 62283 28328 62325 28337
rect 62283 28288 62284 28328
rect 62324 28288 62325 28328
rect 62283 28279 62325 28288
rect 62851 28328 62909 28329
rect 62851 28288 62860 28328
rect 62900 28288 62909 28328
rect 62851 28287 62909 28288
rect 63051 28328 63093 28337
rect 63051 28288 63052 28328
rect 63092 28288 63093 28328
rect 63051 28279 63093 28288
rect 63427 28328 63485 28329
rect 63427 28288 63436 28328
rect 63476 28288 63485 28328
rect 63427 28287 63485 28288
rect 64291 28328 64349 28329
rect 64291 28288 64300 28328
rect 64340 28288 64349 28328
rect 64291 28287 64349 28288
rect 65635 28328 65693 28329
rect 65635 28288 65644 28328
rect 65684 28288 65693 28328
rect 65635 28287 65693 28288
rect 66307 28328 66365 28329
rect 66307 28288 66316 28328
rect 66356 28288 66365 28328
rect 66307 28287 66365 28288
rect 67171 28328 67229 28329
rect 67171 28288 67180 28328
rect 67220 28288 67229 28328
rect 67171 28287 67229 28288
rect 70435 28328 70493 28329
rect 70435 28288 70444 28328
rect 70484 28288 70493 28328
rect 70531 28302 70540 28342
rect 70580 28302 70589 28342
rect 70531 28301 70589 28302
rect 70731 28339 70773 28348
rect 70731 28299 70732 28339
rect 70772 28299 70773 28339
rect 70731 28290 70773 28299
rect 70915 28328 70973 28329
rect 70435 28287 70493 28288
rect 70915 28288 70924 28328
rect 70964 28288 70973 28328
rect 70915 28287 70973 28288
rect 71307 28328 71349 28337
rect 71307 28288 71308 28328
rect 71348 28288 71349 28328
rect 71307 28279 71349 28288
rect 71787 28328 71829 28337
rect 71787 28288 71788 28328
rect 71828 28288 71829 28328
rect 71787 28279 71829 28288
rect 71883 28328 71925 28337
rect 71883 28288 71884 28328
rect 71924 28288 71925 28328
rect 71883 28279 71925 28288
rect 71979 28328 72021 28337
rect 71979 28288 71980 28328
rect 72020 28288 72021 28328
rect 71979 28279 72021 28288
rect 72075 28328 72117 28337
rect 72075 28288 72076 28328
rect 72116 28288 72117 28328
rect 72075 28279 72117 28288
rect 72747 28328 72789 28337
rect 72747 28288 72748 28328
rect 72788 28288 72789 28328
rect 72747 28279 72789 28288
rect 72843 28328 72885 28337
rect 72843 28288 72844 28328
rect 72884 28288 72885 28328
rect 72843 28279 72885 28288
rect 72939 28328 72981 28337
rect 72939 28288 72940 28328
rect 72980 28288 72981 28328
rect 72939 28279 72981 28288
rect 73035 28328 73077 28337
rect 73035 28288 73036 28328
rect 73076 28288 73077 28328
rect 73035 28279 73077 28288
rect 73699 28328 73757 28329
rect 73699 28288 73708 28328
rect 73748 28288 73757 28328
rect 73699 28287 73757 28288
rect 74851 28328 74909 28329
rect 74851 28288 74860 28328
rect 74900 28288 74909 28328
rect 74851 28287 74909 28288
rect 75715 28328 75773 28329
rect 75715 28288 75724 28328
rect 75764 28288 75773 28328
rect 75715 28287 75773 28288
rect 77355 28328 77397 28337
rect 77355 28288 77356 28328
rect 77396 28288 77397 28328
rect 77355 28279 77397 28288
rect 77443 28328 77501 28329
rect 77443 28288 77452 28328
rect 77492 28288 77501 28328
rect 77443 28287 77501 28288
rect 77731 28328 77789 28329
rect 77731 28288 77740 28328
rect 77780 28288 77789 28328
rect 77731 28287 77789 28288
rect 52107 28244 52149 28253
rect 52107 28204 52108 28244
rect 52148 28204 52149 28244
rect 52107 28195 52149 28204
rect 56427 28244 56469 28253
rect 56427 28204 56428 28244
rect 56468 28204 56469 28244
rect 56427 28195 56469 28204
rect 56619 28244 56661 28253
rect 56619 28204 56620 28244
rect 56660 28204 56661 28244
rect 56619 28195 56661 28204
rect 65931 28244 65973 28253
rect 65931 28204 65932 28244
rect 65972 28204 65973 28244
rect 65931 28195 65973 28204
rect 74475 28244 74517 28253
rect 74475 28204 74476 28244
rect 74516 28204 74517 28244
rect 74475 28195 74517 28204
rect 39619 28160 39677 28161
rect 39619 28120 39628 28160
rect 39668 28120 39677 28160
rect 39619 28119 39677 28120
rect 45187 28160 45245 28161
rect 45187 28120 45196 28160
rect 45236 28120 45245 28160
rect 45187 28119 45245 28120
rect 47779 28160 47837 28161
rect 47779 28120 47788 28160
rect 47828 28120 47837 28160
rect 47779 28119 47837 28120
rect 52299 28156 52341 28165
rect 52299 28116 52300 28156
rect 52340 28116 52341 28156
rect 52963 28160 53021 28161
rect 52963 28120 52972 28160
rect 53012 28120 53021 28160
rect 52963 28119 53021 28120
rect 55179 28160 55221 28169
rect 55179 28120 55180 28160
rect 55220 28120 55221 28160
rect 52299 28107 52341 28116
rect 55179 28111 55221 28120
rect 59011 28160 59069 28161
rect 59011 28120 59020 28160
rect 59060 28120 59069 28160
rect 59011 28119 59069 28120
rect 60843 28156 60885 28165
rect 60843 28116 60844 28156
rect 60884 28116 60885 28156
rect 60843 28107 60885 28116
rect 62763 28160 62805 28169
rect 62763 28120 62764 28160
rect 62804 28120 62805 28160
rect 62763 28111 62805 28120
rect 65739 28160 65781 28169
rect 65739 28120 65740 28160
rect 65780 28120 65781 28160
rect 65739 28111 65781 28120
rect 68323 28160 68381 28161
rect 68323 28120 68332 28160
rect 68372 28120 68381 28160
rect 68323 28119 68381 28120
rect 68907 28160 68949 28169
rect 68907 28120 68908 28160
rect 68948 28120 68949 28160
rect 68907 28111 68949 28120
rect 73611 28160 73653 28169
rect 73611 28120 73612 28160
rect 73652 28120 73653 28160
rect 73611 28111 73653 28120
rect 77835 28160 77877 28169
rect 77835 28120 77836 28160
rect 77876 28120 77877 28160
rect 77835 28111 77877 28120
rect 77547 28102 77589 28111
rect 77547 28062 77548 28102
rect 77588 28062 77589 28102
rect 77547 28053 77589 28062
rect 576 27992 79584 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 76352 27992
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76720 27952 79584 27992
rect 576 27928 79584 27952
rect 65547 27882 65589 27891
rect 65547 27842 65548 27882
rect 65588 27842 65589 27882
rect 42219 27824 42261 27833
rect 42219 27784 42220 27824
rect 42260 27784 42261 27824
rect 42219 27775 42261 27784
rect 42507 27828 42549 27837
rect 42507 27788 42508 27828
rect 42548 27788 42549 27828
rect 42507 27779 42549 27788
rect 46059 27824 46101 27833
rect 46059 27784 46060 27824
rect 46100 27784 46101 27824
rect 46059 27775 46101 27784
rect 47307 27824 47349 27833
rect 47307 27784 47308 27824
rect 47348 27784 47349 27824
rect 47307 27775 47349 27784
rect 47595 27828 47637 27837
rect 65547 27833 65589 27842
rect 47595 27788 47596 27828
rect 47636 27788 47637 27828
rect 47595 27779 47637 27788
rect 57475 27824 57533 27825
rect 57475 27784 57484 27824
rect 57524 27784 57533 27824
rect 57475 27783 57533 27784
rect 59403 27824 59445 27833
rect 59403 27784 59404 27824
rect 59444 27784 59445 27824
rect 47971 27782 48029 27783
rect 47971 27742 47980 27782
rect 48020 27742 48029 27782
rect 59403 27775 59445 27784
rect 66019 27824 66077 27825
rect 66019 27784 66028 27824
rect 66068 27784 66077 27824
rect 66019 27783 66077 27784
rect 71115 27824 71157 27833
rect 71115 27784 71116 27824
rect 71156 27784 71157 27824
rect 71115 27775 71157 27784
rect 71499 27828 71541 27837
rect 71499 27788 71500 27828
rect 71540 27788 71541 27828
rect 71499 27779 71541 27788
rect 47971 27741 48029 27742
rect 53163 27740 53205 27749
rect 43179 27698 43221 27707
rect 40587 27656 40629 27665
rect 40587 27616 40588 27656
rect 40628 27616 40629 27656
rect 40587 27607 40629 27616
rect 40779 27656 40821 27665
rect 40779 27616 40780 27656
rect 40820 27616 40821 27656
rect 40779 27607 40821 27616
rect 40867 27656 40925 27657
rect 40867 27616 40876 27656
rect 40916 27616 40925 27656
rect 40867 27615 40925 27616
rect 42115 27656 42173 27657
rect 42115 27616 42124 27656
rect 42164 27616 42173 27656
rect 42115 27615 42173 27616
rect 42595 27656 42653 27657
rect 42595 27616 42604 27656
rect 42644 27616 42653 27656
rect 42595 27615 42653 27616
rect 42699 27656 42741 27665
rect 42699 27616 42700 27656
rect 42740 27616 42741 27656
rect 43179 27658 43180 27698
rect 43220 27658 43221 27698
rect 53163 27700 53164 27740
rect 53204 27700 53205 27740
rect 53163 27691 53205 27700
rect 43179 27649 43221 27658
rect 43371 27656 43413 27665
rect 42699 27607 42741 27616
rect 43371 27616 43372 27656
rect 43412 27616 43413 27656
rect 43371 27607 43413 27616
rect 43459 27656 43517 27657
rect 43459 27616 43468 27656
rect 43508 27616 43517 27656
rect 43459 27615 43517 27616
rect 43651 27656 43709 27657
rect 43651 27616 43660 27656
rect 43700 27616 43709 27656
rect 43651 27615 43709 27616
rect 44035 27656 44093 27657
rect 44035 27616 44044 27656
rect 44084 27616 44093 27656
rect 44035 27615 44093 27616
rect 47395 27656 47453 27657
rect 47395 27616 47404 27656
rect 47444 27616 47453 27656
rect 47395 27615 47453 27616
rect 47683 27656 47741 27657
rect 47683 27616 47692 27656
rect 47732 27616 47741 27656
rect 47683 27615 47741 27616
rect 47787 27656 47829 27665
rect 47787 27616 47788 27656
rect 47828 27616 47829 27656
rect 47787 27607 47829 27616
rect 48267 27656 48309 27665
rect 48267 27616 48268 27656
rect 48308 27616 48309 27656
rect 48267 27607 48309 27616
rect 48363 27656 48405 27665
rect 48363 27616 48364 27656
rect 48404 27616 48405 27656
rect 48363 27607 48405 27616
rect 48459 27656 48501 27665
rect 48459 27616 48460 27656
rect 48500 27616 48501 27656
rect 48459 27607 48501 27616
rect 48555 27656 48597 27665
rect 48555 27616 48556 27656
rect 48596 27616 48597 27656
rect 48555 27607 48597 27616
rect 48747 27656 48789 27665
rect 48747 27616 48748 27656
rect 48788 27616 48789 27656
rect 48747 27607 48789 27616
rect 49123 27656 49181 27657
rect 49123 27616 49132 27656
rect 49172 27616 49181 27656
rect 49123 27615 49181 27616
rect 49987 27656 50045 27657
rect 49987 27616 49996 27656
rect 50036 27616 50045 27656
rect 49987 27615 50045 27616
rect 52011 27656 52053 27665
rect 52011 27616 52012 27656
rect 52052 27616 52053 27656
rect 52011 27607 52053 27616
rect 52387 27656 52445 27657
rect 52387 27616 52396 27656
rect 52436 27616 52445 27656
rect 52779 27656 52821 27665
rect 52387 27615 52445 27616
rect 52587 27645 52629 27654
rect 52587 27605 52588 27645
rect 52628 27605 52629 27645
rect 52779 27616 52780 27656
rect 52820 27616 52821 27656
rect 52779 27607 52821 27616
rect 52867 27656 52925 27657
rect 52867 27616 52876 27656
rect 52916 27616 52925 27656
rect 52867 27615 52925 27616
rect 53539 27656 53597 27657
rect 53539 27616 53548 27656
rect 53588 27616 53597 27656
rect 53539 27615 53597 27616
rect 54403 27656 54461 27657
rect 54403 27616 54412 27656
rect 54452 27616 54461 27656
rect 54403 27615 54461 27616
rect 57579 27656 57621 27665
rect 57579 27616 57580 27656
rect 57620 27616 57621 27656
rect 57579 27607 57621 27616
rect 57675 27656 57717 27665
rect 57675 27616 57676 27656
rect 57716 27616 57717 27656
rect 57675 27607 57717 27616
rect 57771 27656 57813 27665
rect 57771 27616 57772 27656
rect 57812 27616 57813 27656
rect 57771 27607 57813 27616
rect 58051 27656 58109 27657
rect 58051 27616 58060 27656
rect 58100 27616 58109 27656
rect 58051 27615 58109 27616
rect 60651 27656 60693 27665
rect 60651 27616 60652 27656
rect 60692 27616 60693 27656
rect 60651 27607 60693 27616
rect 61027 27656 61085 27657
rect 61027 27616 61036 27656
rect 61076 27616 61085 27656
rect 61027 27615 61085 27616
rect 61227 27656 61269 27665
rect 61227 27616 61228 27656
rect 61268 27616 61269 27656
rect 61227 27607 61269 27616
rect 61419 27656 61461 27665
rect 61419 27616 61420 27656
rect 61460 27616 61461 27656
rect 61419 27607 61461 27616
rect 61507 27656 61565 27657
rect 61507 27616 61516 27656
rect 61556 27616 61565 27656
rect 61507 27615 61565 27616
rect 62379 27656 62421 27665
rect 62379 27616 62380 27656
rect 62420 27616 62421 27656
rect 62379 27607 62421 27616
rect 62755 27656 62813 27657
rect 62755 27616 62764 27656
rect 62804 27616 62813 27656
rect 62755 27615 62813 27616
rect 63619 27656 63677 27657
rect 63619 27616 63628 27656
rect 63668 27616 63677 27656
rect 63619 27615 63677 27616
rect 65355 27656 65397 27665
rect 65355 27616 65356 27656
rect 65396 27616 65397 27656
rect 65355 27607 65397 27616
rect 65443 27656 65501 27657
rect 65443 27616 65452 27656
rect 65492 27616 65501 27656
rect 65443 27615 65501 27616
rect 65739 27656 65781 27665
rect 65739 27616 65740 27656
rect 65780 27616 65781 27656
rect 65739 27607 65781 27616
rect 65835 27656 65877 27665
rect 65835 27616 65836 27656
rect 65876 27616 65877 27656
rect 65835 27607 65877 27616
rect 65931 27656 65973 27665
rect 65931 27616 65932 27656
rect 65972 27616 65973 27656
rect 65931 27607 65973 27616
rect 66499 27656 66557 27657
rect 66499 27616 66508 27656
rect 66548 27616 66557 27656
rect 66499 27615 66557 27616
rect 69571 27656 69629 27657
rect 69571 27616 69580 27656
rect 69620 27616 69629 27656
rect 69571 27615 69629 27616
rect 70435 27656 70493 27657
rect 70435 27616 70444 27656
rect 70484 27616 70493 27656
rect 70435 27615 70493 27616
rect 70827 27656 70869 27665
rect 70827 27616 70828 27656
rect 70868 27616 70869 27656
rect 70827 27607 70869 27616
rect 71203 27656 71261 27657
rect 71203 27616 71212 27656
rect 71252 27616 71261 27656
rect 71203 27615 71261 27616
rect 71587 27656 71645 27657
rect 71587 27616 71596 27656
rect 71636 27616 71645 27656
rect 71587 27615 71645 27616
rect 71691 27656 71733 27665
rect 71691 27616 71692 27656
rect 71732 27616 71733 27656
rect 71691 27607 71733 27616
rect 75723 27656 75765 27665
rect 75723 27616 75724 27656
rect 75764 27616 75765 27656
rect 75723 27607 75765 27616
rect 75915 27656 75957 27665
rect 75915 27616 75916 27656
rect 75956 27616 75957 27656
rect 75915 27607 75957 27616
rect 76003 27656 76061 27657
rect 76003 27616 76012 27656
rect 76052 27616 76061 27656
rect 76003 27615 76061 27616
rect 76203 27656 76245 27665
rect 76203 27616 76204 27656
rect 76244 27616 76245 27656
rect 76203 27607 76245 27616
rect 76579 27656 76637 27657
rect 76579 27616 76588 27656
rect 76628 27616 76637 27656
rect 76579 27615 76637 27616
rect 76867 27656 76925 27657
rect 76867 27616 76876 27656
rect 76916 27616 76925 27656
rect 76867 27615 76925 27616
rect 77067 27656 77109 27665
rect 77067 27616 77068 27656
rect 77108 27616 77109 27656
rect 77067 27607 77109 27616
rect 77443 27656 77501 27657
rect 77443 27616 77452 27656
rect 77492 27616 77501 27656
rect 77443 27615 77501 27616
rect 78307 27656 78365 27657
rect 78307 27616 78316 27656
rect 78356 27616 78365 27656
rect 78307 27615 78365 27616
rect 52587 27596 52629 27605
rect 40387 27572 40445 27573
rect 40387 27532 40396 27572
rect 40436 27532 40445 27572
rect 40387 27531 40445 27532
rect 44227 27572 44285 27573
rect 44227 27532 44236 27572
rect 44276 27532 44285 27572
rect 44227 27531 44285 27532
rect 45859 27572 45917 27573
rect 45859 27532 45868 27572
rect 45908 27532 45917 27572
rect 45859 27531 45917 27532
rect 52107 27572 52149 27581
rect 52107 27532 52108 27572
rect 52148 27532 52149 27572
rect 52107 27523 52149 27532
rect 52299 27572 52341 27581
rect 52299 27532 52300 27572
rect 52340 27532 52341 27572
rect 52299 27523 52341 27532
rect 58819 27572 58877 27573
rect 58819 27532 58828 27572
rect 58868 27532 58877 27572
rect 58819 27531 58877 27532
rect 59203 27572 59261 27573
rect 59203 27532 59212 27572
rect 59252 27532 59261 27572
rect 59203 27531 59261 27532
rect 59587 27572 59645 27573
rect 59587 27532 59596 27572
rect 59636 27532 59645 27572
rect 59587 27531 59645 27532
rect 59971 27572 60029 27573
rect 59971 27532 59980 27572
rect 60020 27532 60029 27572
rect 59971 27531 60029 27532
rect 60747 27572 60789 27581
rect 60747 27532 60748 27572
rect 60788 27532 60789 27572
rect 60747 27523 60789 27532
rect 60939 27572 60981 27581
rect 60939 27532 60940 27572
rect 60980 27532 60981 27572
rect 60939 27523 60981 27532
rect 68427 27572 68469 27581
rect 68427 27532 68428 27572
rect 68468 27532 68469 27572
rect 68427 27523 68469 27532
rect 76299 27572 76341 27581
rect 76299 27532 76300 27572
rect 76340 27532 76341 27572
rect 76299 27523 76341 27532
rect 76491 27572 76533 27581
rect 76491 27532 76492 27572
rect 76532 27532 76533 27572
rect 76491 27523 76533 27532
rect 42987 27488 43029 27497
rect 42987 27448 42988 27488
rect 43028 27448 43029 27488
rect 42987 27439 43029 27448
rect 43179 27488 43221 27497
rect 43179 27448 43180 27488
rect 43220 27448 43221 27488
rect 43179 27439 43221 27448
rect 43755 27488 43797 27497
rect 43755 27448 43756 27488
rect 43796 27448 43797 27488
rect 43755 27439 43797 27448
rect 52203 27488 52245 27497
rect 52203 27448 52204 27488
rect 52244 27448 52245 27488
rect 52203 27439 52245 27448
rect 52587 27488 52629 27497
rect 52587 27448 52588 27488
rect 52628 27448 52629 27488
rect 52587 27439 52629 27448
rect 60843 27488 60885 27497
rect 60843 27448 60844 27488
rect 60884 27448 60885 27488
rect 60843 27439 60885 27448
rect 65067 27488 65109 27497
rect 65067 27448 65068 27488
rect 65108 27448 65109 27488
rect 65067 27439 65109 27448
rect 76395 27488 76437 27497
rect 76395 27448 76396 27488
rect 76436 27448 76437 27488
rect 76395 27439 76437 27448
rect 40203 27404 40245 27413
rect 40203 27364 40204 27404
rect 40244 27364 40245 27404
rect 40203 27355 40245 27364
rect 40587 27404 40629 27413
rect 40587 27364 40588 27404
rect 40628 27364 40629 27404
rect 40587 27355 40629 27364
rect 43947 27404 43989 27413
rect 43947 27364 43948 27404
rect 43988 27364 43989 27404
rect 43947 27355 43989 27364
rect 44427 27404 44469 27413
rect 44427 27364 44428 27404
rect 44468 27364 44469 27404
rect 44427 27355 44469 27364
rect 46059 27404 46101 27413
rect 46059 27364 46060 27404
rect 46100 27364 46101 27404
rect 46059 27355 46101 27364
rect 51139 27404 51197 27405
rect 51139 27364 51148 27404
rect 51188 27364 51197 27404
rect 51139 27363 51197 27364
rect 55555 27404 55613 27405
rect 55555 27364 55564 27404
rect 55604 27364 55613 27404
rect 55555 27363 55613 27364
rect 58155 27404 58197 27413
rect 58155 27364 58156 27404
rect 58196 27364 58197 27404
rect 58155 27355 58197 27364
rect 59019 27404 59061 27413
rect 59019 27364 59020 27404
rect 59060 27364 59061 27404
rect 59019 27355 59061 27364
rect 59787 27404 59829 27413
rect 59787 27364 59788 27404
rect 59828 27364 59829 27404
rect 59787 27355 59829 27364
rect 60171 27404 60213 27413
rect 60171 27364 60172 27404
rect 60212 27364 60213 27404
rect 60171 27355 60213 27364
rect 61227 27404 61269 27413
rect 61227 27364 61228 27404
rect 61268 27364 61269 27404
rect 61227 27355 61269 27364
rect 64771 27404 64829 27405
rect 64771 27364 64780 27404
rect 64820 27364 64829 27404
rect 64771 27363 64829 27364
rect 66603 27404 66645 27413
rect 66603 27364 66604 27404
rect 66644 27364 66645 27404
rect 66603 27355 66645 27364
rect 71115 27404 71157 27413
rect 71115 27364 71116 27404
rect 71156 27364 71157 27404
rect 71115 27355 71157 27364
rect 71979 27404 72021 27413
rect 71979 27364 71980 27404
rect 72020 27364 72021 27404
rect 71979 27355 72021 27364
rect 75723 27404 75765 27413
rect 75723 27364 75724 27404
rect 75764 27364 75765 27404
rect 75723 27355 75765 27364
rect 76779 27404 76821 27413
rect 76779 27364 76780 27404
rect 76820 27364 76821 27404
rect 76779 27355 76821 27364
rect 79459 27404 79517 27405
rect 79459 27364 79468 27404
rect 79508 27364 79517 27404
rect 79459 27363 79517 27364
rect 576 27236 79584 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 75112 27236
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75480 27196 79584 27236
rect 576 27172 79584 27196
rect 44515 27068 44573 27069
rect 44515 27028 44524 27068
rect 44564 27028 44573 27068
rect 44515 27027 44573 27028
rect 49131 27068 49173 27077
rect 49131 27028 49132 27068
rect 49172 27028 49173 27068
rect 49131 27019 49173 27028
rect 50851 27068 50909 27069
rect 50851 27028 50860 27068
rect 50900 27028 50909 27068
rect 50851 27027 50909 27028
rect 61419 27068 61461 27077
rect 61419 27028 61420 27068
rect 61460 27028 61461 27068
rect 61419 27019 61461 27028
rect 61899 27068 61941 27077
rect 61899 27028 61900 27068
rect 61940 27028 61941 27068
rect 61899 27019 61941 27028
rect 64395 27068 64437 27077
rect 64395 27028 64396 27068
rect 64436 27028 64437 27068
rect 64395 27019 64437 27028
rect 76963 27068 77021 27069
rect 76963 27028 76972 27068
rect 77012 27028 77021 27068
rect 76963 27027 77021 27028
rect 78123 27068 78165 27077
rect 78123 27028 78124 27068
rect 78164 27028 78165 27068
rect 78123 27019 78165 27028
rect 39915 26984 39957 26993
rect 39915 26944 39916 26984
rect 39956 26944 39957 26984
rect 39915 26935 39957 26944
rect 47787 26984 47829 26993
rect 47787 26944 47788 26984
rect 47828 26944 47829 26984
rect 47787 26935 47829 26944
rect 63915 26984 63957 26993
rect 63915 26944 63916 26984
rect 63956 26944 63957 26984
rect 63915 26935 63957 26944
rect 71019 26984 71061 26993
rect 71019 26944 71020 26984
rect 71060 26944 71061 26984
rect 71019 26935 71061 26944
rect 39819 26900 39861 26909
rect 39819 26860 39820 26900
rect 39860 26860 39861 26900
rect 39819 26851 39861 26860
rect 40011 26900 40053 26909
rect 40011 26860 40012 26900
rect 40052 26860 40053 26900
rect 40011 26851 40053 26860
rect 40771 26900 40829 26901
rect 40771 26860 40780 26900
rect 40820 26860 40829 26900
rect 40771 26859 40829 26860
rect 44899 26900 44957 26901
rect 44899 26860 44908 26900
rect 44948 26860 44957 26900
rect 44899 26859 44957 26860
rect 47691 26900 47733 26909
rect 47691 26860 47692 26900
rect 47732 26860 47733 26900
rect 47691 26851 47733 26860
rect 47883 26900 47925 26909
rect 47883 26860 47884 26900
rect 47924 26860 47925 26900
rect 47883 26851 47925 26860
rect 58435 26900 58493 26901
rect 58435 26860 58444 26900
rect 58484 26860 58493 26900
rect 58435 26859 58493 26860
rect 61603 26900 61661 26901
rect 61603 26860 61612 26900
rect 61652 26860 61661 26900
rect 61603 26859 61661 26860
rect 63819 26900 63861 26909
rect 63819 26860 63820 26900
rect 63860 26860 63861 26900
rect 63819 26851 63861 26860
rect 64011 26900 64053 26909
rect 64011 26860 64012 26900
rect 64052 26860 64053 26900
rect 64011 26851 64053 26860
rect 70923 26900 70965 26909
rect 70923 26860 70924 26900
rect 70964 26860 70965 26900
rect 70923 26851 70965 26860
rect 71115 26900 71157 26909
rect 71115 26860 71116 26900
rect 71156 26860 71157 26900
rect 71115 26851 71157 26860
rect 78307 26900 78365 26901
rect 78307 26860 78316 26900
rect 78356 26860 78365 26900
rect 78307 26859 78365 26860
rect 39427 26816 39485 26817
rect 39427 26776 39436 26816
rect 39476 26776 39485 26816
rect 39427 26775 39485 26776
rect 39531 26816 39573 26825
rect 39531 26776 39532 26816
rect 39572 26776 39573 26816
rect 39531 26767 39573 26776
rect 39715 26816 39773 26817
rect 39715 26776 39724 26816
rect 39764 26776 39773 26816
rect 39715 26775 39773 26776
rect 40107 26816 40149 26825
rect 40107 26776 40108 26816
rect 40148 26776 40149 26816
rect 40395 26816 40437 26825
rect 40107 26767 40149 26776
rect 40299 26795 40341 26804
rect 40299 26755 40300 26795
rect 40340 26755 40341 26795
rect 40395 26776 40396 26816
rect 40436 26776 40437 26816
rect 40395 26767 40437 26776
rect 40491 26816 40533 26825
rect 40491 26776 40492 26816
rect 40532 26776 40533 26816
rect 40491 26767 40533 26776
rect 42499 26816 42557 26817
rect 42499 26776 42508 26816
rect 42548 26776 42557 26816
rect 42499 26775 42557 26776
rect 43363 26816 43421 26817
rect 43363 26776 43372 26816
rect 43412 26776 43421 26816
rect 43363 26775 43421 26776
rect 47115 26816 47157 26825
rect 47115 26776 47116 26816
rect 47156 26776 47157 26816
rect 47115 26767 47157 26776
rect 47307 26816 47349 26825
rect 47307 26776 47308 26816
rect 47348 26776 47349 26816
rect 47307 26767 47349 26776
rect 47395 26816 47453 26817
rect 47395 26776 47404 26816
rect 47444 26776 47453 26816
rect 47395 26775 47453 26776
rect 47595 26816 47637 26825
rect 47595 26776 47596 26816
rect 47636 26776 47637 26816
rect 47595 26767 47637 26776
rect 47971 26816 48029 26817
rect 47971 26776 47980 26816
rect 48020 26776 48029 26816
rect 47971 26775 48029 26776
rect 48171 26816 48213 26825
rect 48171 26776 48172 26816
rect 48212 26776 48213 26816
rect 48171 26767 48213 26776
rect 48267 26816 48309 26825
rect 48267 26776 48268 26816
rect 48308 26776 48309 26816
rect 48267 26767 48309 26776
rect 48363 26816 48405 26825
rect 48363 26776 48364 26816
rect 48404 26776 48405 26816
rect 48363 26767 48405 26776
rect 48459 26816 48501 26825
rect 48459 26776 48460 26816
rect 48500 26776 48501 26816
rect 48459 26767 48501 26776
rect 49027 26816 49085 26817
rect 49027 26776 49036 26816
rect 49076 26776 49085 26816
rect 49027 26775 49085 26776
rect 52003 26816 52061 26817
rect 52003 26776 52012 26816
rect 52052 26776 52061 26816
rect 52003 26775 52061 26776
rect 52867 26816 52925 26817
rect 52867 26776 52876 26816
rect 52916 26776 52925 26816
rect 52867 26775 52925 26776
rect 53451 26816 53493 26825
rect 53451 26776 53452 26816
rect 53492 26776 53493 26816
rect 53451 26767 53493 26776
rect 53547 26816 53589 26825
rect 53547 26776 53548 26816
rect 53588 26776 53589 26816
rect 53547 26767 53589 26776
rect 53643 26816 53685 26825
rect 53643 26776 53644 26816
rect 53684 26776 53685 26816
rect 53643 26767 53685 26776
rect 53739 26816 53781 26825
rect 53739 26776 53740 26816
rect 53780 26776 53781 26816
rect 53739 26767 53781 26776
rect 55171 26816 55229 26817
rect 55171 26776 55180 26816
rect 55220 26776 55229 26816
rect 55171 26775 55229 26776
rect 56035 26816 56093 26817
rect 56035 26776 56044 26816
rect 56084 26776 56093 26816
rect 56035 26775 56093 26776
rect 59971 26816 60029 26817
rect 59971 26776 59980 26816
rect 60020 26776 60029 26816
rect 59971 26775 60029 26776
rect 60835 26816 60893 26817
rect 60835 26776 60844 26816
rect 60884 26776 60893 26816
rect 60835 26775 60893 26776
rect 61227 26816 61269 26825
rect 61227 26776 61228 26816
rect 61268 26776 61269 26816
rect 61227 26767 61269 26776
rect 61795 26816 61853 26817
rect 61795 26776 61804 26816
rect 61844 26776 61853 26816
rect 61795 26775 61853 26776
rect 63715 26816 63773 26817
rect 63715 26776 63724 26816
rect 63764 26776 63773 26816
rect 63715 26775 63773 26776
rect 64107 26816 64149 26825
rect 64107 26776 64108 26816
rect 64148 26776 64149 26816
rect 64107 26767 64149 26776
rect 64395 26816 64437 26825
rect 64395 26776 64396 26816
rect 64436 26776 64437 26816
rect 64395 26767 64437 26776
rect 64587 26816 64629 26825
rect 64587 26776 64588 26816
rect 64628 26776 64629 26816
rect 64587 26767 64629 26776
rect 64675 26816 64733 26817
rect 64675 26776 64684 26816
rect 64724 26776 64733 26816
rect 64675 26775 64733 26776
rect 64867 26816 64925 26817
rect 64867 26776 64876 26816
rect 64916 26776 64925 26816
rect 64867 26775 64925 26776
rect 64971 26816 65013 26825
rect 64971 26776 64972 26816
rect 65012 26776 65013 26816
rect 64971 26767 65013 26776
rect 69187 26816 69245 26817
rect 69187 26776 69196 26816
rect 69236 26776 69245 26816
rect 69187 26775 69245 26776
rect 70051 26816 70109 26817
rect 70051 26776 70060 26816
rect 70100 26776 70109 26816
rect 70051 26775 70109 26776
rect 70827 26816 70869 26825
rect 70827 26776 70828 26816
rect 70868 26776 70869 26816
rect 70827 26767 70869 26776
rect 71203 26816 71261 26817
rect 71203 26776 71212 26816
rect 71252 26776 71261 26816
rect 71203 26775 71261 26776
rect 71395 26816 71453 26817
rect 71395 26776 71404 26816
rect 71444 26776 71453 26816
rect 71395 26775 71453 26776
rect 71499 26816 71541 26825
rect 71499 26776 71500 26816
rect 71540 26776 71541 26816
rect 71499 26767 71541 26776
rect 71691 26816 71733 26825
rect 71691 26776 71692 26816
rect 71732 26776 71733 26816
rect 71691 26767 71733 26776
rect 72355 26816 72413 26817
rect 72355 26776 72364 26816
rect 72404 26776 72413 26816
rect 72355 26775 72413 26776
rect 73219 26816 73277 26817
rect 73219 26776 73228 26816
rect 73268 26776 73277 26816
rect 73219 26775 73277 26776
rect 74947 26816 75005 26817
rect 74947 26776 74956 26816
rect 74996 26776 75005 26816
rect 74947 26775 75005 26776
rect 75811 26816 75869 26817
rect 75811 26776 75820 26816
rect 75860 26776 75869 26816
rect 75811 26775 75869 26776
rect 77163 26816 77205 26825
rect 77163 26776 77164 26816
rect 77204 26776 77205 26816
rect 77163 26767 77205 26776
rect 77259 26816 77301 26825
rect 77259 26776 77260 26816
rect 77300 26776 77301 26816
rect 77259 26767 77301 26776
rect 77355 26816 77397 26825
rect 77355 26776 77356 26816
rect 77396 26776 77397 26816
rect 77355 26767 77397 26776
rect 77451 26816 77493 26825
rect 77451 26776 77452 26816
rect 77492 26776 77493 26816
rect 77451 26767 77493 26776
rect 77643 26816 77685 26825
rect 77643 26776 77644 26816
rect 77684 26776 77685 26816
rect 77643 26767 77685 26776
rect 77739 26816 77781 26825
rect 77739 26776 77740 26816
rect 77780 26776 77781 26816
rect 77739 26767 77781 26776
rect 77835 26816 77877 26825
rect 77835 26776 77836 26816
rect 77876 26776 77877 26816
rect 77835 26767 77877 26776
rect 77931 26816 77973 26825
rect 77931 26776 77932 26816
rect 77972 26776 77973 26816
rect 77931 26767 77973 26776
rect 78595 26816 78653 26817
rect 78595 26776 78604 26816
rect 78644 26776 78653 26816
rect 78595 26775 78653 26776
rect 40299 26746 40341 26755
rect 42123 26732 42165 26741
rect 42123 26692 42124 26732
rect 42164 26692 42165 26732
rect 42123 26683 42165 26692
rect 47211 26732 47253 26741
rect 47211 26692 47212 26732
rect 47252 26692 47253 26732
rect 47211 26683 47253 26692
rect 53259 26732 53301 26741
rect 53259 26692 53260 26732
rect 53300 26692 53301 26732
rect 53259 26683 53301 26692
rect 56427 26732 56469 26741
rect 56427 26692 56428 26732
rect 56468 26692 56469 26732
rect 56427 26683 56469 26692
rect 70443 26732 70485 26741
rect 70443 26692 70444 26732
rect 70484 26692 70485 26732
rect 70443 26683 70485 26692
rect 71979 26732 72021 26741
rect 71979 26692 71980 26732
rect 72020 26692 72021 26732
rect 71979 26683 72021 26692
rect 74571 26732 74613 26741
rect 74571 26692 74572 26732
rect 74612 26692 74613 26732
rect 74571 26683 74613 26692
rect 40579 26648 40637 26649
rect 40579 26608 40588 26648
rect 40628 26608 40637 26648
rect 40579 26607 40637 26608
rect 40971 26648 41013 26657
rect 40971 26608 40972 26648
rect 41012 26608 41013 26648
rect 40971 26599 41013 26608
rect 44715 26648 44757 26657
rect 44715 26608 44716 26648
rect 44756 26608 44757 26648
rect 44715 26599 44757 26608
rect 49131 26648 49173 26657
rect 49131 26608 49132 26648
rect 49172 26608 49173 26648
rect 49131 26599 49173 26608
rect 54019 26648 54077 26649
rect 54019 26608 54028 26648
rect 54068 26608 54077 26648
rect 54019 26607 54077 26608
rect 58635 26648 58677 26657
rect 58635 26608 58636 26648
rect 58676 26608 58677 26648
rect 58635 26599 58677 26608
rect 58819 26648 58877 26649
rect 58819 26608 58828 26648
rect 58868 26608 58877 26648
rect 58819 26607 58877 26608
rect 61899 26648 61941 26657
rect 61899 26608 61900 26648
rect 61940 26608 61941 26648
rect 61899 26599 61941 26608
rect 68035 26648 68093 26649
rect 68035 26608 68044 26648
rect 68084 26608 68093 26648
rect 68035 26607 68093 26608
rect 71587 26648 71645 26649
rect 71587 26608 71596 26648
rect 71636 26608 71645 26648
rect 71587 26607 71645 26608
rect 74371 26648 74429 26649
rect 74371 26608 74380 26648
rect 74420 26608 74429 26648
rect 74371 26607 74429 26608
rect 78507 26648 78549 26657
rect 78507 26608 78508 26648
rect 78548 26608 78549 26648
rect 78507 26599 78549 26608
rect 576 26480 79584 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 76352 26480
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76720 26440 79584 26480
rect 576 26416 79584 26440
rect 61419 26370 61461 26379
rect 61419 26330 61420 26370
rect 61460 26330 61461 26370
rect 843 26312 885 26321
rect 44139 26316 44181 26325
rect 61419 26321 61461 26330
rect 843 26272 844 26312
rect 884 26272 885 26312
rect 843 26263 885 26272
rect 42403 26312 42461 26313
rect 42403 26272 42412 26312
rect 42452 26272 42461 26312
rect 42403 26271 42461 26272
rect 44139 26276 44140 26316
rect 44180 26276 44181 26316
rect 44139 26267 44181 26276
rect 54603 26312 54645 26321
rect 54603 26272 54604 26312
rect 54644 26272 54645 26312
rect 54603 26263 54645 26272
rect 69963 26312 70005 26321
rect 69963 26272 69964 26312
rect 70004 26272 70005 26312
rect 69963 26263 70005 26272
rect 71211 26312 71253 26321
rect 76683 26316 76725 26325
rect 71211 26272 71212 26312
rect 71252 26272 71253 26312
rect 71211 26263 71253 26272
rect 71779 26312 71837 26313
rect 71779 26272 71788 26312
rect 71828 26272 71837 26312
rect 71779 26271 71837 26272
rect 72643 26312 72701 26313
rect 72643 26272 72652 26312
rect 72692 26272 72701 26312
rect 72643 26271 72701 26272
rect 76683 26276 76684 26316
rect 76724 26276 76725 26316
rect 76683 26267 76725 26276
rect 39339 26228 39381 26237
rect 39339 26188 39340 26228
rect 39380 26188 39381 26228
rect 39339 26179 39381 26188
rect 43083 26228 43125 26237
rect 43083 26188 43084 26228
rect 43124 26188 43125 26228
rect 47787 26228 47829 26237
rect 43083 26179 43125 26188
rect 43179 26186 43221 26195
rect 38083 26144 38141 26145
rect 38083 26104 38092 26144
rect 38132 26104 38141 26144
rect 38083 26103 38141 26104
rect 38947 26144 39005 26145
rect 38947 26104 38956 26144
rect 38996 26104 39005 26144
rect 38947 26103 39005 26104
rect 39531 26144 39573 26153
rect 39531 26104 39532 26144
rect 39572 26104 39573 26144
rect 39531 26095 39573 26104
rect 39627 26144 39669 26153
rect 39627 26104 39628 26144
rect 39668 26104 39669 26144
rect 39627 26095 39669 26104
rect 39723 26144 39765 26153
rect 39723 26104 39724 26144
rect 39764 26104 39765 26144
rect 39723 26095 39765 26104
rect 39819 26144 39861 26153
rect 39819 26104 39820 26144
rect 39860 26104 39861 26144
rect 39819 26095 39861 26104
rect 40011 26144 40053 26153
rect 40011 26104 40012 26144
rect 40052 26104 40053 26144
rect 40011 26095 40053 26104
rect 40387 26144 40445 26145
rect 40387 26104 40396 26144
rect 40436 26104 40445 26144
rect 40387 26103 40445 26104
rect 41251 26144 41309 26145
rect 41251 26104 41260 26144
rect 41300 26104 41309 26144
rect 41251 26103 41309 26104
rect 42987 26144 43029 26153
rect 42987 26104 42988 26144
rect 43028 26104 43029 26144
rect 43179 26146 43180 26186
rect 43220 26146 43221 26186
rect 47787 26188 47788 26228
rect 47828 26188 47829 26228
rect 47787 26179 47829 26188
rect 59115 26228 59157 26237
rect 59115 26188 59116 26228
rect 59156 26188 59157 26228
rect 59115 26179 59157 26188
rect 70539 26186 70581 26195
rect 43179 26137 43221 26146
rect 43267 26144 43325 26145
rect 42987 26095 43029 26104
rect 43267 26104 43276 26144
rect 43316 26104 43325 26144
rect 43267 26103 43325 26104
rect 43467 26144 43509 26153
rect 43467 26104 43468 26144
rect 43508 26104 43509 26144
rect 43467 26095 43509 26104
rect 43843 26144 43901 26145
rect 43843 26104 43852 26144
rect 43892 26104 43901 26144
rect 43843 26103 43901 26104
rect 44227 26144 44285 26145
rect 44227 26104 44236 26144
rect 44276 26104 44285 26144
rect 44227 26103 44285 26104
rect 44331 26144 44373 26153
rect 44331 26104 44332 26144
rect 44372 26104 44373 26144
rect 44331 26095 44373 26104
rect 44811 26144 44853 26153
rect 44811 26104 44812 26144
rect 44852 26104 44853 26144
rect 44811 26095 44853 26104
rect 45187 26144 45245 26145
rect 45187 26104 45196 26144
rect 45236 26104 45245 26144
rect 45187 26103 45245 26104
rect 46051 26144 46109 26145
rect 46051 26104 46060 26144
rect 46100 26104 46109 26144
rect 46051 26103 46109 26104
rect 48163 26144 48221 26145
rect 48163 26104 48172 26144
rect 48212 26104 48221 26144
rect 48163 26103 48221 26104
rect 49027 26144 49085 26145
rect 49027 26104 49036 26144
rect 49076 26104 49085 26144
rect 49027 26103 49085 26104
rect 53155 26144 53213 26145
rect 53155 26104 53164 26144
rect 53204 26104 53213 26144
rect 53155 26103 53213 26104
rect 53347 26144 53405 26145
rect 53347 26104 53356 26144
rect 53396 26104 53405 26144
rect 53347 26103 53405 26104
rect 53451 26144 53493 26153
rect 53451 26104 53452 26144
rect 53492 26104 53493 26144
rect 53451 26095 53493 26104
rect 53635 26144 53693 26145
rect 53635 26104 53644 26144
rect 53684 26104 53693 26144
rect 53635 26103 53693 26104
rect 54027 26144 54069 26153
rect 54027 26104 54028 26144
rect 54068 26104 54069 26144
rect 54027 26095 54069 26104
rect 54795 26144 54837 26153
rect 54795 26104 54796 26144
rect 54836 26104 54837 26144
rect 54795 26095 54837 26104
rect 54987 26144 55029 26153
rect 54987 26104 54988 26144
rect 55028 26104 55029 26144
rect 54987 26095 55029 26104
rect 55075 26144 55133 26145
rect 55075 26104 55084 26144
rect 55124 26104 55133 26144
rect 55075 26103 55133 26104
rect 55843 26144 55901 26145
rect 55843 26104 55852 26144
rect 55892 26104 55901 26144
rect 55843 26103 55901 26104
rect 56131 26144 56189 26145
rect 56131 26104 56140 26144
rect 56180 26104 56189 26144
rect 56131 26103 56189 26104
rect 56523 26144 56565 26153
rect 56523 26104 56524 26144
rect 56564 26104 56565 26144
rect 56523 26095 56565 26104
rect 57859 26144 57917 26145
rect 57859 26104 57868 26144
rect 57908 26104 57917 26144
rect 57859 26103 57917 26104
rect 58723 26144 58781 26145
rect 58723 26104 58732 26144
rect 58772 26104 58781 26144
rect 58723 26103 58781 26104
rect 59299 26144 59357 26145
rect 59299 26104 59308 26144
rect 59348 26104 59357 26144
rect 59299 26103 59357 26104
rect 59691 26144 59733 26153
rect 59691 26104 59692 26144
rect 59732 26104 59733 26144
rect 59691 26095 59733 26104
rect 59979 26144 60021 26153
rect 59979 26104 59980 26144
rect 60020 26104 60021 26144
rect 59979 26095 60021 26104
rect 60171 26144 60213 26153
rect 60171 26104 60172 26144
rect 60212 26104 60213 26144
rect 60171 26095 60213 26104
rect 60259 26144 60317 26145
rect 60259 26104 60268 26144
rect 60308 26104 60317 26144
rect 60259 26103 60317 26104
rect 61227 26144 61269 26153
rect 61227 26104 61228 26144
rect 61268 26104 61269 26144
rect 61227 26095 61269 26104
rect 61315 26144 61373 26145
rect 61315 26104 61324 26144
rect 61364 26104 61373 26144
rect 61315 26103 61373 26104
rect 61707 26144 61749 26153
rect 61707 26104 61708 26144
rect 61748 26104 61749 26144
rect 61707 26095 61749 26104
rect 61803 26144 61845 26153
rect 61803 26104 61804 26144
rect 61844 26104 61845 26144
rect 61803 26095 61845 26104
rect 61899 26144 61941 26153
rect 61899 26104 61900 26144
rect 61940 26104 61941 26144
rect 61899 26095 61941 26104
rect 61995 26144 62037 26153
rect 61995 26104 61996 26144
rect 62036 26104 62037 26144
rect 61995 26095 62037 26104
rect 64387 26144 64445 26145
rect 64387 26104 64396 26144
rect 64436 26104 64445 26144
rect 64387 26103 64445 26104
rect 65251 26144 65309 26145
rect 65251 26104 65260 26144
rect 65300 26104 65309 26144
rect 65251 26103 65309 26104
rect 65643 26144 65685 26153
rect 65643 26104 65644 26144
rect 65684 26104 65685 26144
rect 65643 26095 65685 26104
rect 66123 26144 66165 26153
rect 66123 26104 66124 26144
rect 66164 26104 66165 26144
rect 66123 26095 66165 26104
rect 66499 26144 66557 26145
rect 66499 26104 66508 26144
rect 66548 26104 66557 26144
rect 66499 26103 66557 26104
rect 67363 26144 67421 26145
rect 67363 26104 67372 26144
rect 67412 26104 67421 26144
rect 67363 26103 67421 26104
rect 68803 26144 68861 26145
rect 68803 26104 68812 26144
rect 68852 26104 68861 26144
rect 68803 26103 68861 26104
rect 69195 26144 69237 26153
rect 69195 26104 69196 26144
rect 69236 26104 69237 26144
rect 69195 26095 69237 26104
rect 69483 26144 69525 26153
rect 69483 26104 69484 26144
rect 69524 26104 69525 26144
rect 69483 26095 69525 26104
rect 69675 26144 69717 26153
rect 70539 26146 70540 26186
rect 70580 26146 70581 26186
rect 69675 26104 69676 26144
rect 69716 26104 69717 26144
rect 69675 26095 69717 26104
rect 69763 26144 69821 26145
rect 69763 26104 69772 26144
rect 69812 26104 69821 26144
rect 70539 26137 70581 26146
rect 70915 26144 70973 26145
rect 69763 26103 69821 26104
rect 70915 26104 70924 26144
rect 70964 26104 70973 26144
rect 70915 26103 70973 26104
rect 71107 26144 71165 26145
rect 71107 26104 71116 26144
rect 71156 26104 71165 26144
rect 71107 26103 71165 26104
rect 71883 26144 71925 26153
rect 71883 26104 71884 26144
rect 71924 26104 71925 26144
rect 71883 26095 71925 26104
rect 71979 26144 72021 26153
rect 71979 26104 71980 26144
rect 72020 26104 72021 26144
rect 71979 26095 72021 26104
rect 72075 26144 72117 26153
rect 72075 26104 72076 26144
rect 72116 26104 72117 26144
rect 72075 26095 72117 26104
rect 72747 26144 72789 26153
rect 72747 26104 72748 26144
rect 72788 26104 72789 26144
rect 72747 26095 72789 26104
rect 72843 26144 72885 26153
rect 72843 26104 72844 26144
rect 72884 26104 72885 26144
rect 72843 26095 72885 26104
rect 72939 26144 72981 26153
rect 72939 26104 72940 26144
rect 72980 26104 72981 26144
rect 72939 26095 72981 26104
rect 73315 26144 73373 26145
rect 73315 26104 73324 26144
rect 73364 26104 73373 26144
rect 73315 26103 73373 26104
rect 75627 26144 75669 26153
rect 75627 26104 75628 26144
rect 75668 26104 75669 26144
rect 75627 26095 75669 26104
rect 76003 26144 76061 26145
rect 76003 26104 76012 26144
rect 76052 26104 76061 26144
rect 76003 26103 76061 26104
rect 76491 26144 76533 26153
rect 76491 26104 76492 26144
rect 76532 26104 76533 26144
rect 76491 26095 76533 26104
rect 76579 26144 76637 26145
rect 76579 26104 76588 26144
rect 76628 26104 76637 26144
rect 76579 26103 76637 26104
rect 76875 26144 76917 26153
rect 76875 26104 76876 26144
rect 76916 26104 76917 26144
rect 76875 26095 76917 26104
rect 77251 26144 77309 26145
rect 77251 26104 77260 26144
rect 77300 26104 77309 26144
rect 77251 26103 77309 26104
rect 78115 26144 78173 26145
rect 78115 26104 78124 26144
rect 78164 26104 78173 26144
rect 78115 26103 78173 26104
rect 643 26060 701 26061
rect 643 26020 652 26060
rect 692 26020 701 26060
rect 643 26019 701 26020
rect 42787 26060 42845 26061
rect 42787 26020 42796 26060
rect 42836 26020 42845 26060
rect 42787 26019 42845 26020
rect 43563 26060 43605 26069
rect 43563 26020 43564 26060
rect 43604 26020 43605 26060
rect 43563 26011 43605 26020
rect 43755 26060 43797 26069
rect 43755 26020 43756 26060
rect 43796 26020 43797 26060
rect 43755 26011 43797 26020
rect 53739 26060 53781 26069
rect 53739 26020 53740 26060
rect 53780 26020 53781 26060
rect 53739 26011 53781 26020
rect 53931 26060 53973 26069
rect 53931 26020 53932 26060
rect 53972 26020 53973 26060
rect 53931 26011 53973 26020
rect 54403 26060 54461 26061
rect 54403 26020 54412 26060
rect 54452 26020 54461 26060
rect 54403 26019 54461 26020
rect 56235 26060 56277 26069
rect 56235 26020 56236 26060
rect 56276 26020 56277 26060
rect 56235 26011 56277 26020
rect 56427 26060 56469 26069
rect 56427 26020 56428 26060
rect 56468 26020 56469 26060
rect 56427 26011 56469 26020
rect 59403 26060 59445 26069
rect 59403 26020 59404 26060
rect 59444 26020 59445 26060
rect 59403 26011 59445 26020
rect 59595 26060 59637 26069
rect 59595 26020 59596 26060
rect 59636 26020 59637 26060
rect 59595 26011 59637 26020
rect 60451 26060 60509 26061
rect 60451 26020 60460 26060
rect 60500 26020 60509 26060
rect 60451 26019 60509 26020
rect 68907 26060 68949 26069
rect 68907 26020 68908 26060
rect 68948 26020 68949 26060
rect 68907 26011 68949 26020
rect 69099 26060 69141 26069
rect 69099 26020 69100 26060
rect 69140 26020 69141 26060
rect 69099 26011 69141 26020
rect 70147 26060 70205 26061
rect 70147 26020 70156 26060
rect 70196 26020 70205 26060
rect 70147 26019 70205 26020
rect 70635 26060 70677 26069
rect 70635 26020 70636 26060
rect 70676 26020 70677 26060
rect 70635 26011 70677 26020
rect 70827 26060 70869 26069
rect 70827 26020 70828 26060
rect 70868 26020 70869 26060
rect 70827 26011 70869 26020
rect 75235 26060 75293 26061
rect 75235 26020 75244 26060
rect 75284 26020 75293 26060
rect 75235 26019 75293 26020
rect 75723 26060 75765 26069
rect 75723 26020 75724 26060
rect 75764 26020 75765 26060
rect 75723 26011 75765 26020
rect 75915 26060 75957 26069
rect 75915 26020 75916 26060
rect 75956 26020 75957 26060
rect 75915 26011 75957 26020
rect 36931 25976 36989 25977
rect 36931 25936 36940 25976
rect 36980 25936 36989 25976
rect 36931 25935 36989 25936
rect 43659 25976 43701 25985
rect 43659 25936 43660 25976
rect 43700 25936 43701 25976
rect 43659 25927 43701 25936
rect 47203 25976 47261 25977
rect 47203 25936 47212 25976
rect 47252 25936 47261 25976
rect 47203 25935 47261 25936
rect 53835 25976 53877 25985
rect 53835 25936 53836 25976
rect 53876 25936 53877 25976
rect 53835 25927 53877 25936
rect 54795 25976 54837 25985
rect 54795 25936 54796 25976
rect 54836 25936 54837 25976
rect 54795 25927 54837 25936
rect 55947 25976 55989 25985
rect 55947 25936 55948 25976
rect 55988 25936 55989 25976
rect 55947 25927 55989 25936
rect 56331 25976 56373 25985
rect 56331 25936 56332 25976
rect 56372 25936 56373 25976
rect 56331 25927 56373 25936
rect 59499 25976 59541 25985
rect 59499 25936 59500 25976
rect 59540 25936 59541 25976
rect 59499 25927 59541 25936
rect 59979 25976 60021 25985
rect 59979 25936 59980 25976
rect 60020 25936 60021 25976
rect 59979 25927 60021 25936
rect 60651 25976 60693 25985
rect 60651 25936 60652 25976
rect 60692 25936 60693 25976
rect 60651 25927 60693 25936
rect 60939 25976 60981 25985
rect 60939 25936 60940 25976
rect 60980 25936 60981 25976
rect 60939 25927 60981 25936
rect 63235 25976 63293 25977
rect 63235 25936 63244 25976
rect 63284 25936 63293 25976
rect 63235 25935 63293 25936
rect 69003 25976 69045 25985
rect 69003 25936 69004 25976
rect 69044 25936 69045 25976
rect 69003 25927 69045 25936
rect 69483 25976 69525 25985
rect 69483 25936 69484 25976
rect 69524 25936 69525 25976
rect 69483 25927 69525 25936
rect 70731 25976 70773 25985
rect 70731 25936 70732 25976
rect 70772 25936 70773 25976
rect 70731 25927 70773 25936
rect 73419 25976 73461 25985
rect 73419 25936 73420 25976
rect 73460 25936 73461 25976
rect 73419 25927 73461 25936
rect 75435 25976 75477 25985
rect 75435 25936 75436 25976
rect 75476 25936 75477 25976
rect 75435 25927 75477 25936
rect 75819 25976 75861 25985
rect 75819 25936 75820 25976
rect 75860 25936 75861 25976
rect 75819 25927 75861 25936
rect 76203 25976 76245 25985
rect 76203 25936 76204 25976
rect 76244 25936 76245 25976
rect 76203 25927 76245 25936
rect 42603 25892 42645 25901
rect 42603 25852 42604 25892
rect 42644 25852 42645 25892
rect 42603 25843 42645 25852
rect 44619 25892 44661 25901
rect 44619 25852 44620 25892
rect 44660 25852 44661 25892
rect 44619 25843 44661 25852
rect 50179 25892 50237 25893
rect 50179 25852 50188 25892
rect 50228 25852 50237 25892
rect 50179 25851 50237 25852
rect 53067 25892 53109 25901
rect 53067 25852 53068 25892
rect 53108 25852 53109 25892
rect 53067 25843 53109 25852
rect 54603 25892 54645 25901
rect 54603 25852 54604 25892
rect 54644 25852 54645 25892
rect 54603 25843 54645 25852
rect 56707 25892 56765 25893
rect 56707 25852 56716 25892
rect 56756 25852 56765 25892
rect 56707 25851 56765 25852
rect 68515 25892 68573 25893
rect 68515 25852 68524 25892
rect 68564 25852 68573 25892
rect 68515 25851 68573 25852
rect 79267 25892 79325 25893
rect 79267 25852 79276 25892
rect 79316 25852 79325 25892
rect 79267 25851 79325 25852
rect 576 25724 79584 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 75112 25724
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75480 25684 79584 25724
rect 576 25660 79584 25684
rect 39723 25556 39765 25565
rect 39723 25516 39724 25556
rect 39764 25516 39765 25556
rect 39723 25507 39765 25516
rect 40779 25556 40821 25565
rect 40779 25516 40780 25556
rect 40820 25516 40821 25556
rect 40779 25507 40821 25516
rect 41931 25556 41973 25565
rect 41931 25516 41932 25556
rect 41972 25516 41973 25556
rect 41931 25507 41973 25516
rect 42315 25556 42357 25565
rect 42315 25516 42316 25556
rect 42356 25516 42357 25556
rect 42315 25507 42357 25516
rect 49131 25556 49173 25565
rect 49131 25516 49132 25556
rect 49172 25516 49173 25556
rect 49131 25507 49173 25516
rect 50763 25556 50805 25565
rect 50763 25516 50764 25556
rect 50804 25516 50805 25556
rect 50763 25507 50805 25516
rect 52299 25556 52341 25565
rect 52299 25516 52300 25556
rect 52340 25516 52341 25556
rect 52299 25507 52341 25516
rect 54123 25556 54165 25565
rect 54123 25516 54124 25556
rect 54164 25516 54165 25556
rect 54123 25507 54165 25516
rect 57003 25556 57045 25565
rect 57003 25516 57004 25556
rect 57044 25516 57045 25556
rect 57003 25507 57045 25516
rect 57483 25556 57525 25565
rect 57483 25516 57484 25556
rect 57524 25516 57525 25556
rect 57483 25507 57525 25516
rect 60363 25556 60405 25565
rect 60363 25516 60364 25556
rect 60404 25516 60405 25556
rect 60363 25507 60405 25516
rect 60555 25556 60597 25565
rect 60555 25516 60556 25556
rect 60596 25516 60597 25556
rect 60555 25507 60597 25516
rect 64587 25556 64629 25565
rect 64587 25516 64588 25556
rect 64628 25516 64629 25556
rect 64587 25507 64629 25516
rect 68715 25556 68757 25565
rect 68715 25516 68716 25556
rect 68756 25516 68757 25556
rect 68715 25507 68757 25516
rect 70251 25556 70293 25565
rect 70251 25516 70252 25556
rect 70292 25516 70293 25556
rect 70251 25507 70293 25516
rect 76107 25556 76149 25565
rect 76107 25516 76108 25556
rect 76148 25516 76149 25556
rect 76107 25507 76149 25516
rect 43275 25472 43317 25481
rect 43275 25432 43276 25472
rect 43316 25432 43317 25472
rect 43275 25423 43317 25432
rect 43659 25472 43701 25481
rect 43659 25432 43660 25472
rect 43700 25432 43701 25472
rect 43659 25423 43701 25432
rect 47787 25472 47829 25481
rect 47787 25432 47788 25472
rect 47828 25432 47829 25472
rect 47787 25423 47829 25432
rect 58923 25472 58965 25481
rect 58923 25432 58924 25472
rect 58964 25432 58965 25472
rect 58923 25423 58965 25432
rect 59115 25472 59157 25481
rect 59115 25432 59116 25472
rect 59156 25432 59157 25472
rect 59115 25423 59157 25432
rect 63723 25472 63765 25481
rect 63723 25432 63724 25472
rect 63764 25432 63765 25472
rect 63723 25423 63765 25432
rect 65931 25472 65973 25481
rect 65931 25432 65932 25472
rect 65972 25432 65973 25472
rect 65931 25423 65973 25432
rect 66315 25472 66357 25481
rect 66315 25432 66316 25472
rect 66356 25432 66357 25472
rect 66315 25423 66357 25432
rect 67179 25472 67221 25481
rect 67179 25432 67180 25472
rect 67220 25432 67221 25472
rect 67179 25423 67221 25432
rect 69003 25472 69045 25481
rect 69003 25432 69004 25472
rect 69044 25432 69045 25472
rect 69003 25423 69045 25432
rect 71499 25472 71541 25481
rect 71499 25432 71500 25472
rect 71540 25432 71541 25472
rect 71499 25423 71541 25432
rect 643 25388 701 25389
rect 643 25348 652 25388
rect 692 25348 701 25388
rect 643 25347 701 25348
rect 39523 25388 39581 25389
rect 39523 25348 39532 25388
rect 39572 25348 39581 25388
rect 39523 25347 39581 25348
rect 40579 25388 40637 25389
rect 40579 25348 40588 25388
rect 40628 25348 40637 25388
rect 40579 25347 40637 25348
rect 41731 25388 41789 25389
rect 41731 25348 41740 25388
rect 41780 25348 41789 25388
rect 41731 25347 41789 25348
rect 42115 25388 42173 25389
rect 42115 25348 42124 25388
rect 42164 25348 42173 25388
rect 42115 25347 42173 25348
rect 42499 25388 42557 25389
rect 42499 25348 42508 25388
rect 42548 25348 42557 25388
rect 42499 25347 42557 25348
rect 43075 25388 43133 25389
rect 43075 25348 43084 25388
rect 43124 25348 43133 25388
rect 43075 25347 43133 25348
rect 43459 25388 43517 25389
rect 43459 25348 43468 25388
rect 43508 25348 43517 25388
rect 43459 25347 43517 25348
rect 43843 25388 43901 25389
rect 43843 25348 43852 25388
rect 43892 25348 43901 25388
rect 43843 25347 43901 25348
rect 50563 25388 50621 25389
rect 50563 25348 50572 25388
rect 50612 25348 50621 25388
rect 50563 25347 50621 25348
rect 51235 25388 51293 25389
rect 51235 25348 51244 25388
rect 51284 25348 51293 25388
rect 51235 25347 51293 25348
rect 52099 25388 52157 25389
rect 52099 25348 52108 25388
rect 52148 25348 52157 25388
rect 52099 25347 52157 25348
rect 58723 25388 58781 25389
rect 58723 25348 58732 25388
rect 58772 25348 58781 25388
rect 58723 25347 58781 25348
rect 59971 25388 60029 25389
rect 59971 25348 59980 25388
rect 60020 25348 60029 25388
rect 59971 25347 60029 25348
rect 60163 25388 60221 25389
rect 60163 25348 60172 25388
rect 60212 25348 60221 25388
rect 60163 25347 60221 25348
rect 60739 25388 60797 25389
rect 60739 25348 60748 25388
rect 60788 25348 60797 25388
rect 60739 25347 60797 25348
rect 65835 25388 65877 25397
rect 65835 25348 65836 25388
rect 65876 25348 65877 25388
rect 65835 25339 65877 25348
rect 66027 25388 66069 25397
rect 66027 25348 66028 25388
rect 66068 25348 66069 25388
rect 66027 25339 66069 25348
rect 69859 25388 69917 25389
rect 69859 25348 69868 25388
rect 69908 25348 69917 25388
rect 69859 25347 69917 25348
rect 70051 25388 70109 25389
rect 70051 25348 70060 25388
rect 70100 25348 70109 25388
rect 70051 25347 70109 25348
rect 37699 25304 37757 25305
rect 37699 25264 37708 25304
rect 37748 25264 37757 25304
rect 37699 25263 37757 25264
rect 38379 25304 38421 25313
rect 38379 25264 38380 25304
rect 38420 25264 38421 25304
rect 38379 25255 38421 25264
rect 38571 25304 38613 25313
rect 38571 25264 38572 25304
rect 38612 25264 38613 25304
rect 38571 25255 38613 25264
rect 38659 25304 38717 25305
rect 38659 25264 38668 25304
rect 38708 25264 38717 25304
rect 38659 25263 38717 25264
rect 40011 25304 40053 25313
rect 40011 25264 40012 25304
rect 40052 25264 40053 25304
rect 40011 25255 40053 25264
rect 40099 25304 40157 25305
rect 40099 25264 40108 25304
rect 40148 25264 40157 25304
rect 40099 25263 40157 25264
rect 40963 25304 41021 25305
rect 40963 25264 40972 25304
rect 41012 25264 41021 25304
rect 40963 25263 41021 25264
rect 44427 25304 44469 25313
rect 44427 25264 44428 25304
rect 44468 25264 44469 25304
rect 44427 25255 44469 25264
rect 44523 25304 44565 25313
rect 44523 25264 44524 25304
rect 44564 25264 44565 25304
rect 44523 25255 44565 25264
rect 44619 25304 44661 25313
rect 44619 25264 44620 25304
rect 44660 25264 44661 25304
rect 44619 25255 44661 25264
rect 44715 25304 44757 25313
rect 44715 25264 44716 25304
rect 44756 25264 44757 25304
rect 44715 25255 44757 25264
rect 44907 25304 44949 25313
rect 44907 25264 44908 25304
rect 44948 25264 44949 25304
rect 44907 25255 44949 25264
rect 45003 25304 45045 25313
rect 45003 25264 45004 25304
rect 45044 25264 45045 25304
rect 45003 25255 45045 25264
rect 45099 25304 45141 25313
rect 45099 25264 45100 25304
rect 45140 25264 45141 25304
rect 45099 25255 45141 25264
rect 45195 25304 45237 25313
rect 45195 25264 45196 25304
rect 45236 25264 45237 25304
rect 45195 25255 45237 25264
rect 45667 25304 45725 25305
rect 45667 25264 45676 25304
rect 45716 25264 45725 25304
rect 45667 25263 45725 25264
rect 48075 25304 48117 25313
rect 48075 25264 48076 25304
rect 48116 25264 48117 25304
rect 48075 25255 48117 25264
rect 48163 25304 48221 25305
rect 48163 25264 48172 25304
rect 48212 25264 48221 25304
rect 48163 25263 48221 25264
rect 49219 25304 49277 25305
rect 49219 25264 49228 25304
rect 49268 25264 49277 25304
rect 49219 25263 49277 25264
rect 50083 25304 50141 25305
rect 50083 25264 50092 25304
rect 50132 25264 50141 25304
rect 50083 25263 50141 25264
rect 50187 25304 50229 25313
rect 50187 25264 50188 25304
rect 50228 25264 50229 25304
rect 50187 25255 50229 25264
rect 50379 25304 50421 25313
rect 50379 25264 50380 25304
rect 50420 25264 50421 25304
rect 50379 25255 50421 25264
rect 51043 25304 51101 25305
rect 51043 25264 51052 25304
rect 51092 25264 51101 25304
rect 51043 25263 51101 25264
rect 51723 25304 51765 25313
rect 51723 25264 51724 25304
rect 51764 25264 51765 25304
rect 51723 25255 51765 25264
rect 51819 25304 51861 25313
rect 51819 25264 51820 25304
rect 51860 25264 51861 25304
rect 51819 25255 51861 25264
rect 51915 25304 51957 25313
rect 51915 25264 51916 25304
rect 51956 25264 51957 25304
rect 51915 25255 51957 25264
rect 53731 25304 53789 25305
rect 53731 25264 53740 25304
rect 53780 25264 53789 25304
rect 53731 25263 53789 25264
rect 53835 25304 53877 25313
rect 53835 25264 53836 25304
rect 53876 25264 53877 25304
rect 53835 25255 53877 25264
rect 54315 25304 54357 25313
rect 54315 25264 54316 25304
rect 54356 25264 54357 25304
rect 54315 25255 54357 25264
rect 54411 25304 54453 25313
rect 54411 25264 54412 25304
rect 54452 25264 54453 25304
rect 54411 25255 54453 25264
rect 54507 25304 54549 25313
rect 54507 25264 54508 25304
rect 54548 25264 54549 25304
rect 54507 25255 54549 25264
rect 54603 25304 54645 25313
rect 54603 25264 54604 25304
rect 54644 25264 54645 25304
rect 54603 25255 54645 25264
rect 56611 25304 56669 25305
rect 56611 25264 56620 25304
rect 56660 25264 56669 25304
rect 56611 25263 56669 25264
rect 56715 25304 56757 25313
rect 56715 25264 56716 25304
rect 56756 25264 56757 25304
rect 56715 25255 56757 25264
rect 57483 25304 57525 25313
rect 57483 25264 57484 25304
rect 57524 25264 57525 25304
rect 57483 25255 57525 25264
rect 57675 25304 57717 25313
rect 57675 25264 57676 25304
rect 57716 25264 57717 25304
rect 57675 25255 57717 25264
rect 57763 25304 57821 25305
rect 57763 25264 57772 25304
rect 57812 25264 57821 25304
rect 57763 25263 57821 25264
rect 58435 25304 58493 25305
rect 58435 25264 58444 25304
rect 58484 25264 58493 25304
rect 58435 25263 58493 25264
rect 59403 25304 59445 25313
rect 59403 25264 59404 25304
rect 59444 25264 59445 25304
rect 59403 25255 59445 25264
rect 59491 25304 59549 25305
rect 59491 25264 59500 25304
rect 59540 25264 59549 25304
rect 59491 25263 59549 25264
rect 61315 25304 61373 25305
rect 61315 25264 61324 25304
rect 61364 25264 61373 25304
rect 61315 25263 61373 25264
rect 62179 25304 62237 25305
rect 62179 25264 62188 25304
rect 62228 25264 62237 25304
rect 62179 25263 62237 25264
rect 64011 25304 64053 25313
rect 64011 25264 64012 25304
rect 64052 25264 64053 25304
rect 64011 25255 64053 25264
rect 64099 25304 64157 25305
rect 64099 25264 64108 25304
rect 64148 25264 64157 25304
rect 64779 25304 64821 25313
rect 64099 25263 64157 25264
rect 64587 25262 64629 25271
rect 45579 25220 45621 25229
rect 45579 25180 45580 25220
rect 45620 25180 45621 25220
rect 60939 25220 60981 25229
rect 45579 25171 45621 25180
rect 54123 25178 54165 25187
rect 843 25136 885 25145
rect 843 25096 844 25136
rect 884 25096 885 25136
rect 843 25087 885 25096
rect 37803 25136 37845 25145
rect 37803 25096 37804 25136
rect 37844 25096 37845 25136
rect 37803 25087 37845 25096
rect 38467 25136 38525 25137
rect 38467 25096 38476 25136
rect 38516 25096 38525 25136
rect 38467 25095 38525 25096
rect 39339 25136 39381 25145
rect 39339 25096 39340 25136
rect 39380 25096 39381 25136
rect 39339 25087 39381 25096
rect 40203 25132 40245 25141
rect 40203 25092 40204 25132
rect 40244 25092 40245 25132
rect 40203 25083 40245 25092
rect 41067 25136 41109 25145
rect 41067 25096 41068 25136
rect 41108 25096 41109 25136
rect 41067 25087 41109 25096
rect 42699 25136 42741 25145
rect 42699 25096 42700 25136
rect 42740 25096 42741 25136
rect 42699 25087 42741 25096
rect 44043 25136 44085 25145
rect 44043 25096 44044 25136
rect 44084 25096 44085 25136
rect 44043 25087 44085 25096
rect 48267 25132 48309 25141
rect 48267 25092 48268 25132
rect 48308 25092 48309 25132
rect 50275 25136 50333 25137
rect 50275 25096 50284 25136
rect 50324 25096 50333 25136
rect 50275 25095 50333 25096
rect 50763 25136 50805 25145
rect 50763 25096 50764 25136
rect 50804 25096 50805 25136
rect 48267 25083 48309 25092
rect 50763 25087 50805 25096
rect 50955 25136 50997 25145
rect 50955 25096 50956 25136
rect 50996 25096 50997 25136
rect 50955 25087 50997 25096
rect 51435 25136 51477 25145
rect 51435 25096 51436 25136
rect 51476 25096 51477 25136
rect 51435 25087 51477 25096
rect 51619 25136 51677 25137
rect 51619 25096 51628 25136
rect 51668 25096 51677 25136
rect 51619 25095 51677 25096
rect 53643 25132 53685 25141
rect 53643 25092 53644 25132
rect 53684 25092 53685 25132
rect 54123 25138 54124 25178
rect 54164 25138 54165 25178
rect 60939 25180 60940 25220
rect 60980 25180 60981 25220
rect 64587 25222 64588 25262
rect 64628 25222 64629 25262
rect 64779 25264 64780 25304
rect 64820 25264 64821 25304
rect 64779 25255 64821 25264
rect 64867 25304 64925 25305
rect 64867 25264 64876 25304
rect 64916 25264 64925 25304
rect 64867 25263 64925 25264
rect 65443 25304 65501 25305
rect 65443 25264 65452 25304
rect 65492 25264 65501 25304
rect 65443 25263 65501 25264
rect 65547 25304 65589 25313
rect 65547 25264 65548 25304
rect 65588 25264 65589 25304
rect 65547 25255 65589 25264
rect 65739 25304 65781 25313
rect 65739 25264 65740 25304
rect 65780 25264 65781 25304
rect 65739 25255 65781 25264
rect 66115 25304 66173 25305
rect 66115 25264 66124 25304
rect 66164 25264 66173 25304
rect 66115 25263 66173 25264
rect 66603 25304 66645 25313
rect 66603 25264 66604 25304
rect 66644 25264 66645 25304
rect 66603 25255 66645 25264
rect 66691 25304 66749 25305
rect 66691 25264 66700 25304
rect 66740 25264 66749 25304
rect 66691 25263 66749 25264
rect 67179 25304 67221 25313
rect 67179 25264 67180 25304
rect 67220 25264 67221 25304
rect 67179 25255 67221 25264
rect 67371 25304 67413 25313
rect 67371 25264 67372 25304
rect 67412 25264 67413 25304
rect 67371 25255 67413 25264
rect 67459 25304 67517 25305
rect 67459 25264 67468 25304
rect 67508 25264 67517 25304
rect 67459 25263 67517 25264
rect 68611 25304 68669 25305
rect 68611 25264 68620 25304
rect 68660 25264 68669 25304
rect 68611 25263 68669 25264
rect 69291 25304 69333 25313
rect 69291 25264 69292 25304
rect 69332 25264 69333 25304
rect 69291 25255 69333 25264
rect 69379 25304 69437 25305
rect 69379 25264 69388 25304
rect 69428 25264 69437 25304
rect 69379 25263 69437 25264
rect 71107 25304 71165 25305
rect 71107 25264 71116 25304
rect 71156 25264 71165 25304
rect 71107 25263 71165 25264
rect 71211 25304 71253 25313
rect 71211 25264 71212 25304
rect 71252 25264 71253 25304
rect 71211 25255 71253 25264
rect 71979 25304 72021 25313
rect 71979 25264 71980 25304
rect 72020 25264 72021 25304
rect 71979 25255 72021 25264
rect 72075 25304 72117 25313
rect 72075 25264 72076 25304
rect 72116 25264 72117 25304
rect 72075 25255 72117 25264
rect 72171 25304 72213 25313
rect 72171 25264 72172 25304
rect 72212 25264 72213 25304
rect 72171 25255 72213 25264
rect 72267 25304 72309 25313
rect 72267 25264 72268 25304
rect 72308 25264 72309 25304
rect 72267 25255 72309 25264
rect 73603 25304 73661 25305
rect 73603 25264 73612 25304
rect 73652 25264 73661 25304
rect 73603 25263 73661 25264
rect 74467 25304 74525 25305
rect 74467 25264 74476 25304
rect 74516 25264 74525 25304
rect 74467 25263 74525 25264
rect 75811 25304 75869 25305
rect 75811 25264 75820 25304
rect 75860 25264 75869 25304
rect 75811 25263 75869 25264
rect 75915 25304 75957 25313
rect 75915 25264 75916 25304
rect 75956 25264 75957 25304
rect 75915 25255 75957 25264
rect 76107 25304 76149 25313
rect 76107 25264 76108 25304
rect 76148 25264 76149 25304
rect 76107 25255 76149 25264
rect 76779 25304 76821 25313
rect 76779 25264 76780 25304
rect 76820 25264 76821 25304
rect 76779 25255 76821 25264
rect 76875 25304 76917 25313
rect 76875 25264 76876 25304
rect 76916 25264 76917 25304
rect 76875 25255 76917 25264
rect 76971 25304 77013 25313
rect 76971 25264 76972 25304
rect 77012 25264 77013 25304
rect 76971 25255 77013 25264
rect 77067 25304 77109 25313
rect 77067 25264 77068 25304
rect 77108 25264 77109 25304
rect 77067 25255 77109 25264
rect 77355 25304 77397 25313
rect 77355 25264 77356 25304
rect 77396 25264 77397 25304
rect 77355 25255 77397 25264
rect 77451 25304 77493 25313
rect 77451 25264 77452 25304
rect 77492 25264 77493 25304
rect 77451 25255 77493 25264
rect 77547 25304 77589 25313
rect 77547 25264 77548 25304
rect 77588 25264 77589 25304
rect 77547 25255 77589 25264
rect 77643 25304 77685 25313
rect 77643 25264 77644 25304
rect 77684 25264 77685 25304
rect 77643 25255 77685 25264
rect 78211 25304 78269 25305
rect 78211 25264 78220 25304
rect 78260 25264 78269 25304
rect 78211 25263 78269 25264
rect 64587 25213 64629 25222
rect 73227 25220 73269 25229
rect 60939 25171 60981 25180
rect 73227 25180 73228 25220
rect 73268 25180 73269 25220
rect 73227 25171 73269 25180
rect 54123 25129 54165 25138
rect 56523 25132 56565 25141
rect 53643 25083 53685 25092
rect 56523 25092 56524 25132
rect 56564 25092 56565 25132
rect 56523 25083 56565 25092
rect 58539 25136 58581 25145
rect 58539 25096 58540 25136
rect 58580 25096 58581 25136
rect 58539 25087 58581 25096
rect 59595 25132 59637 25141
rect 59595 25092 59596 25132
rect 59636 25092 59637 25132
rect 59595 25083 59637 25092
rect 59787 25136 59829 25145
rect 59787 25096 59788 25136
rect 59828 25096 59829 25136
rect 59787 25087 59829 25096
rect 63331 25136 63389 25137
rect 63331 25096 63340 25136
rect 63380 25096 63389 25136
rect 63331 25095 63389 25096
rect 64203 25132 64245 25141
rect 64203 25092 64204 25132
rect 64244 25092 64245 25132
rect 64203 25083 64245 25092
rect 66795 25132 66837 25141
rect 66795 25092 66796 25132
rect 66836 25092 66837 25132
rect 66795 25083 66837 25092
rect 69483 25132 69525 25141
rect 69483 25092 69484 25132
rect 69524 25092 69525 25132
rect 69483 25083 69525 25092
rect 69675 25136 69717 25145
rect 69675 25096 69676 25136
rect 69716 25096 69717 25136
rect 69675 25087 69717 25096
rect 71019 25132 71061 25141
rect 71019 25092 71020 25132
rect 71060 25092 71061 25132
rect 75619 25136 75677 25137
rect 75619 25096 75628 25136
rect 75668 25096 75677 25136
rect 75619 25095 75677 25096
rect 78123 25136 78165 25145
rect 78123 25096 78124 25136
rect 78164 25096 78165 25136
rect 71019 25083 71061 25092
rect 78123 25087 78165 25096
rect 576 24968 79584 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 76352 24968
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76720 24928 79584 24968
rect 576 24904 79584 24928
rect 37803 24858 37845 24867
rect 37803 24818 37804 24858
rect 37844 24818 37845 24858
rect 37803 24809 37845 24818
rect 843 24800 885 24809
rect 843 24760 844 24800
rect 884 24760 885 24800
rect 843 24751 885 24760
rect 2379 24800 2421 24809
rect 75435 24804 75477 24813
rect 2379 24760 2380 24800
rect 2420 24760 2421 24800
rect 2379 24751 2421 24760
rect 40867 24800 40925 24801
rect 40867 24760 40876 24800
rect 40916 24760 40925 24800
rect 40867 24759 40925 24760
rect 43459 24800 43517 24801
rect 43459 24760 43468 24800
rect 43508 24760 43517 24800
rect 43459 24759 43517 24760
rect 75435 24764 75436 24804
rect 75476 24764 75477 24804
rect 75435 24755 75477 24764
rect 38475 24716 38517 24725
rect 38475 24676 38476 24716
rect 38516 24676 38517 24716
rect 38475 24667 38517 24676
rect 41067 24716 41109 24725
rect 41067 24676 41068 24716
rect 41108 24676 41109 24716
rect 41067 24667 41109 24676
rect 36355 24632 36413 24633
rect 36355 24592 36364 24632
rect 36404 24592 36413 24632
rect 36355 24591 36413 24592
rect 37219 24632 37277 24633
rect 37219 24592 37228 24632
rect 37268 24592 37277 24632
rect 37219 24591 37277 24592
rect 37611 24632 37653 24641
rect 37611 24592 37612 24632
rect 37652 24592 37653 24632
rect 37611 24583 37653 24592
rect 37891 24632 37949 24633
rect 37891 24592 37900 24632
rect 37940 24592 37949 24632
rect 37891 24591 37949 24592
rect 37995 24632 38037 24641
rect 37995 24592 37996 24632
rect 38036 24592 38037 24632
rect 37995 24583 38037 24592
rect 38851 24632 38909 24633
rect 38851 24592 38860 24632
rect 38900 24592 38909 24632
rect 38851 24591 38909 24592
rect 39715 24632 39773 24633
rect 39715 24592 39724 24632
rect 39764 24592 39773 24632
rect 39715 24591 39773 24592
rect 41443 24632 41501 24633
rect 41443 24592 41452 24632
rect 41492 24592 41501 24632
rect 41443 24591 41501 24592
rect 42307 24632 42365 24633
rect 42307 24592 42316 24632
rect 42356 24592 42365 24632
rect 42307 24591 42365 24592
rect 43659 24632 43701 24641
rect 43659 24592 43660 24632
rect 43700 24592 43701 24632
rect 43659 24583 43701 24592
rect 44035 24632 44093 24633
rect 44035 24592 44044 24632
rect 44084 24592 44093 24632
rect 44035 24591 44093 24592
rect 44899 24632 44957 24633
rect 44899 24592 44908 24632
rect 44948 24592 44957 24632
rect 44899 24591 44957 24592
rect 46251 24632 46293 24641
rect 46251 24592 46252 24632
rect 46292 24592 46293 24632
rect 46251 24583 46293 24592
rect 46627 24632 46685 24633
rect 46627 24592 46636 24632
rect 46676 24592 46685 24632
rect 46627 24591 46685 24592
rect 47491 24632 47549 24633
rect 47491 24592 47500 24632
rect 47540 24592 47549 24632
rect 47491 24591 47549 24592
rect 48843 24632 48885 24641
rect 48843 24592 48844 24632
rect 48884 24592 48885 24632
rect 48843 24583 48885 24592
rect 49219 24632 49277 24633
rect 49219 24592 49228 24632
rect 49268 24592 49277 24632
rect 49219 24591 49277 24592
rect 50083 24632 50141 24633
rect 50083 24592 50092 24632
rect 50132 24592 50141 24632
rect 50083 24591 50141 24592
rect 51435 24632 51477 24641
rect 51435 24592 51436 24632
rect 51476 24592 51477 24632
rect 51435 24583 51477 24592
rect 51811 24632 51869 24633
rect 51811 24592 51820 24632
rect 51860 24592 51869 24632
rect 51811 24591 51869 24592
rect 52675 24632 52733 24633
rect 52675 24592 52684 24632
rect 52724 24592 52733 24632
rect 52675 24591 52733 24592
rect 54027 24632 54069 24641
rect 54027 24592 54028 24632
rect 54068 24592 54069 24632
rect 54027 24583 54069 24592
rect 54403 24632 54461 24633
rect 54403 24592 54412 24632
rect 54452 24592 54461 24632
rect 54403 24591 54461 24592
rect 55267 24632 55325 24633
rect 55267 24592 55276 24632
rect 55316 24592 55325 24632
rect 55267 24591 55325 24592
rect 56619 24632 56661 24641
rect 56619 24592 56620 24632
rect 56660 24592 56661 24632
rect 56619 24583 56661 24592
rect 56995 24632 57053 24633
rect 56995 24592 57004 24632
rect 57044 24592 57053 24632
rect 56995 24591 57053 24592
rect 57859 24632 57917 24633
rect 57859 24592 57868 24632
rect 57908 24592 57917 24632
rect 57859 24591 57917 24592
rect 59499 24632 59541 24641
rect 59499 24592 59500 24632
rect 59540 24592 59541 24632
rect 59499 24583 59541 24592
rect 59875 24632 59933 24633
rect 59875 24592 59884 24632
rect 59924 24592 59933 24632
rect 59875 24591 59933 24592
rect 60739 24632 60797 24633
rect 60739 24592 60748 24632
rect 60788 24592 60797 24632
rect 60739 24591 60797 24592
rect 62859 24632 62901 24641
rect 62859 24592 62860 24632
rect 62900 24592 62901 24632
rect 62859 24583 62901 24592
rect 62955 24632 62997 24641
rect 62955 24592 62956 24632
rect 62996 24592 62997 24632
rect 62955 24583 62997 24592
rect 63051 24632 63093 24641
rect 63051 24592 63052 24632
rect 63092 24592 63093 24632
rect 63051 24583 63093 24592
rect 63147 24632 63189 24641
rect 63147 24592 63148 24632
rect 63188 24592 63189 24632
rect 63147 24583 63189 24592
rect 63339 24632 63381 24641
rect 63339 24592 63340 24632
rect 63380 24592 63381 24632
rect 63339 24583 63381 24592
rect 63715 24632 63773 24633
rect 63715 24592 63724 24632
rect 63764 24592 63773 24632
rect 63715 24591 63773 24592
rect 64579 24632 64637 24633
rect 64579 24592 64588 24632
rect 64628 24592 64637 24632
rect 64579 24591 64637 24592
rect 66987 24632 67029 24641
rect 66987 24592 66988 24632
rect 67028 24592 67029 24632
rect 66987 24583 67029 24592
rect 67083 24632 67125 24641
rect 67083 24592 67084 24632
rect 67124 24592 67125 24632
rect 67083 24583 67125 24592
rect 67179 24632 67221 24641
rect 67179 24592 67180 24632
rect 67220 24592 67221 24632
rect 67179 24583 67221 24592
rect 67275 24632 67317 24641
rect 67275 24592 67276 24632
rect 67316 24592 67317 24632
rect 67275 24583 67317 24592
rect 69099 24632 69141 24641
rect 69099 24592 69100 24632
rect 69140 24592 69141 24632
rect 69099 24583 69141 24592
rect 69475 24632 69533 24633
rect 69475 24592 69484 24632
rect 69524 24592 69533 24632
rect 69475 24591 69533 24592
rect 70339 24632 70397 24633
rect 70339 24592 70348 24632
rect 70388 24592 70397 24632
rect 70339 24591 70397 24592
rect 71691 24632 71733 24641
rect 71691 24592 71692 24632
rect 71732 24592 71733 24632
rect 71691 24583 71733 24592
rect 72067 24632 72125 24633
rect 72067 24592 72076 24632
rect 72116 24592 72125 24632
rect 72067 24591 72125 24592
rect 72931 24632 72989 24633
rect 72931 24592 72940 24632
rect 72980 24592 72989 24632
rect 72931 24591 72989 24592
rect 74859 24632 74901 24641
rect 74859 24592 74860 24632
rect 74900 24592 74901 24632
rect 74859 24583 74901 24592
rect 75235 24632 75293 24633
rect 75235 24592 75244 24632
rect 75284 24592 75293 24632
rect 75235 24591 75293 24592
rect 75523 24632 75581 24633
rect 75523 24592 75532 24632
rect 75572 24592 75581 24632
rect 75523 24591 75581 24592
rect 75627 24632 75669 24641
rect 75627 24592 75628 24632
rect 75668 24592 75669 24632
rect 75627 24583 75669 24592
rect 76587 24632 76629 24641
rect 76587 24592 76588 24632
rect 76628 24592 76629 24632
rect 76587 24583 76629 24592
rect 76963 24632 77021 24633
rect 76963 24592 76972 24632
rect 77012 24592 77021 24632
rect 76963 24591 77021 24592
rect 77827 24632 77885 24633
rect 77827 24592 77836 24632
rect 77876 24592 77885 24632
rect 77827 24591 77885 24592
rect 643 24548 701 24549
rect 643 24508 652 24548
rect 692 24508 701 24548
rect 643 24507 701 24508
rect 1795 24548 1853 24549
rect 1795 24508 1804 24548
rect 1844 24508 1853 24548
rect 1795 24507 1853 24508
rect 2179 24548 2237 24549
rect 2179 24508 2188 24548
rect 2228 24508 2237 24548
rect 2179 24507 2237 24508
rect 35211 24548 35253 24557
rect 35211 24508 35212 24548
rect 35252 24508 35253 24548
rect 35211 24499 35253 24508
rect 51243 24548 51285 24557
rect 51243 24508 51244 24548
rect 51284 24508 51285 24548
rect 51243 24499 51285 24508
rect 53835 24548 53877 24557
rect 53835 24508 53836 24548
rect 53876 24508 53877 24548
rect 53835 24499 53877 24508
rect 56427 24548 56469 24557
rect 56427 24508 56428 24548
rect 56468 24508 56469 24548
rect 56427 24499 56469 24508
rect 61899 24548 61941 24557
rect 61899 24508 61900 24548
rect 61940 24508 61941 24548
rect 61899 24499 61941 24508
rect 65739 24548 65781 24557
rect 65739 24508 65740 24548
rect 65780 24508 65781 24548
rect 65739 24499 65781 24508
rect 68707 24548 68765 24549
rect 68707 24508 68716 24548
rect 68756 24508 68765 24548
rect 68707 24507 68765 24508
rect 74091 24548 74133 24557
rect 74091 24508 74092 24548
rect 74132 24508 74133 24548
rect 74091 24499 74133 24508
rect 74955 24548 74997 24557
rect 74955 24508 74956 24548
rect 74996 24508 74997 24548
rect 74955 24499 74997 24508
rect 75147 24548 75189 24557
rect 75147 24508 75148 24548
rect 75188 24508 75189 24548
rect 75147 24499 75189 24508
rect 76195 24548 76253 24549
rect 76195 24508 76204 24548
rect 76244 24508 76253 24548
rect 76195 24507 76253 24508
rect 78987 24548 79029 24557
rect 78987 24508 78988 24548
rect 79028 24508 79029 24548
rect 78987 24499 79029 24508
rect 75051 24464 75093 24473
rect 75051 24424 75052 24464
rect 75092 24424 75093 24464
rect 75051 24415 75093 24424
rect 75915 24464 75957 24473
rect 75915 24424 75916 24464
rect 75956 24424 75957 24464
rect 75915 24415 75957 24424
rect 1995 24380 2037 24389
rect 1995 24340 1996 24380
rect 2036 24340 2037 24380
rect 1995 24331 2037 24340
rect 38283 24380 38325 24389
rect 38283 24340 38284 24380
rect 38324 24340 38325 24380
rect 38283 24331 38325 24340
rect 40867 24380 40925 24381
rect 40867 24340 40876 24380
rect 40916 24340 40925 24380
rect 40867 24339 40925 24340
rect 46051 24380 46109 24381
rect 46051 24340 46060 24380
rect 46100 24340 46109 24380
rect 46051 24339 46109 24340
rect 48643 24380 48701 24381
rect 48643 24340 48652 24380
rect 48692 24340 48701 24380
rect 48643 24339 48701 24340
rect 59011 24380 59069 24381
rect 59011 24340 59020 24380
rect 59060 24340 59069 24380
rect 59011 24339 59069 24340
rect 68907 24380 68949 24389
rect 68907 24340 68908 24380
rect 68948 24340 68949 24380
rect 68907 24331 68949 24340
rect 71491 24380 71549 24381
rect 71491 24340 71500 24380
rect 71540 24340 71549 24380
rect 71491 24339 71549 24340
rect 76395 24380 76437 24389
rect 76395 24340 76396 24380
rect 76436 24340 76437 24380
rect 76395 24331 76437 24340
rect 576 24212 79584 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 79584 24212
rect 576 24148 79584 24172
rect 41739 24044 41781 24053
rect 41739 24004 41740 24044
rect 41780 24004 41781 24044
rect 51339 24044 51381 24053
rect 41739 23995 41781 24004
rect 50475 24002 50517 24011
rect 37995 23960 38037 23969
rect 37995 23920 37996 23960
rect 38036 23920 38037 23960
rect 37995 23911 38037 23920
rect 42795 23960 42837 23969
rect 42795 23920 42796 23960
rect 42836 23920 42837 23960
rect 42795 23911 42837 23920
rect 43851 23960 43893 23969
rect 43851 23920 43852 23960
rect 43892 23920 43893 23960
rect 50475 23962 50476 24002
rect 50516 23962 50517 24002
rect 51339 24004 51340 24044
rect 51380 24004 51381 24044
rect 51339 23995 51381 24004
rect 52203 24044 52245 24053
rect 52203 24004 52204 24044
rect 52244 24004 52245 24044
rect 52203 23995 52245 24004
rect 53067 24044 53109 24053
rect 53067 24004 53068 24044
rect 53108 24004 53109 24044
rect 53067 23995 53109 24004
rect 54987 24044 55029 24053
rect 54987 24004 54988 24044
rect 55028 24004 55029 24044
rect 54987 23995 55029 24004
rect 55947 24044 55989 24053
rect 55947 24004 55948 24044
rect 55988 24004 55989 24044
rect 55947 23995 55989 24004
rect 56427 24044 56469 24053
rect 56427 24004 56428 24044
rect 56468 24004 56469 24044
rect 56427 23995 56469 24004
rect 62187 24044 62229 24053
rect 62187 24004 62188 24044
rect 62228 24004 62229 24044
rect 62187 23995 62229 24004
rect 64011 24044 64053 24053
rect 64011 24004 64012 24044
rect 64052 24004 64053 24044
rect 64011 23995 64053 24004
rect 65259 24044 65301 24053
rect 65259 24004 65260 24044
rect 65300 24004 65301 24044
rect 65259 23995 65301 24004
rect 68803 24044 68861 24045
rect 68803 24004 68812 24044
rect 68852 24004 68861 24044
rect 68803 24003 68861 24004
rect 74859 24044 74901 24053
rect 74859 24004 74860 24044
rect 74900 24004 74901 24044
rect 74859 23995 74901 24004
rect 75531 24044 75573 24053
rect 75531 24004 75532 24044
rect 75572 24004 75573 24044
rect 75531 23995 75573 24004
rect 50475 23953 50517 23962
rect 57771 23960 57813 23969
rect 43851 23911 43893 23920
rect 57771 23920 57772 23960
rect 57812 23920 57813 23960
rect 57771 23911 57813 23920
rect 65451 23960 65493 23969
rect 65451 23920 65452 23960
rect 65492 23920 65493 23960
rect 65451 23911 65493 23920
rect 71979 23960 72021 23969
rect 71979 23920 71980 23960
rect 72020 23920 72021 23960
rect 71979 23911 72021 23920
rect 643 23876 701 23877
rect 643 23836 652 23876
rect 692 23836 701 23876
rect 643 23835 701 23836
rect 1795 23876 1853 23877
rect 1795 23836 1804 23876
rect 1844 23836 1853 23876
rect 1795 23835 1853 23836
rect 2179 23876 2237 23877
rect 2179 23836 2188 23876
rect 2228 23836 2237 23876
rect 2179 23835 2237 23836
rect 37899 23876 37941 23885
rect 37899 23836 37900 23876
rect 37940 23836 37941 23876
rect 37899 23827 37941 23836
rect 38091 23876 38133 23885
rect 38091 23836 38092 23876
rect 38132 23836 38133 23876
rect 38091 23827 38133 23836
rect 40483 23876 40541 23877
rect 40483 23836 40492 23876
rect 40532 23836 40541 23876
rect 40483 23835 40541 23836
rect 42699 23876 42741 23885
rect 42699 23836 42700 23876
rect 42740 23836 42741 23876
rect 42699 23827 42741 23836
rect 42891 23876 42933 23885
rect 42891 23836 42892 23876
rect 42932 23836 42933 23876
rect 50379 23876 50421 23885
rect 50379 23836 50380 23876
rect 50420 23836 50421 23876
rect 42891 23827 42933 23836
rect 43459 23835 43517 23836
rect 36363 23792 36405 23801
rect 36171 23750 36213 23759
rect 36171 23710 36172 23750
rect 36212 23710 36213 23750
rect 36363 23752 36364 23792
rect 36404 23752 36405 23792
rect 36363 23743 36405 23752
rect 36451 23792 36509 23793
rect 36451 23752 36460 23792
rect 36500 23752 36509 23792
rect 36451 23751 36509 23752
rect 36747 23792 36789 23801
rect 36747 23752 36748 23792
rect 36788 23752 36789 23792
rect 36747 23743 36789 23752
rect 36843 23792 36885 23801
rect 36843 23752 36844 23792
rect 36884 23752 36885 23792
rect 36843 23743 36885 23752
rect 36939 23792 36981 23801
rect 36939 23752 36940 23792
rect 36980 23752 36981 23792
rect 36939 23743 36981 23752
rect 37803 23792 37845 23801
rect 37803 23752 37804 23792
rect 37844 23752 37845 23792
rect 37803 23743 37845 23752
rect 38179 23792 38237 23793
rect 38179 23752 38188 23792
rect 38228 23752 38237 23792
rect 38179 23751 38237 23752
rect 38667 23792 38709 23801
rect 38667 23752 38668 23792
rect 38708 23752 38709 23792
rect 38667 23743 38709 23752
rect 38763 23792 38805 23801
rect 38763 23752 38764 23792
rect 38804 23752 38805 23792
rect 38763 23743 38805 23752
rect 38859 23792 38901 23801
rect 38859 23752 38860 23792
rect 38900 23752 38901 23792
rect 38859 23743 38901 23752
rect 38955 23792 38997 23801
rect 38955 23752 38956 23792
rect 38996 23752 38997 23792
rect 38955 23743 38997 23752
rect 39147 23792 39189 23801
rect 39147 23752 39148 23792
rect 39188 23752 39189 23792
rect 39147 23743 39189 23752
rect 39243 23792 39285 23801
rect 39243 23752 39244 23792
rect 39284 23752 39285 23792
rect 39243 23743 39285 23752
rect 39339 23792 39381 23801
rect 39339 23752 39340 23792
rect 39380 23752 39381 23792
rect 39339 23743 39381 23752
rect 39435 23792 39477 23801
rect 39435 23752 39436 23792
rect 39476 23752 39477 23792
rect 39435 23743 39477 23752
rect 40875 23792 40917 23801
rect 40875 23752 40876 23792
rect 40916 23752 40917 23792
rect 40875 23743 40917 23752
rect 41067 23792 41109 23801
rect 41067 23752 41068 23792
rect 41108 23752 41109 23792
rect 41067 23743 41109 23752
rect 41155 23792 41213 23793
rect 41155 23752 41164 23792
rect 41204 23752 41213 23792
rect 41155 23751 41213 23752
rect 41443 23792 41501 23793
rect 41443 23752 41452 23792
rect 41492 23752 41501 23792
rect 41443 23751 41501 23752
rect 42603 23792 42645 23801
rect 43459 23795 43468 23835
rect 43508 23795 43517 23835
rect 50379 23827 50421 23836
rect 50571 23876 50613 23885
rect 50571 23836 50572 23876
rect 50612 23836 50613 23876
rect 50571 23827 50613 23836
rect 52003 23876 52061 23877
rect 52003 23836 52012 23876
rect 52052 23836 52061 23876
rect 52003 23835 52061 23836
rect 63243 23876 63285 23885
rect 63243 23836 63244 23876
rect 63284 23836 63285 23876
rect 51619 23834 51677 23835
rect 43459 23794 43517 23795
rect 42603 23752 42604 23792
rect 42644 23752 42645 23792
rect 42603 23743 42645 23752
rect 42979 23792 43037 23793
rect 42979 23752 42988 23792
rect 43028 23752 43037 23792
rect 42979 23751 43037 23752
rect 43563 23792 43605 23801
rect 43563 23752 43564 23792
rect 43604 23752 43605 23792
rect 43563 23743 43605 23752
rect 44139 23792 44181 23801
rect 44139 23752 44140 23792
rect 44180 23752 44181 23792
rect 44139 23743 44181 23752
rect 44235 23792 44277 23801
rect 44235 23752 44236 23792
rect 44276 23752 44277 23792
rect 44235 23743 44277 23752
rect 44331 23792 44373 23801
rect 44331 23752 44332 23792
rect 44372 23752 44373 23792
rect 44331 23743 44373 23752
rect 44427 23792 44469 23801
rect 44427 23752 44428 23792
rect 44468 23752 44469 23792
rect 44427 23743 44469 23752
rect 47307 23792 47349 23801
rect 47307 23752 47308 23792
rect 47348 23752 47349 23792
rect 47307 23743 47349 23752
rect 47403 23792 47445 23801
rect 47403 23752 47404 23792
rect 47444 23752 47445 23792
rect 47403 23743 47445 23752
rect 47499 23792 47541 23801
rect 47499 23752 47500 23792
rect 47540 23752 47541 23792
rect 47499 23743 47541 23752
rect 47595 23792 47637 23801
rect 47595 23752 47596 23792
rect 47636 23752 47637 23792
rect 47595 23743 47637 23752
rect 48171 23792 48213 23801
rect 48171 23752 48172 23792
rect 48212 23752 48213 23792
rect 48171 23743 48213 23752
rect 48267 23792 48309 23801
rect 48267 23752 48268 23792
rect 48308 23752 48309 23792
rect 48267 23743 48309 23752
rect 48363 23792 48405 23801
rect 48363 23752 48364 23792
rect 48404 23752 48405 23792
rect 48363 23743 48405 23752
rect 48459 23792 48501 23801
rect 48459 23752 48460 23792
rect 48500 23752 48501 23792
rect 48459 23743 48501 23752
rect 48747 23792 48789 23801
rect 48747 23752 48748 23792
rect 48788 23752 48789 23792
rect 48747 23743 48789 23752
rect 48835 23792 48893 23793
rect 48835 23752 48844 23792
rect 48884 23752 48893 23792
rect 48835 23751 48893 23752
rect 49795 23792 49853 23793
rect 49795 23752 49804 23792
rect 49844 23752 49853 23792
rect 49795 23751 49853 23752
rect 49899 23792 49941 23801
rect 49899 23752 49900 23792
rect 49940 23752 49941 23792
rect 49899 23743 49941 23752
rect 50091 23792 50133 23801
rect 50091 23752 50092 23792
rect 50132 23752 50133 23792
rect 50091 23743 50133 23752
rect 50283 23792 50325 23801
rect 50283 23752 50284 23792
rect 50324 23752 50325 23792
rect 50283 23743 50325 23752
rect 50947 23792 51005 23793
rect 50947 23752 50956 23792
rect 50996 23752 51005 23792
rect 50947 23751 51005 23752
rect 51051 23792 51093 23801
rect 51051 23752 51052 23792
rect 51092 23752 51093 23792
rect 50659 23750 50717 23751
rect 36171 23701 36213 23710
rect 40971 23708 41013 23717
rect 50659 23710 50668 23750
rect 50708 23710 50717 23750
rect 51051 23743 51093 23752
rect 51531 23792 51573 23801
rect 51619 23794 51628 23834
rect 51668 23794 51677 23834
rect 63243 23827 63285 23836
rect 51619 23793 51677 23794
rect 51531 23752 51532 23792
rect 51572 23752 51573 23792
rect 51531 23743 51573 23752
rect 51723 23792 51765 23801
rect 51723 23752 51724 23792
rect 51764 23752 51765 23792
rect 51723 23743 51765 23752
rect 51819 23800 51861 23809
rect 51819 23760 51820 23800
rect 51860 23760 51861 23800
rect 51819 23751 51861 23760
rect 53155 23792 53213 23793
rect 53155 23752 53164 23792
rect 53204 23752 53213 23792
rect 53155 23751 53213 23752
rect 53835 23792 53877 23801
rect 53835 23752 53836 23792
rect 53876 23752 53877 23792
rect 53835 23743 53877 23752
rect 53931 23792 53973 23801
rect 53931 23752 53932 23792
rect 53972 23752 53973 23792
rect 53931 23743 53973 23752
rect 54027 23792 54069 23801
rect 54027 23752 54028 23792
rect 54068 23752 54069 23792
rect 54027 23743 54069 23752
rect 54123 23792 54165 23801
rect 54123 23752 54124 23792
rect 54164 23752 54165 23792
rect 54123 23743 54165 23752
rect 55075 23792 55133 23793
rect 55075 23752 55084 23792
rect 55124 23752 55133 23792
rect 55075 23751 55133 23752
rect 55651 23792 55709 23793
rect 55651 23752 55660 23792
rect 55700 23752 55709 23792
rect 55651 23751 55709 23752
rect 56035 23792 56093 23793
rect 56035 23752 56044 23792
rect 56084 23752 56093 23792
rect 56035 23751 56093 23752
rect 56323 23792 56381 23793
rect 56323 23752 56332 23792
rect 56372 23752 56381 23792
rect 56323 23751 56381 23752
rect 56619 23792 56661 23801
rect 56619 23752 56620 23792
rect 56660 23752 56661 23792
rect 56619 23743 56661 23752
rect 56715 23792 56757 23801
rect 56715 23752 56716 23792
rect 56756 23752 56757 23792
rect 56715 23743 56757 23752
rect 56811 23792 56853 23801
rect 56811 23752 56812 23792
rect 56852 23752 56853 23792
rect 56811 23743 56853 23752
rect 56907 23792 56949 23801
rect 56907 23752 56908 23792
rect 56948 23752 56949 23792
rect 56907 23743 56949 23752
rect 57099 23792 57141 23801
rect 57099 23752 57100 23792
rect 57140 23752 57141 23792
rect 57099 23743 57141 23752
rect 57195 23792 57237 23801
rect 57195 23752 57196 23792
rect 57236 23752 57237 23792
rect 57195 23743 57237 23752
rect 57291 23792 57333 23801
rect 57291 23752 57292 23792
rect 57332 23752 57333 23792
rect 57291 23743 57333 23752
rect 57387 23792 57429 23801
rect 57387 23752 57388 23792
rect 57428 23752 57429 23792
rect 57387 23743 57429 23752
rect 57859 23792 57917 23793
rect 57859 23752 57868 23792
rect 57908 23752 57917 23792
rect 57859 23751 57917 23752
rect 59307 23792 59349 23801
rect 59307 23752 59308 23792
rect 59348 23752 59349 23792
rect 59307 23743 59349 23752
rect 59403 23792 59445 23801
rect 59403 23752 59404 23792
rect 59444 23752 59445 23792
rect 59403 23743 59445 23752
rect 59499 23792 59541 23801
rect 59499 23752 59500 23792
rect 59540 23752 59541 23792
rect 59499 23743 59541 23752
rect 59595 23792 59637 23801
rect 59595 23752 59596 23792
rect 59636 23752 59637 23792
rect 59595 23743 59637 23752
rect 59787 23792 59829 23801
rect 59787 23752 59788 23792
rect 59828 23752 59829 23792
rect 59787 23743 59829 23752
rect 59883 23792 59925 23801
rect 59883 23752 59884 23792
rect 59924 23752 59925 23792
rect 59883 23743 59925 23752
rect 59979 23792 60021 23801
rect 59979 23752 59980 23792
rect 60020 23752 60021 23792
rect 59979 23743 60021 23752
rect 60075 23792 60117 23801
rect 60075 23752 60076 23792
rect 60116 23752 60117 23792
rect 60075 23743 60117 23752
rect 60355 23792 60413 23793
rect 60355 23752 60364 23792
rect 60404 23752 60413 23792
rect 60355 23751 60413 23752
rect 60939 23792 60981 23801
rect 60939 23752 60940 23792
rect 60980 23752 60981 23792
rect 60939 23743 60981 23752
rect 61035 23792 61077 23801
rect 61035 23752 61036 23792
rect 61076 23752 61077 23792
rect 61035 23743 61077 23752
rect 61131 23792 61173 23801
rect 61131 23752 61132 23792
rect 61172 23752 61173 23792
rect 61131 23743 61173 23752
rect 61227 23792 61269 23801
rect 61227 23752 61228 23792
rect 61268 23752 61269 23792
rect 61227 23743 61269 23752
rect 62083 23792 62141 23793
rect 62083 23752 62092 23792
rect 62132 23752 62141 23792
rect 62083 23751 62141 23752
rect 62571 23792 62613 23801
rect 62571 23752 62572 23792
rect 62612 23752 62613 23792
rect 62571 23743 62613 23752
rect 62659 23792 62717 23793
rect 62659 23752 62668 23792
rect 62708 23752 62717 23792
rect 62659 23751 62717 23752
rect 63907 23792 63965 23793
rect 63907 23752 63916 23792
rect 63956 23752 63965 23792
rect 63907 23751 63965 23752
rect 64203 23792 64245 23801
rect 64203 23752 64204 23792
rect 64244 23752 64245 23792
rect 64203 23743 64245 23752
rect 64299 23792 64341 23801
rect 64299 23752 64300 23792
rect 64340 23752 64341 23792
rect 64299 23743 64341 23752
rect 64395 23792 64437 23801
rect 64395 23752 64396 23792
rect 64436 23752 64437 23792
rect 64395 23743 64437 23752
rect 64491 23792 64533 23801
rect 64491 23752 64492 23792
rect 64532 23752 64533 23792
rect 64491 23743 64533 23752
rect 64771 23792 64829 23793
rect 64771 23752 64780 23792
rect 64820 23752 64829 23792
rect 64771 23751 64829 23752
rect 65155 23792 65213 23793
rect 65155 23752 65164 23792
rect 65204 23752 65213 23792
rect 65155 23751 65213 23752
rect 65931 23792 65973 23801
rect 65931 23752 65932 23792
rect 65972 23752 65973 23792
rect 65931 23743 65973 23752
rect 66027 23792 66069 23801
rect 66027 23752 66028 23792
rect 66068 23752 66069 23792
rect 66027 23743 66069 23752
rect 66123 23792 66165 23801
rect 66123 23752 66124 23792
rect 66164 23752 66165 23792
rect 66123 23743 66165 23752
rect 66787 23792 66845 23793
rect 66787 23752 66796 23792
rect 66836 23752 66845 23792
rect 66787 23751 66845 23752
rect 67651 23792 67709 23793
rect 67651 23752 67660 23792
rect 67700 23752 67709 23792
rect 67651 23751 67709 23752
rect 69099 23792 69141 23801
rect 69099 23752 69100 23792
rect 69140 23752 69141 23792
rect 69099 23743 69141 23752
rect 69195 23792 69237 23801
rect 69195 23752 69196 23792
rect 69236 23752 69237 23792
rect 69195 23743 69237 23752
rect 69291 23792 69333 23801
rect 69291 23752 69292 23792
rect 69332 23752 69333 23792
rect 69291 23743 69333 23752
rect 69387 23792 69429 23801
rect 69387 23752 69388 23792
rect 69428 23752 69429 23792
rect 69387 23743 69429 23752
rect 69963 23792 70005 23801
rect 69963 23752 69964 23792
rect 70004 23752 70005 23792
rect 69963 23743 70005 23752
rect 70059 23792 70101 23801
rect 70059 23752 70060 23792
rect 70100 23752 70101 23792
rect 70059 23743 70101 23752
rect 70155 23792 70197 23801
rect 70155 23752 70156 23792
rect 70196 23752 70197 23792
rect 70155 23743 70197 23752
rect 70251 23792 70293 23801
rect 70251 23752 70252 23792
rect 70292 23752 70293 23792
rect 70251 23743 70293 23752
rect 71211 23792 71253 23801
rect 71211 23752 71212 23792
rect 71252 23752 71253 23792
rect 71211 23743 71253 23752
rect 71307 23792 71349 23801
rect 71307 23752 71308 23792
rect 71348 23752 71349 23792
rect 71307 23743 71349 23752
rect 71403 23792 71445 23801
rect 71403 23752 71404 23792
rect 71444 23752 71445 23792
rect 71403 23743 71445 23752
rect 71499 23792 71541 23801
rect 71499 23752 71500 23792
rect 71540 23752 71541 23792
rect 71499 23743 71541 23752
rect 72067 23792 72125 23793
rect 72067 23752 72076 23792
rect 72116 23752 72125 23792
rect 72067 23751 72125 23752
rect 72451 23792 72509 23793
rect 72451 23752 72460 23792
rect 72500 23752 72509 23792
rect 72451 23751 72509 23752
rect 72747 23792 72789 23801
rect 72747 23752 72748 23792
rect 72788 23752 72789 23792
rect 72747 23743 72789 23752
rect 72835 23792 72893 23793
rect 72835 23752 72844 23792
rect 72884 23752 72893 23792
rect 72835 23751 72893 23752
rect 74859 23792 74901 23801
rect 74859 23752 74860 23792
rect 74900 23752 74901 23792
rect 74859 23743 74901 23752
rect 75051 23792 75093 23801
rect 75051 23752 75052 23792
rect 75092 23752 75093 23792
rect 75051 23743 75093 23752
rect 75139 23792 75197 23793
rect 75139 23752 75148 23792
rect 75188 23752 75197 23792
rect 75139 23751 75197 23752
rect 75619 23792 75677 23793
rect 75619 23752 75628 23792
rect 75668 23752 75677 23792
rect 75619 23751 75677 23752
rect 76203 23792 76245 23801
rect 76203 23752 76204 23792
rect 76244 23752 76245 23792
rect 76203 23743 76245 23752
rect 76299 23792 76341 23801
rect 76299 23752 76300 23792
rect 76340 23752 76341 23792
rect 76299 23743 76341 23752
rect 76395 23792 76437 23801
rect 76395 23752 76396 23792
rect 76436 23752 76437 23792
rect 76395 23743 76437 23752
rect 76587 23792 76629 23801
rect 76587 23752 76588 23792
rect 76628 23752 76629 23792
rect 76587 23743 76629 23752
rect 76683 23792 76725 23801
rect 76683 23752 76684 23792
rect 76724 23752 76725 23792
rect 76683 23743 76725 23752
rect 76779 23792 76821 23801
rect 76779 23752 76780 23792
rect 76820 23752 76821 23792
rect 76779 23743 76821 23752
rect 77251 23792 77309 23793
rect 77251 23752 77260 23792
rect 77300 23752 77309 23792
rect 77251 23751 77309 23752
rect 78787 23792 78845 23793
rect 78787 23752 78796 23792
rect 78836 23752 78845 23792
rect 78787 23751 78845 23752
rect 78979 23792 79037 23793
rect 78979 23752 78988 23792
rect 79028 23752 79037 23792
rect 78979 23751 79037 23752
rect 50659 23709 50717 23710
rect 40971 23668 40972 23708
rect 41012 23668 41013 23708
rect 40971 23659 41013 23668
rect 55563 23708 55605 23717
rect 55563 23668 55564 23708
rect 55604 23668 55605 23708
rect 55563 23659 55605 23668
rect 66219 23708 66261 23717
rect 66219 23668 66220 23708
rect 66260 23668 66261 23708
rect 66219 23659 66261 23668
rect 66411 23708 66453 23717
rect 66411 23668 66412 23708
rect 66452 23668 66453 23708
rect 66411 23659 66453 23668
rect 843 23624 885 23633
rect 843 23584 844 23624
rect 884 23584 885 23624
rect 843 23575 885 23584
rect 1611 23624 1653 23633
rect 1611 23584 1612 23624
rect 1652 23584 1653 23624
rect 1611 23575 1653 23584
rect 1995 23624 2037 23633
rect 1995 23584 1996 23624
rect 2036 23584 2037 23624
rect 1995 23575 2037 23584
rect 36259 23624 36317 23625
rect 36259 23584 36268 23624
rect 36308 23584 36317 23624
rect 36259 23583 36317 23584
rect 36643 23624 36701 23625
rect 36643 23584 36652 23624
rect 36692 23584 36701 23624
rect 36643 23583 36701 23584
rect 40683 23624 40725 23633
rect 40683 23584 40684 23624
rect 40724 23584 40725 23624
rect 40683 23575 40725 23584
rect 49987 23624 50045 23625
rect 49987 23584 49996 23624
rect 50036 23584 50045 23624
rect 49987 23583 50045 23584
rect 50859 23620 50901 23629
rect 50859 23580 50860 23620
rect 50900 23580 50901 23620
rect 43371 23566 43413 23575
rect 50859 23571 50901 23580
rect 55947 23624 55989 23633
rect 55947 23584 55948 23624
rect 55988 23584 55989 23624
rect 55947 23575 55989 23584
rect 60267 23624 60309 23633
rect 60267 23584 60268 23624
rect 60308 23584 60309 23624
rect 60267 23575 60309 23584
rect 64875 23624 64917 23633
rect 64875 23584 64876 23624
rect 64916 23584 64917 23624
rect 64875 23575 64917 23584
rect 65259 23624 65301 23633
rect 65259 23584 65260 23624
rect 65300 23584 65301 23624
rect 65259 23575 65301 23584
rect 72363 23624 72405 23633
rect 72363 23584 72364 23624
rect 72404 23584 72405 23624
rect 72363 23575 72405 23584
rect 76099 23624 76157 23625
rect 76099 23584 76108 23624
rect 76148 23584 76157 23624
rect 76099 23583 76157 23584
rect 76867 23624 76925 23625
rect 76867 23584 76876 23624
rect 76916 23584 76925 23624
rect 76867 23583 76925 23584
rect 77163 23624 77205 23633
rect 77163 23584 77164 23624
rect 77204 23584 77205 23624
rect 77163 23575 77205 23584
rect 78699 23624 78741 23633
rect 78699 23584 78700 23624
rect 78740 23584 78741 23624
rect 78699 23575 78741 23584
rect 79083 23624 79125 23633
rect 79083 23584 79084 23624
rect 79124 23584 79125 23624
rect 79083 23575 79125 23584
rect 43371 23526 43372 23566
rect 43412 23526 43413 23566
rect 43371 23517 43413 23526
rect 576 23456 79584 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 79584 23456
rect 576 23392 79584 23416
rect 36843 23292 36885 23301
rect 33763 23288 33821 23289
rect 33763 23248 33772 23288
rect 33812 23248 33821 23288
rect 33763 23247 33821 23248
rect 36843 23252 36844 23292
rect 36884 23252 36885 23292
rect 36843 23243 36885 23252
rect 39811 23288 39869 23289
rect 39811 23248 39820 23288
rect 39860 23248 39869 23288
rect 39811 23247 39869 23248
rect 42403 23288 42461 23289
rect 42403 23248 42412 23288
rect 42452 23248 42461 23288
rect 42403 23247 42461 23248
rect 43371 23288 43413 23297
rect 43371 23248 43372 23288
rect 43412 23248 43413 23288
rect 43371 23239 43413 23248
rect 43843 23288 43901 23289
rect 43843 23248 43852 23288
rect 43892 23248 43901 23288
rect 43843 23247 43901 23248
rect 45003 23288 45045 23297
rect 45003 23248 45004 23288
rect 45044 23248 45045 23288
rect 45003 23239 45045 23248
rect 48835 23288 48893 23289
rect 48835 23248 48844 23288
rect 48884 23248 48893 23288
rect 48835 23247 48893 23248
rect 50283 23288 50325 23297
rect 50283 23248 50284 23288
rect 50324 23248 50325 23288
rect 50283 23239 50325 23248
rect 50859 23288 50901 23297
rect 50859 23248 50860 23288
rect 50900 23248 50901 23288
rect 50859 23239 50901 23248
rect 52395 23204 52437 23213
rect 52395 23164 52396 23204
rect 52436 23164 52437 23204
rect 52395 23155 52437 23164
rect 42795 23141 42837 23150
rect 1515 23120 1557 23129
rect 1515 23080 1516 23120
rect 1556 23080 1557 23120
rect 1515 23071 1557 23080
rect 1707 23120 1749 23129
rect 1707 23080 1708 23120
rect 1748 23080 1749 23120
rect 1707 23071 1749 23080
rect 34915 23120 34973 23121
rect 34915 23080 34924 23120
rect 34964 23080 34973 23120
rect 34915 23079 34973 23080
rect 35779 23120 35837 23121
rect 35779 23080 35788 23120
rect 35828 23080 35837 23120
rect 35779 23079 35837 23080
rect 36171 23120 36213 23129
rect 36171 23080 36172 23120
rect 36212 23080 36213 23120
rect 36171 23071 36213 23080
rect 36651 23120 36693 23129
rect 36651 23080 36652 23120
rect 36692 23080 36693 23120
rect 36651 23071 36693 23080
rect 36739 23120 36797 23121
rect 36739 23080 36748 23120
rect 36788 23080 36797 23120
rect 36739 23079 36797 23080
rect 37027 23120 37085 23121
rect 37027 23080 37036 23120
rect 37076 23080 37085 23120
rect 37027 23079 37085 23080
rect 37419 23120 37461 23129
rect 37419 23080 37420 23120
rect 37460 23080 37461 23120
rect 37419 23071 37461 23080
rect 37795 23120 37853 23121
rect 37795 23080 37804 23120
rect 37844 23080 37853 23120
rect 37795 23079 37853 23080
rect 38659 23120 38717 23121
rect 38659 23080 38668 23120
rect 38708 23080 38717 23120
rect 38659 23079 38717 23080
rect 40011 23120 40053 23129
rect 40011 23080 40012 23120
rect 40052 23080 40053 23120
rect 40011 23071 40053 23080
rect 40387 23120 40445 23121
rect 40387 23080 40396 23120
rect 40436 23080 40445 23120
rect 40387 23079 40445 23080
rect 41251 23120 41309 23121
rect 41251 23080 41260 23120
rect 41300 23080 41309 23120
rect 41251 23079 41309 23080
rect 42603 23120 42645 23129
rect 42603 23080 42604 23120
rect 42644 23080 42645 23120
rect 42603 23071 42645 23080
rect 42699 23120 42741 23129
rect 42699 23080 42700 23120
rect 42740 23080 42741 23120
rect 42795 23101 42796 23141
rect 42836 23101 42837 23141
rect 42795 23092 42837 23101
rect 42891 23120 42933 23129
rect 42699 23071 42741 23080
rect 42891 23080 42892 23120
rect 42932 23080 42933 23120
rect 42891 23071 42933 23080
rect 43075 23120 43133 23121
rect 43075 23080 43084 23120
rect 43124 23080 43133 23120
rect 43075 23079 43133 23080
rect 43459 23120 43517 23121
rect 43459 23080 43468 23120
rect 43508 23080 43517 23120
rect 43459 23079 43517 23080
rect 43947 23120 43989 23129
rect 43947 23080 43948 23120
rect 43988 23080 43989 23120
rect 43947 23071 43989 23080
rect 44043 23120 44085 23129
rect 44043 23080 44044 23120
rect 44084 23080 44085 23120
rect 44043 23071 44085 23080
rect 44139 23120 44181 23129
rect 44139 23080 44140 23120
rect 44180 23080 44181 23120
rect 44139 23071 44181 23080
rect 44899 23120 44957 23121
rect 44899 23080 44908 23120
rect 44948 23080 44957 23120
rect 44899 23079 44957 23080
rect 45963 23120 46005 23129
rect 45963 23080 45964 23120
rect 46004 23080 46005 23120
rect 45963 23071 46005 23080
rect 46059 23120 46101 23129
rect 46059 23080 46060 23120
rect 46100 23080 46101 23120
rect 46059 23071 46101 23080
rect 46155 23120 46197 23129
rect 46155 23080 46156 23120
rect 46196 23080 46197 23120
rect 46155 23071 46197 23080
rect 46251 23120 46293 23129
rect 46251 23080 46252 23120
rect 46292 23080 46293 23120
rect 46251 23071 46293 23080
rect 46443 23120 46485 23129
rect 46443 23080 46444 23120
rect 46484 23080 46485 23120
rect 46443 23071 46485 23080
rect 46819 23120 46877 23121
rect 46819 23080 46828 23120
rect 46868 23080 46877 23120
rect 46819 23079 46877 23080
rect 47683 23120 47741 23121
rect 47683 23080 47692 23120
rect 47732 23080 47741 23120
rect 47683 23079 47741 23080
rect 49219 23120 49277 23121
rect 49219 23080 49228 23120
rect 49268 23080 49277 23120
rect 49219 23079 49277 23080
rect 49699 23120 49757 23121
rect 49699 23080 49708 23120
rect 49748 23080 49757 23120
rect 49699 23079 49757 23080
rect 50091 23120 50133 23129
rect 50091 23080 50092 23120
rect 50132 23080 50133 23120
rect 50091 23071 50133 23080
rect 52003 23120 52061 23121
rect 52003 23080 52012 23120
rect 52052 23080 52061 23120
rect 52003 23079 52061 23080
rect 52107 23120 52149 23129
rect 52107 23080 52108 23120
rect 52148 23080 52149 23120
rect 52107 23071 52149 23080
rect 52291 23120 52349 23121
rect 52291 23080 52300 23120
rect 52340 23080 52349 23120
rect 52291 23079 52349 23080
rect 52675 23120 52733 23121
rect 52675 23080 52684 23120
rect 52724 23080 52733 23120
rect 52675 23079 52733 23080
rect 643 23036 701 23037
rect 643 22996 652 23036
rect 692 22996 701 23036
rect 643 22995 701 22996
rect 1611 23036 1653 23045
rect 1611 22996 1612 23036
rect 1652 22996 1653 23036
rect 1611 22987 1653 22996
rect 49323 23036 49365 23045
rect 49323 22996 49324 23036
rect 49364 22996 49365 23036
rect 49323 22987 49365 22996
rect 49803 23036 49845 23045
rect 49803 22996 49804 23036
rect 49844 22996 49845 23036
rect 49803 22987 49845 22996
rect 49995 23036 50037 23045
rect 49995 22996 49996 23036
rect 50036 22996 50037 23036
rect 49995 22987 50037 22996
rect 50467 23036 50525 23037
rect 50467 22996 50476 23036
rect 50516 22996 50525 23036
rect 50467 22995 50525 22996
rect 50659 23036 50717 23037
rect 50659 22996 50668 23036
rect 50708 22996 50717 23036
rect 50659 22995 50717 22996
rect 51523 23036 51581 23037
rect 51523 22996 51532 23036
rect 51572 22996 51581 23036
rect 51523 22995 51581 22996
rect 843 22952 885 22961
rect 843 22912 844 22952
rect 884 22912 885 22952
rect 843 22903 885 22912
rect 49899 22952 49941 22961
rect 49899 22912 49900 22952
rect 49940 22912 49941 22952
rect 49899 22903 49941 22912
rect 36363 22868 36405 22877
rect 36363 22828 36364 22868
rect 36404 22828 36405 22868
rect 36363 22819 36405 22828
rect 37131 22868 37173 22877
rect 37131 22828 37132 22868
rect 37172 22828 37173 22868
rect 37131 22819 37173 22828
rect 43179 22868 43221 22877
rect 43179 22828 43180 22868
rect 43220 22828 43221 22868
rect 43179 22819 43221 22828
rect 48835 22868 48893 22869
rect 48835 22828 48844 22868
rect 48884 22828 48893 22868
rect 48835 22827 48893 22828
rect 51339 22868 51381 22877
rect 51339 22828 51340 22868
rect 51380 22828 51381 22868
rect 51339 22819 51381 22828
rect 52587 22868 52629 22877
rect 52587 22828 52588 22868
rect 52628 22828 52629 22868
rect 52587 22819 52629 22828
rect 576 22700 52800 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 52800 22700
rect 576 22636 52800 22660
rect 42027 22574 42069 22583
rect 31083 22532 31125 22541
rect 31083 22492 31084 22532
rect 31124 22492 31125 22532
rect 31083 22483 31125 22492
rect 32043 22532 32085 22541
rect 32043 22492 32044 22532
rect 32084 22492 32085 22532
rect 32043 22483 32085 22492
rect 37803 22532 37845 22541
rect 37803 22492 37804 22532
rect 37844 22492 37845 22532
rect 37803 22483 37845 22492
rect 39435 22532 39477 22541
rect 39435 22492 39436 22532
rect 39476 22492 39477 22532
rect 42027 22534 42028 22574
rect 42068 22534 42069 22574
rect 42027 22525 42069 22534
rect 43467 22532 43509 22541
rect 39435 22483 39477 22492
rect 43467 22492 43468 22532
rect 43508 22492 43509 22532
rect 43467 22483 43509 22492
rect 46443 22532 46485 22541
rect 46443 22492 46444 22532
rect 46484 22492 46485 22532
rect 46443 22483 46485 22492
rect 47115 22532 47157 22541
rect 47115 22492 47116 22532
rect 47156 22492 47157 22532
rect 47115 22483 47157 22492
rect 52387 22532 52445 22533
rect 52387 22492 52396 22532
rect 52436 22492 52445 22532
rect 52387 22491 52445 22492
rect 52683 22532 52725 22541
rect 52683 22492 52684 22532
rect 52724 22492 52725 22532
rect 52683 22483 52725 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 36171 22448 36213 22457
rect 36171 22408 36172 22448
rect 36212 22408 36213 22448
rect 36171 22399 36213 22408
rect 41643 22448 41685 22457
rect 41643 22408 41644 22448
rect 41684 22408 41685 22448
rect 41643 22399 41685 22408
rect 42891 22448 42933 22457
rect 42891 22408 42892 22448
rect 42932 22408 42933 22448
rect 42891 22399 42933 22408
rect 49323 22448 49365 22457
rect 49323 22408 49324 22448
rect 49364 22408 49365 22448
rect 49323 22399 49365 22408
rect 31267 22364 31325 22365
rect 31267 22324 31276 22364
rect 31316 22324 31325 22364
rect 31267 22323 31325 22324
rect 32227 22364 32285 22365
rect 32227 22324 32236 22364
rect 32276 22324 32285 22364
rect 32227 22323 32285 22324
rect 33283 22364 33341 22365
rect 33283 22324 33292 22364
rect 33332 22324 33341 22364
rect 33283 22323 33341 22324
rect 36075 22364 36117 22373
rect 36075 22324 36076 22364
rect 36116 22324 36117 22364
rect 36075 22315 36117 22324
rect 36267 22364 36309 22373
rect 36267 22324 36268 22364
rect 36308 22324 36309 22364
rect 36267 22315 36309 22324
rect 41547 22364 41589 22373
rect 41547 22324 41548 22364
rect 41588 22324 41589 22364
rect 41547 22315 41589 22324
rect 41739 22364 41781 22373
rect 41739 22324 41740 22364
rect 41780 22324 41781 22364
rect 41739 22315 41781 22324
rect 7939 22280 7997 22281
rect 7939 22240 7948 22280
rect 7988 22240 7997 22280
rect 7939 22239 7997 22240
rect 31563 22280 31605 22289
rect 31563 22240 31564 22280
rect 31604 22240 31605 22280
rect 31563 22231 31605 22240
rect 31659 22280 31701 22289
rect 31659 22240 31660 22280
rect 31700 22240 31701 22280
rect 31659 22231 31701 22240
rect 31755 22280 31797 22289
rect 31755 22240 31756 22280
rect 31796 22240 31797 22280
rect 31755 22231 31797 22240
rect 35499 22280 35541 22289
rect 35499 22240 35500 22280
rect 35540 22240 35541 22280
rect 35499 22231 35541 22240
rect 35691 22280 35733 22289
rect 35691 22240 35692 22280
rect 35732 22240 35733 22280
rect 35691 22231 35733 22240
rect 35779 22280 35837 22281
rect 35779 22240 35788 22280
rect 35828 22240 35837 22280
rect 35779 22239 35837 22240
rect 35979 22280 36021 22289
rect 35979 22240 35980 22280
rect 36020 22240 36021 22280
rect 35979 22231 36021 22240
rect 36355 22280 36413 22281
rect 36355 22240 36364 22280
rect 36404 22240 36413 22280
rect 36355 22239 36413 22240
rect 36939 22280 36981 22289
rect 36939 22240 36940 22280
rect 36980 22240 36981 22280
rect 36939 22231 36981 22240
rect 37035 22280 37077 22289
rect 37035 22240 37036 22280
rect 37076 22240 37077 22280
rect 37035 22231 37077 22240
rect 37131 22280 37173 22289
rect 37131 22240 37132 22280
rect 37172 22240 37173 22280
rect 37131 22231 37173 22240
rect 37227 22280 37269 22289
rect 37227 22240 37228 22280
rect 37268 22240 37269 22280
rect 37227 22231 37269 22240
rect 37507 22280 37565 22281
rect 37507 22240 37516 22280
rect 37556 22240 37565 22280
rect 37507 22239 37565 22240
rect 37699 22280 37757 22281
rect 37699 22240 37708 22280
rect 37748 22240 37757 22280
rect 37699 22239 37757 22240
rect 39523 22280 39581 22281
rect 39523 22240 39532 22280
rect 39572 22240 39581 22280
rect 39523 22239 39581 22240
rect 41451 22280 41493 22289
rect 41451 22240 41452 22280
rect 41492 22240 41493 22280
rect 41451 22231 41493 22240
rect 41827 22280 41885 22281
rect 41827 22240 41836 22280
rect 41876 22240 41885 22280
rect 41827 22239 41885 22240
rect 42315 22280 42357 22289
rect 42315 22240 42316 22280
rect 42356 22240 42357 22280
rect 42315 22231 42357 22240
rect 42403 22280 42461 22281
rect 42403 22240 42412 22280
rect 42452 22240 42461 22280
rect 42403 22239 42461 22240
rect 42891 22280 42933 22289
rect 42891 22240 42892 22280
rect 42932 22240 42933 22280
rect 42891 22231 42933 22240
rect 43083 22280 43125 22289
rect 43083 22240 43084 22280
rect 43124 22240 43125 22280
rect 43083 22231 43125 22240
rect 43197 22273 43239 22282
rect 43197 22233 43198 22273
rect 43238 22233 43239 22273
rect 43363 22280 43421 22281
rect 43363 22240 43372 22280
rect 43412 22240 43421 22280
rect 43363 22239 43421 22240
rect 44995 22280 45053 22281
rect 44995 22240 45004 22280
rect 45044 22240 45053 22280
rect 44995 22239 45053 22240
rect 45859 22280 45917 22281
rect 45859 22240 45868 22280
rect 45908 22240 45917 22280
rect 45859 22239 45917 22240
rect 46731 22280 46773 22289
rect 46731 22240 46732 22280
rect 46772 22240 46773 22280
rect 43197 22224 43239 22233
rect 46731 22231 46773 22240
rect 46819 22280 46877 22281
rect 46819 22240 46828 22280
rect 46868 22240 46877 22280
rect 46819 22239 46877 22240
rect 47203 22280 47261 22281
rect 47203 22240 47212 22280
rect 47252 22240 47261 22280
rect 47203 22239 47261 22240
rect 47403 22280 47445 22289
rect 47403 22240 47404 22280
rect 47444 22240 47445 22280
rect 47403 22231 47445 22240
rect 47595 22280 47637 22289
rect 47595 22240 47596 22280
rect 47636 22240 47637 22280
rect 47595 22231 47637 22240
rect 47683 22280 47741 22281
rect 47683 22240 47692 22280
rect 47732 22240 47741 22280
rect 47683 22239 47741 22240
rect 49611 22280 49653 22289
rect 49611 22240 49612 22280
rect 49652 22240 49653 22280
rect 49611 22231 49653 22240
rect 49699 22280 49757 22281
rect 49699 22240 49708 22280
rect 49748 22240 49757 22280
rect 49699 22239 49757 22240
rect 50371 22280 50429 22281
rect 50371 22240 50380 22280
rect 50420 22240 50429 22280
rect 50371 22239 50429 22240
rect 51235 22280 51293 22281
rect 51235 22240 51244 22280
rect 51284 22240 51293 22280
rect 51235 22239 51293 22240
rect 52579 22280 52637 22281
rect 52579 22240 52588 22280
rect 52628 22240 52637 22280
rect 52579 22239 52637 22240
rect 46251 22196 46293 22205
rect 46251 22156 46252 22196
rect 46292 22156 46293 22196
rect 46251 22147 46293 22156
rect 49995 22196 50037 22205
rect 49995 22156 49996 22196
rect 50036 22156 50037 22196
rect 49995 22147 50037 22156
rect 31083 22112 31125 22121
rect 31083 22072 31084 22112
rect 31124 22072 31125 22112
rect 31083 22063 31125 22072
rect 31459 22112 31517 22113
rect 31459 22072 31468 22112
rect 31508 22072 31517 22112
rect 31459 22071 31517 22072
rect 32043 22112 32085 22121
rect 32043 22072 32044 22112
rect 32084 22072 32085 22112
rect 32043 22063 32085 22072
rect 33483 22112 33525 22121
rect 33483 22072 33484 22112
rect 33524 22072 33525 22112
rect 33483 22063 33525 22072
rect 35587 22112 35645 22113
rect 35587 22072 35596 22112
rect 35636 22072 35645 22112
rect 35587 22071 35645 22072
rect 37419 22112 37461 22121
rect 37419 22072 37420 22112
rect 37460 22072 37461 22112
rect 37419 22063 37461 22072
rect 37803 22112 37845 22121
rect 37803 22072 37804 22112
rect 37844 22072 37845 22112
rect 37803 22063 37845 22072
rect 39435 22112 39477 22121
rect 39435 22072 39436 22112
rect 39476 22072 39477 22112
rect 39435 22063 39477 22072
rect 42507 22108 42549 22117
rect 42507 22068 42508 22108
rect 42548 22068 42549 22108
rect 43843 22112 43901 22113
rect 43843 22072 43852 22112
rect 43892 22072 43901 22112
rect 43843 22071 43901 22072
rect 47491 22112 47549 22113
rect 47491 22072 47500 22112
rect 47540 22072 47549 22112
rect 47491 22071 47549 22072
rect 52387 22112 52445 22113
rect 52387 22072 52396 22112
rect 52436 22072 52445 22112
rect 52387 22071 52445 22072
rect 42507 22059 42549 22068
rect 46923 22054 46965 22063
rect 46923 22014 46924 22054
rect 46964 22014 46965 22054
rect 46923 22005 46965 22014
rect 49803 22054 49845 22063
rect 49803 22014 49804 22054
rect 49844 22014 49845 22054
rect 49803 22005 49845 22014
rect 576 21944 52800 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 52800 21944
rect 576 21880 52800 21904
rect 36075 21780 36117 21789
rect 36075 21740 36076 21780
rect 36116 21740 36117 21780
rect 36075 21731 36117 21740
rect 42115 21776 42173 21777
rect 42115 21736 42124 21776
rect 42164 21736 42173 21776
rect 42115 21735 42173 21736
rect 44995 21776 45053 21777
rect 44995 21736 45004 21776
rect 45044 21736 45053 21776
rect 44995 21735 45053 21736
rect 46723 21776 46781 21777
rect 46723 21736 46732 21776
rect 46772 21736 46781 21776
rect 46723 21735 46781 21736
rect 49987 21776 50045 21777
rect 49987 21736 49996 21776
rect 50036 21736 50045 21776
rect 49987 21735 50045 21736
rect 30891 21692 30933 21701
rect 30891 21652 30892 21692
rect 30932 21652 30933 21692
rect 30891 21643 30933 21652
rect 37227 21692 37269 21701
rect 37227 21652 37228 21692
rect 37268 21652 37269 21692
rect 37227 21643 37269 21652
rect 37419 21692 37461 21701
rect 37419 21652 37420 21692
rect 37460 21652 37461 21692
rect 42603 21692 42645 21701
rect 37419 21643 37461 21652
rect 40299 21650 40341 21659
rect 3723 21608 3765 21617
rect 3723 21568 3724 21608
rect 3764 21568 3765 21608
rect 3723 21559 3765 21568
rect 3819 21608 3861 21617
rect 3819 21568 3820 21608
rect 3860 21568 3861 21608
rect 3819 21559 3861 21568
rect 3915 21608 3957 21617
rect 3915 21568 3916 21608
rect 3956 21568 3957 21608
rect 3915 21559 3957 21568
rect 4011 21608 4053 21617
rect 4011 21568 4012 21608
rect 4052 21568 4053 21608
rect 4011 21559 4053 21568
rect 4491 21608 4533 21617
rect 4491 21568 4492 21608
rect 4532 21568 4533 21608
rect 4491 21559 4533 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 4683 21608 4725 21617
rect 4683 21568 4684 21608
rect 4724 21568 4725 21608
rect 4683 21559 4725 21568
rect 4779 21608 4821 21617
rect 4779 21568 4780 21608
rect 4820 21568 4821 21608
rect 4779 21559 4821 21568
rect 4971 21608 5013 21617
rect 4971 21568 4972 21608
rect 5012 21568 5013 21608
rect 4971 21559 5013 21568
rect 5347 21608 5405 21609
rect 5347 21568 5356 21608
rect 5396 21568 5405 21608
rect 5347 21567 5405 21568
rect 6211 21608 6269 21609
rect 6211 21568 6220 21608
rect 6260 21568 6269 21608
rect 6211 21567 6269 21568
rect 7755 21608 7797 21617
rect 7755 21568 7756 21608
rect 7796 21568 7797 21608
rect 7755 21559 7797 21568
rect 8131 21608 8189 21609
rect 8131 21568 8140 21608
rect 8180 21568 8189 21608
rect 8131 21567 8189 21568
rect 8995 21608 9053 21609
rect 8995 21568 9004 21608
rect 9044 21568 9053 21608
rect 8995 21567 9053 21568
rect 11211 21608 11253 21617
rect 11211 21568 11212 21608
rect 11252 21568 11253 21608
rect 11211 21559 11253 21568
rect 11587 21608 11645 21609
rect 11587 21568 11596 21608
rect 11636 21568 11645 21608
rect 11587 21567 11645 21568
rect 12451 21608 12509 21609
rect 12451 21568 12460 21608
rect 12500 21568 12509 21608
rect 12451 21567 12509 21568
rect 31267 21608 31325 21609
rect 31267 21568 31276 21608
rect 31316 21568 31325 21608
rect 31267 21567 31325 21568
rect 32131 21608 32189 21609
rect 32131 21568 32140 21608
rect 32180 21568 32189 21608
rect 32131 21567 32189 21568
rect 34627 21608 34685 21609
rect 34627 21568 34636 21608
rect 34676 21568 34685 21608
rect 34627 21567 34685 21568
rect 35491 21608 35549 21609
rect 35491 21568 35500 21608
rect 35540 21568 35549 21608
rect 35491 21567 35549 21568
rect 35883 21608 35925 21617
rect 35883 21568 35884 21608
rect 35924 21568 35925 21608
rect 35883 21559 35925 21568
rect 36163 21608 36221 21609
rect 36163 21568 36172 21608
rect 36212 21568 36221 21608
rect 36163 21567 36221 21568
rect 36267 21608 36309 21617
rect 36267 21568 36268 21608
rect 36308 21568 36309 21608
rect 36267 21559 36309 21568
rect 36939 21608 36981 21617
rect 36939 21568 36940 21608
rect 36980 21568 36981 21608
rect 36939 21559 36981 21568
rect 37035 21608 37077 21617
rect 37035 21568 37036 21608
rect 37076 21568 37077 21608
rect 37035 21559 37077 21568
rect 37131 21608 37173 21617
rect 37131 21568 37132 21608
rect 37172 21568 37173 21608
rect 37131 21559 37173 21568
rect 37795 21608 37853 21609
rect 37795 21568 37804 21608
rect 37844 21568 37853 21608
rect 37795 21567 37853 21568
rect 38659 21608 38717 21609
rect 38659 21568 38668 21608
rect 38708 21568 38717 21608
rect 38659 21567 38717 21568
rect 40003 21608 40061 21609
rect 40003 21568 40012 21608
rect 40052 21568 40061 21608
rect 40003 21567 40061 21568
rect 40107 21608 40149 21617
rect 40107 21568 40108 21608
rect 40148 21568 40149 21608
rect 40299 21610 40300 21650
rect 40340 21610 40341 21650
rect 42603 21652 42604 21692
rect 42644 21652 42645 21692
rect 42603 21643 42645 21652
rect 49803 21692 49845 21701
rect 49803 21652 49804 21692
rect 49844 21652 49845 21692
rect 49803 21643 49845 21652
rect 40299 21601 40341 21610
rect 42219 21608 42261 21617
rect 40107 21559 40149 21568
rect 42219 21568 42220 21608
rect 42260 21568 42261 21608
rect 42219 21559 42261 21568
rect 42315 21608 42357 21617
rect 42315 21568 42316 21608
rect 42356 21568 42357 21608
rect 42315 21559 42357 21568
rect 42411 21608 42453 21617
rect 42411 21568 42412 21608
rect 42452 21568 42453 21608
rect 42411 21559 42453 21568
rect 42979 21608 43037 21609
rect 42979 21568 42988 21608
rect 43028 21568 43037 21608
rect 42979 21567 43037 21568
rect 43843 21608 43901 21609
rect 43843 21568 43852 21608
rect 43892 21568 43901 21608
rect 43843 21567 43901 21568
rect 45859 21608 45917 21609
rect 45859 21568 45868 21608
rect 45908 21568 45917 21608
rect 45859 21567 45917 21568
rect 45963 21608 46005 21617
rect 45963 21568 45964 21608
rect 46004 21568 46005 21608
rect 45963 21559 46005 21568
rect 46147 21608 46205 21609
rect 46147 21568 46156 21608
rect 46196 21568 46205 21608
rect 46147 21567 46205 21568
rect 46539 21608 46581 21617
rect 46539 21568 46540 21608
rect 46580 21568 46581 21608
rect 46539 21559 46581 21568
rect 46827 21608 46869 21617
rect 46827 21568 46828 21608
rect 46868 21568 46869 21608
rect 46827 21559 46869 21568
rect 46923 21608 46965 21617
rect 46923 21568 46924 21608
rect 46964 21568 46965 21608
rect 46923 21559 46965 21568
rect 47019 21608 47061 21617
rect 47019 21568 47020 21608
rect 47060 21568 47061 21608
rect 47019 21559 47061 21568
rect 48547 21608 48605 21609
rect 48547 21568 48556 21608
rect 48596 21568 48605 21608
rect 48547 21567 48605 21568
rect 49411 21608 49469 21609
rect 49411 21568 49420 21608
rect 49460 21568 49469 21608
rect 49411 21567 49469 21568
rect 50091 21608 50133 21617
rect 50091 21568 50092 21608
rect 50132 21568 50133 21608
rect 50091 21559 50133 21568
rect 50187 21608 50229 21617
rect 50187 21568 50188 21608
rect 50228 21568 50229 21608
rect 50187 21559 50229 21568
rect 50283 21608 50325 21617
rect 50283 21568 50284 21608
rect 50324 21568 50325 21608
rect 50283 21559 50325 21568
rect 50475 21608 50517 21617
rect 50475 21568 50476 21608
rect 50516 21568 50517 21608
rect 50475 21559 50517 21568
rect 50571 21608 50613 21617
rect 50571 21568 50572 21608
rect 50612 21568 50613 21608
rect 50571 21559 50613 21568
rect 50667 21608 50709 21617
rect 50667 21568 50668 21608
rect 50708 21568 50709 21608
rect 50667 21559 50709 21568
rect 50763 21608 50805 21617
rect 50763 21568 50764 21608
rect 50804 21568 50805 21608
rect 50763 21559 50805 21568
rect 51235 21608 51293 21609
rect 51235 21568 51244 21608
rect 51284 21568 51293 21608
rect 51235 21567 51293 21568
rect 51523 21608 51581 21609
rect 51523 21568 51532 21608
rect 51572 21568 51581 21608
rect 51523 21567 51581 21568
rect 51811 21608 51869 21609
rect 51811 21568 51820 21608
rect 51860 21568 51869 21608
rect 51811 21567 51869 21568
rect 52195 21608 52253 21609
rect 52195 21568 52204 21608
rect 52244 21568 52253 21608
rect 52195 21567 52253 21568
rect 52483 21608 52541 21609
rect 52483 21568 52492 21608
rect 52532 21568 52541 21608
rect 52483 21567 52541 21568
rect 3331 21524 3389 21525
rect 3331 21484 3340 21524
rect 3380 21484 3389 21524
rect 3331 21483 3389 21484
rect 7371 21524 7413 21533
rect 7371 21484 7372 21524
rect 7412 21484 7413 21524
rect 7371 21475 7413 21484
rect 29731 21524 29789 21525
rect 29731 21484 29740 21524
rect 29780 21484 29789 21524
rect 29731 21483 29789 21484
rect 30115 21524 30173 21525
rect 30115 21484 30124 21524
rect 30164 21484 30173 21524
rect 30115 21483 30173 21484
rect 30499 21524 30557 21525
rect 30499 21484 30508 21524
rect 30548 21484 30557 21524
rect 30499 21483 30557 21484
rect 39819 21524 39861 21533
rect 39819 21484 39820 21524
rect 39860 21484 39861 21524
rect 39819 21475 39861 21484
rect 46251 21524 46293 21533
rect 46251 21484 46252 21524
rect 46292 21484 46293 21524
rect 46251 21475 46293 21484
rect 46443 21524 46485 21533
rect 46443 21484 46444 21524
rect 46484 21484 46485 21524
rect 46443 21475 46485 21484
rect 51147 21524 51189 21533
rect 51147 21484 51148 21524
rect 51188 21484 51189 21524
rect 51147 21475 51189 21484
rect 46347 21440 46389 21449
rect 46347 21400 46348 21440
rect 46388 21400 46389 21440
rect 46347 21391 46389 21400
rect 52587 21440 52629 21449
rect 52587 21400 52588 21440
rect 52628 21400 52629 21440
rect 52587 21391 52629 21400
rect 3531 21356 3573 21365
rect 3531 21316 3532 21356
rect 3572 21316 3573 21356
rect 3531 21307 3573 21316
rect 10147 21356 10205 21357
rect 10147 21316 10156 21356
rect 10196 21316 10205 21356
rect 10147 21315 10205 21316
rect 13603 21356 13661 21357
rect 13603 21316 13612 21356
rect 13652 21316 13661 21356
rect 13603 21315 13661 21316
rect 29931 21356 29973 21365
rect 29931 21316 29932 21356
rect 29972 21316 29973 21356
rect 29931 21307 29973 21316
rect 30315 21356 30357 21365
rect 30315 21316 30316 21356
rect 30356 21316 30357 21356
rect 30315 21307 30357 21316
rect 30699 21356 30741 21365
rect 30699 21316 30700 21356
rect 30740 21316 30741 21356
rect 30699 21307 30741 21316
rect 33283 21356 33341 21357
rect 33283 21316 33292 21356
rect 33332 21316 33341 21356
rect 33283 21315 33341 21316
rect 33475 21356 33533 21357
rect 33475 21316 33484 21356
rect 33524 21316 33533 21356
rect 33475 21315 33533 21316
rect 36555 21356 36597 21365
rect 36555 21316 36556 21356
rect 36596 21316 36597 21356
rect 36555 21307 36597 21316
rect 40299 21356 40341 21365
rect 40299 21316 40300 21356
rect 40340 21316 40341 21356
rect 40299 21307 40341 21316
rect 47395 21356 47453 21357
rect 47395 21316 47404 21356
rect 47444 21316 47453 21356
rect 47395 21315 47453 21316
rect 51627 21356 51669 21365
rect 51627 21316 51628 21356
rect 51668 21316 51669 21356
rect 51627 21307 51669 21316
rect 51915 21356 51957 21365
rect 51915 21316 51916 21356
rect 51956 21316 51957 21356
rect 51915 21307 51957 21316
rect 52299 21356 52341 21365
rect 52299 21316 52300 21356
rect 52340 21316 52341 21356
rect 52299 21307 52341 21316
rect 576 21188 52800 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 52800 21188
rect 576 21124 52800 21148
rect 7947 21020 7989 21029
rect 7947 20980 7948 21020
rect 7988 20980 7989 21020
rect 7947 20971 7989 20980
rect 33003 21020 33045 21029
rect 33003 20980 33004 21020
rect 33044 20980 33045 21020
rect 33003 20971 33045 20980
rect 43659 21020 43701 21029
rect 43659 20980 43660 21020
rect 43700 20980 43701 21020
rect 43659 20971 43701 20980
rect 49611 21020 49653 21029
rect 49611 20980 49612 21020
rect 49652 20980 49653 21020
rect 49611 20971 49653 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 3819 20936 3861 20945
rect 3819 20896 3820 20936
rect 3860 20896 3861 20936
rect 3819 20887 3861 20896
rect 6795 20936 6837 20945
rect 6795 20896 6796 20936
rect 6836 20896 6837 20936
rect 6795 20887 6837 20896
rect 10251 20936 10293 20945
rect 10251 20896 10252 20936
rect 10292 20896 10293 20936
rect 10251 20887 10293 20896
rect 32619 20936 32661 20945
rect 32619 20896 32620 20936
rect 32660 20896 32661 20936
rect 35691 20936 35733 20945
rect 32619 20887 32661 20896
rect 32715 20894 32757 20903
rect 1315 20852 1373 20853
rect 1315 20812 1324 20852
rect 1364 20812 1373 20852
rect 1315 20811 1373 20812
rect 2755 20852 2813 20853
rect 2755 20812 2764 20852
rect 2804 20812 2813 20852
rect 2755 20811 2813 20812
rect 3619 20852 3677 20853
rect 3619 20812 3628 20852
rect 3668 20812 3677 20852
rect 3619 20811 3677 20812
rect 6411 20852 6453 20861
rect 6411 20812 6412 20852
rect 6452 20812 6453 20852
rect 6411 20803 6453 20812
rect 6699 20852 6741 20861
rect 6699 20812 6700 20852
rect 6740 20812 6741 20852
rect 6699 20803 6741 20812
rect 6891 20852 6933 20861
rect 6891 20812 6892 20852
rect 6932 20812 6933 20852
rect 6891 20803 6933 20812
rect 10155 20852 10197 20861
rect 10155 20812 10156 20852
rect 10196 20812 10197 20852
rect 10155 20803 10197 20812
rect 10347 20852 10389 20861
rect 10347 20812 10348 20852
rect 10388 20812 10389 20852
rect 10347 20803 10389 20812
rect 16299 20852 16341 20861
rect 16299 20812 16300 20852
rect 16340 20812 16341 20852
rect 16299 20803 16341 20812
rect 29635 20852 29693 20853
rect 29635 20812 29644 20852
rect 29684 20812 29693 20852
rect 29635 20811 29693 20812
rect 32523 20852 32565 20861
rect 32523 20812 32524 20852
rect 32564 20812 32565 20852
rect 32715 20854 32716 20894
rect 32756 20854 32757 20894
rect 35691 20896 35692 20936
rect 35732 20896 35733 20936
rect 35691 20887 35733 20896
rect 52491 20936 52533 20945
rect 52491 20896 52492 20936
rect 52532 20896 52533 20936
rect 52491 20887 52533 20896
rect 32715 20845 32757 20854
rect 35595 20852 35637 20861
rect 32523 20803 32565 20812
rect 35595 20812 35596 20852
rect 35636 20812 35637 20852
rect 35595 20803 35637 20812
rect 35787 20852 35829 20861
rect 35787 20812 35788 20852
rect 35828 20812 35829 20852
rect 35787 20803 35829 20812
rect 37411 20852 37469 20853
rect 37411 20812 37420 20852
rect 37460 20812 37469 20852
rect 37411 20811 37469 20812
rect 40003 20852 40061 20853
rect 40003 20812 40012 20852
rect 40052 20812 40061 20852
rect 40003 20811 40061 20812
rect 42603 20852 42645 20861
rect 42603 20812 42604 20852
rect 42644 20812 42645 20852
rect 42603 20803 42645 20812
rect 43843 20852 43901 20853
rect 43843 20812 43852 20852
rect 43892 20812 43901 20852
rect 43843 20811 43901 20812
rect 46819 20852 46877 20853
rect 46819 20812 46828 20852
rect 46868 20812 46877 20852
rect 46819 20811 46877 20812
rect 49987 20852 50045 20853
rect 49987 20812 49996 20852
rect 50036 20812 50045 20852
rect 49987 20811 50045 20812
rect 50371 20852 50429 20853
rect 50371 20812 50380 20852
rect 50420 20812 50429 20852
rect 50371 20811 50429 20812
rect 50563 20852 50621 20853
rect 50563 20812 50572 20852
rect 50612 20812 50621 20852
rect 50563 20811 50621 20812
rect 3147 20768 3189 20777
rect 3147 20728 3148 20768
rect 3188 20728 3189 20768
rect 3147 20719 3189 20728
rect 3243 20768 3285 20777
rect 3243 20728 3244 20768
rect 3284 20728 3285 20768
rect 3243 20719 3285 20728
rect 3339 20768 3381 20777
rect 3339 20728 3340 20768
rect 3380 20728 3381 20768
rect 3339 20719 3381 20728
rect 4387 20768 4445 20769
rect 4387 20728 4396 20768
rect 4436 20728 4445 20768
rect 4387 20727 4445 20728
rect 5251 20768 5309 20769
rect 5251 20728 5260 20768
rect 5300 20728 5309 20768
rect 5251 20727 5309 20728
rect 6595 20768 6653 20769
rect 6595 20728 6604 20768
rect 6644 20728 6653 20768
rect 6595 20727 6653 20728
rect 6987 20768 7029 20777
rect 6987 20728 6988 20768
rect 7028 20728 7029 20768
rect 6987 20719 7029 20728
rect 7459 20768 7517 20769
rect 7459 20728 7468 20768
rect 7508 20728 7517 20768
rect 7459 20727 7517 20728
rect 8419 20768 8477 20769
rect 8419 20728 8428 20768
rect 8468 20728 8477 20768
rect 8419 20727 8477 20728
rect 9763 20768 9821 20769
rect 9763 20728 9772 20768
rect 9812 20728 9821 20768
rect 9763 20727 9821 20728
rect 10051 20768 10109 20769
rect 10051 20728 10060 20768
rect 10100 20728 10109 20768
rect 10051 20727 10109 20728
rect 10443 20768 10485 20777
rect 10443 20728 10444 20768
rect 10484 20728 10485 20768
rect 10443 20719 10485 20728
rect 10827 20768 10869 20777
rect 10827 20728 10828 20768
rect 10868 20728 10869 20768
rect 10827 20719 10869 20728
rect 10923 20768 10965 20777
rect 10923 20728 10924 20768
rect 10964 20728 10965 20768
rect 10923 20719 10965 20728
rect 11019 20768 11061 20777
rect 11019 20728 11020 20768
rect 11060 20728 11061 20768
rect 11019 20719 11061 20728
rect 11115 20768 11157 20777
rect 11115 20728 11116 20768
rect 11156 20728 11157 20768
rect 11115 20719 11157 20728
rect 13515 20768 13557 20777
rect 13515 20728 13516 20768
rect 13556 20728 13557 20768
rect 13515 20719 13557 20728
rect 13611 20768 13653 20777
rect 13611 20728 13612 20768
rect 13652 20728 13653 20768
rect 13611 20719 13653 20728
rect 13707 20768 13749 20777
rect 13707 20728 13708 20768
rect 13748 20728 13749 20768
rect 13707 20719 13749 20728
rect 14275 20768 14333 20769
rect 14275 20728 14284 20768
rect 14324 20728 14333 20768
rect 14275 20727 14333 20728
rect 15139 20768 15197 20769
rect 15139 20728 15148 20768
rect 15188 20728 15197 20768
rect 15139 20727 15197 20728
rect 30979 20768 31037 20769
rect 30979 20728 30988 20768
rect 31028 20728 31037 20768
rect 30979 20727 31037 20728
rect 31843 20768 31901 20769
rect 31843 20728 31852 20768
rect 31892 20728 31901 20768
rect 31843 20727 31901 20728
rect 32235 20768 32277 20777
rect 32235 20728 32236 20768
rect 32276 20728 32277 20768
rect 32235 20719 32277 20728
rect 32419 20768 32477 20769
rect 32419 20728 32428 20768
rect 32468 20728 32477 20768
rect 32419 20727 32477 20728
rect 32811 20768 32853 20777
rect 32811 20728 32812 20768
rect 32852 20728 32853 20768
rect 32811 20719 32853 20728
rect 33003 20768 33045 20777
rect 33003 20728 33004 20768
rect 33044 20728 33045 20768
rect 33003 20719 33045 20728
rect 33195 20768 33237 20777
rect 33195 20728 33196 20768
rect 33236 20728 33237 20768
rect 33195 20719 33237 20728
rect 33283 20768 33341 20769
rect 33283 20728 33292 20768
rect 33332 20728 33341 20768
rect 33283 20727 33341 20728
rect 35203 20768 35261 20769
rect 35203 20728 35212 20768
rect 35252 20728 35261 20768
rect 35203 20727 35261 20728
rect 35499 20768 35541 20777
rect 35499 20728 35500 20768
rect 35540 20728 35541 20768
rect 35499 20719 35541 20728
rect 35875 20768 35933 20769
rect 35875 20728 35884 20768
rect 35924 20728 35933 20768
rect 35875 20727 35933 20728
rect 36747 20768 36789 20777
rect 36747 20728 36748 20768
rect 36788 20728 36789 20768
rect 36747 20719 36789 20728
rect 36843 20768 36885 20777
rect 36843 20728 36844 20768
rect 36884 20728 36885 20768
rect 36843 20719 36885 20728
rect 36939 20768 36981 20777
rect 36939 20728 36940 20768
rect 36980 20728 36981 20768
rect 36939 20719 36981 20728
rect 37035 20768 37077 20777
rect 37035 20728 37036 20768
rect 37076 20728 37077 20768
rect 37035 20719 37077 20728
rect 40579 20768 40637 20769
rect 40579 20728 40588 20768
rect 40628 20728 40637 20768
rect 40579 20727 40637 20728
rect 41443 20768 41501 20769
rect 41443 20728 41452 20768
rect 41492 20728 41501 20768
rect 41443 20727 41501 20728
rect 42883 20768 42941 20769
rect 42883 20728 42892 20768
rect 42932 20728 42941 20768
rect 42883 20727 42941 20728
rect 47203 20768 47261 20769
rect 47203 20728 47212 20768
rect 47252 20728 47261 20768
rect 47203 20727 47261 20728
rect 48843 20768 48885 20777
rect 48843 20728 48844 20768
rect 48884 20728 48885 20768
rect 48843 20719 48885 20728
rect 49131 20768 49173 20777
rect 49131 20728 49132 20768
rect 49172 20728 49173 20768
rect 49131 20719 49173 20728
rect 49507 20768 49565 20769
rect 49507 20728 49516 20768
rect 49556 20728 49565 20768
rect 49507 20727 49565 20728
rect 52195 20768 52253 20769
rect 52195 20728 52204 20768
rect 52244 20728 52253 20768
rect 52195 20727 52253 20728
rect 52579 20768 52637 20769
rect 52579 20728 52588 20768
rect 52628 20728 52637 20768
rect 52579 20727 52637 20728
rect 4011 20684 4053 20693
rect 4011 20644 4012 20684
rect 4052 20644 4053 20684
rect 4011 20635 4053 20644
rect 13899 20684 13941 20693
rect 13899 20644 13900 20684
rect 13940 20644 13941 20684
rect 13899 20635 13941 20644
rect 40203 20684 40245 20693
rect 40203 20644 40204 20684
rect 40244 20644 40245 20684
rect 40203 20635 40245 20644
rect 1515 20600 1557 20609
rect 1515 20560 1516 20600
rect 1556 20560 1557 20600
rect 1515 20551 1557 20560
rect 2955 20600 2997 20609
rect 2955 20560 2956 20600
rect 2996 20560 2997 20600
rect 2955 20551 2997 20560
rect 3427 20600 3485 20601
rect 3427 20560 3436 20600
rect 3476 20560 3485 20600
rect 3427 20559 3485 20560
rect 9867 20600 9909 20609
rect 9867 20560 9868 20600
rect 9908 20560 9909 20600
rect 9867 20551 9909 20560
rect 13411 20600 13469 20601
rect 13411 20560 13420 20600
rect 13460 20560 13469 20600
rect 13411 20559 13469 20560
rect 29451 20600 29493 20609
rect 29451 20560 29452 20600
rect 29492 20560 29493 20600
rect 29451 20551 29493 20560
rect 29827 20600 29885 20601
rect 29827 20560 29836 20600
rect 29876 20560 29885 20600
rect 29827 20559 29885 20560
rect 35307 20600 35349 20609
rect 35307 20560 35308 20600
rect 35348 20560 35349 20600
rect 35307 20551 35349 20560
rect 37611 20600 37653 20609
rect 37611 20560 37612 20600
rect 37652 20560 37653 20600
rect 37611 20551 37653 20560
rect 39819 20600 39861 20609
rect 39819 20560 39820 20600
rect 39860 20560 39861 20600
rect 39819 20551 39861 20560
rect 42795 20600 42837 20609
rect 42795 20560 42796 20600
rect 42836 20560 42837 20600
rect 42795 20551 42837 20560
rect 43659 20600 43701 20609
rect 43659 20560 43660 20600
rect 43700 20560 43701 20600
rect 43659 20551 43701 20560
rect 46635 20600 46677 20609
rect 46635 20560 46636 20600
rect 46676 20560 46677 20600
rect 46635 20551 46677 20560
rect 47115 20600 47157 20609
rect 47115 20560 47116 20600
rect 47156 20560 47157 20600
rect 47115 20551 47157 20560
rect 49803 20600 49845 20609
rect 49803 20560 49804 20600
rect 49844 20560 49845 20600
rect 49803 20551 49845 20560
rect 50187 20600 50229 20609
rect 50187 20560 50188 20600
rect 50228 20560 50229 20600
rect 50187 20551 50229 20560
rect 50763 20600 50805 20609
rect 50763 20560 50764 20600
rect 50804 20560 50805 20600
rect 50763 20551 50805 20560
rect 52299 20600 52341 20609
rect 52299 20560 52300 20600
rect 52340 20560 52341 20600
rect 52299 20551 52341 20560
rect 576 20432 52800 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 52800 20432
rect 576 20368 52800 20392
rect 31659 20322 31701 20331
rect 31659 20282 31660 20322
rect 31700 20282 31701 20322
rect 3339 20268 3381 20277
rect 31659 20273 31701 20282
rect 3339 20228 3340 20268
rect 3380 20228 3381 20268
rect 3339 20219 3381 20228
rect 9283 20264 9341 20265
rect 9283 20224 9292 20264
rect 9332 20224 9341 20264
rect 9283 20223 9341 20224
rect 30507 20264 30549 20273
rect 42411 20268 42453 20277
rect 30507 20224 30508 20264
rect 30548 20224 30549 20264
rect 30507 20215 30549 20224
rect 41731 20264 41789 20265
rect 41731 20224 41740 20264
rect 41780 20224 41789 20264
rect 41731 20223 41789 20224
rect 42411 20228 42412 20268
rect 42452 20228 42453 20268
rect 42411 20219 42453 20228
rect 7659 20180 7701 20189
rect 7659 20140 7660 20180
rect 7700 20140 7701 20180
rect 7659 20131 7701 20140
rect 7851 20180 7893 20189
rect 7851 20140 7852 20180
rect 7892 20140 7893 20180
rect 7851 20131 7893 20140
rect 11691 20180 11733 20189
rect 11691 20140 11692 20180
rect 11732 20140 11733 20180
rect 11691 20131 11733 20140
rect 28483 20180 28541 20181
rect 28483 20140 28492 20180
rect 28532 20140 28541 20180
rect 28483 20139 28541 20140
rect 42795 20180 42837 20189
rect 42795 20140 42796 20180
rect 42836 20140 42837 20180
rect 42795 20131 42837 20140
rect 41643 20117 41685 20126
rect 1891 20096 1949 20097
rect 1891 20056 1900 20096
rect 1940 20056 1949 20096
rect 1891 20055 1949 20056
rect 2755 20096 2813 20097
rect 2755 20056 2764 20096
rect 2804 20056 2813 20096
rect 2755 20055 2813 20056
rect 3147 20096 3189 20105
rect 3147 20056 3148 20096
rect 3188 20056 3189 20096
rect 3147 20047 3189 20056
rect 3427 20096 3485 20097
rect 3427 20056 3436 20096
rect 3476 20056 3485 20096
rect 3427 20055 3485 20056
rect 3531 20096 3573 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 4011 20096 4053 20105
rect 4011 20056 4012 20096
rect 4052 20056 4053 20096
rect 4011 20047 4053 20056
rect 4203 20096 4245 20105
rect 4203 20056 4204 20096
rect 4244 20056 4245 20096
rect 4203 20047 4245 20056
rect 4291 20096 4349 20097
rect 4291 20056 4300 20096
rect 4340 20056 4349 20096
rect 4291 20055 4349 20056
rect 6403 20096 6461 20097
rect 6403 20056 6412 20096
rect 6452 20056 6461 20096
rect 6403 20055 6461 20056
rect 7267 20096 7325 20097
rect 7267 20056 7276 20096
rect 7316 20056 7325 20096
rect 7267 20055 7325 20056
rect 7947 20096 7989 20105
rect 7947 20056 7948 20096
rect 7988 20056 7989 20096
rect 7947 20047 7989 20056
rect 8043 20096 8085 20105
rect 8043 20056 8044 20096
rect 8084 20056 8085 20096
rect 8043 20047 8085 20056
rect 8139 20096 8181 20105
rect 8139 20056 8140 20096
rect 8180 20056 8181 20096
rect 8139 20047 8181 20056
rect 8331 20096 8373 20105
rect 8331 20056 8332 20096
rect 8372 20056 8373 20096
rect 8331 20047 8373 20056
rect 8427 20096 8469 20105
rect 8427 20056 8428 20096
rect 8468 20056 8469 20096
rect 8427 20047 8469 20056
rect 8523 20096 8565 20105
rect 8523 20056 8524 20096
rect 8564 20056 8565 20096
rect 8523 20047 8565 20056
rect 8619 20096 8661 20105
rect 8619 20056 8620 20096
rect 8660 20056 8661 20096
rect 8619 20047 8661 20056
rect 10435 20096 10493 20097
rect 10435 20056 10444 20096
rect 10484 20056 10493 20096
rect 10435 20055 10493 20056
rect 11299 20096 11357 20097
rect 11299 20056 11308 20096
rect 11348 20056 11357 20096
rect 11299 20055 11357 20056
rect 26955 20096 26997 20105
rect 26955 20056 26956 20096
rect 26996 20056 26997 20096
rect 26955 20047 26997 20056
rect 27619 20096 27677 20097
rect 27619 20056 27628 20096
rect 27668 20056 27677 20096
rect 27619 20055 27677 20056
rect 30699 20096 30741 20105
rect 30699 20056 30700 20096
rect 30740 20056 30741 20096
rect 30699 20047 30741 20056
rect 30795 20096 30837 20105
rect 30795 20056 30796 20096
rect 30836 20056 30837 20096
rect 30795 20047 30837 20056
rect 30891 20096 30933 20105
rect 30891 20056 30892 20096
rect 30932 20056 30933 20096
rect 30891 20047 30933 20056
rect 30987 20096 31029 20105
rect 30987 20056 30988 20096
rect 31028 20056 31029 20096
rect 30987 20047 31029 20056
rect 31467 20096 31509 20105
rect 31467 20056 31468 20096
rect 31508 20056 31509 20096
rect 31467 20047 31509 20056
rect 31555 20096 31613 20097
rect 31555 20056 31564 20096
rect 31604 20056 31613 20096
rect 31555 20055 31613 20056
rect 35683 20096 35741 20097
rect 35683 20056 35692 20096
rect 35732 20056 35741 20096
rect 35683 20055 35741 20056
rect 36547 20096 36605 20097
rect 36547 20056 36556 20096
rect 36596 20056 36605 20096
rect 36547 20055 36605 20056
rect 36939 20096 36981 20105
rect 36939 20056 36940 20096
rect 36980 20056 36981 20096
rect 36939 20047 36981 20056
rect 38563 20096 38621 20097
rect 38563 20056 38572 20096
rect 38612 20056 38621 20096
rect 38563 20055 38621 20056
rect 39427 20096 39485 20097
rect 39427 20056 39436 20096
rect 39476 20056 39485 20096
rect 39427 20055 39485 20056
rect 39819 20096 39861 20105
rect 39819 20056 39820 20096
rect 39860 20056 39861 20096
rect 39819 20047 39861 20056
rect 40483 20096 40541 20097
rect 40483 20056 40492 20096
rect 40532 20056 40541 20096
rect 40483 20055 40541 20056
rect 40875 20096 40917 20105
rect 40875 20056 40876 20096
rect 40916 20056 40917 20096
rect 41643 20077 41644 20117
rect 41684 20077 41685 20117
rect 43171 20109 43229 20110
rect 41643 20068 41685 20077
rect 42219 20096 42261 20105
rect 40875 20047 40917 20056
rect 41451 20051 41493 20060
rect 42219 20056 42220 20096
rect 42260 20056 42261 20096
rect 43171 20069 43180 20109
rect 43220 20069 43229 20109
rect 43171 20068 43229 20069
rect 44035 20096 44093 20097
rect 4675 20012 4733 20013
rect 4675 19972 4684 20012
rect 4724 19972 4733 20012
rect 4675 19971 4733 19972
rect 5259 20012 5301 20021
rect 5259 19972 5260 20012
rect 5300 19972 5301 20012
rect 5259 19963 5301 19972
rect 30307 20012 30365 20013
rect 30307 19972 30316 20012
rect 30356 19972 30365 20012
rect 30307 19971 30365 19972
rect 31939 20012 31997 20013
rect 31939 19972 31948 20012
rect 31988 19972 31997 20012
rect 31939 19971 31997 19972
rect 33187 20012 33245 20013
rect 33187 19972 33196 20012
rect 33236 19972 33245 20012
rect 33187 19971 33245 19972
rect 33571 20012 33629 20013
rect 33571 19972 33580 20012
rect 33620 19972 33629 20012
rect 33571 19971 33629 19972
rect 33955 20012 34013 20013
rect 33955 19972 33964 20012
rect 34004 19972 34013 20012
rect 33955 19971 34013 19972
rect 40099 20012 40157 20013
rect 40099 19972 40108 20012
rect 40148 19972 40157 20012
rect 40099 19971 40157 19972
rect 40587 20012 40629 20021
rect 40587 19972 40588 20012
rect 40628 19972 40629 20012
rect 40587 19963 40629 19972
rect 40779 20012 40821 20021
rect 40779 19972 40780 20012
rect 40820 19972 40821 20012
rect 40779 19963 40821 19972
rect 41059 20012 41117 20013
rect 41059 19972 41068 20012
rect 41108 19972 41117 20012
rect 41451 20011 41452 20051
rect 41492 20011 41493 20051
rect 41539 20054 41597 20055
rect 41539 20014 41548 20054
rect 41588 20014 41597 20054
rect 42219 20047 42261 20056
rect 44035 20056 44044 20096
rect 44084 20056 44093 20096
rect 44035 20055 44093 20056
rect 45387 20096 45429 20105
rect 45387 20056 45388 20096
rect 45428 20056 45429 20096
rect 42307 20054 42365 20055
rect 41539 20013 41597 20014
rect 42307 20014 42316 20054
rect 42356 20014 42365 20054
rect 45387 20047 45429 20056
rect 45763 20096 45821 20097
rect 45763 20056 45772 20096
rect 45812 20056 45821 20096
rect 45763 20055 45821 20056
rect 46627 20096 46685 20097
rect 46627 20056 46636 20096
rect 46676 20056 46685 20096
rect 46627 20055 46685 20056
rect 48363 20096 48405 20105
rect 48363 20056 48364 20096
rect 48404 20056 48405 20096
rect 48363 20047 48405 20056
rect 48739 20096 48797 20097
rect 48739 20056 48748 20096
rect 48788 20056 48797 20096
rect 48739 20055 48797 20056
rect 49603 20096 49661 20097
rect 49603 20056 49612 20096
rect 49652 20056 49661 20096
rect 49603 20055 49661 20056
rect 42307 20013 42365 20014
rect 41451 20002 41493 20011
rect 47787 20012 47829 20021
rect 41059 19971 41117 19972
rect 47787 19972 47788 20012
rect 47828 19972 47829 20012
rect 47787 19963 47829 19972
rect 50947 20012 51005 20013
rect 50947 19972 50956 20012
rect 50996 19972 51005 20012
rect 50947 19971 51005 19972
rect 51331 20012 51389 20013
rect 51331 19972 51340 20012
rect 51380 19972 51389 20012
rect 51331 19971 51389 19972
rect 51907 20012 51965 20013
rect 51907 19972 51916 20012
rect 51956 19972 51965 20012
rect 51907 19971 51965 19972
rect 3819 19928 3861 19937
rect 3819 19888 3820 19928
rect 3860 19888 3861 19928
rect 3819 19879 3861 19888
rect 27915 19928 27957 19937
rect 27915 19888 27916 19928
rect 27956 19888 27957 19928
rect 27915 19879 27957 19888
rect 31179 19928 31221 19937
rect 31179 19888 31180 19928
rect 31220 19888 31221 19928
rect 31179 19879 31221 19888
rect 32139 19928 32181 19937
rect 32139 19888 32140 19928
rect 32180 19888 32181 19928
rect 32139 19879 32181 19888
rect 40683 19928 40725 19937
rect 40683 19888 40684 19928
rect 40724 19888 40725 19928
rect 40683 19879 40725 19888
rect 41931 19928 41973 19937
rect 41931 19888 41932 19928
rect 41972 19888 41973 19928
rect 41931 19879 41973 19888
rect 51147 19928 51189 19937
rect 51147 19888 51148 19928
rect 51188 19888 51189 19928
rect 51147 19879 51189 19888
rect 739 19844 797 19845
rect 739 19804 748 19844
rect 788 19804 797 19844
rect 739 19803 797 19804
rect 4011 19844 4053 19853
rect 4011 19804 4012 19844
rect 4052 19804 4053 19844
rect 4011 19795 4053 19804
rect 4491 19844 4533 19853
rect 4491 19804 4492 19844
rect 4532 19804 4533 19844
rect 4491 19795 4533 19804
rect 33003 19844 33045 19853
rect 33003 19804 33004 19844
rect 33044 19804 33045 19844
rect 33003 19795 33045 19804
rect 33387 19844 33429 19853
rect 33387 19804 33388 19844
rect 33428 19804 33429 19844
rect 33387 19795 33429 19804
rect 33771 19844 33813 19853
rect 33771 19804 33772 19844
rect 33812 19804 33813 19844
rect 33771 19795 33813 19804
rect 34531 19844 34589 19845
rect 34531 19804 34540 19844
rect 34580 19804 34589 19844
rect 34531 19803 34589 19804
rect 37411 19844 37469 19845
rect 37411 19804 37420 19844
rect 37460 19804 37469 19844
rect 37411 19803 37469 19804
rect 40299 19844 40341 19853
rect 40299 19804 40300 19844
rect 40340 19804 40341 19844
rect 40299 19795 40341 19804
rect 41259 19844 41301 19853
rect 41259 19804 41260 19844
rect 41300 19804 41301 19844
rect 41259 19795 41301 19804
rect 45187 19844 45245 19845
rect 45187 19804 45196 19844
rect 45236 19804 45245 19844
rect 45187 19803 45245 19804
rect 50755 19844 50813 19845
rect 50755 19804 50764 19844
rect 50804 19804 50813 19844
rect 50755 19803 50813 19804
rect 51531 19844 51573 19853
rect 51531 19804 51532 19844
rect 51572 19804 51573 19844
rect 51531 19795 51573 19804
rect 51723 19844 51765 19853
rect 51723 19804 51724 19844
rect 51764 19804 51765 19844
rect 51723 19795 51765 19804
rect 576 19676 52800 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 52800 19676
rect 576 19612 52800 19636
rect 1227 19508 1269 19517
rect 1227 19468 1228 19508
rect 1268 19468 1269 19508
rect 1227 19459 1269 19468
rect 3051 19508 3093 19517
rect 3051 19468 3052 19508
rect 3092 19468 3093 19508
rect 3051 19459 3093 19468
rect 6411 19508 6453 19517
rect 6411 19468 6412 19508
rect 6452 19468 6453 19508
rect 6411 19459 6453 19468
rect 7083 19508 7125 19517
rect 7083 19468 7084 19508
rect 7124 19468 7125 19508
rect 7083 19459 7125 19468
rect 7275 19508 7317 19517
rect 7275 19468 7276 19508
rect 7316 19468 7317 19508
rect 7275 19459 7317 19468
rect 10731 19508 10773 19517
rect 10731 19468 10732 19508
rect 10772 19468 10773 19508
rect 10731 19459 10773 19468
rect 31659 19508 31701 19517
rect 31659 19468 31660 19508
rect 31700 19468 31701 19508
rect 31659 19459 31701 19468
rect 38859 19508 38901 19517
rect 38859 19468 38860 19508
rect 38900 19468 38901 19508
rect 38859 19459 38901 19468
rect 48075 19508 48117 19517
rect 48075 19468 48076 19508
rect 48116 19468 48117 19508
rect 48075 19459 48117 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 3435 19424 3477 19433
rect 3435 19384 3436 19424
rect 3476 19384 3477 19424
rect 3435 19375 3477 19384
rect 4587 19424 4629 19433
rect 4587 19384 4588 19424
rect 4628 19384 4629 19424
rect 4587 19375 4629 19384
rect 13419 19424 13461 19433
rect 13419 19384 13420 19424
rect 13460 19384 13461 19424
rect 13419 19375 13461 19384
rect 32811 19424 32853 19433
rect 32811 19384 32812 19424
rect 32852 19384 32853 19424
rect 32811 19375 32853 19384
rect 36459 19424 36501 19433
rect 36459 19384 36460 19424
rect 36500 19384 36501 19424
rect 36459 19375 36501 19384
rect 36843 19424 36885 19433
rect 36843 19384 36844 19424
rect 36884 19384 36885 19424
rect 36843 19375 36885 19384
rect 38091 19424 38133 19433
rect 38091 19384 38092 19424
rect 38132 19384 38133 19424
rect 38091 19375 38133 19384
rect 39243 19424 39285 19433
rect 39243 19384 39244 19424
rect 39284 19384 39285 19424
rect 39243 19375 39285 19384
rect 39627 19424 39669 19433
rect 39627 19384 39628 19424
rect 39668 19384 39669 19424
rect 39627 19375 39669 19384
rect 40011 19424 40053 19433
rect 40011 19384 40012 19424
rect 40052 19384 40053 19424
rect 40011 19375 40053 19384
rect 41163 19424 41205 19433
rect 41163 19384 41164 19424
rect 41204 19384 41205 19424
rect 41163 19375 41205 19384
rect 44331 19424 44373 19433
rect 44331 19384 44332 19424
rect 44372 19384 44373 19424
rect 44331 19375 44373 19384
rect 45675 19424 45717 19433
rect 45675 19384 45676 19424
rect 45716 19384 45717 19424
rect 45675 19375 45717 19384
rect 46155 19424 46197 19433
rect 46155 19384 46156 19424
rect 46196 19384 46197 19424
rect 46155 19375 46197 19384
rect 48459 19424 48501 19433
rect 48459 19384 48460 19424
rect 48500 19384 48501 19424
rect 48459 19375 48501 19384
rect 1411 19340 1469 19341
rect 1411 19300 1420 19340
rect 1460 19300 1469 19340
rect 1411 19299 1469 19300
rect 1795 19340 1853 19341
rect 1795 19300 1804 19340
rect 1844 19300 1853 19340
rect 1795 19299 1853 19300
rect 2179 19340 2237 19341
rect 2179 19300 2188 19340
rect 2228 19300 2237 19340
rect 2179 19299 2237 19300
rect 3339 19340 3381 19349
rect 3339 19300 3340 19340
rect 3380 19300 3381 19340
rect 3339 19291 3381 19300
rect 3531 19340 3573 19349
rect 3531 19300 3532 19340
rect 3572 19300 3573 19340
rect 3531 19291 3573 19300
rect 4099 19340 4157 19341
rect 4099 19300 4108 19340
rect 4148 19300 4157 19340
rect 4099 19299 4157 19300
rect 5923 19340 5981 19341
rect 5923 19300 5932 19340
rect 5972 19300 5981 19340
rect 5923 19299 5981 19300
rect 30691 19340 30749 19341
rect 30691 19300 30700 19340
rect 30740 19300 30749 19340
rect 30691 19299 30749 19300
rect 32419 19340 32477 19341
rect 32419 19300 32428 19340
rect 32468 19300 32477 19340
rect 32419 19299 32477 19300
rect 36363 19340 36405 19349
rect 36363 19300 36364 19340
rect 36404 19300 36405 19340
rect 36363 19291 36405 19300
rect 36555 19340 36597 19349
rect 36555 19300 36556 19340
rect 36596 19300 36597 19340
rect 36555 19291 36597 19300
rect 38659 19340 38717 19341
rect 38659 19300 38668 19340
rect 38708 19300 38717 19340
rect 38659 19299 38717 19300
rect 39043 19340 39101 19341
rect 39043 19300 39052 19340
rect 39092 19300 39101 19340
rect 39043 19299 39101 19300
rect 39531 19340 39573 19349
rect 39531 19300 39532 19340
rect 39572 19300 39573 19340
rect 39531 19291 39573 19300
rect 39723 19340 39765 19349
rect 39723 19300 39724 19340
rect 39764 19300 39765 19340
rect 45091 19340 45149 19341
rect 39723 19291 39765 19300
rect 40971 19301 41013 19310
rect 2947 19256 3005 19257
rect 2947 19216 2956 19256
rect 2996 19216 3005 19256
rect 2947 19215 3005 19216
rect 3235 19256 3293 19257
rect 3235 19216 3244 19256
rect 3284 19216 3293 19256
rect 3235 19215 3293 19216
rect 3627 19256 3669 19265
rect 3627 19216 3628 19256
rect 3668 19216 3669 19256
rect 4395 19256 4437 19265
rect 3627 19207 3669 19216
rect 4281 19241 4339 19242
rect 4281 19201 4290 19241
rect 4330 19201 4339 19241
rect 4395 19216 4396 19256
rect 4436 19216 4437 19256
rect 4395 19207 4437 19216
rect 4587 19256 4629 19265
rect 4587 19216 4588 19256
rect 4628 19216 4629 19256
rect 4587 19207 4629 19216
rect 6307 19256 6365 19257
rect 6307 19216 6316 19256
rect 6356 19216 6365 19256
rect 6307 19215 6365 19216
rect 6691 19256 6749 19257
rect 6691 19216 6700 19256
rect 6740 19216 6749 19256
rect 6691 19215 6749 19216
rect 6795 19256 6837 19265
rect 6795 19216 6796 19256
rect 6836 19216 6837 19256
rect 6795 19207 6837 19216
rect 7275 19256 7317 19265
rect 7275 19216 7276 19256
rect 7316 19216 7317 19256
rect 7275 19207 7317 19216
rect 7467 19256 7509 19265
rect 7467 19216 7468 19256
rect 7508 19216 7509 19256
rect 7467 19207 7509 19216
rect 7555 19256 7613 19257
rect 7555 19216 7564 19256
rect 7604 19216 7613 19256
rect 7555 19215 7613 19216
rect 9771 19256 9813 19265
rect 9771 19216 9772 19256
rect 9812 19216 9813 19256
rect 9771 19207 9813 19216
rect 9867 19256 9909 19265
rect 9867 19216 9868 19256
rect 9908 19216 9909 19256
rect 9867 19207 9909 19216
rect 9963 19256 10005 19265
rect 9963 19216 9964 19256
rect 10004 19216 10005 19256
rect 9963 19207 10005 19216
rect 10059 19256 10101 19265
rect 10059 19216 10060 19256
rect 10100 19216 10101 19256
rect 10059 19207 10101 19216
rect 10339 19256 10397 19257
rect 10339 19216 10348 19256
rect 10388 19216 10397 19256
rect 10339 19215 10397 19216
rect 10443 19256 10485 19265
rect 10443 19216 10444 19256
rect 10484 19216 10485 19256
rect 10443 19207 10485 19216
rect 10923 19256 10965 19265
rect 10923 19216 10924 19256
rect 10964 19216 10965 19256
rect 10923 19207 10965 19216
rect 11115 19256 11157 19265
rect 11115 19216 11116 19256
rect 11156 19216 11157 19256
rect 11115 19207 11157 19216
rect 11203 19256 11261 19257
rect 11203 19216 11212 19256
rect 11252 19216 11261 19256
rect 11203 19215 11261 19216
rect 12459 19256 12501 19265
rect 12459 19216 12460 19256
rect 12500 19216 12501 19256
rect 12459 19207 12501 19216
rect 12555 19256 12597 19265
rect 12555 19216 12556 19256
rect 12596 19216 12597 19256
rect 12555 19207 12597 19216
rect 12651 19256 12693 19265
rect 12651 19216 12652 19256
rect 12692 19216 12693 19256
rect 12651 19207 12693 19216
rect 12747 19256 12789 19265
rect 12747 19216 12748 19256
rect 12788 19216 12789 19256
rect 12747 19207 12789 19216
rect 13027 19256 13085 19257
rect 13027 19216 13036 19256
rect 13076 19216 13085 19256
rect 13027 19215 13085 19216
rect 13131 19256 13173 19265
rect 13131 19216 13132 19256
rect 13172 19216 13173 19256
rect 13131 19207 13173 19216
rect 31555 19256 31613 19257
rect 31555 19216 31564 19256
rect 31604 19216 31613 19256
rect 31555 19215 31613 19216
rect 33099 19254 33141 19263
rect 33099 19214 33100 19254
rect 33140 19214 33141 19254
rect 33187 19256 33245 19257
rect 33187 19216 33196 19256
rect 33236 19216 33245 19256
rect 33187 19215 33245 19216
rect 33579 19256 33621 19265
rect 33579 19216 33580 19256
rect 33620 19216 33621 19256
rect 33099 19205 33141 19214
rect 33579 19207 33621 19216
rect 33955 19256 34013 19257
rect 33955 19216 33964 19256
rect 34004 19216 34013 19256
rect 33955 19215 34013 19216
rect 34819 19256 34877 19257
rect 34819 19216 34828 19256
rect 34868 19216 34877 19256
rect 34819 19215 34877 19216
rect 36259 19256 36317 19257
rect 36259 19216 36268 19256
rect 36308 19216 36317 19256
rect 36259 19215 36317 19216
rect 36651 19256 36693 19265
rect 36651 19216 36652 19256
rect 36692 19216 36693 19256
rect 36651 19207 36693 19216
rect 37131 19256 37173 19265
rect 37131 19216 37132 19256
rect 37172 19216 37173 19256
rect 37131 19207 37173 19216
rect 37219 19256 37277 19257
rect 37219 19216 37228 19256
rect 37268 19216 37277 19256
rect 37219 19215 37277 19216
rect 37507 19256 37565 19257
rect 37507 19216 37516 19256
rect 37556 19216 37565 19256
rect 37507 19215 37565 19216
rect 37611 19256 37653 19265
rect 37611 19216 37612 19256
rect 37652 19216 37653 19256
rect 37611 19207 37653 19216
rect 38091 19256 38133 19265
rect 38091 19216 38092 19256
rect 38132 19216 38133 19256
rect 38091 19207 38133 19216
rect 38283 19256 38325 19265
rect 38283 19216 38284 19256
rect 38324 19216 38325 19256
rect 38283 19207 38325 19216
rect 38371 19256 38429 19257
rect 38371 19216 38380 19256
rect 38420 19216 38429 19256
rect 38371 19215 38429 19216
rect 39435 19256 39477 19265
rect 39435 19216 39436 19256
rect 39476 19216 39477 19256
rect 39435 19207 39477 19216
rect 39811 19256 39869 19257
rect 39811 19216 39820 19256
rect 39860 19216 39869 19256
rect 39811 19215 39869 19216
rect 40299 19256 40341 19265
rect 40299 19216 40300 19256
rect 40340 19216 40341 19256
rect 40299 19207 40341 19216
rect 40387 19256 40445 19257
rect 40387 19216 40396 19256
rect 40436 19216 40445 19256
rect 40387 19215 40445 19216
rect 40683 19256 40725 19265
rect 40683 19216 40684 19256
rect 40724 19216 40725 19256
rect 40683 19207 40725 19216
rect 40779 19256 40821 19265
rect 40779 19216 40780 19256
rect 40820 19216 40821 19256
rect 40779 19207 40821 19216
rect 40875 19256 40917 19265
rect 40875 19216 40876 19256
rect 40916 19216 40917 19256
rect 40971 19261 40972 19301
rect 41012 19261 41013 19301
rect 45091 19300 45100 19340
rect 45140 19300 45149 19340
rect 45091 19299 45149 19300
rect 45579 19340 45621 19349
rect 45579 19300 45580 19340
rect 45620 19300 45621 19340
rect 45579 19291 45621 19300
rect 45771 19340 45813 19349
rect 45771 19300 45772 19340
rect 45812 19300 45813 19340
rect 45771 19291 45813 19300
rect 47491 19340 47549 19341
rect 47491 19300 47500 19340
rect 47540 19300 47549 19340
rect 47491 19299 47549 19300
rect 48363 19340 48405 19349
rect 48363 19300 48364 19340
rect 48404 19300 48405 19340
rect 48363 19291 48405 19300
rect 48555 19340 48597 19349
rect 48555 19300 48556 19340
rect 48596 19300 48597 19340
rect 48555 19291 48597 19300
rect 40971 19252 41013 19261
rect 41163 19256 41205 19265
rect 40875 19207 40917 19216
rect 41163 19216 41164 19256
rect 41204 19216 41205 19256
rect 41163 19207 41205 19216
rect 41355 19256 41397 19265
rect 41355 19216 41356 19256
rect 41396 19216 41397 19256
rect 41355 19207 41397 19216
rect 41443 19256 41501 19257
rect 41443 19216 41452 19256
rect 41492 19216 41501 19256
rect 41443 19215 41501 19216
rect 41731 19256 41789 19257
rect 41731 19216 41740 19256
rect 41780 19216 41789 19256
rect 41731 19215 41789 19216
rect 43179 19256 43221 19265
rect 43179 19216 43180 19256
rect 43220 19216 43221 19256
rect 43179 19207 43221 19216
rect 44035 19256 44093 19257
rect 44035 19216 44044 19256
rect 44084 19216 44093 19256
rect 44035 19215 44093 19216
rect 44139 19256 44181 19265
rect 44139 19216 44140 19256
rect 44180 19216 44181 19256
rect 44139 19207 44181 19216
rect 44331 19256 44373 19265
rect 44331 19216 44332 19256
rect 44372 19216 44373 19256
rect 44331 19207 44373 19216
rect 45483 19256 45525 19265
rect 45483 19216 45484 19256
rect 45524 19216 45525 19256
rect 45483 19207 45525 19216
rect 45859 19256 45917 19257
rect 45859 19216 45868 19256
rect 45908 19216 45917 19256
rect 45859 19215 45917 19216
rect 46443 19256 46485 19265
rect 46443 19216 46444 19256
rect 46484 19216 46485 19256
rect 46443 19207 46485 19216
rect 46531 19256 46589 19257
rect 46531 19216 46540 19256
rect 46580 19216 46589 19256
rect 46531 19215 46589 19216
rect 46923 19256 46965 19265
rect 46923 19216 46924 19256
rect 46964 19216 46965 19256
rect 46923 19207 46965 19216
rect 47019 19256 47061 19265
rect 47019 19216 47020 19256
rect 47060 19216 47061 19256
rect 47019 19207 47061 19216
rect 47115 19256 47157 19265
rect 47115 19216 47116 19256
rect 47156 19216 47157 19256
rect 47115 19207 47157 19216
rect 47779 19256 47837 19257
rect 47779 19216 47788 19256
rect 47828 19216 47837 19256
rect 47779 19215 47837 19216
rect 47883 19256 47925 19265
rect 47883 19216 47884 19256
rect 47924 19216 47925 19256
rect 48267 19256 48309 19265
rect 47883 19207 47925 19216
rect 48075 19242 48117 19251
rect 4281 19200 4339 19201
rect 48075 19202 48076 19242
rect 48116 19202 48117 19242
rect 48267 19216 48268 19256
rect 48308 19216 48309 19256
rect 48267 19207 48309 19216
rect 48643 19256 48701 19257
rect 48643 19216 48652 19256
rect 48692 19216 48701 19256
rect 48643 19215 48701 19216
rect 49035 19256 49077 19265
rect 49035 19216 49036 19256
rect 49076 19216 49077 19256
rect 49035 19207 49077 19216
rect 49891 19256 49949 19257
rect 49891 19216 49900 19256
rect 49940 19216 49949 19256
rect 49891 19215 49949 19216
rect 50659 19256 50717 19257
rect 50659 19216 50668 19256
rect 50708 19216 50717 19256
rect 50659 19215 50717 19216
rect 51523 19256 51581 19257
rect 51523 19216 51532 19256
rect 51572 19216 51581 19256
rect 51523 19215 51581 19216
rect 48075 19193 48117 19202
rect 11019 19172 11061 19181
rect 11019 19132 11020 19172
rect 11060 19132 11061 19172
rect 11019 19123 11061 19132
rect 50283 19172 50325 19181
rect 50283 19132 50284 19172
rect 50324 19132 50325 19172
rect 50283 19123 50325 19132
rect 1611 19088 1653 19097
rect 1611 19048 1612 19088
rect 1652 19048 1653 19088
rect 1611 19039 1653 19048
rect 1995 19088 2037 19097
rect 1995 19048 1996 19088
rect 2036 19048 2037 19088
rect 1995 19039 2037 19048
rect 3915 19088 3957 19097
rect 3915 19048 3916 19088
rect 3956 19048 3957 19088
rect 3915 19039 3957 19048
rect 5739 19088 5781 19097
rect 5739 19048 5740 19088
rect 5780 19048 5781 19088
rect 5739 19039 5781 19048
rect 6603 19084 6645 19093
rect 6603 19044 6604 19084
rect 6644 19044 6645 19084
rect 6603 19035 6645 19044
rect 10251 19084 10293 19093
rect 10251 19044 10252 19084
rect 10292 19044 10293 19084
rect 10251 19035 10293 19044
rect 30891 19088 30933 19097
rect 30891 19048 30892 19088
rect 30932 19048 30933 19088
rect 30891 19039 30933 19048
rect 32619 19088 32661 19097
rect 32619 19048 32620 19088
rect 32660 19048 32661 19088
rect 32619 19039 32661 19048
rect 35971 19088 36029 19089
rect 35971 19048 35980 19088
rect 36020 19048 36029 19088
rect 35971 19047 36029 19048
rect 37323 19084 37365 19093
rect 37323 19044 37324 19084
rect 37364 19044 37365 19084
rect 12939 19030 12981 19039
rect 12939 18990 12940 19030
rect 12980 18990 12981 19030
rect 12939 18981 12981 18990
rect 33291 19030 33333 19039
rect 37323 19035 37365 19044
rect 40491 19084 40533 19093
rect 40491 19044 40492 19084
rect 40532 19044 40533 19084
rect 40491 19035 40533 19044
rect 45291 19088 45333 19097
rect 45291 19048 45292 19088
rect 45332 19048 45333 19088
rect 45291 19039 45333 19048
rect 46819 19088 46877 19089
rect 46819 19048 46828 19088
rect 46868 19048 46877 19088
rect 46819 19047 46877 19048
rect 47307 19088 47349 19097
rect 47307 19048 47308 19088
rect 47348 19048 47349 19088
rect 47307 19039 47349 19048
rect 49419 19088 49461 19097
rect 49419 19048 49420 19088
rect 49460 19048 49461 19088
rect 49419 19039 49461 19048
rect 52675 19088 52733 19089
rect 52675 19048 52684 19088
rect 52724 19048 52733 19088
rect 52675 19047 52733 19048
rect 33291 18990 33292 19030
rect 33332 18990 33333 19030
rect 33291 18981 33333 18990
rect 46635 19030 46677 19039
rect 46635 18990 46636 19030
rect 46676 18990 46677 19030
rect 46635 18981 46677 18990
rect 576 18920 52800 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 52800 18920
rect 576 18856 52800 18880
rect 50091 18810 50133 18819
rect 50091 18770 50092 18810
rect 50132 18770 50133 18810
rect 3915 18756 3957 18765
rect 50091 18761 50133 18770
rect 3915 18716 3916 18756
rect 3956 18716 3957 18756
rect 3915 18707 3957 18716
rect 33483 18752 33525 18761
rect 33483 18712 33484 18752
rect 33524 18712 33525 18752
rect 33483 18703 33525 18712
rect 34147 18752 34205 18753
rect 34147 18712 34156 18752
rect 34196 18712 34205 18752
rect 34147 18711 34205 18712
rect 42595 18752 42653 18753
rect 42595 18712 42604 18752
rect 42644 18712 42653 18752
rect 42595 18711 42653 18712
rect 43563 18752 43605 18761
rect 43563 18712 43564 18752
rect 43604 18712 43605 18752
rect 43563 18703 43605 18712
rect 50275 18752 50333 18753
rect 50275 18712 50284 18752
rect 50324 18712 50333 18752
rect 50275 18711 50333 18712
rect 51627 18752 51669 18761
rect 51627 18712 51628 18752
rect 51668 18712 51669 18752
rect 51627 18703 51669 18712
rect 32803 18626 32861 18627
rect 3435 18584 3477 18593
rect 3435 18544 3436 18584
rect 3476 18544 3477 18584
rect 3435 18535 3477 18544
rect 3531 18584 3573 18593
rect 3531 18544 3532 18584
rect 3572 18544 3573 18584
rect 3531 18535 3573 18544
rect 3627 18584 3669 18593
rect 3627 18544 3628 18584
rect 3668 18544 3669 18584
rect 3627 18535 3669 18544
rect 3723 18584 3765 18593
rect 3723 18544 3724 18584
rect 3764 18544 3765 18584
rect 3723 18535 3765 18544
rect 4003 18584 4061 18585
rect 4003 18544 4012 18584
rect 4052 18544 4061 18584
rect 4003 18543 4061 18544
rect 4107 18584 4149 18593
rect 4107 18544 4108 18584
rect 4148 18544 4149 18584
rect 4107 18535 4149 18544
rect 4579 18584 4637 18585
rect 4579 18544 4588 18584
rect 4628 18544 4637 18584
rect 4579 18543 4637 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 7275 18584 7317 18593
rect 7275 18544 7276 18584
rect 7316 18544 7317 18584
rect 7275 18535 7317 18544
rect 7371 18584 7413 18593
rect 7371 18544 7372 18584
rect 7412 18544 7413 18584
rect 7371 18535 7413 18544
rect 7467 18584 7509 18593
rect 7467 18544 7468 18584
rect 7508 18544 7509 18584
rect 7467 18535 7509 18544
rect 7563 18584 7605 18593
rect 7563 18544 7564 18584
rect 7604 18544 7605 18584
rect 7563 18535 7605 18544
rect 7755 18584 7797 18593
rect 7755 18544 7756 18584
rect 7796 18544 7797 18584
rect 7755 18535 7797 18544
rect 8131 18584 8189 18585
rect 8131 18544 8140 18584
rect 8180 18544 8189 18584
rect 8131 18543 8189 18544
rect 8995 18584 9053 18585
rect 8995 18544 9004 18584
rect 9044 18544 9053 18584
rect 8995 18543 9053 18544
rect 10635 18584 10677 18593
rect 10635 18544 10636 18584
rect 10676 18544 10677 18584
rect 10635 18535 10677 18544
rect 10731 18584 10773 18593
rect 10731 18544 10732 18584
rect 10772 18544 10773 18584
rect 10731 18535 10773 18544
rect 10827 18584 10869 18593
rect 10827 18544 10828 18584
rect 10868 18544 10869 18584
rect 10827 18535 10869 18544
rect 10923 18584 10965 18593
rect 10923 18544 10924 18584
rect 10964 18544 10965 18584
rect 10923 18535 10965 18544
rect 12075 18584 12117 18593
rect 12075 18544 12076 18584
rect 12116 18544 12117 18584
rect 12075 18535 12117 18544
rect 12451 18584 12509 18585
rect 12451 18544 12460 18584
rect 12500 18544 12509 18584
rect 12451 18543 12509 18544
rect 12651 18584 12693 18593
rect 12651 18544 12652 18584
rect 12692 18544 12693 18584
rect 12651 18535 12693 18544
rect 13027 18584 13085 18585
rect 13027 18544 13036 18584
rect 13076 18544 13085 18584
rect 13027 18543 13085 18544
rect 13891 18584 13949 18585
rect 13891 18544 13900 18584
rect 13940 18544 13949 18584
rect 13891 18543 13949 18544
rect 15243 18584 15285 18593
rect 15243 18544 15244 18584
rect 15284 18544 15285 18584
rect 15243 18535 15285 18544
rect 15339 18584 15381 18593
rect 15339 18544 15340 18584
rect 15380 18544 15381 18584
rect 15339 18535 15381 18544
rect 15435 18584 15477 18593
rect 15435 18544 15436 18584
rect 15476 18544 15477 18584
rect 15435 18535 15477 18544
rect 15531 18584 15573 18593
rect 15531 18544 15532 18584
rect 15572 18544 15573 18584
rect 15531 18535 15573 18544
rect 15723 18584 15765 18593
rect 15723 18544 15724 18584
rect 15764 18544 15765 18584
rect 15723 18535 15765 18544
rect 16099 18584 16157 18585
rect 16099 18544 16108 18584
rect 16148 18544 16157 18584
rect 16099 18543 16157 18544
rect 16963 18584 17021 18585
rect 16963 18544 16972 18584
rect 17012 18544 17021 18584
rect 16963 18543 17021 18544
rect 31363 18584 31421 18585
rect 31363 18544 31372 18584
rect 31412 18544 31421 18584
rect 31363 18543 31421 18544
rect 32227 18584 32285 18585
rect 32227 18544 32236 18584
rect 32276 18544 32285 18584
rect 32227 18543 32285 18544
rect 32619 18584 32661 18593
rect 32803 18586 32812 18626
rect 32852 18586 32861 18626
rect 32803 18585 32861 18586
rect 32619 18544 32620 18584
rect 32660 18544 32661 18584
rect 32619 18535 32661 18544
rect 33195 18584 33237 18593
rect 33195 18544 33196 18584
rect 33236 18544 33237 18584
rect 32926 18542 32984 18543
rect 1315 18500 1373 18501
rect 1315 18460 1324 18500
rect 1364 18460 1373 18500
rect 1315 18459 1373 18460
rect 1699 18500 1757 18501
rect 1699 18460 1708 18500
rect 1748 18460 1757 18500
rect 1699 18459 1757 18460
rect 4683 18500 4725 18509
rect 4683 18460 4684 18500
rect 4724 18460 4725 18500
rect 4683 18451 4725 18460
rect 4875 18500 4917 18509
rect 4875 18460 4876 18500
rect 4916 18460 4917 18500
rect 4875 18451 4917 18460
rect 5347 18500 5405 18501
rect 5347 18460 5356 18500
rect 5396 18460 5405 18500
rect 5347 18459 5405 18460
rect 6787 18500 6845 18501
rect 6787 18460 6796 18500
rect 6836 18460 6845 18500
rect 6787 18459 6845 18460
rect 12171 18500 12213 18509
rect 12171 18460 12172 18500
rect 12212 18460 12213 18500
rect 12171 18451 12213 18460
rect 12363 18500 12405 18509
rect 32926 18502 32935 18542
rect 32975 18502 32984 18542
rect 33195 18535 33237 18544
rect 33379 18584 33437 18585
rect 33379 18544 33388 18584
rect 33428 18544 33437 18584
rect 33379 18543 33437 18544
rect 33675 18584 33717 18593
rect 33675 18544 33676 18584
rect 33716 18544 33717 18584
rect 33675 18535 33717 18544
rect 33867 18584 33909 18593
rect 33867 18544 33868 18584
rect 33908 18544 33909 18584
rect 33867 18535 33909 18544
rect 33955 18584 34013 18585
rect 33955 18544 33964 18584
rect 34004 18544 34013 18584
rect 33955 18543 34013 18544
rect 34251 18584 34293 18593
rect 34251 18544 34252 18584
rect 34292 18544 34293 18584
rect 34251 18535 34293 18544
rect 34347 18584 34389 18593
rect 34347 18544 34348 18584
rect 34388 18544 34389 18584
rect 34347 18535 34389 18544
rect 34443 18584 34485 18593
rect 34443 18544 34444 18584
rect 34484 18544 34485 18584
rect 34443 18535 34485 18544
rect 34627 18584 34685 18585
rect 34627 18544 34636 18584
rect 34676 18544 34685 18584
rect 34627 18543 34685 18544
rect 36459 18584 36501 18593
rect 36459 18544 36460 18584
rect 36500 18544 36501 18584
rect 36459 18535 36501 18544
rect 36555 18584 36597 18593
rect 36555 18544 36556 18584
rect 36596 18544 36597 18584
rect 36555 18535 36597 18544
rect 36651 18584 36693 18593
rect 36651 18544 36652 18584
rect 36692 18544 36693 18584
rect 36651 18535 36693 18544
rect 36747 18584 36789 18593
rect 36747 18544 36748 18584
rect 36788 18544 36789 18584
rect 36747 18535 36789 18544
rect 36939 18584 36981 18593
rect 36939 18544 36940 18584
rect 36980 18544 36981 18584
rect 36939 18535 36981 18544
rect 37315 18584 37373 18585
rect 37315 18544 37324 18584
rect 37364 18544 37373 18584
rect 37315 18543 37373 18544
rect 38179 18584 38237 18585
rect 38179 18544 38188 18584
rect 38228 18544 38237 18584
rect 38179 18543 38237 18544
rect 39531 18584 39573 18593
rect 39531 18544 39532 18584
rect 39572 18544 39573 18584
rect 39531 18535 39573 18544
rect 39627 18584 39669 18593
rect 39627 18544 39628 18584
rect 39668 18544 39669 18584
rect 39627 18535 39669 18544
rect 39723 18584 39765 18593
rect 39723 18544 39724 18584
rect 39764 18544 39765 18584
rect 39723 18535 39765 18544
rect 39819 18584 39861 18593
rect 39819 18544 39820 18584
rect 39860 18544 39861 18584
rect 39819 18535 39861 18544
rect 40011 18584 40053 18593
rect 40011 18544 40012 18584
rect 40052 18544 40053 18584
rect 40011 18535 40053 18544
rect 40387 18584 40445 18585
rect 40387 18544 40396 18584
rect 40436 18544 40445 18584
rect 40387 18543 40445 18544
rect 41251 18584 41309 18585
rect 41251 18544 41260 18584
rect 41300 18544 41309 18584
rect 41251 18543 41309 18544
rect 42699 18584 42741 18593
rect 42699 18544 42700 18584
rect 42740 18544 42741 18584
rect 42699 18535 42741 18544
rect 42795 18584 42837 18593
rect 42795 18544 42796 18584
rect 42836 18544 42837 18584
rect 42795 18535 42837 18544
rect 42891 18584 42933 18593
rect 42891 18544 42892 18584
rect 42932 18544 42933 18584
rect 42891 18535 42933 18544
rect 43459 18584 43517 18585
rect 43459 18544 43468 18584
rect 43508 18544 43517 18584
rect 43459 18543 43517 18544
rect 43755 18584 43797 18593
rect 43755 18544 43756 18584
rect 43796 18544 43797 18584
rect 43755 18535 43797 18544
rect 44131 18584 44189 18585
rect 44131 18544 44140 18584
rect 44180 18544 44189 18584
rect 44131 18543 44189 18544
rect 44995 18584 45053 18585
rect 44995 18544 45004 18584
rect 45044 18544 45053 18584
rect 44995 18543 45053 18544
rect 46347 18584 46389 18593
rect 46347 18544 46348 18584
rect 46388 18544 46389 18584
rect 46347 18535 46389 18544
rect 46723 18584 46781 18585
rect 46723 18544 46732 18584
rect 46772 18544 46781 18584
rect 46723 18543 46781 18544
rect 47587 18584 47645 18585
rect 47587 18544 47596 18584
rect 47636 18544 47645 18584
rect 47587 18543 47645 18544
rect 49131 18584 49173 18593
rect 49131 18544 49132 18584
rect 49172 18544 49173 18584
rect 49131 18535 49173 18544
rect 49323 18584 49365 18593
rect 49323 18544 49324 18584
rect 49364 18544 49365 18584
rect 49323 18535 49365 18544
rect 49411 18584 49469 18585
rect 49411 18544 49420 18584
rect 49460 18544 49469 18584
rect 49411 18543 49469 18544
rect 49899 18584 49941 18593
rect 49899 18544 49900 18584
rect 49940 18544 49941 18584
rect 49899 18535 49941 18544
rect 49987 18584 50045 18585
rect 49987 18544 49996 18584
rect 50036 18544 50045 18584
rect 49987 18543 50045 18544
rect 50379 18584 50421 18593
rect 50379 18544 50380 18584
rect 50420 18544 50421 18584
rect 50379 18535 50421 18544
rect 50475 18584 50517 18593
rect 50475 18544 50476 18584
rect 50516 18544 50517 18584
rect 50475 18535 50517 18544
rect 50571 18584 50613 18593
rect 50571 18544 50572 18584
rect 50612 18544 50613 18584
rect 50571 18535 50613 18544
rect 50955 18584 50997 18593
rect 50955 18544 50956 18584
rect 50996 18544 50997 18584
rect 50955 18535 50997 18544
rect 51051 18584 51093 18593
rect 51051 18544 51052 18584
rect 51092 18544 51093 18584
rect 51051 18535 51093 18544
rect 51147 18584 51189 18593
rect 51147 18544 51148 18584
rect 51188 18544 51189 18584
rect 51147 18535 51189 18544
rect 51243 18584 51285 18593
rect 51243 18544 51244 18584
rect 51284 18544 51285 18584
rect 51243 18535 51285 18544
rect 51811 18584 51869 18585
rect 51811 18544 51820 18584
rect 51860 18544 51869 18584
rect 51811 18543 51869 18544
rect 32926 18501 32984 18502
rect 12363 18460 12364 18500
rect 12404 18460 12405 18500
rect 42411 18500 42453 18509
rect 12363 18451 12405 18460
rect 33099 18458 33141 18467
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 4779 18416 4821 18425
rect 4779 18376 4780 18416
rect 4820 18376 4821 18416
rect 4779 18367 4821 18376
rect 6603 18416 6645 18425
rect 6603 18376 6604 18416
rect 6644 18376 6645 18416
rect 6603 18367 6645 18376
rect 12267 18416 12309 18425
rect 12267 18376 12268 18416
rect 12308 18376 12309 18416
rect 12267 18367 12309 18376
rect 18115 18416 18173 18417
rect 18115 18376 18124 18416
rect 18164 18376 18173 18416
rect 18115 18375 18173 18376
rect 33003 18416 33045 18425
rect 33003 18376 33004 18416
rect 33044 18376 33045 18416
rect 33099 18418 33100 18458
rect 33140 18418 33141 18458
rect 42411 18460 42412 18500
rect 42452 18460 42453 18500
rect 42411 18451 42453 18460
rect 43075 18500 43133 18501
rect 43075 18460 43084 18500
rect 43124 18460 43133 18500
rect 43075 18459 43133 18460
rect 51427 18500 51485 18501
rect 51427 18460 51436 18500
rect 51476 18460 51485 18500
rect 51427 18459 51485 18460
rect 33099 18409 33141 18418
rect 43275 18416 43317 18425
rect 33003 18367 33045 18376
rect 43275 18376 43276 18416
rect 43316 18376 43317 18416
rect 43275 18367 43317 18376
rect 49611 18416 49653 18425
rect 49611 18376 49612 18416
rect 49652 18376 49653 18416
rect 49611 18367 49653 18376
rect 1131 18332 1173 18341
rect 1131 18292 1132 18332
rect 1172 18292 1173 18332
rect 1131 18283 1173 18292
rect 1515 18332 1557 18341
rect 1515 18292 1516 18332
rect 1556 18292 1557 18332
rect 1515 18283 1557 18292
rect 4395 18332 4437 18341
rect 4395 18292 4396 18332
rect 4436 18292 4437 18332
rect 4395 18283 4437 18292
rect 5163 18332 5205 18341
rect 5163 18292 5164 18332
rect 5204 18292 5205 18332
rect 5163 18283 5205 18292
rect 10147 18332 10205 18333
rect 10147 18292 10156 18332
rect 10196 18292 10205 18332
rect 10147 18291 10205 18292
rect 15043 18332 15101 18333
rect 15043 18292 15052 18332
rect 15092 18292 15101 18332
rect 15043 18291 15101 18292
rect 30211 18332 30269 18333
rect 30211 18292 30220 18332
rect 30260 18292 30269 18332
rect 30211 18291 30269 18292
rect 33675 18332 33717 18341
rect 33675 18292 33676 18332
rect 33716 18292 33717 18332
rect 33675 18283 33717 18292
rect 34731 18332 34773 18341
rect 34731 18292 34732 18332
rect 34772 18292 34773 18332
rect 34731 18283 34773 18292
rect 39331 18332 39389 18333
rect 39331 18292 39340 18332
rect 39380 18292 39389 18332
rect 39331 18291 39389 18292
rect 46147 18332 46205 18333
rect 46147 18292 46156 18332
rect 46196 18292 46205 18332
rect 46147 18291 46205 18292
rect 48739 18332 48797 18333
rect 48739 18292 48748 18332
rect 48788 18292 48797 18332
rect 48739 18291 48797 18292
rect 49131 18332 49173 18341
rect 49131 18292 49132 18332
rect 49172 18292 49173 18332
rect 49131 18283 49173 18292
rect 51627 18332 51669 18341
rect 51627 18292 51628 18332
rect 51668 18292 51669 18332
rect 51627 18283 51669 18292
rect 51915 18332 51957 18341
rect 51915 18292 51916 18332
rect 51956 18292 51957 18332
rect 51915 18283 51957 18292
rect 576 18164 52800 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 52800 18164
rect 576 18100 52800 18124
rect 3819 17996 3861 18005
rect 3819 17956 3820 17996
rect 3860 17956 3861 17996
rect 3819 17947 3861 17956
rect 7179 17996 7221 18005
rect 7179 17956 7180 17996
rect 7220 17956 7221 17996
rect 7179 17947 7221 17956
rect 10347 17996 10389 18005
rect 10347 17956 10348 17996
rect 10388 17956 10389 17996
rect 10347 17947 10389 17956
rect 13131 17996 13173 18005
rect 13131 17956 13132 17996
rect 13172 17956 13173 17996
rect 13131 17947 13173 17956
rect 13611 17996 13653 18005
rect 13611 17956 13612 17996
rect 13652 17956 13653 17996
rect 13611 17947 13653 17956
rect 31947 17996 31989 18005
rect 31947 17956 31948 17996
rect 31988 17956 31989 17996
rect 31947 17947 31989 17956
rect 39723 17996 39765 18005
rect 39723 17956 39724 17996
rect 39764 17956 39765 17996
rect 39723 17947 39765 17956
rect 48747 17996 48789 18005
rect 48747 17956 48748 17996
rect 48788 17956 48789 17996
rect 48747 17947 48789 17956
rect 51051 17996 51093 18005
rect 51051 17956 51052 17996
rect 51092 17956 51093 17996
rect 51051 17947 51093 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 49899 17912 49941 17921
rect 49899 17872 49900 17912
rect 49940 17872 49941 17912
rect 49899 17863 49941 17872
rect 1315 17828 1373 17829
rect 1315 17788 1324 17828
rect 1364 17788 1373 17828
rect 1315 17787 1373 17788
rect 1699 17828 1757 17829
rect 1699 17788 1708 17828
rect 1748 17788 1757 17828
rect 1699 17787 1757 17788
rect 4011 17828 4053 17837
rect 4011 17788 4012 17828
rect 4052 17788 4053 17828
rect 4011 17779 4053 17788
rect 7363 17828 7421 17829
rect 7363 17788 7372 17828
rect 7412 17788 7421 17828
rect 7363 17787 7421 17788
rect 31747 17828 31805 17829
rect 31747 17788 31756 17828
rect 31796 17788 31805 17828
rect 31747 17787 31805 17788
rect 39907 17828 39965 17829
rect 39907 17788 39916 17828
rect 39956 17788 39965 17828
rect 39907 17787 39965 17788
rect 40291 17828 40349 17829
rect 40291 17788 40300 17828
rect 40340 17788 40349 17828
rect 40291 17787 40349 17788
rect 40491 17828 40533 17837
rect 40491 17788 40492 17828
rect 40532 17788 40533 17828
rect 40491 17779 40533 17788
rect 48547 17828 48605 17829
rect 48547 17788 48556 17828
rect 48596 17788 48605 17828
rect 48547 17787 48605 17788
rect 49123 17828 49181 17829
rect 49123 17788 49132 17828
rect 49172 17788 49181 17828
rect 49123 17787 49181 17788
rect 49315 17828 49373 17829
rect 49315 17788 49324 17828
rect 49364 17788 49373 17828
rect 49315 17787 49373 17788
rect 49803 17828 49845 17837
rect 49803 17788 49804 17828
rect 49844 17788 49845 17828
rect 49803 17779 49845 17788
rect 49995 17828 50037 17837
rect 49995 17788 49996 17828
rect 50036 17788 50037 17828
rect 49995 17779 50037 17788
rect 3715 17744 3773 17745
rect 3715 17704 3724 17744
rect 3764 17704 3773 17744
rect 3715 17703 3773 17704
rect 5155 17744 5213 17745
rect 5155 17704 5164 17744
rect 5204 17704 5213 17744
rect 5155 17703 5213 17704
rect 6019 17744 6077 17745
rect 6019 17704 6028 17744
rect 6068 17704 6077 17744
rect 6019 17703 6077 17704
rect 6411 17744 6453 17753
rect 6411 17704 6412 17744
rect 6452 17704 6453 17744
rect 6411 17695 6453 17704
rect 6787 17744 6845 17745
rect 6787 17704 6796 17744
rect 6836 17704 6845 17744
rect 6787 17703 6845 17704
rect 6891 17744 6933 17753
rect 6891 17704 6892 17744
rect 6932 17704 6933 17744
rect 6891 17695 6933 17704
rect 9955 17744 10013 17745
rect 9955 17704 9964 17744
rect 10004 17704 10013 17744
rect 9955 17703 10013 17704
rect 10059 17744 10101 17753
rect 10059 17704 10060 17744
rect 10100 17704 10101 17744
rect 10059 17695 10101 17704
rect 10915 17744 10973 17745
rect 10915 17704 10924 17744
rect 10964 17704 10973 17744
rect 10915 17703 10973 17704
rect 11779 17744 11837 17745
rect 11779 17704 11788 17744
rect 11828 17704 11837 17744
rect 11779 17703 11837 17704
rect 13131 17744 13173 17753
rect 13131 17704 13132 17744
rect 13172 17704 13173 17744
rect 13131 17695 13173 17704
rect 13323 17744 13365 17753
rect 13323 17704 13324 17744
rect 13364 17704 13365 17744
rect 13323 17695 13365 17704
rect 13411 17744 13469 17745
rect 13411 17704 13420 17744
rect 13460 17704 13469 17744
rect 13411 17703 13469 17704
rect 13699 17744 13757 17745
rect 13699 17704 13708 17744
rect 13748 17704 13757 17744
rect 13699 17703 13757 17704
rect 32131 17744 32189 17745
rect 32131 17704 32140 17744
rect 32180 17704 32189 17744
rect 32131 17703 32189 17704
rect 32235 17744 32277 17753
rect 32235 17704 32236 17744
rect 32276 17704 32277 17744
rect 32235 17695 32277 17704
rect 32427 17744 32469 17753
rect 32427 17704 32428 17744
rect 32468 17704 32469 17744
rect 32427 17695 32469 17704
rect 32715 17744 32757 17753
rect 32715 17704 32716 17744
rect 32756 17704 32757 17744
rect 32715 17695 32757 17704
rect 32811 17744 32853 17753
rect 32811 17704 32812 17744
rect 32852 17704 32853 17744
rect 32811 17695 32853 17704
rect 32907 17744 32949 17753
rect 32907 17704 32908 17744
rect 32948 17704 32949 17744
rect 32907 17695 32949 17704
rect 33099 17744 33141 17753
rect 33099 17704 33100 17744
rect 33140 17704 33141 17744
rect 33099 17695 33141 17704
rect 33187 17744 33245 17745
rect 33187 17704 33196 17744
rect 33236 17704 33245 17744
rect 33187 17703 33245 17704
rect 33387 17744 33429 17753
rect 33387 17704 33388 17744
rect 33428 17704 33429 17744
rect 33579 17744 33621 17753
rect 33387 17695 33429 17704
rect 33483 17723 33525 17732
rect 33483 17683 33484 17723
rect 33524 17683 33525 17723
rect 33579 17704 33580 17744
rect 33620 17704 33621 17744
rect 33579 17695 33621 17704
rect 33675 17744 33717 17753
rect 33675 17704 33676 17744
rect 33716 17704 33717 17744
rect 33675 17695 33717 17704
rect 37419 17744 37461 17753
rect 37419 17704 37420 17744
rect 37460 17704 37461 17744
rect 37419 17695 37461 17704
rect 37515 17744 37557 17753
rect 37515 17704 37516 17744
rect 37556 17704 37557 17744
rect 37515 17695 37557 17704
rect 37611 17744 37653 17753
rect 37611 17704 37612 17744
rect 37652 17704 37653 17744
rect 37611 17695 37653 17704
rect 37707 17744 37749 17753
rect 37707 17704 37708 17744
rect 37748 17704 37749 17744
rect 37707 17695 37749 17704
rect 38179 17744 38237 17745
rect 38179 17704 38188 17744
rect 38228 17704 38237 17744
rect 38179 17703 38237 17704
rect 41635 17744 41693 17745
rect 41635 17704 41644 17744
rect 41684 17704 41693 17744
rect 41635 17703 41693 17704
rect 42499 17744 42557 17745
rect 42499 17704 42508 17744
rect 42548 17704 42557 17744
rect 42499 17703 42557 17704
rect 43075 17744 43133 17745
rect 43075 17704 43084 17744
rect 43124 17704 43133 17744
rect 43075 17703 43133 17704
rect 43459 17744 43517 17745
rect 43459 17704 43468 17744
rect 43508 17704 43517 17744
rect 43459 17703 43517 17704
rect 43563 17744 43605 17753
rect 43563 17704 43564 17744
rect 43604 17704 43605 17744
rect 43563 17695 43605 17704
rect 44043 17744 44085 17753
rect 44043 17704 44044 17744
rect 44084 17704 44085 17744
rect 44043 17695 44085 17704
rect 44139 17744 44181 17753
rect 44139 17704 44140 17744
rect 44180 17704 44181 17744
rect 44139 17695 44181 17704
rect 44235 17744 44277 17753
rect 44235 17704 44236 17744
rect 44276 17704 44277 17744
rect 44235 17695 44277 17704
rect 44523 17744 44565 17753
rect 44523 17704 44524 17744
rect 44564 17704 44565 17744
rect 44523 17695 44565 17704
rect 44619 17744 44661 17753
rect 44619 17704 44620 17744
rect 44660 17704 44661 17744
rect 44619 17695 44661 17704
rect 44715 17744 44757 17753
rect 44715 17704 44716 17744
rect 44756 17704 44757 17744
rect 44715 17695 44757 17704
rect 44811 17744 44853 17753
rect 44811 17704 44812 17744
rect 44852 17704 44853 17744
rect 44811 17695 44853 17704
rect 45091 17744 45149 17745
rect 45091 17704 45100 17744
rect 45140 17704 45149 17744
rect 45091 17703 45149 17704
rect 46155 17744 46197 17753
rect 46155 17704 46156 17744
rect 46196 17704 46197 17744
rect 46155 17695 46197 17704
rect 46251 17744 46293 17753
rect 46251 17704 46252 17744
rect 46292 17704 46293 17744
rect 46251 17695 46293 17704
rect 46347 17744 46389 17753
rect 46347 17704 46348 17744
rect 46388 17704 46389 17744
rect 46347 17695 46389 17704
rect 46443 17744 46485 17753
rect 46443 17704 46444 17744
rect 46484 17704 46485 17744
rect 46443 17695 46485 17704
rect 47491 17744 47549 17745
rect 47491 17704 47500 17744
rect 47540 17704 47549 17744
rect 47491 17703 47549 17704
rect 49707 17744 49749 17753
rect 49707 17704 49708 17744
rect 49748 17704 49749 17744
rect 49707 17695 49749 17704
rect 50083 17744 50141 17745
rect 50083 17704 50092 17744
rect 50132 17704 50141 17744
rect 50083 17703 50141 17704
rect 50571 17744 50613 17753
rect 50571 17704 50572 17744
rect 50612 17704 50613 17744
rect 50571 17695 50613 17704
rect 50667 17744 50709 17753
rect 50667 17704 50668 17744
rect 50708 17704 50709 17744
rect 50667 17695 50709 17704
rect 50763 17744 50805 17753
rect 50763 17704 50764 17744
rect 50804 17704 50805 17744
rect 50763 17695 50805 17704
rect 50947 17744 51005 17745
rect 50947 17704 50956 17744
rect 50996 17704 51005 17744
rect 50947 17703 51005 17704
rect 51331 17744 51389 17745
rect 51331 17704 51340 17744
rect 51380 17704 51389 17744
rect 51331 17703 51389 17704
rect 52387 17744 52445 17745
rect 52387 17704 52396 17744
rect 52436 17704 52445 17744
rect 52387 17703 52445 17704
rect 52675 17744 52733 17745
rect 52675 17704 52684 17744
rect 52724 17704 52733 17744
rect 52675 17703 52733 17704
rect 33483 17674 33525 17683
rect 10539 17660 10581 17669
rect 10539 17620 10540 17660
rect 10580 17620 10581 17660
rect 10539 17611 10581 17620
rect 42891 17660 42933 17669
rect 42891 17620 42892 17660
rect 42932 17620 42933 17660
rect 42891 17611 42933 17620
rect 43747 17618 43805 17619
rect 1131 17576 1173 17585
rect 1131 17536 1132 17576
rect 1172 17536 1173 17576
rect 1131 17527 1173 17536
rect 1515 17576 1557 17585
rect 1515 17536 1516 17576
rect 1556 17536 1557 17576
rect 1515 17527 1557 17536
rect 7563 17576 7605 17585
rect 7563 17536 7564 17576
rect 7604 17536 7605 17576
rect 7563 17527 7605 17536
rect 9867 17572 9909 17581
rect 9867 17532 9868 17572
rect 9908 17532 9909 17572
rect 12931 17576 12989 17577
rect 12931 17536 12940 17576
rect 12980 17536 12989 17576
rect 12931 17535 12989 17536
rect 32323 17576 32381 17577
rect 32323 17536 32332 17576
rect 32372 17536 32381 17576
rect 32323 17535 32381 17536
rect 32611 17576 32669 17577
rect 32611 17536 32620 17576
rect 32660 17536 32669 17576
rect 32611 17535 32669 17536
rect 38283 17576 38325 17585
rect 38283 17536 38284 17576
rect 38324 17536 38325 17576
rect 6699 17518 6741 17527
rect 9867 17523 9909 17532
rect 38283 17527 38325 17536
rect 40107 17576 40149 17585
rect 40107 17536 40108 17576
rect 40148 17536 40149 17576
rect 40107 17527 40149 17536
rect 43179 17576 43221 17585
rect 43179 17536 43180 17576
rect 43220 17536 43221 17576
rect 43179 17527 43221 17536
rect 43371 17572 43413 17581
rect 43747 17578 43756 17618
rect 43796 17578 43805 17618
rect 43747 17577 43805 17578
rect 43371 17532 43372 17572
rect 43412 17532 43413 17572
rect 44323 17576 44381 17577
rect 44323 17536 44332 17576
rect 44372 17536 44381 17576
rect 44323 17535 44381 17536
rect 45003 17576 45045 17585
rect 45003 17536 45004 17576
rect 45044 17536 45045 17576
rect 43371 17523 43413 17532
rect 45003 17527 45045 17536
rect 47403 17576 47445 17585
rect 47403 17536 47404 17576
rect 47444 17536 47445 17576
rect 47403 17527 47445 17536
rect 48939 17576 48981 17585
rect 48939 17536 48940 17576
rect 48980 17536 48981 17576
rect 48939 17527 48981 17536
rect 49515 17576 49557 17585
rect 49515 17536 49516 17576
rect 49556 17536 49557 17576
rect 49515 17527 49557 17536
rect 50467 17576 50525 17577
rect 50467 17536 50476 17576
rect 50516 17536 50525 17576
rect 50467 17535 50525 17536
rect 51243 17576 51285 17585
rect 51243 17536 51244 17576
rect 51284 17536 51285 17576
rect 51243 17527 51285 17536
rect 52299 17576 52341 17585
rect 52299 17536 52300 17576
rect 52340 17536 52341 17576
rect 52299 17527 52341 17536
rect 52587 17576 52629 17585
rect 52587 17536 52588 17576
rect 52628 17536 52629 17576
rect 52587 17527 52629 17536
rect 6699 17478 6700 17518
rect 6740 17478 6741 17518
rect 6699 17469 6741 17478
rect 576 17408 52800 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 52800 17408
rect 576 17344 52800 17368
rect 6307 17240 6365 17241
rect 6307 17200 6316 17240
rect 6356 17200 6365 17240
rect 6307 17199 6365 17200
rect 29163 17240 29205 17249
rect 29163 17200 29164 17240
rect 29204 17200 29205 17240
rect 29163 17191 29205 17200
rect 32715 17244 32757 17253
rect 32715 17204 32716 17244
rect 32756 17204 32757 17244
rect 32715 17195 32757 17204
rect 41259 17240 41301 17249
rect 41259 17200 41260 17240
rect 41300 17200 41301 17240
rect 41259 17191 41301 17200
rect 32907 17156 32949 17165
rect 32907 17116 32908 17156
rect 32948 17116 32949 17156
rect 32907 17107 32949 17116
rect 50091 17156 50133 17165
rect 50091 17116 50092 17156
rect 50132 17116 50133 17156
rect 50091 17107 50133 17116
rect 40963 17083 41021 17084
rect 6027 17072 6069 17081
rect 6027 17032 6028 17072
rect 6068 17032 6069 17072
rect 6027 17023 6069 17032
rect 6123 17072 6165 17081
rect 6123 17032 6124 17072
rect 6164 17032 6165 17072
rect 6123 17023 6165 17032
rect 6219 17072 6261 17081
rect 6219 17032 6220 17072
rect 6260 17032 6261 17072
rect 6219 17023 6261 17032
rect 6507 17072 6549 17081
rect 6507 17032 6508 17072
rect 6548 17032 6549 17072
rect 6507 17023 6549 17032
rect 6883 17072 6941 17073
rect 6883 17032 6892 17072
rect 6932 17032 6941 17072
rect 6883 17031 6941 17032
rect 7083 17072 7125 17081
rect 7083 17032 7084 17072
rect 7124 17032 7125 17072
rect 7083 17023 7125 17032
rect 7459 17072 7517 17073
rect 7459 17032 7468 17072
rect 7508 17032 7517 17072
rect 7459 17031 7517 17032
rect 8323 17072 8381 17073
rect 8323 17032 8332 17072
rect 8372 17032 8381 17072
rect 8323 17031 8381 17032
rect 9763 17072 9821 17073
rect 9763 17032 9772 17072
rect 9812 17032 9821 17072
rect 9763 17031 9821 17032
rect 9867 17072 9909 17081
rect 9867 17032 9868 17072
rect 9908 17032 9909 17072
rect 9867 17023 9909 17032
rect 10059 17072 10101 17081
rect 10059 17032 10060 17072
rect 10100 17032 10101 17072
rect 10059 17023 10101 17032
rect 10347 17072 10389 17081
rect 10347 17032 10348 17072
rect 10388 17032 10389 17072
rect 10347 17023 10389 17032
rect 10723 17072 10781 17073
rect 10723 17032 10732 17072
rect 10772 17032 10781 17072
rect 10723 17031 10781 17032
rect 10923 17072 10965 17081
rect 10923 17032 10924 17072
rect 10964 17032 10965 17072
rect 10923 17023 10965 17032
rect 11011 17072 11069 17073
rect 11011 17032 11020 17072
rect 11060 17032 11069 17072
rect 11011 17031 11069 17032
rect 31171 17072 31229 17073
rect 31171 17032 31180 17072
rect 31220 17032 31229 17072
rect 31171 17031 31229 17032
rect 32523 17072 32565 17081
rect 32523 17032 32524 17072
rect 32564 17032 32565 17072
rect 32523 17023 32565 17032
rect 32611 17072 32669 17073
rect 32611 17032 32620 17072
rect 32660 17032 32669 17072
rect 32611 17031 32669 17032
rect 33283 17072 33341 17073
rect 33283 17032 33292 17072
rect 33332 17032 33341 17072
rect 33283 17031 33341 17032
rect 34147 17072 34205 17073
rect 34147 17032 34156 17072
rect 34196 17032 34205 17072
rect 34147 17031 34205 17032
rect 35595 17072 35637 17081
rect 35595 17032 35596 17072
rect 35636 17032 35637 17072
rect 35595 17023 35637 17032
rect 35971 17072 36029 17073
rect 35971 17032 35980 17072
rect 36020 17032 36029 17072
rect 35971 17031 36029 17032
rect 36835 17072 36893 17073
rect 36835 17032 36844 17072
rect 36884 17032 36893 17072
rect 36835 17031 36893 17032
rect 39043 17072 39101 17073
rect 39043 17032 39052 17072
rect 39092 17032 39101 17072
rect 40963 17043 40972 17083
rect 41012 17043 41021 17083
rect 40963 17042 41021 17043
rect 41155 17072 41213 17073
rect 39043 17031 39101 17032
rect 41155 17032 41164 17072
rect 41204 17032 41213 17072
rect 41155 17031 41213 17032
rect 43267 17072 43325 17073
rect 43267 17032 43276 17072
rect 43316 17032 43325 17072
rect 43267 17031 43325 17032
rect 43659 17072 43701 17081
rect 43659 17032 43660 17072
rect 43700 17032 43701 17072
rect 43659 17023 43701 17032
rect 44139 17072 44181 17081
rect 44139 17032 44140 17072
rect 44180 17032 44181 17072
rect 44139 17023 44181 17032
rect 44331 17072 44373 17081
rect 44331 17032 44332 17072
rect 44372 17032 44373 17072
rect 44331 17023 44373 17032
rect 44419 17072 44477 17073
rect 44419 17032 44428 17072
rect 44468 17032 44477 17072
rect 44419 17031 44477 17032
rect 45475 17072 45533 17073
rect 45475 17032 45484 17072
rect 45524 17032 45533 17072
rect 45475 17031 45533 17032
rect 46155 17072 46197 17081
rect 46155 17032 46156 17072
rect 46196 17032 46197 17072
rect 46155 17023 46197 17032
rect 46251 17072 46293 17081
rect 46251 17032 46252 17072
rect 46292 17032 46293 17072
rect 46251 17023 46293 17032
rect 46347 17072 46389 17081
rect 46347 17032 46348 17072
rect 46388 17032 46389 17072
rect 46347 17023 46389 17032
rect 46443 17072 46485 17081
rect 46443 17032 46444 17072
rect 46484 17032 46485 17072
rect 46443 17023 46485 17032
rect 46635 17072 46677 17081
rect 46635 17032 46636 17072
rect 46676 17032 46677 17072
rect 46635 17023 46677 17032
rect 46731 17072 46773 17081
rect 46731 17032 46732 17072
rect 46772 17032 46773 17072
rect 46731 17023 46773 17032
rect 46827 17072 46869 17081
rect 46827 17032 46828 17072
rect 46868 17032 46869 17072
rect 46827 17023 46869 17032
rect 46923 17072 46965 17081
rect 46923 17032 46924 17072
rect 46964 17032 46965 17072
rect 46923 17023 46965 17032
rect 47395 17072 47453 17073
rect 47395 17032 47404 17072
rect 47444 17032 47453 17072
rect 47395 17031 47453 17032
rect 48835 17072 48893 17073
rect 48835 17032 48844 17072
rect 48884 17032 48893 17072
rect 48835 17031 48893 17032
rect 49699 17072 49757 17073
rect 49699 17032 49708 17072
rect 49748 17032 49757 17072
rect 49699 17031 49757 17032
rect 50283 17072 50325 17081
rect 50283 17032 50284 17072
rect 50324 17032 50325 17072
rect 50283 17023 50325 17032
rect 50659 17072 50717 17073
rect 50659 17032 50668 17072
rect 50708 17032 50717 17072
rect 50659 17031 50717 17032
rect 51523 17072 51581 17073
rect 51523 17032 51532 17072
rect 51572 17032 51581 17072
rect 51523 17031 51581 17032
rect 2659 16988 2717 16989
rect 2659 16948 2668 16988
rect 2708 16948 2717 16988
rect 2659 16947 2717 16948
rect 6603 16988 6645 16997
rect 6603 16948 6604 16988
rect 6644 16948 6645 16988
rect 6603 16939 6645 16948
rect 6795 16988 6837 16997
rect 6795 16948 6796 16988
rect 6836 16948 6837 16988
rect 6795 16939 6837 16948
rect 10443 16988 10485 16997
rect 10443 16948 10444 16988
rect 10484 16948 10485 16988
rect 10443 16939 10485 16948
rect 10635 16988 10677 16997
rect 10635 16948 10636 16988
rect 10676 16948 10677 16988
rect 10635 16939 10677 16948
rect 29731 16988 29789 16989
rect 29731 16948 29740 16988
rect 29780 16948 29789 16988
rect 29731 16947 29789 16948
rect 35307 16988 35349 16997
rect 35307 16948 35308 16988
rect 35348 16948 35349 16988
rect 35307 16939 35349 16948
rect 37995 16988 38037 16997
rect 37995 16948 37996 16988
rect 38036 16948 38037 16988
rect 37995 16939 38037 16948
rect 39147 16988 39189 16997
rect 39147 16948 39148 16988
rect 39188 16948 39189 16988
rect 39147 16939 39189 16948
rect 40483 16988 40541 16989
rect 40483 16948 40492 16988
rect 40532 16948 40541 16988
rect 40483 16947 40541 16948
rect 43371 16988 43413 16997
rect 43371 16948 43372 16988
rect 43412 16948 43413 16988
rect 45763 16988 45821 16989
rect 43371 16939 43413 16948
rect 43563 16946 43605 16955
rect 45763 16948 45772 16988
rect 45812 16948 45821 16988
rect 45763 16947 45821 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 1035 16904 1077 16913
rect 1035 16864 1036 16904
rect 1076 16864 1077 16904
rect 1035 16855 1077 16864
rect 6699 16904 6741 16913
rect 6699 16864 6700 16904
rect 6740 16864 6741 16904
rect 6699 16855 6741 16864
rect 10059 16904 10101 16913
rect 10059 16864 10060 16904
rect 10100 16864 10101 16904
rect 10059 16855 10101 16864
rect 10539 16904 10581 16913
rect 10539 16864 10540 16904
rect 10580 16864 10581 16904
rect 10539 16855 10581 16864
rect 32235 16904 32277 16913
rect 32235 16864 32236 16904
rect 32276 16864 32277 16904
rect 43563 16906 43564 16946
rect 43604 16906 43605 16946
rect 43563 16897 43605 16906
rect 44139 16904 44181 16913
rect 32235 16855 32277 16864
rect 43467 16862 43509 16871
rect 2475 16820 2517 16829
rect 2475 16780 2476 16820
rect 2516 16780 2517 16820
rect 2475 16771 2517 16780
rect 9475 16820 9533 16821
rect 9475 16780 9484 16820
rect 9524 16780 9533 16820
rect 9475 16779 9533 16780
rect 40683 16820 40725 16829
rect 40683 16780 40684 16820
rect 40724 16780 40725 16820
rect 40683 16771 40725 16780
rect 40875 16820 40917 16829
rect 40875 16780 40876 16820
rect 40916 16780 40917 16820
rect 43467 16822 43468 16862
rect 43508 16822 43509 16862
rect 44139 16864 44140 16904
rect 44180 16864 44181 16904
rect 44139 16855 44181 16864
rect 43467 16813 43509 16822
rect 45579 16820 45621 16829
rect 40875 16771 40917 16780
rect 45579 16780 45580 16820
rect 45620 16780 45621 16820
rect 45579 16771 45621 16780
rect 45963 16820 46005 16829
rect 45963 16780 45964 16820
rect 46004 16780 46005 16820
rect 45963 16771 46005 16780
rect 47307 16820 47349 16829
rect 47307 16780 47308 16820
rect 47348 16780 47349 16820
rect 47307 16771 47349 16780
rect 47683 16820 47741 16821
rect 47683 16780 47692 16820
rect 47732 16780 47741 16820
rect 47683 16779 47741 16780
rect 52675 16820 52733 16821
rect 52675 16780 52684 16820
rect 52724 16780 52733 16820
rect 52675 16779 52733 16780
rect 576 16652 79584 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 79584 16652
rect 576 16588 79584 16612
rect 6603 16484 6645 16493
rect 6603 16444 6604 16484
rect 6644 16444 6645 16484
rect 6603 16435 6645 16444
rect 6891 16484 6933 16493
rect 6891 16444 6892 16484
rect 6932 16444 6933 16484
rect 6891 16435 6933 16444
rect 27627 16484 27669 16493
rect 27627 16444 27628 16484
rect 27668 16444 27669 16484
rect 27627 16435 27669 16444
rect 40483 16484 40541 16485
rect 40483 16444 40492 16484
rect 40532 16444 40541 16484
rect 40483 16443 40541 16444
rect 45475 16484 45533 16485
rect 45475 16444 45484 16484
rect 45524 16444 45533 16484
rect 45475 16443 45533 16444
rect 50379 16484 50421 16493
rect 50379 16444 50380 16484
rect 50420 16444 50421 16484
rect 50379 16435 50421 16444
rect 54883 16484 54941 16485
rect 54883 16444 54892 16484
rect 54932 16444 54941 16484
rect 54883 16443 54941 16444
rect 56331 16484 56373 16493
rect 56331 16444 56332 16484
rect 56372 16444 56373 16484
rect 56331 16435 56373 16444
rect 57003 16484 57045 16493
rect 57003 16444 57004 16484
rect 57044 16444 57045 16484
rect 57003 16435 57045 16444
rect 57291 16484 57333 16493
rect 57291 16444 57292 16484
rect 57332 16444 57333 16484
rect 57291 16435 57333 16444
rect 59595 16484 59637 16493
rect 59595 16444 59596 16484
rect 59636 16444 59637 16484
rect 59595 16435 59637 16444
rect 63915 16484 63957 16493
rect 63915 16444 63916 16484
rect 63956 16444 63957 16484
rect 63915 16435 63957 16444
rect 65739 16484 65781 16493
rect 65739 16444 65740 16484
rect 65780 16444 65781 16484
rect 65739 16435 65781 16444
rect 66123 16484 66165 16493
rect 66123 16444 66124 16484
rect 66164 16444 66165 16484
rect 66123 16435 66165 16444
rect 66699 16484 66741 16493
rect 66699 16444 66700 16484
rect 66740 16444 66741 16484
rect 66699 16435 66741 16444
rect 69283 16484 69341 16485
rect 69283 16444 69292 16484
rect 69332 16444 69341 16484
rect 69283 16443 69341 16444
rect 69963 16484 70005 16493
rect 69963 16444 69964 16484
rect 70004 16444 70005 16484
rect 69963 16435 70005 16444
rect 73419 16484 73461 16493
rect 73419 16444 73420 16484
rect 73460 16444 73461 16484
rect 73419 16435 73461 16444
rect 74187 16484 74229 16493
rect 74187 16444 74188 16484
rect 74228 16444 74229 16484
rect 74187 16435 74229 16444
rect 77835 16484 77877 16493
rect 77835 16444 77836 16484
rect 77876 16444 77877 16484
rect 77835 16435 77877 16444
rect 79467 16484 79509 16493
rect 79467 16444 79468 16484
rect 79508 16444 79509 16484
rect 79467 16435 79509 16444
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 32235 16400 32277 16409
rect 32235 16360 32236 16400
rect 32276 16360 32277 16400
rect 32235 16351 32277 16360
rect 46347 16400 46389 16409
rect 46347 16360 46348 16400
rect 46388 16360 46389 16400
rect 46347 16351 46389 16360
rect 71787 16400 71829 16409
rect 71787 16360 71788 16400
rect 71828 16360 71829 16400
rect 71787 16351 71829 16360
rect 60739 16327 60797 16328
rect 1699 16316 1757 16317
rect 1699 16276 1708 16316
rect 1748 16276 1757 16316
rect 1699 16275 1757 16276
rect 10531 16316 10589 16317
rect 10531 16276 10540 16316
rect 10580 16276 10589 16316
rect 10531 16275 10589 16276
rect 32139 16316 32181 16325
rect 32139 16276 32140 16316
rect 32180 16276 32181 16316
rect 32139 16267 32181 16276
rect 32331 16316 32373 16325
rect 32331 16276 32332 16316
rect 32372 16276 32373 16316
rect 32331 16267 32373 16276
rect 49707 16316 49749 16325
rect 49707 16276 49708 16316
rect 49748 16276 49749 16316
rect 49707 16267 49749 16276
rect 56035 16316 56093 16317
rect 56035 16276 56044 16316
rect 56084 16276 56093 16316
rect 56035 16275 56093 16276
rect 59107 16316 59165 16317
rect 59107 16276 59116 16316
rect 59156 16276 59165 16316
rect 60739 16287 60748 16327
rect 60788 16287 60797 16327
rect 60739 16286 60797 16287
rect 70339 16316 70397 16317
rect 59107 16275 59165 16276
rect 70339 16276 70348 16316
rect 70388 16276 70397 16316
rect 70339 16275 70397 16276
rect 70723 16316 70781 16317
rect 70723 16276 70732 16316
rect 70772 16276 70781 16316
rect 70723 16275 70781 16276
rect 70915 16316 70973 16317
rect 70915 16276 70924 16316
rect 70964 16276 70973 16316
rect 70915 16275 70973 16276
rect 75619 16316 75677 16317
rect 75619 16276 75628 16316
rect 75668 16276 75677 16316
rect 75619 16275 75677 16276
rect 76003 16316 76061 16317
rect 76003 16276 76012 16316
rect 76052 16276 76061 16316
rect 76003 16275 76061 16276
rect 78603 16316 78645 16325
rect 78603 16276 78604 16316
rect 78644 16276 78645 16316
rect 78603 16267 78645 16276
rect 6307 16232 6365 16233
rect 6307 16192 6316 16232
rect 6356 16192 6365 16232
rect 6307 16191 6365 16192
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 6603 16232 6645 16241
rect 6603 16192 6604 16232
rect 6644 16192 6645 16232
rect 6603 16183 6645 16192
rect 6979 16232 7037 16233
rect 6979 16192 6988 16232
rect 7028 16192 7037 16232
rect 6979 16191 7037 16192
rect 28291 16232 28349 16233
rect 28291 16192 28300 16232
rect 28340 16192 28349 16232
rect 28291 16191 28349 16192
rect 29931 16232 29973 16241
rect 29931 16192 29932 16232
rect 29972 16192 29973 16232
rect 29931 16183 29973 16192
rect 32035 16232 32093 16233
rect 32035 16192 32044 16232
rect 32084 16192 32093 16232
rect 32035 16191 32093 16192
rect 32427 16232 32469 16241
rect 32427 16192 32428 16232
rect 32468 16192 32469 16232
rect 32427 16183 32469 16192
rect 32811 16232 32853 16241
rect 32811 16192 32812 16232
rect 32852 16192 32853 16232
rect 32811 16183 32853 16192
rect 32907 16232 32949 16241
rect 32907 16192 32908 16232
rect 32948 16192 32949 16232
rect 32907 16183 32949 16192
rect 33003 16232 33045 16241
rect 33003 16192 33004 16232
rect 33044 16192 33045 16232
rect 33003 16183 33045 16192
rect 33099 16232 33141 16241
rect 33099 16192 33100 16232
rect 33140 16192 33141 16232
rect 33099 16183 33141 16192
rect 33387 16232 33429 16241
rect 33387 16192 33388 16232
rect 33428 16192 33429 16232
rect 33387 16183 33429 16192
rect 33475 16232 33533 16233
rect 33475 16192 33484 16232
rect 33524 16192 33533 16232
rect 33475 16191 33533 16192
rect 35499 16232 35541 16241
rect 35499 16192 35500 16232
rect 35540 16192 35541 16232
rect 35499 16183 35541 16192
rect 35595 16232 35637 16241
rect 35595 16192 35596 16232
rect 35636 16192 35637 16232
rect 35595 16183 35637 16192
rect 35691 16232 35733 16241
rect 35691 16192 35692 16232
rect 35732 16192 35733 16232
rect 35691 16183 35733 16192
rect 35787 16232 35829 16241
rect 35787 16192 35788 16232
rect 35828 16192 35829 16232
rect 35787 16183 35829 16192
rect 36171 16232 36213 16241
rect 36171 16192 36172 16232
rect 36212 16192 36213 16232
rect 36171 16183 36213 16192
rect 36267 16232 36309 16241
rect 36267 16192 36268 16232
rect 36308 16192 36309 16232
rect 36267 16183 36309 16192
rect 36363 16232 36405 16241
rect 36363 16192 36364 16232
rect 36404 16192 36405 16232
rect 36363 16183 36405 16192
rect 36835 16232 36893 16233
rect 36835 16192 36844 16232
rect 36884 16192 36893 16232
rect 36835 16191 36893 16192
rect 37707 16232 37749 16241
rect 37707 16192 37708 16232
rect 37748 16192 37749 16232
rect 37707 16183 37749 16192
rect 37803 16232 37845 16241
rect 37803 16192 37804 16232
rect 37844 16192 37845 16232
rect 37803 16183 37845 16192
rect 37899 16232 37941 16241
rect 37899 16192 37900 16232
rect 37940 16192 37941 16232
rect 37899 16183 37941 16192
rect 38467 16232 38525 16233
rect 38467 16192 38476 16232
rect 38516 16192 38525 16232
rect 38467 16191 38525 16192
rect 39331 16232 39389 16233
rect 39331 16192 39340 16232
rect 39380 16192 39389 16232
rect 39331 16191 39389 16192
rect 41059 16232 41117 16233
rect 41059 16192 41068 16232
rect 41108 16192 41117 16232
rect 41059 16191 41117 16192
rect 42883 16232 42941 16233
rect 42883 16192 42892 16232
rect 42932 16192 42941 16232
rect 42883 16191 42941 16192
rect 43459 16232 43517 16233
rect 43459 16192 43468 16232
rect 43508 16192 43517 16232
rect 43459 16191 43517 16192
rect 44323 16232 44381 16233
rect 44323 16192 44332 16232
rect 44372 16192 44381 16232
rect 44323 16191 44381 16192
rect 45955 16232 46013 16233
rect 45955 16192 45964 16232
rect 46004 16192 46013 16232
rect 45955 16191 46013 16192
rect 46059 16232 46101 16241
rect 46059 16192 46060 16232
rect 46100 16192 46101 16232
rect 46059 16183 46101 16192
rect 46539 16232 46581 16241
rect 46539 16192 46540 16232
rect 46580 16192 46581 16232
rect 46539 16183 46581 16192
rect 46915 16232 46973 16233
rect 46915 16192 46924 16232
rect 46964 16192 46973 16232
rect 46915 16191 46973 16192
rect 47779 16232 47837 16233
rect 47779 16192 47788 16232
rect 47828 16192 47837 16232
rect 47779 16191 47837 16192
rect 49603 16232 49661 16233
rect 49603 16192 49612 16232
rect 49652 16192 49661 16232
rect 49603 16191 49661 16192
rect 49987 16232 50045 16233
rect 49987 16192 49996 16232
rect 50036 16192 50045 16232
rect 49987 16191 50045 16192
rect 50091 16232 50133 16241
rect 50091 16192 50092 16232
rect 50132 16192 50133 16232
rect 50091 16183 50133 16192
rect 50571 16232 50613 16241
rect 50571 16192 50572 16232
rect 50612 16192 50613 16232
rect 50571 16183 50613 16192
rect 50667 16232 50709 16241
rect 50667 16192 50668 16232
rect 50708 16192 50709 16232
rect 50667 16183 50709 16192
rect 50763 16232 50805 16241
rect 50763 16192 50764 16232
rect 50804 16192 50805 16232
rect 50763 16183 50805 16192
rect 50859 16232 50901 16241
rect 50859 16192 50860 16232
rect 50900 16192 50901 16232
rect 50859 16183 50901 16192
rect 51043 16232 51101 16233
rect 51043 16192 51052 16232
rect 51092 16192 51101 16232
rect 51043 16191 51101 16192
rect 52195 16232 52253 16233
rect 52195 16192 52204 16232
rect 52244 16192 52253 16232
rect 52195 16191 52253 16192
rect 52867 16232 52925 16233
rect 52867 16192 52876 16232
rect 52916 16192 52925 16232
rect 52867 16191 52925 16192
rect 53731 16232 53789 16233
rect 53731 16192 53740 16232
rect 53780 16192 53789 16232
rect 53731 16191 53789 16192
rect 55179 16232 55221 16241
rect 55179 16192 55180 16232
rect 55220 16192 55221 16232
rect 55179 16183 55221 16192
rect 55275 16232 55317 16241
rect 55275 16192 55276 16232
rect 55316 16192 55317 16232
rect 55275 16183 55317 16192
rect 55371 16232 55413 16241
rect 55371 16192 55372 16232
rect 55412 16192 55413 16232
rect 55371 16183 55413 16192
rect 56227 16232 56285 16233
rect 56227 16192 56236 16232
rect 56276 16192 56285 16232
rect 56227 16191 56285 16192
rect 56611 16232 56669 16233
rect 56611 16192 56620 16232
rect 56660 16192 56669 16232
rect 56611 16191 56669 16192
rect 56899 16232 56957 16233
rect 56899 16192 56908 16232
rect 56948 16192 56957 16232
rect 56899 16191 56957 16192
rect 57187 16232 57245 16233
rect 57187 16192 57196 16232
rect 57236 16192 57245 16232
rect 57187 16191 57245 16192
rect 58059 16232 58101 16241
rect 58059 16192 58060 16232
rect 58100 16192 58101 16232
rect 58059 16183 58101 16192
rect 58155 16232 58197 16241
rect 58155 16192 58156 16232
rect 58196 16192 58197 16232
rect 58155 16183 58197 16192
rect 58251 16232 58293 16241
rect 58251 16192 58252 16232
rect 58292 16192 58293 16232
rect 58251 16183 58293 16192
rect 58635 16232 58677 16241
rect 58635 16192 58636 16232
rect 58676 16192 58677 16232
rect 58635 16183 58677 16192
rect 58731 16232 58773 16241
rect 58731 16192 58732 16232
rect 58772 16192 58773 16232
rect 58731 16183 58773 16192
rect 58827 16232 58869 16241
rect 58827 16192 58828 16232
rect 58868 16192 58869 16232
rect 58827 16183 58869 16192
rect 59491 16232 59549 16233
rect 59491 16192 59500 16232
rect 59540 16192 59549 16232
rect 59491 16191 59549 16192
rect 60067 16232 60125 16233
rect 60067 16192 60076 16232
rect 60116 16192 60125 16232
rect 60067 16191 60125 16192
rect 60459 16232 60501 16241
rect 60459 16192 60460 16232
rect 60500 16192 60501 16232
rect 60459 16183 60501 16192
rect 60547 16232 60605 16233
rect 60547 16192 60556 16232
rect 60596 16192 60605 16232
rect 60547 16191 60605 16192
rect 61507 16232 61565 16233
rect 61507 16192 61516 16232
rect 61556 16192 61565 16232
rect 61507 16191 61565 16192
rect 62371 16232 62429 16233
rect 62371 16192 62380 16232
rect 62420 16192 62429 16232
rect 62371 16191 62429 16192
rect 63811 16232 63869 16233
rect 63811 16192 63820 16232
rect 63860 16192 63869 16232
rect 63811 16191 63869 16192
rect 65635 16232 65693 16233
rect 65635 16192 65644 16232
rect 65684 16192 65693 16232
rect 65635 16191 65693 16192
rect 66019 16232 66077 16233
rect 66019 16192 66028 16232
rect 66068 16192 66077 16232
rect 66019 16191 66077 16192
rect 66315 16232 66357 16241
rect 66315 16192 66316 16232
rect 66356 16192 66357 16232
rect 66315 16183 66357 16192
rect 66595 16232 66653 16233
rect 66595 16192 66604 16232
rect 66644 16192 66653 16232
rect 66595 16191 66653 16192
rect 67267 16232 67325 16233
rect 67267 16192 67276 16232
rect 67316 16192 67325 16232
rect 67267 16191 67325 16192
rect 68131 16232 68189 16233
rect 68131 16192 68140 16232
rect 68180 16192 68189 16232
rect 68131 16191 68189 16192
rect 69571 16232 69629 16233
rect 69571 16192 69580 16232
rect 69620 16192 69629 16232
rect 69571 16191 69629 16192
rect 69675 16232 69717 16241
rect 69675 16192 69676 16232
rect 69716 16192 69717 16232
rect 69675 16183 69717 16192
rect 69859 16232 69917 16233
rect 69859 16192 69868 16232
rect 69908 16192 69917 16232
rect 69859 16191 69917 16192
rect 72163 16232 72221 16233
rect 72163 16192 72172 16232
rect 72212 16192 72221 16232
rect 72163 16191 72221 16192
rect 72451 16232 72509 16233
rect 72451 16192 72460 16232
rect 72500 16192 72509 16232
rect 72451 16191 72509 16192
rect 73315 16232 73373 16233
rect 73315 16192 73324 16232
rect 73364 16192 73373 16232
rect 73315 16191 73373 16192
rect 74083 16232 74141 16233
rect 74083 16192 74092 16232
rect 74132 16192 74141 16232
rect 74083 16191 74141 16192
rect 75331 16232 75389 16233
rect 75331 16192 75340 16232
rect 75380 16192 75389 16232
rect 75331 16191 75389 16192
rect 77731 16232 77789 16233
rect 77731 16192 77740 16232
rect 77780 16192 77789 16232
rect 77731 16191 77789 16192
rect 78499 16232 78557 16233
rect 78499 16192 78508 16232
rect 78548 16192 78557 16232
rect 78499 16191 78557 16192
rect 79363 16232 79421 16233
rect 79363 16192 79372 16232
rect 79412 16192 79421 16232
rect 79363 16191 79421 16192
rect 37611 16148 37653 16157
rect 37611 16108 37612 16148
rect 37652 16108 37653 16148
rect 37611 16099 37653 16108
rect 38091 16148 38133 16157
rect 38091 16108 38092 16148
rect 38132 16108 38133 16148
rect 38091 16099 38133 16108
rect 42795 16148 42837 16157
rect 42795 16108 42796 16148
rect 42836 16108 42837 16148
rect 42795 16099 42837 16108
rect 43083 16148 43125 16157
rect 43083 16108 43084 16148
rect 43124 16108 43125 16148
rect 43083 16099 43125 16108
rect 52491 16148 52533 16157
rect 52491 16108 52492 16148
rect 52532 16108 52533 16148
rect 52491 16099 52533 16108
rect 61131 16148 61173 16157
rect 61131 16108 61132 16148
rect 61172 16108 61173 16148
rect 61131 16099 61173 16108
rect 66891 16148 66933 16157
rect 66891 16108 66892 16148
rect 66932 16108 66933 16148
rect 66891 16099 66933 16108
rect 1515 16064 1557 16073
rect 1515 16024 1516 16064
rect 1556 16024 1557 16064
rect 1515 16015 1557 16024
rect 10347 16064 10389 16073
rect 10347 16024 10348 16064
rect 10388 16024 10389 16064
rect 10347 16015 10389 16024
rect 36067 16064 36125 16065
rect 36067 16024 36076 16064
rect 36116 16024 36125 16064
rect 36067 16023 36125 16024
rect 36747 16064 36789 16073
rect 36747 16024 36748 16064
rect 36788 16024 36789 16064
rect 36747 16015 36789 16024
rect 41163 16064 41205 16073
rect 41163 16024 41164 16064
rect 41204 16024 41205 16064
rect 41163 16015 41205 16024
rect 45867 16060 45909 16069
rect 45867 16020 45868 16060
rect 45908 16020 45909 16060
rect 48931 16064 48989 16065
rect 48931 16024 48940 16064
rect 48980 16024 48989 16064
rect 48931 16023 48989 16024
rect 49899 16060 49941 16069
rect 45867 16011 45909 16020
rect 49899 16020 49900 16060
rect 49940 16020 49941 16060
rect 49899 16011 49941 16020
rect 51147 16064 51189 16073
rect 51147 16024 51148 16064
rect 51188 16024 51189 16064
rect 51147 16015 51189 16024
rect 52299 16064 52341 16073
rect 52299 16024 52300 16064
rect 52340 16024 52341 16064
rect 52299 16015 52341 16024
rect 55075 16064 55133 16065
rect 55075 16024 55084 16064
rect 55124 16024 55133 16064
rect 55075 16023 55133 16024
rect 55851 16064 55893 16073
rect 55851 16024 55852 16064
rect 55892 16024 55893 16064
rect 55851 16015 55893 16024
rect 56715 16064 56757 16073
rect 56715 16024 56716 16064
rect 56756 16024 56757 16064
rect 56715 16015 56757 16024
rect 57291 16064 57333 16073
rect 57291 16024 57292 16064
rect 57332 16024 57333 16064
rect 57291 16015 57333 16024
rect 58339 16064 58397 16065
rect 58339 16024 58348 16064
rect 58388 16024 58397 16064
rect 58339 16023 58397 16024
rect 58915 16064 58973 16065
rect 58915 16024 58924 16064
rect 58964 16024 58973 16064
rect 58915 16023 58973 16024
rect 59307 16064 59349 16073
rect 59307 16024 59308 16064
rect 59348 16024 59349 16064
rect 59307 16015 59349 16024
rect 60171 16064 60213 16073
rect 60171 16024 60172 16064
rect 60212 16024 60213 16064
rect 60171 16015 60213 16024
rect 60939 16064 60981 16073
rect 60939 16024 60940 16064
rect 60980 16024 60981 16064
rect 60939 16015 60981 16024
rect 63523 16064 63581 16065
rect 63523 16024 63532 16064
rect 63572 16024 63581 16064
rect 63523 16023 63581 16024
rect 66123 16064 66165 16073
rect 66123 16024 66124 16064
rect 66164 16024 66165 16064
rect 66123 16015 66165 16024
rect 66699 16064 66741 16073
rect 66699 16024 66700 16064
rect 66740 16024 66741 16064
rect 66699 16015 66741 16024
rect 69283 16064 69341 16065
rect 69283 16024 69292 16064
rect 69332 16024 69341 16064
rect 69283 16023 69341 16024
rect 69963 16064 70005 16073
rect 69963 16024 69964 16064
rect 70004 16024 70005 16064
rect 69963 16015 70005 16024
rect 70155 16064 70197 16073
rect 70155 16024 70156 16064
rect 70196 16024 70197 16064
rect 70155 16015 70197 16024
rect 70539 16064 70581 16073
rect 70539 16024 70540 16064
rect 70580 16024 70581 16064
rect 70539 16015 70581 16024
rect 71115 16064 71157 16073
rect 71115 16024 71116 16064
rect 71156 16024 71157 16064
rect 71115 16015 71157 16024
rect 72267 16064 72309 16073
rect 72267 16024 72268 16064
rect 72308 16024 72309 16064
rect 72267 16015 72309 16024
rect 72555 16064 72597 16073
rect 72555 16024 72556 16064
rect 72596 16024 72597 16064
rect 72555 16015 72597 16024
rect 73419 16064 73461 16073
rect 73419 16024 73420 16064
rect 73460 16024 73461 16064
rect 73419 16015 73461 16024
rect 74187 16064 74229 16073
rect 74187 16024 74188 16064
rect 74228 16024 74229 16064
rect 74187 16015 74229 16024
rect 75435 16064 75477 16073
rect 75435 16024 75436 16064
rect 75476 16024 75477 16064
rect 75435 16015 75477 16024
rect 75819 16064 75861 16073
rect 75819 16024 75820 16064
rect 75860 16024 75861 16064
rect 75819 16015 75861 16024
rect 76203 16064 76245 16073
rect 76203 16024 76204 16064
rect 76244 16024 76245 16064
rect 76203 16015 76245 16024
rect 76387 16064 76445 16065
rect 76387 16024 76396 16064
rect 76436 16024 76445 16064
rect 76387 16023 76445 16024
rect 77835 16064 77877 16073
rect 77835 16024 77836 16064
rect 77876 16024 77877 16064
rect 77835 16015 77877 16024
rect 576 15896 79584 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 79584 15896
rect 576 15832 79584 15856
rect 75531 15786 75573 15795
rect 75531 15746 75532 15786
rect 75572 15746 75573 15786
rect 35979 15732 36021 15741
rect 34051 15728 34109 15729
rect 34051 15688 34060 15728
rect 34100 15688 34109 15728
rect 34051 15687 34109 15688
rect 35979 15692 35980 15732
rect 36020 15692 36021 15732
rect 35979 15683 36021 15692
rect 36171 15728 36213 15737
rect 36171 15688 36172 15728
rect 36212 15688 36213 15728
rect 36171 15679 36213 15688
rect 38187 15732 38229 15741
rect 75531 15737 75573 15746
rect 38187 15692 38188 15732
rect 38228 15692 38229 15732
rect 38187 15683 38229 15692
rect 39811 15728 39869 15729
rect 39811 15688 39820 15728
rect 39860 15688 39869 15728
rect 39811 15687 39869 15688
rect 42403 15728 42461 15729
rect 42403 15688 42412 15728
rect 42452 15688 42461 15728
rect 42403 15687 42461 15688
rect 52291 15728 52349 15729
rect 52291 15688 52300 15728
rect 52340 15688 52349 15728
rect 52291 15687 52349 15688
rect 57763 15728 57821 15729
rect 57763 15688 57772 15728
rect 57812 15688 57821 15728
rect 57763 15687 57821 15688
rect 60355 15728 60413 15729
rect 60355 15688 60364 15728
rect 60404 15688 60413 15728
rect 60355 15687 60413 15688
rect 60931 15728 60989 15729
rect 60931 15688 60940 15728
rect 60980 15688 60989 15728
rect 60931 15687 60989 15688
rect 61611 15728 61653 15737
rect 61611 15688 61612 15728
rect 61652 15688 61653 15728
rect 61611 15679 61653 15688
rect 66883 15728 66941 15729
rect 66883 15688 66892 15728
rect 66932 15688 66941 15728
rect 66883 15687 66941 15688
rect 69859 15728 69917 15729
rect 69859 15688 69868 15728
rect 69908 15688 69917 15728
rect 69859 15687 69917 15688
rect 72739 15728 72797 15729
rect 72739 15688 72748 15728
rect 72788 15688 72797 15728
rect 72739 15687 72797 15688
rect 72931 15728 72989 15729
rect 72931 15688 72940 15728
rect 72980 15688 72989 15728
rect 72931 15687 72989 15688
rect 78787 15728 78845 15729
rect 78787 15688 78796 15728
rect 78836 15688 78845 15728
rect 78787 15687 78845 15688
rect 31659 15644 31701 15653
rect 31659 15604 31660 15644
rect 31700 15604 31701 15644
rect 31659 15595 31701 15604
rect 38379 15644 38421 15653
rect 38379 15604 38380 15644
rect 38420 15604 38421 15644
rect 38379 15595 38421 15604
rect 40011 15644 40053 15653
rect 40011 15604 40012 15644
rect 40052 15604 40053 15644
rect 40011 15595 40053 15604
rect 55371 15644 55413 15653
rect 55371 15604 55372 15644
rect 55412 15604 55413 15644
rect 55371 15595 55413 15604
rect 57963 15644 58005 15653
rect 57963 15604 57964 15644
rect 58004 15604 58005 15644
rect 57963 15595 58005 15604
rect 67467 15644 67509 15653
rect 67467 15604 67468 15644
rect 67508 15604 67509 15644
rect 67467 15595 67509 15604
rect 70347 15644 70389 15653
rect 70347 15604 70348 15644
rect 70388 15604 70389 15644
rect 70347 15595 70389 15604
rect 61995 15581 62037 15590
rect 27619 15560 27677 15561
rect 27619 15520 27628 15560
rect 27668 15520 27677 15560
rect 27619 15519 27677 15520
rect 32035 15560 32093 15561
rect 32035 15520 32044 15560
rect 32084 15520 32093 15560
rect 32035 15519 32093 15520
rect 32899 15560 32957 15561
rect 32899 15520 32908 15560
rect 32948 15520 32957 15560
rect 32899 15519 32957 15520
rect 34243 15560 34301 15561
rect 34243 15520 34252 15560
rect 34292 15520 34301 15560
rect 34243 15519 34301 15520
rect 34347 15560 34389 15569
rect 34347 15520 34348 15560
rect 34388 15520 34389 15560
rect 34347 15511 34389 15520
rect 34539 15560 34581 15569
rect 34539 15520 34540 15560
rect 34580 15520 34581 15560
rect 34539 15511 34581 15520
rect 34731 15560 34773 15569
rect 34731 15520 34732 15560
rect 34772 15520 34773 15560
rect 34731 15511 34773 15520
rect 35107 15560 35165 15561
rect 35107 15520 35116 15560
rect 35156 15520 35165 15560
rect 35107 15519 35165 15520
rect 35787 15560 35829 15569
rect 35787 15520 35788 15560
rect 35828 15520 35829 15560
rect 35787 15511 35829 15520
rect 35875 15560 35933 15561
rect 35875 15520 35884 15560
rect 35924 15520 35933 15560
rect 35875 15519 35933 15520
rect 36259 15560 36317 15561
rect 36259 15520 36268 15560
rect 36308 15520 36317 15560
rect 36259 15519 36317 15520
rect 36643 15560 36701 15561
rect 36643 15520 36652 15560
rect 36692 15520 36701 15560
rect 36643 15519 36701 15520
rect 36747 15560 36789 15569
rect 36747 15520 36748 15560
rect 36788 15520 36789 15560
rect 37995 15560 38037 15569
rect 36747 15511 36789 15520
rect 36939 15549 36981 15558
rect 36939 15509 36940 15549
rect 36980 15509 36981 15549
rect 37995 15520 37996 15560
rect 38036 15520 38037 15560
rect 37995 15511 38037 15520
rect 38083 15560 38141 15561
rect 38083 15520 38092 15560
rect 38132 15520 38141 15560
rect 38083 15519 38141 15520
rect 38475 15560 38517 15569
rect 38475 15520 38476 15560
rect 38516 15520 38517 15560
rect 38475 15511 38517 15520
rect 38571 15560 38613 15569
rect 38571 15520 38572 15560
rect 38612 15520 38613 15560
rect 38571 15511 38613 15520
rect 38667 15560 38709 15569
rect 38667 15520 38668 15560
rect 38708 15520 38709 15560
rect 38667 15511 38709 15520
rect 39531 15560 39573 15569
rect 39531 15520 39532 15560
rect 39572 15520 39573 15560
rect 39531 15511 39573 15520
rect 39627 15560 39669 15569
rect 39627 15520 39628 15560
rect 39668 15520 39669 15560
rect 39627 15511 39669 15520
rect 39723 15560 39765 15569
rect 39723 15520 39724 15560
rect 39764 15520 39765 15560
rect 39723 15511 39765 15520
rect 40387 15560 40445 15561
rect 40387 15520 40396 15560
rect 40436 15520 40445 15560
rect 40387 15519 40445 15520
rect 41251 15560 41309 15561
rect 41251 15520 41260 15560
rect 41300 15520 41309 15560
rect 41251 15519 41309 15520
rect 42603 15560 42645 15569
rect 42603 15520 42604 15560
rect 42644 15520 42645 15560
rect 42603 15511 42645 15520
rect 42979 15560 43037 15561
rect 42979 15520 42988 15560
rect 43028 15520 43037 15560
rect 42979 15519 43037 15520
rect 43843 15560 43901 15561
rect 43843 15520 43852 15560
rect 43892 15520 43901 15560
rect 43843 15519 43901 15520
rect 45675 15560 45717 15569
rect 45675 15520 45676 15560
rect 45716 15520 45717 15560
rect 45675 15511 45717 15520
rect 46723 15560 46781 15561
rect 46723 15520 46732 15560
rect 46772 15520 46781 15560
rect 46723 15519 46781 15520
rect 47115 15560 47157 15569
rect 47115 15520 47116 15560
rect 47156 15520 47157 15560
rect 47115 15511 47157 15520
rect 47307 15560 47349 15569
rect 47307 15520 47308 15560
rect 47348 15520 47349 15560
rect 47307 15511 47349 15520
rect 47499 15560 47541 15569
rect 47499 15520 47500 15560
rect 47540 15520 47541 15560
rect 47499 15511 47541 15520
rect 47587 15560 47645 15561
rect 47587 15520 47596 15560
rect 47636 15520 47645 15560
rect 47587 15519 47645 15520
rect 47779 15560 47837 15561
rect 47779 15520 47788 15560
rect 47828 15520 47837 15560
rect 47779 15519 47837 15520
rect 49035 15560 49077 15569
rect 49035 15520 49036 15560
rect 49076 15520 49077 15560
rect 49035 15511 49077 15520
rect 49131 15560 49173 15569
rect 49131 15520 49132 15560
rect 49172 15520 49173 15560
rect 49131 15511 49173 15520
rect 49227 15560 49269 15569
rect 49227 15520 49228 15560
rect 49268 15520 49269 15560
rect 49227 15511 49269 15520
rect 49323 15560 49365 15569
rect 49323 15520 49324 15560
rect 49364 15520 49365 15560
rect 49323 15511 49365 15520
rect 49707 15560 49749 15569
rect 49707 15520 49708 15560
rect 49748 15520 49749 15560
rect 49707 15511 49749 15520
rect 49803 15560 49845 15569
rect 49803 15520 49804 15560
rect 49844 15520 49845 15560
rect 49803 15511 49845 15520
rect 49899 15560 49941 15569
rect 49899 15520 49900 15560
rect 49940 15520 49941 15560
rect 49899 15511 49941 15520
rect 49995 15560 50037 15569
rect 49995 15520 49996 15560
rect 50036 15520 50037 15560
rect 49995 15511 50037 15520
rect 52395 15560 52437 15569
rect 52395 15520 52396 15560
rect 52436 15520 52437 15560
rect 52395 15511 52437 15520
rect 52491 15560 52533 15569
rect 52491 15520 52492 15560
rect 52532 15520 52533 15560
rect 52491 15511 52533 15520
rect 52587 15560 52629 15569
rect 52587 15520 52588 15560
rect 52628 15520 52629 15560
rect 52587 15511 52629 15520
rect 53059 15560 53117 15561
rect 53059 15520 53068 15560
rect 53108 15520 53117 15560
rect 53059 15519 53117 15520
rect 55747 15560 55805 15561
rect 55747 15520 55756 15560
rect 55796 15520 55805 15560
rect 55747 15519 55805 15520
rect 56611 15560 56669 15561
rect 56611 15520 56620 15560
rect 56660 15520 56669 15560
rect 56611 15519 56669 15520
rect 58339 15560 58397 15561
rect 58339 15520 58348 15560
rect 58388 15520 58397 15560
rect 58339 15519 58397 15520
rect 59203 15560 59261 15561
rect 59203 15520 59212 15560
rect 59252 15520 59261 15560
rect 59203 15519 59261 15520
rect 61035 15560 61077 15569
rect 61035 15520 61036 15560
rect 61076 15520 61077 15560
rect 61035 15511 61077 15520
rect 61131 15560 61173 15569
rect 61131 15520 61132 15560
rect 61172 15520 61173 15560
rect 61131 15511 61173 15520
rect 61227 15560 61269 15569
rect 61227 15520 61228 15560
rect 61268 15520 61269 15560
rect 61227 15511 61269 15520
rect 61803 15560 61845 15569
rect 61803 15520 61804 15560
rect 61844 15520 61845 15560
rect 61803 15511 61845 15520
rect 61899 15560 61941 15569
rect 61899 15520 61900 15560
rect 61940 15520 61941 15560
rect 61995 15541 61996 15581
rect 62036 15541 62037 15581
rect 61995 15532 62037 15541
rect 62091 15560 62133 15569
rect 61899 15511 61941 15520
rect 62091 15520 62092 15560
rect 62132 15520 62133 15560
rect 62091 15511 62133 15520
rect 66987 15560 67029 15569
rect 66987 15520 66988 15560
rect 67028 15520 67029 15560
rect 66987 15511 67029 15520
rect 67083 15560 67125 15569
rect 67083 15520 67084 15560
rect 67124 15520 67125 15560
rect 67083 15511 67125 15520
rect 67179 15560 67221 15569
rect 67179 15520 67180 15560
rect 67220 15520 67221 15560
rect 67179 15511 67221 15520
rect 67555 15560 67613 15561
rect 67555 15520 67564 15560
rect 67604 15520 67613 15560
rect 67555 15519 67613 15520
rect 67947 15560 67989 15569
rect 67947 15520 67948 15560
rect 67988 15520 67989 15560
rect 67947 15511 67989 15520
rect 68043 15560 68085 15569
rect 68043 15520 68044 15560
rect 68084 15520 68085 15560
rect 68043 15511 68085 15520
rect 68139 15560 68181 15569
rect 68139 15520 68140 15560
rect 68180 15520 68181 15560
rect 68139 15511 68181 15520
rect 68235 15560 68277 15569
rect 68235 15520 68236 15560
rect 68276 15520 68277 15560
rect 68235 15511 68277 15520
rect 68419 15560 68477 15561
rect 68419 15520 68428 15560
rect 68468 15520 68477 15560
rect 68419 15519 68477 15520
rect 69963 15560 70005 15569
rect 69963 15520 69964 15560
rect 70004 15520 70005 15560
rect 69963 15511 70005 15520
rect 70059 15560 70101 15569
rect 70059 15520 70060 15560
rect 70100 15520 70101 15560
rect 70059 15511 70101 15520
rect 70155 15560 70197 15569
rect 70155 15520 70156 15560
rect 70196 15520 70197 15560
rect 70155 15511 70197 15520
rect 70723 15560 70781 15561
rect 70723 15520 70732 15560
rect 70772 15520 70781 15560
rect 70723 15519 70781 15520
rect 71587 15560 71645 15561
rect 71587 15520 71596 15560
rect 71636 15520 71645 15560
rect 71587 15519 71645 15520
rect 74083 15560 74141 15561
rect 74083 15520 74092 15560
rect 74132 15520 74141 15560
rect 74083 15519 74141 15520
rect 74947 15560 75005 15561
rect 74947 15520 74956 15560
rect 74996 15520 75005 15560
rect 74947 15519 75005 15520
rect 75339 15560 75381 15569
rect 75339 15520 75340 15560
rect 75380 15520 75381 15560
rect 75339 15511 75381 15520
rect 75619 15560 75677 15561
rect 75619 15520 75628 15560
rect 75668 15520 75677 15560
rect 75619 15519 75677 15520
rect 75723 15560 75765 15569
rect 75723 15520 75724 15560
rect 75764 15520 75765 15560
rect 75723 15511 75765 15520
rect 76395 15560 76437 15569
rect 76395 15520 76396 15560
rect 76436 15520 76437 15560
rect 76395 15511 76437 15520
rect 76771 15560 76829 15561
rect 76771 15520 76780 15560
rect 76820 15520 76829 15560
rect 76771 15519 76829 15520
rect 77635 15560 77693 15561
rect 77635 15520 77644 15560
rect 77684 15520 77693 15560
rect 77635 15519 77693 15520
rect 36939 15500 36981 15509
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 1699 15476 1757 15477
rect 1699 15436 1708 15476
rect 1748 15436 1757 15476
rect 1699 15435 1757 15436
rect 34827 15476 34869 15485
rect 34827 15436 34828 15476
rect 34868 15436 34869 15476
rect 34827 15427 34869 15436
rect 35019 15476 35061 15485
rect 35019 15436 35020 15476
rect 35060 15436 35061 15476
rect 35019 15427 35061 15436
rect 46827 15476 46869 15485
rect 46827 15436 46828 15476
rect 46868 15436 46869 15476
rect 46827 15427 46869 15436
rect 47019 15476 47061 15485
rect 47019 15436 47020 15476
rect 47060 15436 47061 15476
rect 47019 15427 47061 15436
rect 61411 15476 61469 15477
rect 61411 15436 61420 15476
rect 61460 15436 61469 15476
rect 61411 15435 61469 15436
rect 62275 15476 62333 15477
rect 62275 15436 62284 15476
rect 62324 15436 62333 15476
rect 62275 15435 62333 15436
rect 65059 15476 65117 15477
rect 65059 15436 65068 15476
rect 65108 15436 65117 15476
rect 65059 15435 65117 15436
rect 68523 15476 68565 15485
rect 68523 15436 68524 15476
rect 68564 15436 68565 15476
rect 68523 15427 68565 15436
rect 69475 15476 69533 15477
rect 69475 15436 69484 15476
rect 69524 15436 69533 15476
rect 69475 15435 69533 15436
rect 1515 15392 1557 15401
rect 1515 15352 1516 15392
rect 1556 15352 1557 15392
rect 1515 15343 1557 15352
rect 34539 15392 34581 15401
rect 34539 15352 34540 15392
rect 34580 15352 34581 15392
rect 34539 15343 34581 15352
rect 34923 15392 34965 15401
rect 34923 15352 34924 15392
rect 34964 15352 34965 15392
rect 34923 15343 34965 15352
rect 35499 15392 35541 15401
rect 35499 15352 35500 15392
rect 35540 15352 35541 15392
rect 35499 15343 35541 15352
rect 46923 15392 46965 15401
rect 46923 15352 46924 15392
rect 46964 15352 46965 15392
rect 46923 15343 46965 15352
rect 47883 15392 47925 15401
rect 47883 15352 47884 15392
rect 47924 15352 47925 15392
rect 47883 15343 47925 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 36939 15308 36981 15317
rect 36939 15268 36940 15308
rect 36980 15268 36981 15308
rect 36939 15259 36981 15268
rect 37707 15308 37749 15317
rect 37707 15268 37708 15308
rect 37748 15268 37749 15308
rect 37707 15259 37749 15268
rect 42403 15308 42461 15309
rect 42403 15268 42412 15308
rect 42452 15268 42461 15308
rect 42403 15267 42461 15268
rect 44995 15308 45053 15309
rect 44995 15268 45004 15308
rect 45044 15268 45053 15308
rect 44995 15267 45053 15268
rect 47307 15308 47349 15317
rect 47307 15268 47308 15308
rect 47348 15268 47349 15308
rect 47307 15259 47349 15268
rect 54603 15308 54645 15317
rect 54603 15268 54604 15308
rect 54644 15268 54645 15308
rect 54603 15259 54645 15268
rect 61611 15308 61653 15317
rect 61611 15268 61612 15308
rect 61652 15268 61653 15308
rect 61611 15259 61653 15268
rect 62475 15308 62517 15317
rect 62475 15268 62476 15308
rect 62516 15268 62517 15308
rect 62475 15259 62517 15268
rect 65259 15308 65301 15317
rect 65259 15268 65260 15308
rect 65300 15268 65301 15308
rect 65259 15259 65301 15268
rect 69675 15308 69717 15317
rect 69675 15268 69676 15308
rect 69716 15268 69717 15308
rect 69675 15259 69717 15268
rect 76011 15308 76053 15317
rect 76011 15268 76012 15308
rect 76052 15268 76053 15308
rect 76011 15259 76053 15268
rect 576 15140 79584 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 75112 15140
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75480 15100 79584 15140
rect 576 15076 79584 15100
rect 36835 14972 36893 14973
rect 36835 14932 36844 14972
rect 36884 14932 36893 14972
rect 36835 14931 36893 14932
rect 38379 14972 38421 14981
rect 38379 14932 38380 14972
rect 38420 14932 38421 14972
rect 38379 14923 38421 14932
rect 48259 14972 48317 14973
rect 48259 14932 48268 14972
rect 48308 14932 48317 14972
rect 48259 14931 48317 14932
rect 51139 14972 51197 14973
rect 51139 14932 51148 14972
rect 51188 14932 51197 14972
rect 51139 14931 51197 14932
rect 52299 14972 52341 14981
rect 52299 14932 52300 14972
rect 52340 14932 52341 14972
rect 52299 14923 52341 14932
rect 53451 14972 53493 14981
rect 53451 14932 53452 14972
rect 53492 14932 53493 14972
rect 53451 14923 53493 14932
rect 58251 14972 58293 14981
rect 58251 14932 58252 14972
rect 58292 14932 58293 14972
rect 58251 14923 58293 14932
rect 58923 14972 58965 14981
rect 58923 14932 58924 14972
rect 58964 14932 58965 14972
rect 58923 14923 58965 14932
rect 65251 14972 65309 14973
rect 65251 14932 65260 14972
rect 65300 14932 65309 14972
rect 65251 14931 65309 14932
rect 70923 14972 70965 14981
rect 70923 14932 70924 14972
rect 70964 14932 70965 14972
rect 70923 14923 70965 14932
rect 37227 14888 37269 14897
rect 37227 14848 37228 14888
rect 37268 14848 37269 14888
rect 37227 14839 37269 14848
rect 51915 14888 51957 14897
rect 51915 14848 51916 14888
rect 51956 14848 51957 14888
rect 51915 14839 51957 14848
rect 55083 14888 55125 14897
rect 55083 14848 55084 14888
rect 55124 14848 55125 14888
rect 55083 14839 55125 14848
rect 61035 14888 61077 14897
rect 61035 14848 61036 14888
rect 61076 14848 61077 14888
rect 61035 14839 61077 14848
rect 67179 14888 67221 14897
rect 67179 14848 67180 14888
rect 67220 14848 67221 14888
rect 67179 14839 67221 14848
rect 70059 14888 70101 14897
rect 70059 14848 70060 14888
rect 70100 14848 70101 14888
rect 70059 14839 70101 14848
rect 75435 14888 75477 14897
rect 75435 14848 75436 14888
rect 75476 14848 75477 14888
rect 75435 14839 75477 14848
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 37131 14804 37173 14813
rect 37131 14764 37132 14804
rect 37172 14764 37173 14804
rect 37131 14755 37173 14764
rect 37323 14804 37365 14813
rect 37323 14764 37324 14804
rect 37364 14764 37365 14804
rect 37323 14755 37365 14764
rect 51819 14804 51861 14813
rect 51819 14764 51820 14804
rect 51860 14764 51861 14804
rect 51819 14755 51861 14764
rect 52011 14804 52053 14813
rect 52011 14764 52012 14804
rect 52052 14764 52053 14804
rect 52011 14755 52053 14764
rect 59107 14804 59165 14805
rect 59107 14764 59116 14804
rect 59156 14764 59165 14804
rect 59107 14763 59165 14764
rect 60355 14804 60413 14805
rect 60355 14764 60364 14804
rect 60404 14764 60413 14804
rect 60355 14763 60413 14764
rect 61891 14804 61949 14805
rect 61891 14764 61900 14804
rect 61940 14764 61949 14804
rect 61891 14763 61949 14764
rect 68419 14804 68477 14805
rect 68419 14764 68428 14804
rect 68468 14764 68477 14804
rect 68419 14763 68477 14764
rect 69283 14804 69341 14805
rect 69283 14764 69292 14804
rect 69332 14764 69341 14804
rect 69283 14763 69341 14764
rect 70723 14804 70781 14805
rect 70723 14764 70732 14804
rect 70772 14764 70781 14804
rect 70723 14763 70781 14764
rect 73438 14799 73480 14808
rect 73438 14759 73439 14799
rect 73479 14759 73480 14799
rect 73438 14750 73480 14759
rect 75339 14804 75381 14813
rect 75339 14764 75340 14804
rect 75380 14764 75381 14804
rect 75339 14755 75381 14764
rect 75531 14762 75573 14771
rect 34443 14720 34485 14729
rect 34443 14680 34444 14720
rect 34484 14680 34485 14720
rect 34443 14671 34485 14680
rect 34819 14720 34877 14721
rect 34819 14680 34828 14720
rect 34868 14680 34877 14720
rect 34819 14679 34877 14680
rect 35683 14720 35741 14721
rect 35683 14680 35692 14720
rect 35732 14680 35741 14720
rect 35683 14679 35741 14680
rect 37035 14720 37077 14729
rect 37035 14680 37036 14720
rect 37076 14680 37077 14720
rect 37035 14671 37077 14680
rect 37411 14720 37469 14721
rect 37411 14680 37420 14720
rect 37460 14680 37469 14720
rect 37411 14679 37469 14680
rect 38467 14720 38525 14721
rect 38467 14680 38476 14720
rect 38516 14680 38525 14720
rect 38467 14679 38525 14680
rect 38659 14720 38717 14721
rect 38659 14680 38668 14720
rect 38708 14680 38717 14720
rect 38659 14679 38717 14680
rect 38763 14720 38805 14729
rect 38763 14680 38764 14720
rect 38804 14680 38805 14720
rect 38763 14671 38805 14680
rect 38955 14720 38997 14729
rect 38955 14680 38956 14720
rect 38996 14680 38997 14720
rect 38955 14671 38997 14680
rect 39235 14720 39293 14721
rect 39235 14680 39244 14720
rect 39284 14680 39293 14720
rect 39235 14679 39293 14680
rect 42411 14720 42453 14729
rect 42411 14680 42412 14720
rect 42452 14680 42453 14720
rect 42411 14671 42453 14680
rect 42507 14720 42549 14729
rect 42507 14680 42508 14720
rect 42548 14680 42549 14720
rect 42507 14671 42549 14680
rect 42603 14720 42645 14729
rect 42603 14680 42604 14720
rect 42644 14680 42645 14720
rect 42603 14671 42645 14680
rect 42699 14720 42741 14729
rect 42699 14680 42700 14720
rect 42740 14680 42741 14720
rect 42699 14671 42741 14680
rect 43083 14720 43125 14729
rect 43083 14680 43084 14720
rect 43124 14680 43125 14720
rect 43083 14671 43125 14680
rect 43179 14720 43221 14729
rect 43179 14680 43180 14720
rect 43220 14680 43221 14720
rect 43179 14671 43221 14680
rect 43275 14720 43317 14729
rect 43275 14680 43276 14720
rect 43316 14680 43317 14720
rect 43275 14671 43317 14680
rect 45483 14720 45525 14729
rect 45483 14680 45484 14720
rect 45524 14680 45525 14720
rect 45483 14671 45525 14680
rect 45579 14720 45621 14729
rect 45579 14680 45580 14720
rect 45620 14680 45621 14720
rect 45579 14671 45621 14680
rect 45675 14720 45717 14729
rect 45675 14680 45676 14720
rect 45716 14680 45717 14720
rect 45675 14671 45717 14680
rect 46243 14720 46301 14721
rect 46243 14680 46252 14720
rect 46292 14680 46301 14720
rect 46243 14679 46301 14680
rect 47107 14720 47165 14721
rect 47107 14680 47116 14720
rect 47156 14680 47165 14720
rect 47107 14679 47165 14680
rect 48747 14720 48789 14729
rect 48747 14680 48748 14720
rect 48788 14680 48789 14720
rect 48747 14671 48789 14680
rect 49123 14720 49181 14721
rect 49123 14680 49132 14720
rect 49172 14680 49181 14720
rect 49123 14679 49181 14680
rect 49987 14720 50045 14721
rect 49987 14680 49996 14720
rect 50036 14680 50045 14720
rect 49987 14679 50045 14680
rect 51331 14720 51389 14721
rect 51331 14680 51340 14720
rect 51380 14680 51389 14720
rect 51331 14679 51389 14680
rect 51723 14720 51765 14729
rect 51723 14680 51724 14720
rect 51764 14680 51765 14720
rect 51723 14671 51765 14680
rect 52099 14720 52157 14721
rect 52099 14680 52108 14720
rect 52148 14680 52157 14720
rect 52099 14679 52157 14680
rect 52587 14720 52629 14729
rect 52587 14680 52588 14720
rect 52628 14680 52629 14720
rect 52587 14671 52629 14680
rect 52675 14720 52733 14721
rect 52675 14680 52684 14720
rect 52724 14680 52733 14720
rect 52675 14679 52733 14680
rect 52971 14720 53013 14729
rect 52971 14680 52972 14720
rect 53012 14680 53013 14720
rect 52971 14671 53013 14680
rect 53067 14720 53109 14729
rect 53067 14680 53068 14720
rect 53108 14680 53109 14720
rect 53067 14671 53109 14680
rect 53163 14720 53205 14729
rect 53163 14680 53164 14720
rect 53204 14680 53205 14720
rect 53539 14720 53597 14721
rect 53163 14671 53205 14680
rect 53259 14699 53301 14708
rect 53259 14659 53260 14699
rect 53300 14659 53301 14699
rect 53539 14680 53548 14720
rect 53588 14680 53597 14720
rect 53539 14679 53597 14680
rect 53923 14720 53981 14721
rect 53923 14680 53932 14720
rect 53972 14680 53981 14720
rect 53923 14679 53981 14680
rect 54027 14720 54069 14729
rect 54027 14680 54028 14720
rect 54068 14680 54069 14720
rect 54027 14671 54069 14680
rect 54219 14720 54261 14729
rect 54219 14680 54220 14720
rect 54260 14680 54261 14720
rect 54219 14671 54261 14680
rect 54403 14720 54461 14721
rect 54403 14680 54412 14720
rect 54452 14680 54461 14720
rect 54403 14679 54461 14680
rect 55371 14720 55413 14729
rect 55371 14680 55372 14720
rect 55412 14680 55413 14720
rect 55371 14671 55413 14680
rect 55459 14720 55517 14721
rect 55459 14680 55468 14720
rect 55508 14680 55517 14720
rect 55459 14679 55517 14680
rect 55755 14720 55797 14729
rect 55755 14680 55756 14720
rect 55796 14680 55797 14720
rect 55755 14671 55797 14680
rect 55851 14720 55893 14729
rect 55851 14680 55852 14720
rect 55892 14680 55893 14720
rect 55851 14671 55893 14680
rect 55947 14720 55989 14729
rect 55947 14680 55948 14720
rect 55988 14680 55989 14720
rect 55947 14671 55989 14680
rect 56043 14720 56085 14729
rect 56043 14680 56044 14720
rect 56084 14680 56085 14720
rect 56043 14671 56085 14680
rect 58539 14720 58581 14729
rect 58539 14680 58540 14720
rect 58580 14680 58581 14720
rect 58539 14671 58581 14680
rect 58627 14720 58685 14721
rect 58627 14680 58636 14720
rect 58676 14680 58685 14720
rect 58627 14679 58685 14680
rect 61323 14720 61365 14729
rect 61323 14680 61324 14720
rect 61364 14680 61365 14720
rect 61323 14671 61365 14680
rect 61411 14720 61469 14721
rect 61411 14680 61420 14720
rect 61460 14680 61469 14720
rect 61411 14679 61469 14680
rect 62379 14720 62421 14729
rect 62379 14680 62380 14720
rect 62420 14680 62421 14720
rect 62379 14671 62421 14680
rect 62475 14720 62517 14729
rect 62475 14680 62476 14720
rect 62516 14680 62517 14720
rect 62475 14671 62517 14680
rect 62571 14720 62613 14729
rect 62571 14680 62572 14720
rect 62612 14680 62613 14720
rect 62571 14671 62613 14680
rect 63235 14720 63293 14721
rect 63235 14680 63244 14720
rect 63284 14680 63293 14720
rect 63235 14679 63293 14680
rect 64099 14720 64157 14721
rect 64099 14680 64108 14720
rect 64148 14680 64157 14720
rect 64099 14679 64157 14680
rect 65547 14720 65589 14729
rect 65547 14680 65548 14720
rect 65588 14680 65589 14720
rect 65547 14671 65589 14680
rect 65643 14720 65685 14729
rect 65643 14680 65644 14720
rect 65684 14680 65685 14720
rect 65643 14671 65685 14680
rect 65739 14720 65781 14729
rect 65739 14680 65740 14720
rect 65780 14680 65781 14720
rect 65739 14671 65781 14680
rect 67467 14720 67509 14729
rect 67467 14680 67468 14720
rect 67508 14680 67509 14720
rect 67467 14671 67509 14680
rect 67555 14720 67613 14721
rect 67555 14680 67564 14720
rect 67604 14680 67613 14720
rect 67555 14679 67613 14680
rect 68803 14720 68861 14721
rect 68803 14680 68812 14720
rect 68852 14680 68861 14720
rect 68803 14679 68861 14680
rect 68907 14720 68949 14729
rect 68907 14680 68908 14720
rect 68948 14680 68949 14720
rect 68907 14671 68949 14680
rect 69099 14720 69141 14729
rect 69099 14680 69100 14720
rect 69140 14680 69141 14720
rect 69099 14671 69141 14680
rect 70347 14720 70389 14729
rect 70347 14680 70348 14720
rect 70388 14680 70389 14720
rect 70347 14671 70389 14680
rect 70435 14720 70493 14721
rect 70435 14680 70444 14720
rect 70484 14680 70493 14720
rect 70435 14679 70493 14680
rect 71115 14720 71157 14729
rect 71115 14680 71116 14720
rect 71156 14680 71157 14720
rect 71115 14671 71157 14680
rect 71211 14720 71253 14729
rect 71211 14680 71212 14720
rect 71252 14680 71253 14720
rect 71211 14671 71253 14680
rect 71307 14720 71349 14729
rect 71307 14680 71308 14720
rect 71348 14680 71349 14720
rect 71307 14671 71349 14680
rect 71403 14720 71445 14729
rect 71403 14680 71404 14720
rect 71444 14680 71445 14720
rect 71403 14671 71445 14680
rect 71883 14720 71925 14729
rect 71883 14680 71884 14720
rect 71924 14680 71925 14720
rect 71883 14671 71925 14680
rect 71979 14720 72021 14729
rect 71979 14680 71980 14720
rect 72020 14680 72021 14720
rect 71979 14671 72021 14680
rect 72075 14720 72117 14729
rect 72075 14680 72076 14720
rect 72116 14680 72117 14720
rect 72075 14671 72117 14680
rect 75243 14720 75285 14729
rect 75243 14680 75244 14720
rect 75284 14680 75285 14720
rect 75531 14722 75532 14762
rect 75572 14722 75573 14762
rect 75531 14713 75573 14722
rect 75619 14762 75677 14763
rect 75619 14722 75628 14762
rect 75668 14722 75677 14762
rect 75619 14721 75677 14722
rect 75915 14720 75957 14729
rect 75243 14671 75285 14680
rect 75915 14680 75916 14720
rect 75956 14680 75957 14720
rect 75915 14671 75957 14680
rect 76011 14720 76053 14729
rect 76011 14680 76012 14720
rect 76052 14680 76053 14720
rect 76011 14671 76053 14680
rect 76107 14720 76149 14729
rect 76107 14680 76108 14720
rect 76148 14680 76149 14720
rect 76107 14671 76149 14680
rect 76203 14720 76245 14729
rect 76203 14680 76204 14720
rect 76244 14680 76245 14720
rect 76203 14671 76245 14680
rect 76683 14720 76725 14729
rect 76683 14680 76684 14720
rect 76724 14680 76725 14720
rect 76683 14671 76725 14680
rect 76779 14720 76821 14729
rect 76779 14680 76780 14720
rect 76820 14680 76821 14720
rect 76779 14671 76821 14680
rect 76875 14720 76917 14729
rect 76875 14680 76876 14720
rect 76916 14680 76917 14720
rect 76875 14671 76917 14680
rect 76971 14720 77013 14729
rect 76971 14680 76972 14720
rect 77012 14680 77013 14720
rect 76971 14671 77013 14680
rect 53259 14650 53301 14659
rect 45387 14636 45429 14645
rect 45387 14596 45388 14636
rect 45428 14596 45429 14636
rect 45387 14587 45429 14596
rect 45867 14636 45909 14645
rect 45867 14596 45868 14636
rect 45908 14596 45909 14636
rect 45867 14587 45909 14596
rect 62667 14636 62709 14645
rect 62667 14596 62668 14636
rect 62708 14596 62709 14636
rect 62667 14587 62709 14596
rect 62859 14636 62901 14645
rect 62859 14596 62860 14636
rect 62900 14596 62901 14636
rect 62859 14587 62901 14596
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 38851 14552 38909 14553
rect 38851 14512 38860 14552
rect 38900 14512 38909 14552
rect 38851 14511 38909 14512
rect 41259 14552 41301 14561
rect 41259 14512 41260 14552
rect 41300 14512 41301 14552
rect 41259 14503 41301 14512
rect 42979 14552 43037 14553
rect 42979 14512 42988 14552
rect 43028 14512 43037 14552
rect 42979 14511 43037 14512
rect 48259 14552 48317 14553
rect 48259 14512 48268 14552
rect 48308 14512 48317 14552
rect 48259 14511 48317 14512
rect 52779 14548 52821 14557
rect 52779 14508 52780 14548
rect 52820 14508 52821 14548
rect 54115 14552 54173 14553
rect 54115 14512 54124 14552
rect 54164 14512 54173 14552
rect 54115 14511 54173 14512
rect 54507 14552 54549 14561
rect 54507 14512 54508 14552
rect 54548 14512 54549 14552
rect 52779 14499 52821 14508
rect 54507 14503 54549 14512
rect 58923 14552 58965 14561
rect 58923 14512 58924 14552
rect 58964 14512 58965 14552
rect 58923 14503 58965 14512
rect 60171 14552 60213 14561
rect 60171 14512 60172 14552
rect 60212 14512 60213 14552
rect 60171 14503 60213 14512
rect 62091 14552 62133 14561
rect 62091 14512 62092 14552
rect 62132 14512 62133 14552
rect 62091 14503 62133 14512
rect 65443 14552 65501 14553
rect 65443 14512 65452 14552
rect 65492 14512 65501 14552
rect 65443 14511 65501 14512
rect 68619 14552 68661 14561
rect 68619 14512 68620 14552
rect 68660 14512 68661 14552
rect 68619 14503 68661 14512
rect 68995 14552 69053 14553
rect 68995 14512 69004 14552
rect 69044 14512 69053 14552
rect 68995 14511 69053 14512
rect 69483 14552 69525 14561
rect 69483 14512 69484 14552
rect 69524 14512 69525 14552
rect 69483 14503 69525 14512
rect 70923 14552 70965 14561
rect 70923 14512 70924 14552
rect 70964 14512 70965 14552
rect 70923 14503 70965 14512
rect 71779 14552 71837 14553
rect 71779 14512 71788 14552
rect 71828 14512 71837 14552
rect 71779 14511 71837 14512
rect 73611 14552 73653 14561
rect 73611 14512 73612 14552
rect 73652 14512 73653 14552
rect 73611 14503 73653 14512
rect 55563 14494 55605 14503
rect 55563 14454 55564 14494
rect 55604 14454 55605 14494
rect 55563 14445 55605 14454
rect 58731 14494 58773 14503
rect 58731 14454 58732 14494
rect 58772 14454 58773 14494
rect 58731 14445 58773 14454
rect 61515 14494 61557 14503
rect 61515 14454 61516 14494
rect 61556 14454 61557 14494
rect 61515 14445 61557 14454
rect 67659 14494 67701 14503
rect 67659 14454 67660 14494
rect 67700 14454 67701 14494
rect 67659 14445 67701 14454
rect 70539 14494 70581 14503
rect 70539 14454 70540 14494
rect 70580 14454 70581 14494
rect 70539 14445 70581 14454
rect 576 14384 79584 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 76352 14384
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76720 14344 79584 14384
rect 576 14320 79584 14344
rect 40395 14220 40437 14229
rect 39043 14216 39101 14217
rect 39043 14176 39052 14216
rect 39092 14176 39101 14216
rect 39043 14175 39101 14176
rect 40395 14180 40396 14220
rect 40436 14180 40437 14220
rect 40395 14171 40437 14180
rect 41067 14216 41109 14225
rect 41067 14176 41068 14216
rect 41108 14176 41109 14216
rect 41067 14167 41109 14176
rect 42891 14220 42933 14229
rect 42891 14180 42892 14220
rect 42932 14180 42933 14220
rect 42891 14171 42933 14180
rect 45291 14220 45333 14229
rect 45291 14180 45292 14220
rect 45332 14180 45333 14220
rect 45291 14171 45333 14180
rect 53923 14216 53981 14217
rect 53923 14176 53932 14216
rect 53972 14176 53981 14216
rect 53923 14175 53981 14176
rect 66979 14216 67037 14217
rect 66979 14176 66988 14216
rect 67028 14176 67037 14216
rect 66979 14175 67037 14176
rect 70539 14216 70581 14225
rect 70539 14176 70540 14216
rect 70580 14176 70581 14216
rect 70539 14167 70581 14176
rect 74275 14216 74333 14217
rect 74275 14176 74284 14216
rect 74324 14176 74333 14216
rect 74275 14175 74333 14176
rect 75811 14216 75869 14217
rect 75811 14176 75820 14216
rect 75860 14176 75869 14216
rect 75811 14175 75869 14176
rect 79363 14216 79421 14217
rect 79363 14176 79372 14216
rect 79412 14176 79421 14216
rect 79363 14175 79421 14176
rect 36651 14132 36693 14141
rect 36651 14092 36652 14132
rect 36692 14092 36693 14132
rect 36651 14083 36693 14092
rect 46731 14132 46773 14141
rect 46731 14092 46732 14132
rect 46772 14092 46773 14132
rect 46731 14083 46773 14092
rect 51531 14132 51573 14141
rect 51531 14092 51532 14132
rect 51572 14092 51573 14132
rect 51531 14083 51573 14092
rect 64587 14132 64629 14141
rect 64587 14092 64588 14132
rect 64628 14092 64629 14132
rect 64587 14083 64629 14092
rect 71883 14132 71925 14141
rect 71883 14092 71884 14132
rect 71924 14092 71925 14132
rect 71883 14083 71925 14092
rect 63339 14069 63381 14078
rect 37027 14048 37085 14049
rect 37027 14008 37036 14048
rect 37076 14008 37085 14048
rect 37027 14007 37085 14008
rect 37891 14048 37949 14049
rect 37891 14008 37900 14048
rect 37940 14008 37949 14048
rect 37891 14007 37949 14008
rect 39339 14048 39381 14057
rect 39339 14008 39340 14048
rect 39380 14008 39381 14048
rect 39339 13999 39381 14008
rect 39715 14048 39773 14049
rect 39715 14008 39724 14048
rect 39764 14008 39773 14048
rect 39715 14007 39773 14008
rect 40203 14048 40245 14057
rect 40203 14008 40204 14048
rect 40244 14008 40245 14048
rect 40203 13999 40245 14008
rect 40291 14048 40349 14049
rect 40291 14008 40300 14048
rect 40340 14008 40349 14048
rect 40291 14007 40349 14008
rect 40587 14048 40629 14057
rect 40587 14008 40588 14048
rect 40628 14008 40629 14048
rect 40587 13999 40629 14008
rect 40683 14048 40725 14057
rect 40683 14008 40684 14048
rect 40724 14008 40725 14048
rect 40683 13999 40725 14008
rect 40779 14048 40821 14057
rect 40779 14008 40780 14048
rect 40820 14008 40821 14048
rect 40779 13999 40821 14008
rect 40875 14048 40917 14057
rect 40875 14008 40876 14048
rect 40916 14008 40917 14048
rect 40875 13999 40917 14008
rect 41155 14048 41213 14049
rect 41155 14008 41164 14048
rect 41204 14008 41213 14048
rect 41155 14007 41213 14008
rect 41643 14048 41685 14057
rect 41643 14008 41644 14048
rect 41684 14008 41685 14048
rect 41643 13999 41685 14008
rect 42019 14048 42077 14049
rect 42019 14008 42028 14048
rect 42068 14008 42077 14048
rect 42787 14048 42845 14049
rect 42019 14007 42077 14008
rect 42699 14031 42741 14040
rect 42699 13991 42700 14031
rect 42740 13991 42741 14031
rect 42787 14008 42796 14048
rect 42836 14008 42845 14048
rect 42787 14007 42845 14008
rect 45099 14048 45141 14057
rect 45099 14008 45100 14048
rect 45140 14008 45141 14048
rect 45099 13999 45141 14008
rect 45187 14048 45245 14049
rect 45187 14008 45196 14048
rect 45236 14008 45245 14048
rect 45187 14007 45245 14008
rect 45571 14048 45629 14049
rect 45571 14008 45580 14048
rect 45620 14008 45629 14048
rect 45571 14007 45629 14008
rect 46531 14048 46589 14049
rect 46531 14008 46540 14048
rect 46580 14008 46589 14048
rect 46531 14007 46589 14008
rect 46827 14048 46869 14057
rect 46827 14008 46828 14048
rect 46868 14008 46869 14048
rect 46827 13999 46869 14008
rect 46923 14048 46965 14057
rect 46923 14008 46924 14048
rect 46964 14008 46965 14048
rect 46923 13999 46965 14008
rect 47019 14048 47061 14057
rect 47019 14008 47020 14048
rect 47060 14008 47061 14048
rect 47019 13999 47061 14008
rect 48075 14048 48117 14057
rect 48075 14008 48076 14048
rect 48116 14008 48117 14048
rect 48075 13999 48117 14008
rect 48451 14048 48509 14049
rect 48451 14008 48460 14048
rect 48500 14008 48509 14048
rect 48451 14007 48509 14008
rect 48651 14048 48693 14057
rect 48651 14008 48652 14048
rect 48692 14008 48693 14048
rect 48651 13999 48693 14008
rect 49027 14048 49085 14049
rect 49027 14008 49036 14048
rect 49076 14008 49085 14048
rect 49027 14007 49085 14008
rect 49891 14048 49949 14049
rect 49891 14008 49900 14048
rect 49940 14008 49949 14048
rect 49891 14007 49949 14008
rect 51907 14048 51965 14049
rect 51907 14008 51916 14048
rect 51956 14008 51965 14048
rect 51907 14007 51965 14008
rect 52771 14048 52829 14049
rect 52771 14008 52780 14048
rect 52820 14008 52829 14048
rect 52771 14007 52829 14008
rect 54123 14048 54165 14057
rect 54123 14008 54124 14048
rect 54164 14008 54165 14048
rect 54123 13999 54165 14008
rect 54499 14048 54557 14049
rect 54499 14008 54508 14048
rect 54548 14008 54557 14048
rect 54499 14007 54557 14008
rect 55363 14048 55421 14049
rect 55363 14008 55372 14048
rect 55412 14008 55421 14048
rect 55363 14007 55421 14008
rect 58051 14048 58109 14049
rect 58051 14008 58060 14048
rect 58100 14008 58109 14048
rect 58051 14007 58109 14008
rect 58443 14048 58485 14057
rect 58443 14008 58444 14048
rect 58484 14008 58485 14048
rect 58443 13999 58485 14008
rect 59299 14048 59357 14049
rect 59299 14008 59308 14048
rect 59348 14008 59357 14048
rect 59299 14007 59357 14008
rect 59491 14048 59549 14049
rect 59491 14008 59500 14048
rect 59540 14008 59549 14048
rect 59491 14007 59549 14008
rect 59595 14048 59637 14057
rect 59595 14008 59596 14048
rect 59636 14008 59637 14048
rect 59595 13999 59637 14008
rect 59787 14048 59829 14057
rect 59787 14008 59788 14048
rect 59828 14008 59829 14048
rect 59787 13999 59829 14008
rect 59979 14048 60021 14057
rect 59979 14008 59980 14048
rect 60020 14008 60021 14048
rect 59979 13999 60021 14008
rect 60355 14048 60413 14049
rect 60355 14008 60364 14048
rect 60404 14008 60413 14048
rect 60355 14007 60413 14008
rect 61219 14048 61277 14049
rect 61219 14008 61228 14048
rect 61268 14008 61277 14048
rect 61219 14007 61277 14008
rect 62563 14048 62621 14049
rect 62563 14008 62572 14048
rect 62612 14008 62621 14048
rect 62563 14007 62621 14008
rect 63147 14048 63189 14057
rect 63147 14008 63148 14048
rect 63188 14008 63189 14048
rect 63147 13999 63189 14008
rect 63243 14048 63285 14057
rect 63243 14008 63244 14048
rect 63284 14008 63285 14048
rect 63339 14029 63340 14069
rect 63380 14029 63381 14069
rect 63339 14020 63381 14029
rect 63435 14048 63477 14057
rect 63243 13999 63285 14008
rect 63435 14008 63436 14048
rect 63476 14008 63477 14048
rect 63435 13999 63477 14008
rect 64963 14048 65021 14049
rect 64963 14008 64972 14048
rect 65012 14008 65021 14048
rect 64963 14007 65021 14008
rect 65827 14048 65885 14049
rect 65827 14008 65836 14048
rect 65876 14008 65885 14048
rect 65827 14007 65885 14008
rect 67179 14048 67221 14057
rect 67179 14008 67180 14048
rect 67220 14008 67221 14048
rect 67179 13999 67221 14008
rect 67555 14048 67613 14049
rect 67555 14008 67564 14048
rect 67604 14008 67613 14048
rect 67555 14007 67613 14008
rect 68419 14048 68477 14049
rect 68419 14008 68428 14048
rect 68468 14008 68477 14048
rect 68419 14007 68477 14008
rect 69771 14048 69813 14057
rect 69771 14008 69772 14048
rect 69812 14008 69813 14048
rect 69771 13999 69813 14008
rect 70147 14048 70205 14049
rect 70147 14008 70156 14048
rect 70196 14008 70205 14048
rect 70147 14007 70205 14008
rect 70627 14048 70685 14049
rect 70627 14008 70636 14048
rect 70676 14008 70685 14048
rect 70627 14007 70685 14008
rect 70923 14048 70965 14057
rect 70923 14008 70924 14048
rect 70964 14008 70965 14048
rect 70923 13999 70965 14008
rect 71299 14048 71357 14049
rect 71299 14008 71308 14048
rect 71348 14008 71357 14048
rect 71299 14007 71357 14008
rect 72259 14048 72317 14049
rect 72259 14008 72268 14048
rect 72308 14008 72317 14048
rect 72259 14007 72317 14008
rect 73123 14048 73181 14049
rect 73123 14008 73132 14048
rect 73172 14008 73181 14048
rect 73123 14007 73181 14008
rect 75723 14048 75765 14057
rect 75723 14008 75724 14048
rect 75764 14008 75765 14048
rect 75723 13999 75765 14008
rect 75915 14048 75957 14057
rect 75915 14008 75916 14048
rect 75956 14008 75957 14048
rect 75915 13999 75957 14008
rect 76003 14048 76061 14049
rect 76003 14008 76012 14048
rect 76052 14008 76061 14048
rect 76003 14007 76061 14008
rect 76195 14048 76253 14049
rect 76195 14008 76204 14048
rect 76244 14008 76253 14048
rect 76195 14007 76253 14008
rect 76491 14048 76533 14057
rect 76491 14008 76492 14048
rect 76532 14008 76533 14048
rect 76491 13999 76533 14008
rect 76587 14048 76629 14057
rect 76587 14008 76588 14048
rect 76628 14008 76629 14048
rect 76587 13999 76629 14008
rect 76683 14048 76725 14057
rect 76683 14008 76684 14048
rect 76724 14008 76725 14048
rect 76683 13999 76725 14008
rect 76779 14048 76821 14057
rect 76779 14008 76780 14048
rect 76820 14008 76821 14048
rect 76779 13999 76821 14008
rect 76971 14048 77013 14057
rect 76971 14008 76972 14048
rect 77012 14008 77013 14048
rect 76971 13999 77013 14008
rect 77347 14048 77405 14049
rect 77347 14008 77356 14048
rect 77396 14008 77405 14048
rect 77347 14007 77405 14008
rect 78211 14048 78269 14049
rect 78211 14008 78220 14048
rect 78260 14008 78269 14048
rect 78211 14007 78269 14008
rect 42699 13982 42741 13991
rect 1699 13964 1757 13965
rect 1699 13924 1708 13964
rect 1748 13924 1757 13964
rect 1699 13923 1757 13924
rect 39435 13964 39477 13973
rect 39435 13924 39436 13964
rect 39476 13924 39477 13964
rect 39435 13915 39477 13924
rect 39627 13964 39669 13973
rect 39627 13924 39628 13964
rect 39668 13924 39669 13964
rect 39627 13915 39669 13924
rect 41739 13964 41781 13973
rect 41739 13924 41740 13964
rect 41780 13924 41781 13964
rect 41739 13915 41781 13924
rect 41931 13964 41973 13973
rect 41931 13924 41932 13964
rect 41972 13924 41973 13964
rect 41931 13915 41973 13924
rect 48171 13964 48213 13973
rect 48171 13924 48172 13964
rect 48212 13924 48213 13964
rect 48171 13915 48213 13924
rect 48363 13964 48405 13973
rect 48363 13924 48364 13964
rect 48404 13924 48405 13964
rect 48363 13915 48405 13924
rect 58155 13964 58197 13973
rect 58155 13924 58156 13964
rect 58196 13924 58197 13964
rect 58155 13915 58197 13924
rect 58347 13964 58389 13973
rect 58347 13924 58348 13964
rect 58388 13924 58389 13964
rect 58347 13915 58389 13924
rect 69867 13964 69909 13973
rect 69867 13924 69868 13964
rect 69908 13924 69909 13964
rect 69867 13915 69909 13924
rect 70059 13964 70101 13973
rect 70059 13924 70060 13964
rect 70100 13924 70101 13964
rect 70059 13915 70101 13924
rect 71019 13964 71061 13973
rect 71019 13924 71020 13964
rect 71060 13924 71061 13964
rect 71019 13915 71061 13924
rect 71211 13964 71253 13973
rect 71211 13924 71212 13964
rect 71252 13924 71253 13964
rect 71211 13915 71253 13924
rect 39531 13880 39573 13889
rect 39531 13840 39532 13880
rect 39572 13840 39573 13880
rect 39531 13831 39573 13840
rect 39915 13880 39957 13889
rect 39915 13840 39916 13880
rect 39956 13840 39957 13880
rect 39915 13831 39957 13840
rect 41835 13880 41877 13889
rect 41835 13840 41836 13880
rect 41876 13840 41877 13880
rect 41835 13831 41877 13840
rect 42411 13880 42453 13889
rect 42411 13840 42412 13880
rect 42452 13840 42453 13880
rect 42411 13831 42453 13840
rect 44811 13880 44853 13889
rect 44811 13840 44812 13880
rect 44852 13840 44853 13880
rect 44811 13831 44853 13840
rect 48267 13880 48309 13889
rect 48267 13840 48268 13880
rect 48308 13840 48309 13880
rect 48267 13831 48309 13840
rect 58251 13880 58293 13889
rect 58251 13840 58252 13880
rect 58292 13840 58293 13880
rect 58251 13831 58293 13840
rect 59211 13880 59253 13889
rect 59211 13840 59212 13880
rect 59252 13840 59253 13880
rect 59211 13831 59253 13840
rect 62667 13880 62709 13889
rect 62667 13840 62668 13880
rect 62708 13840 62709 13880
rect 62667 13831 62709 13840
rect 69963 13880 70005 13889
rect 69963 13840 69964 13880
rect 70004 13840 70005 13880
rect 69963 13831 70005 13840
rect 71115 13880 71157 13889
rect 71115 13840 71116 13880
rect 71156 13840 71157 13880
rect 71115 13831 71157 13840
rect 1515 13796 1557 13805
rect 1515 13756 1516 13796
rect 1556 13756 1557 13796
rect 1515 13747 1557 13756
rect 45867 13796 45909 13805
rect 45867 13756 45868 13796
rect 45908 13756 45909 13796
rect 45867 13747 45909 13756
rect 51043 13796 51101 13797
rect 51043 13756 51052 13796
rect 51092 13756 51101 13796
rect 51043 13755 51101 13756
rect 56515 13796 56573 13797
rect 56515 13756 56524 13796
rect 56564 13756 56573 13796
rect 56515 13755 56573 13756
rect 59787 13796 59829 13805
rect 59787 13756 59788 13796
rect 59828 13756 59829 13796
rect 59787 13747 59829 13756
rect 62371 13796 62429 13797
rect 62371 13756 62380 13796
rect 62420 13756 62429 13796
rect 62371 13755 62429 13756
rect 69571 13796 69629 13797
rect 69571 13756 69580 13796
rect 69620 13756 69629 13796
rect 69571 13755 69629 13756
rect 76299 13796 76341 13805
rect 76299 13756 76300 13796
rect 76340 13756 76341 13796
rect 76299 13747 76341 13756
rect 576 13628 79584 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 75112 13628
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75480 13588 79584 13628
rect 576 13564 79584 13588
rect 41155 13460 41213 13461
rect 41155 13420 41164 13460
rect 41204 13420 41213 13460
rect 41155 13419 41213 13420
rect 49323 13460 49365 13469
rect 49323 13420 49324 13460
rect 49364 13420 49365 13460
rect 49323 13411 49365 13420
rect 51435 13460 51477 13469
rect 51435 13420 51436 13460
rect 51476 13420 51477 13460
rect 51435 13411 51477 13420
rect 52011 13460 52053 13469
rect 52011 13420 52012 13460
rect 52052 13420 52053 13460
rect 52011 13411 52053 13420
rect 55179 13460 55221 13469
rect 55179 13420 55180 13460
rect 55220 13420 55221 13460
rect 55179 13411 55221 13420
rect 59107 13460 59165 13461
rect 59107 13420 59116 13460
rect 59156 13420 59165 13460
rect 59107 13419 59165 13420
rect 60171 13460 60213 13469
rect 60171 13420 60172 13460
rect 60212 13420 60213 13460
rect 60171 13411 60213 13420
rect 62571 13460 62613 13469
rect 62571 13420 62572 13460
rect 62612 13420 62613 13460
rect 62571 13411 62613 13420
rect 65259 13460 65301 13469
rect 65259 13420 65260 13460
rect 65300 13420 65301 13460
rect 65259 13411 65301 13420
rect 71011 13460 71069 13461
rect 71011 13420 71020 13460
rect 71060 13420 71069 13460
rect 71011 13419 71069 13420
rect 71499 13460 71541 13469
rect 71499 13420 71500 13460
rect 71540 13420 71541 13460
rect 71499 13411 71541 13420
rect 71691 13460 71733 13469
rect 71691 13420 71692 13460
rect 71732 13420 71733 13460
rect 71691 13411 71733 13420
rect 73995 13460 74037 13469
rect 73995 13420 73996 13460
rect 74036 13420 74037 13460
rect 73995 13411 74037 13420
rect 76579 13460 76637 13461
rect 76579 13420 76588 13460
rect 76628 13420 76637 13460
rect 76579 13419 76637 13420
rect 76779 13460 76821 13469
rect 76779 13420 76780 13460
rect 76820 13420 76821 13460
rect 76779 13411 76821 13420
rect 78219 13460 78261 13469
rect 78219 13420 78220 13460
rect 78260 13420 78261 13460
rect 78219 13411 78261 13420
rect 50283 13376 50325 13385
rect 50283 13336 50284 13376
rect 50324 13336 50325 13376
rect 50283 13327 50325 13336
rect 54507 13376 54549 13385
rect 54507 13336 54508 13376
rect 54548 13336 54549 13376
rect 54507 13327 54549 13336
rect 60555 13376 60597 13385
rect 60555 13336 60556 13376
rect 60596 13336 60597 13376
rect 60555 13327 60597 13336
rect 62187 13376 62229 13385
rect 62187 13336 62188 13376
rect 62228 13336 62229 13376
rect 62187 13327 62229 13336
rect 66891 13376 66933 13385
rect 66891 13336 66892 13376
rect 66932 13336 66933 13376
rect 66891 13327 66933 13336
rect 67275 13376 67317 13385
rect 67275 13336 67276 13376
rect 67316 13336 67317 13376
rect 67275 13327 67317 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1699 13292 1757 13293
rect 1699 13252 1708 13292
rect 1748 13252 1757 13292
rect 1699 13251 1757 13252
rect 47787 13292 47829 13301
rect 47787 13252 47788 13292
rect 47828 13252 47829 13292
rect 47787 13243 47829 13252
rect 54411 13292 54453 13301
rect 54411 13252 54412 13292
rect 54452 13252 54453 13292
rect 54411 13243 54453 13252
rect 54603 13292 54645 13301
rect 54603 13252 54604 13292
rect 54644 13252 54645 13292
rect 54603 13243 54645 13252
rect 59971 13292 60029 13293
rect 59971 13252 59980 13292
rect 60020 13252 60029 13292
rect 59971 13251 60029 13252
rect 60459 13292 60501 13301
rect 60459 13252 60460 13292
rect 60500 13252 60501 13292
rect 60459 13243 60501 13252
rect 60651 13292 60693 13301
rect 60651 13252 60652 13292
rect 60692 13252 60693 13292
rect 60651 13243 60693 13252
rect 62091 13292 62133 13301
rect 62091 13252 62092 13292
rect 62132 13252 62133 13292
rect 62091 13243 62133 13252
rect 62283 13292 62325 13301
rect 62283 13252 62284 13292
rect 62324 13252 62325 13292
rect 62283 13243 62325 13252
rect 66795 13292 66837 13301
rect 66795 13252 66796 13292
rect 66836 13252 66837 13292
rect 66795 13243 66837 13252
rect 66987 13292 67029 13301
rect 66987 13252 66988 13292
rect 67028 13252 67029 13292
rect 66987 13243 67029 13252
rect 66499 13221 66557 13222
rect 38763 13208 38805 13217
rect 38763 13168 38764 13208
rect 38804 13168 38805 13208
rect 38763 13159 38805 13168
rect 39139 13208 39197 13209
rect 39139 13168 39148 13208
rect 39188 13168 39197 13208
rect 39139 13167 39197 13168
rect 40003 13208 40061 13209
rect 40003 13168 40012 13208
rect 40052 13168 40061 13208
rect 40003 13167 40061 13168
rect 41355 13208 41397 13217
rect 41355 13168 41356 13208
rect 41396 13168 41397 13208
rect 41355 13159 41397 13168
rect 41731 13208 41789 13209
rect 41731 13168 41740 13208
rect 41780 13168 41789 13208
rect 41731 13167 41789 13168
rect 42595 13208 42653 13209
rect 42595 13168 42604 13208
rect 42644 13168 42653 13208
rect 42595 13167 42653 13168
rect 44419 13208 44477 13209
rect 44419 13168 44428 13208
rect 44468 13168 44477 13208
rect 44419 13167 44477 13168
rect 45283 13208 45341 13209
rect 45283 13168 45292 13208
rect 45332 13168 45341 13208
rect 45283 13167 45341 13168
rect 46731 13208 46773 13217
rect 46731 13168 46732 13208
rect 46772 13168 46773 13208
rect 46731 13159 46773 13168
rect 46827 13208 46869 13217
rect 46827 13168 46828 13208
rect 46868 13168 46869 13208
rect 46827 13159 46869 13168
rect 46923 13208 46965 13217
rect 46923 13168 46924 13208
rect 46964 13168 46965 13208
rect 46923 13159 46965 13168
rect 47683 13208 47741 13209
rect 47683 13168 47692 13208
rect 47732 13168 47741 13208
rect 47683 13167 47741 13168
rect 49611 13208 49653 13217
rect 49611 13168 49612 13208
rect 49652 13168 49653 13208
rect 49611 13159 49653 13168
rect 49699 13208 49757 13209
rect 49699 13168 49708 13208
rect 49748 13168 49757 13208
rect 49699 13167 49757 13168
rect 50371 13208 50429 13209
rect 50371 13168 50380 13208
rect 50420 13168 50429 13208
rect 50371 13167 50429 13168
rect 51139 13208 51197 13209
rect 51139 13168 51148 13208
rect 51188 13168 51197 13208
rect 51139 13167 51197 13168
rect 51243 13208 51285 13217
rect 51243 13168 51244 13208
rect 51284 13168 51285 13208
rect 51243 13159 51285 13168
rect 51435 13208 51477 13217
rect 51435 13168 51436 13208
rect 51476 13168 51477 13208
rect 51435 13159 51477 13168
rect 51715 13208 51773 13209
rect 51715 13168 51724 13208
rect 51764 13168 51773 13208
rect 51715 13167 51773 13168
rect 52675 13208 52733 13209
rect 52675 13168 52684 13208
rect 52724 13168 52733 13208
rect 52675 13167 52733 13168
rect 54315 13208 54357 13217
rect 54315 13168 54316 13208
rect 54356 13168 54357 13208
rect 54315 13159 54357 13168
rect 54691 13208 54749 13209
rect 54691 13168 54700 13208
rect 54740 13168 54749 13208
rect 54691 13167 54749 13168
rect 55267 13208 55325 13209
rect 55267 13168 55276 13208
rect 55316 13168 55325 13208
rect 55267 13167 55325 13168
rect 55467 13208 55509 13217
rect 55467 13168 55468 13208
rect 55508 13168 55509 13208
rect 55467 13159 55509 13168
rect 55659 13208 55701 13217
rect 55659 13168 55660 13208
rect 55700 13168 55701 13208
rect 55659 13159 55701 13168
rect 55747 13208 55805 13209
rect 55747 13168 55756 13208
rect 55796 13168 55805 13208
rect 55747 13167 55805 13168
rect 56235 13208 56277 13217
rect 56235 13168 56236 13208
rect 56276 13168 56277 13208
rect 56235 13159 56277 13168
rect 56331 13208 56373 13217
rect 56331 13168 56332 13208
rect 56372 13168 56373 13208
rect 56331 13159 56373 13168
rect 56427 13208 56469 13217
rect 56427 13168 56428 13208
rect 56468 13168 56469 13208
rect 56427 13159 56469 13168
rect 56523 13208 56565 13217
rect 56523 13168 56524 13208
rect 56564 13168 56565 13208
rect 56523 13159 56565 13168
rect 56715 13208 56757 13217
rect 56715 13168 56716 13208
rect 56756 13168 56757 13208
rect 56715 13159 56757 13168
rect 57091 13208 57149 13209
rect 57091 13168 57100 13208
rect 57140 13168 57149 13208
rect 57091 13167 57149 13168
rect 57955 13208 58013 13209
rect 57955 13168 57964 13208
rect 58004 13168 58013 13208
rect 57955 13167 58013 13168
rect 60363 13208 60405 13217
rect 60363 13168 60364 13208
rect 60404 13168 60405 13208
rect 60363 13159 60405 13168
rect 60739 13208 60797 13209
rect 60739 13168 60748 13208
rect 60788 13168 60797 13208
rect 60739 13167 60797 13168
rect 61515 13208 61557 13217
rect 61515 13168 61516 13208
rect 61556 13168 61557 13208
rect 61515 13159 61557 13168
rect 61707 13208 61749 13217
rect 61707 13168 61708 13208
rect 61748 13168 61749 13208
rect 61707 13159 61749 13168
rect 61795 13208 61853 13209
rect 61795 13168 61804 13208
rect 61844 13168 61853 13208
rect 61795 13167 61853 13168
rect 61995 13208 62037 13217
rect 61995 13168 61996 13208
rect 62036 13168 62037 13208
rect 61995 13159 62037 13168
rect 62371 13208 62429 13209
rect 62371 13168 62380 13208
rect 62420 13168 62429 13208
rect 62371 13167 62429 13168
rect 62859 13208 62901 13217
rect 62859 13168 62860 13208
rect 62900 13168 62901 13208
rect 62859 13159 62901 13168
rect 62947 13208 63005 13209
rect 62947 13168 62956 13208
rect 62996 13168 63005 13208
rect 62947 13167 63005 13168
rect 65547 13208 65589 13217
rect 65547 13168 65548 13208
rect 65588 13168 65589 13208
rect 65547 13159 65589 13168
rect 65635 13208 65693 13209
rect 65635 13168 65644 13208
rect 65684 13168 65693 13208
rect 65635 13167 65693 13168
rect 66027 13208 66069 13217
rect 66027 13168 66028 13208
rect 66068 13168 66069 13208
rect 66027 13159 66069 13168
rect 66123 13208 66165 13217
rect 66123 13168 66124 13208
rect 66164 13168 66165 13208
rect 66123 13159 66165 13168
rect 66219 13208 66261 13217
rect 66219 13168 66220 13208
rect 66260 13168 66261 13208
rect 66499 13181 66508 13221
rect 66548 13181 66557 13221
rect 66499 13180 66557 13181
rect 66699 13208 66741 13217
rect 66219 13159 66261 13168
rect 66699 13168 66700 13208
rect 66740 13168 66741 13208
rect 66699 13159 66741 13168
rect 67075 13208 67133 13209
rect 67075 13168 67084 13208
rect 67124 13168 67133 13208
rect 67075 13167 67133 13168
rect 67275 13208 67317 13217
rect 67275 13168 67276 13208
rect 67316 13168 67317 13208
rect 67275 13159 67317 13168
rect 67467 13208 67509 13217
rect 67467 13168 67468 13208
rect 67508 13168 67509 13208
rect 67467 13159 67509 13168
rect 67555 13208 67613 13209
rect 67555 13168 67564 13208
rect 67604 13168 67613 13208
rect 67555 13167 67613 13168
rect 68139 13208 68181 13217
rect 68139 13168 68140 13208
rect 68180 13168 68181 13208
rect 68139 13159 68181 13168
rect 68227 13208 68285 13209
rect 68227 13168 68236 13208
rect 68276 13168 68285 13208
rect 68227 13167 68285 13168
rect 68619 13208 68661 13217
rect 68619 13168 68620 13208
rect 68660 13168 68661 13208
rect 68619 13159 68661 13168
rect 68995 13208 69053 13209
rect 68995 13168 69004 13208
rect 69044 13168 69053 13208
rect 68995 13167 69053 13168
rect 69859 13208 69917 13209
rect 69859 13168 69868 13208
rect 69908 13168 69917 13208
rect 69859 13167 69917 13168
rect 71203 13208 71261 13209
rect 71203 13168 71212 13208
rect 71252 13168 71261 13208
rect 71203 13167 71261 13168
rect 71307 13208 71349 13217
rect 71307 13168 71308 13208
rect 71348 13168 71349 13208
rect 71307 13159 71349 13168
rect 71499 13208 71541 13217
rect 71499 13168 71500 13208
rect 71540 13168 71541 13208
rect 71499 13159 71541 13168
rect 71979 13208 72021 13217
rect 71979 13168 71980 13208
rect 72020 13168 72021 13208
rect 71979 13159 72021 13168
rect 72067 13208 72125 13209
rect 72067 13168 72076 13208
rect 72116 13168 72125 13208
rect 72067 13167 72125 13168
rect 72651 13208 72693 13217
rect 72651 13168 72652 13208
rect 72692 13168 72693 13208
rect 72651 13159 72693 13168
rect 72747 13208 72789 13217
rect 72747 13168 72748 13208
rect 72788 13168 72789 13208
rect 72747 13159 72789 13168
rect 72843 13208 72885 13217
rect 72843 13168 72844 13208
rect 72884 13168 72885 13208
rect 72843 13159 72885 13168
rect 72939 13208 72981 13217
rect 72939 13168 72940 13208
rect 72980 13168 72981 13208
rect 72939 13159 72981 13168
rect 73891 13208 73949 13209
rect 73891 13168 73900 13208
rect 73940 13168 73949 13208
rect 73891 13167 73949 13168
rect 74187 13208 74229 13217
rect 74187 13168 74188 13208
rect 74228 13168 74229 13208
rect 74187 13159 74229 13168
rect 74563 13208 74621 13209
rect 74563 13168 74572 13208
rect 74612 13168 74621 13208
rect 74563 13167 74621 13168
rect 75427 13208 75485 13209
rect 75427 13168 75436 13208
rect 75476 13168 75485 13208
rect 75427 13167 75485 13168
rect 77067 13208 77109 13217
rect 77067 13168 77068 13208
rect 77108 13168 77109 13208
rect 77067 13159 77109 13168
rect 77155 13208 77213 13209
rect 77155 13168 77164 13208
rect 77204 13168 77213 13208
rect 77155 13167 77213 13168
rect 77547 13208 77589 13217
rect 77547 13168 77548 13208
rect 77588 13168 77589 13208
rect 77547 13159 77589 13168
rect 77643 13208 77685 13217
rect 77643 13168 77644 13208
rect 77684 13168 77685 13208
rect 77643 13159 77685 13168
rect 77739 13208 77781 13217
rect 77739 13168 77740 13208
rect 77780 13168 77781 13208
rect 77739 13159 77781 13168
rect 77835 13208 77877 13217
rect 77835 13168 77836 13208
rect 77876 13168 77877 13208
rect 77835 13159 77877 13168
rect 78307 13208 78365 13209
rect 78307 13168 78316 13208
rect 78356 13168 78365 13208
rect 78307 13167 78365 13168
rect 44043 13124 44085 13133
rect 44043 13084 44044 13124
rect 44084 13084 44085 13124
rect 44043 13075 44085 13084
rect 61611 13124 61653 13133
rect 61611 13084 61612 13124
rect 61652 13084 61653 13124
rect 61611 13075 61653 13084
rect 66411 13124 66453 13133
rect 66411 13084 66412 13124
rect 66452 13084 66453 13124
rect 66411 13075 66453 13084
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 1515 13040 1557 13049
rect 1515 13000 1516 13040
rect 1556 13000 1557 13040
rect 1515 12991 1557 13000
rect 41155 13040 41213 13041
rect 41155 13000 41164 13040
rect 41204 13000 41213 13040
rect 41155 12999 41213 13000
rect 43747 13040 43805 13041
rect 43747 13000 43756 13040
rect 43796 13000 43805 13040
rect 43747 12999 43805 13000
rect 46435 13040 46493 13041
rect 46435 13000 46444 13040
rect 46484 13000 46493 13040
rect 46435 12999 46493 13000
rect 46627 13040 46685 13041
rect 46627 13000 46636 13040
rect 46676 13000 46685 13040
rect 46627 12999 46685 13000
rect 49803 13036 49845 13045
rect 49803 12996 49804 13036
rect 49844 12996 49845 13036
rect 55555 13040 55613 13041
rect 55555 13000 55564 13040
rect 55604 13000 55613 13040
rect 55555 12999 55613 13000
rect 65739 13036 65781 13045
rect 49803 12987 49845 12996
rect 65739 12996 65740 13036
rect 65780 12996 65781 13036
rect 65923 13040 65981 13041
rect 65923 13000 65932 13040
rect 65972 13000 65981 13040
rect 65923 12999 65981 13000
rect 72171 13036 72213 13045
rect 63051 12982 63093 12991
rect 65739 12987 65781 12996
rect 72171 12996 72172 13036
rect 72212 12996 72213 13036
rect 72171 12987 72213 12996
rect 63051 12942 63052 12982
rect 63092 12942 63093 12982
rect 63051 12933 63093 12942
rect 77259 12982 77301 12991
rect 77259 12942 77260 12982
rect 77300 12942 77301 12982
rect 77259 12933 77301 12942
rect 576 12872 79584 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 76352 12872
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76720 12832 79584 12872
rect 576 12808 79584 12832
rect 43179 12704 43221 12713
rect 43179 12664 43180 12704
rect 43220 12664 43221 12704
rect 43179 12655 43221 12664
rect 45579 12704 45621 12713
rect 56235 12708 56277 12717
rect 45579 12664 45580 12704
rect 45620 12664 45621 12704
rect 45579 12655 45621 12664
rect 49219 12704 49277 12705
rect 49219 12664 49228 12704
rect 49268 12664 49277 12704
rect 49219 12663 49277 12664
rect 49795 12704 49853 12705
rect 49795 12664 49804 12704
rect 49844 12664 49853 12704
rect 49795 12663 49853 12664
rect 50851 12704 50909 12705
rect 50851 12664 50860 12704
rect 50900 12664 50909 12704
rect 50851 12663 50909 12664
rect 53731 12704 53789 12705
rect 53731 12664 53740 12704
rect 53780 12664 53789 12704
rect 53731 12663 53789 12664
rect 56235 12668 56236 12708
rect 56276 12668 56277 12708
rect 56235 12659 56277 12668
rect 60067 12704 60125 12705
rect 60067 12664 60076 12704
rect 60116 12664 60125 12704
rect 60067 12663 60125 12664
rect 62955 12704 62997 12713
rect 62955 12664 62956 12704
rect 62996 12664 62997 12704
rect 62955 12655 62997 12664
rect 63723 12704 63765 12713
rect 63723 12664 63724 12704
rect 63764 12664 63765 12704
rect 63723 12655 63765 12664
rect 66787 12704 66845 12705
rect 66787 12664 66796 12704
rect 66836 12664 66845 12704
rect 66787 12663 66845 12664
rect 72171 12704 72213 12713
rect 72171 12664 72172 12704
rect 72212 12664 72213 12704
rect 72171 12655 72213 12664
rect 75043 12704 75101 12705
rect 75043 12664 75052 12704
rect 75092 12664 75101 12704
rect 75043 12663 75101 12664
rect 46827 12620 46869 12629
rect 44043 12578 44085 12587
rect 41251 12536 41309 12537
rect 41251 12496 41260 12536
rect 41300 12496 41309 12536
rect 41251 12495 41309 12496
rect 41355 12536 41397 12545
rect 41355 12496 41356 12536
rect 41396 12496 41397 12536
rect 41355 12487 41397 12496
rect 41547 12536 41589 12545
rect 41547 12496 41548 12536
rect 41588 12496 41589 12536
rect 41547 12487 41589 12496
rect 43267 12536 43325 12537
rect 43267 12496 43276 12536
rect 43316 12496 43325 12536
rect 43267 12495 43325 12496
rect 43555 12536 43613 12537
rect 43555 12496 43564 12536
rect 43604 12496 43613 12536
rect 43555 12495 43613 12496
rect 43747 12536 43805 12537
rect 43747 12496 43756 12536
rect 43796 12496 43805 12536
rect 43747 12495 43805 12496
rect 43851 12536 43893 12545
rect 43851 12496 43852 12536
rect 43892 12496 43893 12536
rect 44043 12538 44044 12578
rect 44084 12538 44085 12578
rect 46827 12580 46828 12620
rect 46868 12580 46869 12620
rect 46827 12571 46869 12580
rect 51339 12620 51381 12629
rect 51339 12580 51340 12620
rect 51380 12580 51381 12620
rect 51339 12571 51381 12580
rect 56427 12620 56469 12629
rect 56427 12580 56428 12620
rect 56468 12580 56469 12620
rect 56427 12571 56469 12580
rect 57675 12620 57717 12629
rect 57675 12580 57676 12620
rect 57716 12580 57717 12620
rect 57675 12571 57717 12580
rect 60267 12620 60309 12629
rect 60267 12580 60268 12620
rect 60308 12580 60309 12620
rect 60267 12571 60309 12580
rect 69483 12620 69525 12629
rect 69483 12580 69484 12620
rect 69524 12580 69525 12620
rect 69483 12571 69525 12580
rect 78211 12547 78269 12548
rect 44043 12529 44085 12538
rect 44427 12536 44469 12545
rect 43851 12487 43893 12496
rect 44427 12496 44428 12536
rect 44468 12496 44469 12536
rect 44427 12487 44469 12496
rect 44803 12536 44861 12537
rect 44803 12496 44812 12536
rect 44852 12496 44861 12536
rect 44803 12495 44861 12496
rect 45667 12536 45725 12537
rect 45667 12496 45676 12536
rect 45716 12496 45725 12536
rect 45667 12495 45725 12496
rect 45859 12536 45917 12537
rect 45859 12496 45868 12536
rect 45908 12496 45917 12536
rect 45859 12495 45917 12496
rect 45963 12536 46005 12545
rect 45963 12496 45964 12536
rect 46004 12496 46005 12536
rect 45963 12487 46005 12496
rect 46155 12536 46197 12545
rect 46155 12496 46156 12536
rect 46196 12496 46197 12536
rect 46155 12487 46197 12496
rect 46347 12536 46389 12545
rect 46347 12496 46348 12536
rect 46388 12496 46389 12536
rect 46347 12487 46389 12496
rect 46443 12536 46485 12545
rect 46443 12496 46444 12536
rect 46484 12496 46485 12536
rect 46443 12487 46485 12496
rect 46539 12536 46581 12545
rect 46539 12496 46540 12536
rect 46580 12496 46581 12536
rect 46539 12487 46581 12496
rect 46635 12536 46677 12545
rect 46635 12496 46636 12536
rect 46676 12496 46677 12536
rect 46635 12487 46677 12496
rect 47203 12536 47261 12537
rect 47203 12496 47212 12536
rect 47252 12496 47261 12536
rect 47203 12495 47261 12496
rect 48067 12536 48125 12537
rect 48067 12496 48076 12536
rect 48116 12496 48125 12536
rect 48067 12495 48125 12496
rect 49707 12536 49749 12545
rect 49707 12496 49708 12536
rect 49748 12496 49749 12536
rect 49707 12487 49749 12496
rect 49899 12536 49941 12545
rect 49899 12496 49900 12536
rect 49940 12496 49941 12536
rect 49899 12487 49941 12496
rect 49987 12536 50045 12537
rect 49987 12496 49996 12536
rect 50036 12496 50045 12536
rect 49987 12495 50045 12496
rect 50563 12536 50621 12537
rect 50563 12496 50572 12536
rect 50612 12496 50621 12536
rect 50563 12495 50621 12496
rect 50955 12536 50997 12545
rect 50955 12496 50956 12536
rect 50996 12496 50997 12536
rect 50955 12487 50997 12496
rect 51051 12536 51093 12545
rect 51051 12496 51052 12536
rect 51092 12496 51093 12536
rect 51051 12487 51093 12496
rect 51147 12536 51189 12545
rect 51147 12496 51148 12536
rect 51188 12496 51189 12536
rect 51147 12487 51189 12496
rect 51715 12536 51773 12537
rect 51715 12496 51724 12536
rect 51764 12496 51773 12536
rect 51715 12495 51773 12496
rect 52579 12536 52637 12537
rect 52579 12496 52588 12536
rect 52628 12496 52637 12536
rect 52579 12495 52637 12496
rect 55179 12536 55221 12545
rect 55179 12496 55180 12536
rect 55220 12496 55221 12536
rect 55179 12487 55221 12496
rect 55555 12536 55613 12537
rect 55555 12496 55564 12536
rect 55604 12496 55613 12536
rect 55555 12495 55613 12496
rect 56043 12536 56085 12545
rect 56043 12496 56044 12536
rect 56084 12496 56085 12536
rect 56043 12487 56085 12496
rect 56131 12536 56189 12537
rect 56131 12496 56140 12536
rect 56180 12496 56189 12536
rect 56131 12495 56189 12496
rect 56523 12536 56565 12545
rect 56523 12496 56524 12536
rect 56564 12496 56565 12536
rect 56523 12487 56565 12496
rect 56619 12536 56661 12545
rect 56619 12496 56620 12536
rect 56660 12496 56661 12536
rect 56619 12487 56661 12496
rect 56715 12536 56757 12545
rect 56715 12496 56716 12536
rect 56756 12496 56757 12536
rect 56715 12487 56757 12496
rect 58051 12536 58109 12537
rect 58051 12496 58060 12536
rect 58100 12496 58109 12536
rect 58051 12495 58109 12496
rect 58915 12536 58973 12537
rect 58915 12496 58924 12536
rect 58964 12496 58973 12536
rect 58915 12495 58973 12496
rect 60643 12536 60701 12537
rect 60643 12496 60652 12536
rect 60692 12496 60701 12536
rect 60643 12495 60701 12496
rect 61507 12536 61565 12537
rect 61507 12496 61516 12536
rect 61556 12496 61565 12536
rect 61507 12495 61565 12496
rect 62851 12536 62909 12537
rect 62851 12496 62860 12536
rect 62900 12496 62909 12536
rect 62851 12495 62909 12496
rect 63619 12536 63677 12537
rect 63619 12496 63628 12536
rect 63668 12496 63677 12536
rect 63619 12495 63677 12496
rect 64395 12536 64437 12545
rect 64395 12496 64396 12536
rect 64436 12496 64437 12536
rect 64395 12487 64437 12496
rect 64771 12536 64829 12537
rect 64771 12496 64780 12536
rect 64820 12496 64829 12536
rect 64771 12495 64829 12496
rect 65635 12536 65693 12537
rect 65635 12496 65644 12536
rect 65684 12496 65693 12536
rect 65635 12495 65693 12496
rect 67851 12536 67893 12545
rect 67851 12496 67852 12536
rect 67892 12496 67893 12536
rect 67851 12487 67893 12496
rect 67947 12536 67989 12545
rect 67947 12496 67948 12536
rect 67988 12496 67989 12536
rect 67947 12487 67989 12496
rect 68043 12536 68085 12545
rect 68043 12496 68044 12536
rect 68084 12496 68085 12536
rect 68043 12487 68085 12496
rect 68139 12536 68181 12545
rect 68139 12496 68140 12536
rect 68180 12496 68181 12536
rect 68139 12487 68181 12496
rect 69859 12536 69917 12537
rect 69859 12496 69868 12536
rect 69908 12496 69917 12536
rect 69859 12495 69917 12496
rect 70723 12536 70781 12537
rect 70723 12496 70732 12536
rect 70772 12496 70781 12536
rect 70723 12495 70781 12496
rect 72067 12536 72125 12537
rect 72067 12496 72076 12536
rect 72116 12496 72125 12536
rect 72067 12495 72125 12496
rect 72651 12536 72693 12545
rect 72651 12496 72652 12536
rect 72692 12496 72693 12536
rect 72651 12487 72693 12496
rect 73027 12536 73085 12537
rect 73027 12496 73036 12536
rect 73076 12496 73085 12536
rect 73027 12495 73085 12496
rect 73891 12536 73949 12537
rect 73891 12496 73900 12536
rect 73940 12496 73949 12536
rect 73891 12495 73949 12496
rect 76395 12536 76437 12545
rect 76395 12496 76396 12536
rect 76436 12496 76437 12536
rect 76395 12487 76437 12496
rect 76771 12536 76829 12537
rect 76771 12496 76780 12536
rect 76820 12496 76829 12536
rect 76771 12495 76829 12496
rect 77163 12536 77205 12545
rect 77163 12496 77164 12536
rect 77204 12496 77205 12536
rect 77163 12487 77205 12496
rect 77259 12536 77301 12545
rect 77259 12496 77260 12536
rect 77300 12496 77301 12536
rect 77259 12487 77301 12496
rect 77451 12536 77493 12545
rect 77451 12496 77452 12536
rect 77492 12496 77493 12536
rect 77347 12494 77405 12495
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1699 12452 1757 12453
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 1699 12411 1757 12412
rect 44523 12452 44565 12461
rect 44523 12412 44524 12452
rect 44564 12412 44565 12452
rect 44523 12403 44565 12412
rect 44715 12452 44757 12461
rect 44715 12412 44716 12452
rect 44756 12412 44757 12452
rect 44715 12403 44757 12412
rect 55275 12452 55317 12461
rect 55275 12412 55276 12452
rect 55316 12412 55317 12452
rect 55275 12403 55317 12412
rect 55467 12452 55509 12461
rect 55467 12412 55468 12452
rect 55508 12412 55509 12452
rect 55467 12403 55509 12412
rect 71883 12452 71925 12461
rect 71883 12412 71884 12452
rect 71924 12412 71925 12452
rect 71883 12403 71925 12412
rect 76491 12452 76533 12461
rect 76491 12412 76492 12452
rect 76532 12412 76533 12452
rect 76491 12403 76533 12412
rect 76683 12452 76725 12461
rect 77347 12454 77356 12494
rect 77396 12454 77405 12494
rect 77451 12487 77493 12496
rect 77643 12536 77685 12545
rect 77643 12496 77644 12536
rect 77684 12496 77685 12536
rect 77643 12487 77685 12496
rect 77739 12536 77781 12545
rect 77739 12496 77740 12536
rect 77780 12496 77781 12536
rect 77739 12487 77781 12496
rect 77835 12536 77877 12545
rect 77835 12496 77836 12536
rect 77876 12496 77877 12536
rect 77835 12487 77877 12496
rect 77931 12536 77973 12545
rect 77931 12496 77932 12536
rect 77972 12496 77973 12536
rect 78211 12507 78220 12547
rect 78260 12507 78269 12547
rect 78211 12506 78269 12507
rect 77931 12487 77973 12496
rect 77347 12453 77405 12454
rect 76683 12412 76684 12452
rect 76724 12412 76725 12452
rect 76683 12403 76725 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 41547 12368 41589 12377
rect 41547 12328 41548 12368
rect 41588 12328 41589 12368
rect 41547 12319 41589 12328
rect 44043 12368 44085 12377
rect 44043 12328 44044 12368
rect 44084 12328 44085 12368
rect 44043 12319 44085 12328
rect 44619 12368 44661 12377
rect 44619 12328 44620 12368
rect 44660 12328 44661 12368
rect 44619 12319 44661 12328
rect 55371 12368 55413 12377
rect 55371 12328 55372 12368
rect 55412 12328 55413 12368
rect 55371 12319 55413 12328
rect 55755 12368 55797 12377
rect 55755 12328 55756 12368
rect 55796 12328 55797 12368
rect 55755 12319 55797 12328
rect 76587 12368 76629 12377
rect 76587 12328 76588 12368
rect 76628 12328 76629 12368
rect 76587 12319 76629 12328
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 43467 12284 43509 12293
rect 43467 12244 43468 12284
rect 43508 12244 43509 12284
rect 43467 12235 43509 12244
rect 46155 12284 46197 12293
rect 46155 12244 46156 12284
rect 46196 12244 46197 12284
rect 46155 12235 46197 12244
rect 50667 12284 50709 12293
rect 50667 12244 50668 12284
rect 50708 12244 50709 12284
rect 50667 12235 50709 12244
rect 53731 12284 53789 12285
rect 53731 12244 53740 12284
rect 53780 12244 53789 12284
rect 53731 12243 53789 12244
rect 62659 12284 62717 12285
rect 62659 12244 62668 12284
rect 62708 12244 62717 12284
rect 62659 12243 62717 12244
rect 63723 12284 63765 12293
rect 63723 12244 63724 12284
rect 63764 12244 63765 12284
rect 63723 12235 63765 12244
rect 78123 12284 78165 12293
rect 78123 12244 78124 12284
rect 78164 12244 78165 12284
rect 78123 12235 78165 12244
rect 576 12116 79584 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 75112 12116
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75480 12076 79584 12116
rect 576 12052 79584 12076
rect 50659 11948 50717 11949
rect 50659 11908 50668 11948
rect 50708 11908 50717 11948
rect 50659 11907 50717 11908
rect 51339 11948 51381 11957
rect 51339 11908 51340 11948
rect 51380 11908 51381 11948
rect 51339 11899 51381 11908
rect 56523 11948 56565 11957
rect 56523 11908 56524 11948
rect 56564 11908 56565 11948
rect 56523 11899 56565 11908
rect 65155 11948 65213 11949
rect 65155 11908 65164 11948
rect 65204 11908 65213 11948
rect 65155 11907 65213 11908
rect 70051 11948 70109 11949
rect 70051 11908 70060 11948
rect 70100 11908 70109 11948
rect 70051 11907 70109 11908
rect 76491 11948 76533 11957
rect 76491 11908 76492 11948
rect 76532 11908 76533 11948
rect 76491 11899 76533 11908
rect 79363 11948 79421 11949
rect 79363 11908 79372 11948
rect 79412 11908 79421 11948
rect 79363 11907 79421 11908
rect 46923 11864 46965 11873
rect 46923 11824 46924 11864
rect 46964 11824 46965 11864
rect 46923 11815 46965 11824
rect 61227 11864 61269 11873
rect 61227 11824 61228 11864
rect 61268 11824 61269 11864
rect 61227 11815 61269 11824
rect 65547 11864 65589 11873
rect 65547 11824 65548 11864
rect 65588 11824 65589 11864
rect 65547 11815 65589 11824
rect 65931 11864 65973 11873
rect 65931 11824 65932 11864
rect 65972 11824 65973 11864
rect 65931 11815 65973 11824
rect 72843 11864 72885 11873
rect 72843 11824 72844 11864
rect 72884 11824 72885 11864
rect 72843 11815 72885 11824
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 1699 11780 1757 11781
rect 1699 11740 1708 11780
rect 1748 11740 1757 11780
rect 1699 11739 1757 11740
rect 43659 11780 43701 11789
rect 43659 11740 43660 11780
rect 43700 11740 43701 11780
rect 43659 11731 43701 11740
rect 53355 11780 53397 11789
rect 53355 11740 53356 11780
rect 53396 11740 53397 11780
rect 59971 11780 60029 11781
rect 53355 11731 53397 11740
rect 55755 11738 55797 11747
rect 59971 11740 59980 11780
rect 60020 11740 60029 11780
rect 59971 11739 60029 11740
rect 61411 11780 61469 11781
rect 61411 11740 61420 11780
rect 61460 11740 61469 11780
rect 61411 11739 61469 11740
rect 65451 11780 65493 11789
rect 65451 11740 65452 11780
rect 65492 11740 65493 11780
rect 41635 11696 41693 11697
rect 41635 11656 41644 11696
rect 41684 11656 41693 11696
rect 41635 11655 41693 11656
rect 42499 11696 42557 11697
rect 42499 11656 42508 11696
rect 42548 11656 42557 11696
rect 42499 11655 42557 11656
rect 44995 11696 45053 11697
rect 44995 11656 45004 11696
rect 45044 11656 45053 11696
rect 44995 11655 45053 11656
rect 45859 11696 45917 11697
rect 45859 11656 45868 11696
rect 45908 11656 45917 11696
rect 45859 11655 45917 11656
rect 46531 11696 46589 11697
rect 46531 11656 46540 11696
rect 46580 11656 46589 11696
rect 46531 11655 46589 11656
rect 46635 11696 46677 11705
rect 46635 11656 46636 11696
rect 46676 11656 46677 11696
rect 46635 11647 46677 11656
rect 48643 11696 48701 11697
rect 48643 11656 48652 11696
rect 48692 11656 48701 11696
rect 48643 11655 48701 11656
rect 49507 11696 49565 11697
rect 49507 11656 49516 11696
rect 49556 11656 49565 11696
rect 49507 11655 49565 11656
rect 50947 11696 51005 11697
rect 50947 11656 50956 11696
rect 50996 11656 51005 11696
rect 50947 11655 51005 11656
rect 51051 11696 51093 11705
rect 51051 11656 51052 11696
rect 51092 11656 51093 11696
rect 51051 11647 51093 11656
rect 51627 11696 51669 11705
rect 51627 11656 51628 11696
rect 51668 11656 51669 11696
rect 51627 11647 51669 11656
rect 51723 11696 51765 11705
rect 51723 11656 51724 11696
rect 51764 11656 51765 11696
rect 51723 11647 51765 11656
rect 51819 11696 51861 11705
rect 55755 11698 55756 11738
rect 55796 11698 55797 11738
rect 56131 11738 56189 11739
rect 51819 11656 51820 11696
rect 51860 11656 51861 11696
rect 51819 11647 51861 11656
rect 54499 11696 54557 11697
rect 54499 11656 54508 11696
rect 54548 11656 54557 11696
rect 54499 11655 54557 11656
rect 55363 11696 55421 11697
rect 55363 11656 55372 11696
rect 55412 11656 55421 11696
rect 55755 11689 55797 11698
rect 56043 11696 56085 11705
rect 56131 11698 56140 11738
rect 56180 11698 56189 11738
rect 65451 11731 65493 11740
rect 65643 11780 65685 11789
rect 65643 11740 65644 11780
rect 65684 11740 65685 11780
rect 65643 11731 65685 11740
rect 56131 11697 56189 11698
rect 55363 11655 55421 11656
rect 56043 11656 56044 11696
rect 56084 11656 56085 11696
rect 56419 11696 56477 11697
rect 56043 11647 56085 11656
rect 56235 11675 56277 11684
rect 56235 11635 56236 11675
rect 56276 11635 56277 11675
rect 56419 11656 56428 11696
rect 56468 11656 56477 11696
rect 56419 11655 56477 11656
rect 59019 11696 59061 11705
rect 59019 11656 59020 11696
rect 59060 11656 59061 11696
rect 59019 11647 59061 11656
rect 59115 11696 59157 11705
rect 59115 11656 59116 11696
rect 59156 11656 59157 11696
rect 59115 11647 59157 11656
rect 59211 11696 59253 11705
rect 59211 11656 59212 11696
rect 59252 11656 59253 11696
rect 59211 11647 59253 11656
rect 59595 11696 59637 11705
rect 59595 11656 59596 11696
rect 59636 11656 59637 11696
rect 59595 11647 59637 11656
rect 59691 11696 59733 11705
rect 59691 11656 59692 11696
rect 59732 11656 59733 11696
rect 59691 11647 59733 11656
rect 59787 11696 59829 11705
rect 59787 11656 59788 11696
rect 59828 11656 59829 11696
rect 59787 11647 59829 11656
rect 62187 11696 62229 11705
rect 62187 11656 62188 11696
rect 62228 11656 62229 11696
rect 62187 11647 62229 11656
rect 62379 11696 62421 11705
rect 62379 11656 62380 11696
rect 62420 11656 62421 11696
rect 62379 11647 62421 11656
rect 62467 11696 62525 11697
rect 62467 11656 62476 11696
rect 62516 11656 62525 11696
rect 62467 11655 62525 11656
rect 63139 11696 63197 11697
rect 63139 11656 63148 11696
rect 63188 11656 63197 11696
rect 63139 11655 63197 11656
rect 64003 11696 64061 11697
rect 64003 11656 64012 11696
rect 64052 11656 64061 11696
rect 64003 11655 64061 11656
rect 65347 11696 65405 11697
rect 65347 11656 65356 11696
rect 65396 11656 65405 11696
rect 65347 11655 65405 11656
rect 65739 11696 65781 11705
rect 65739 11656 65740 11696
rect 65780 11656 65781 11696
rect 65739 11647 65781 11656
rect 65931 11696 65973 11705
rect 65931 11656 65932 11696
rect 65972 11656 65973 11696
rect 65931 11647 65973 11656
rect 66123 11696 66165 11705
rect 66123 11656 66124 11696
rect 66164 11656 66165 11696
rect 66123 11647 66165 11656
rect 66211 11696 66269 11697
rect 66211 11656 66220 11696
rect 66260 11656 66269 11696
rect 66211 11655 66269 11656
rect 66883 11696 66941 11697
rect 66883 11656 66892 11696
rect 66932 11656 66941 11696
rect 66883 11655 66941 11656
rect 67179 11696 67221 11705
rect 67179 11656 67180 11696
rect 67220 11656 67221 11696
rect 67179 11647 67221 11656
rect 67275 11696 67317 11705
rect 67275 11656 67276 11696
rect 67316 11656 67317 11696
rect 67275 11647 67317 11656
rect 67371 11696 67413 11705
rect 67371 11656 67372 11696
rect 67412 11656 67413 11696
rect 67371 11647 67413 11656
rect 68035 11696 68093 11697
rect 68035 11656 68044 11696
rect 68084 11656 68093 11696
rect 68035 11655 68093 11656
rect 68899 11696 68957 11697
rect 68899 11656 68908 11696
rect 68948 11656 68957 11696
rect 68899 11655 68957 11656
rect 71595 11696 71637 11705
rect 71595 11656 71596 11696
rect 71636 11656 71637 11696
rect 71595 11647 71637 11656
rect 71787 11696 71829 11705
rect 71787 11656 71788 11696
rect 71828 11656 71829 11696
rect 71787 11647 71829 11656
rect 71875 11696 71933 11697
rect 71875 11656 71884 11696
rect 71924 11656 71933 11696
rect 71875 11655 71933 11656
rect 72163 11696 72221 11697
rect 72163 11656 72172 11696
rect 72212 11656 72221 11696
rect 72163 11655 72221 11656
rect 72451 11696 72509 11697
rect 72451 11656 72460 11696
rect 72500 11656 72509 11696
rect 72451 11655 72509 11656
rect 72555 11696 72597 11705
rect 72555 11656 72556 11696
rect 72596 11656 72597 11696
rect 72555 11647 72597 11656
rect 73035 11696 73077 11705
rect 73035 11656 73036 11696
rect 73076 11656 73077 11696
rect 73035 11647 73077 11656
rect 73131 11696 73173 11705
rect 73131 11656 73132 11696
rect 73172 11656 73173 11696
rect 73131 11647 73173 11656
rect 73227 11696 73269 11705
rect 73227 11656 73228 11696
rect 73268 11656 73269 11696
rect 73227 11647 73269 11656
rect 73323 11696 73365 11705
rect 73323 11656 73324 11696
rect 73364 11656 73365 11696
rect 73323 11647 73365 11656
rect 73515 11696 73557 11705
rect 73515 11656 73516 11696
rect 73556 11656 73557 11696
rect 73515 11647 73557 11656
rect 73611 11696 73653 11705
rect 73611 11656 73612 11696
rect 73652 11656 73653 11696
rect 73611 11647 73653 11656
rect 73707 11696 73749 11705
rect 73707 11656 73708 11696
rect 73748 11656 73749 11696
rect 73707 11647 73749 11656
rect 73803 11696 73845 11705
rect 73803 11656 73804 11696
rect 73844 11656 73845 11696
rect 73803 11647 73845 11656
rect 76491 11696 76533 11705
rect 76491 11656 76492 11696
rect 76532 11656 76533 11696
rect 76491 11647 76533 11656
rect 76683 11696 76725 11705
rect 76683 11656 76684 11696
rect 76724 11656 76725 11696
rect 76683 11647 76725 11656
rect 76771 11696 76829 11697
rect 76771 11656 76780 11696
rect 76820 11656 76829 11696
rect 76771 11655 76829 11656
rect 76971 11696 77013 11705
rect 76971 11656 76972 11696
rect 77012 11656 77013 11696
rect 76971 11647 77013 11656
rect 77347 11696 77405 11697
rect 77347 11656 77356 11696
rect 77396 11656 77405 11696
rect 77347 11655 77405 11656
rect 78211 11696 78269 11697
rect 78211 11656 78220 11696
rect 78260 11656 78269 11696
rect 78211 11655 78269 11656
rect 56235 11626 56277 11635
rect 41259 11612 41301 11621
rect 41259 11572 41260 11612
rect 41300 11572 41301 11612
rect 41259 11563 41301 11572
rect 46251 11612 46293 11621
rect 46251 11572 46252 11612
rect 46292 11572 46293 11612
rect 46251 11563 46293 11572
rect 48267 11612 48309 11621
rect 48267 11572 48268 11612
rect 48308 11572 48309 11612
rect 48267 11563 48309 11572
rect 51531 11612 51573 11621
rect 51531 11572 51532 11612
rect 51572 11572 51573 11612
rect 51235 11570 51293 11571
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 1515 11528 1557 11537
rect 1515 11488 1516 11528
rect 1556 11488 1557 11528
rect 1515 11479 1557 11488
rect 43843 11528 43901 11529
rect 43843 11488 43852 11528
rect 43892 11488 43901 11528
rect 43843 11487 43901 11488
rect 50859 11524 50901 11533
rect 51235 11530 51244 11570
rect 51284 11530 51293 11570
rect 51531 11563 51573 11572
rect 62283 11612 62325 11621
rect 62283 11572 62284 11612
rect 62324 11572 62325 11612
rect 62283 11563 62325 11572
rect 62763 11612 62805 11621
rect 62763 11572 62764 11612
rect 62804 11572 62805 11612
rect 62763 11563 62805 11572
rect 67467 11612 67509 11621
rect 67467 11572 67468 11612
rect 67508 11572 67509 11612
rect 67467 11563 67509 11572
rect 67659 11612 67701 11621
rect 67659 11572 67660 11612
rect 67700 11572 67701 11612
rect 67659 11563 67701 11572
rect 51235 11529 51293 11530
rect 50859 11484 50860 11524
rect 50900 11484 50901 11524
rect 55939 11528 55997 11529
rect 55939 11488 55948 11528
rect 55988 11488 55997 11528
rect 55939 11487 55997 11488
rect 58915 11528 58973 11529
rect 58915 11488 58924 11528
rect 58964 11488 58973 11528
rect 58915 11487 58973 11488
rect 59491 11528 59549 11529
rect 59491 11488 59500 11528
rect 59540 11488 59549 11528
rect 59491 11487 59549 11488
rect 60171 11528 60213 11537
rect 60171 11488 60172 11528
rect 60212 11488 60213 11528
rect 46443 11470 46485 11479
rect 50859 11475 50901 11484
rect 60171 11479 60213 11488
rect 66987 11528 67029 11537
rect 66987 11488 66988 11528
rect 67028 11488 67029 11528
rect 66987 11479 67029 11488
rect 71683 11528 71741 11529
rect 71683 11488 71692 11528
rect 71732 11488 71741 11528
rect 71683 11487 71741 11488
rect 72075 11528 72117 11537
rect 72075 11488 72076 11528
rect 72116 11488 72117 11528
rect 72075 11479 72117 11488
rect 72363 11524 72405 11533
rect 72363 11484 72364 11524
rect 72404 11484 72405 11524
rect 72363 11475 72405 11484
rect 46443 11430 46444 11470
rect 46484 11430 46485 11470
rect 46443 11421 46485 11430
rect 576 11360 79584 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 76352 11360
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76720 11320 79584 11360
rect 576 11296 79584 11320
rect 67851 11250 67893 11259
rect 67851 11210 67852 11250
rect 67892 11210 67893 11250
rect 43467 11196 43509 11205
rect 42499 11192 42557 11193
rect 42499 11152 42508 11192
rect 42548 11152 42557 11192
rect 42499 11151 42557 11152
rect 43467 11156 43468 11196
rect 43508 11156 43509 11196
rect 43467 11147 43509 11156
rect 46347 11192 46389 11201
rect 46347 11152 46348 11192
rect 46388 11152 46389 11192
rect 46347 11143 46389 11152
rect 49419 11192 49461 11201
rect 49419 11152 49420 11192
rect 49460 11152 49461 11192
rect 49419 11143 49461 11152
rect 52779 11192 52821 11201
rect 62763 11196 62805 11205
rect 67851 11201 67893 11210
rect 52779 11152 52780 11192
rect 52820 11152 52821 11192
rect 52779 11143 52821 11152
rect 58627 11192 58685 11193
rect 58627 11152 58636 11192
rect 58676 11152 58685 11192
rect 58627 11151 58685 11152
rect 61315 11192 61373 11193
rect 61315 11152 61324 11192
rect 61364 11152 61373 11192
rect 61315 11151 61373 11152
rect 62763 11156 62764 11196
rect 62804 11156 62805 11196
rect 62763 11147 62805 11156
rect 62947 11192 63005 11193
rect 62947 11152 62956 11192
rect 62996 11152 63005 11192
rect 62947 11151 63005 11152
rect 64771 11192 64829 11193
rect 64771 11152 64780 11192
rect 64820 11152 64829 11192
rect 64771 11151 64829 11152
rect 72355 11192 72413 11193
rect 72355 11152 72364 11192
rect 72404 11152 72413 11192
rect 72355 11151 72413 11152
rect 74091 11192 74133 11201
rect 77739 11196 77781 11205
rect 74091 11152 74092 11192
rect 74132 11152 74133 11192
rect 74091 11143 74133 11152
rect 77059 11192 77117 11193
rect 77059 11152 77068 11192
rect 77108 11152 77117 11192
rect 77059 11151 77117 11152
rect 77739 11156 77740 11196
rect 77780 11156 77781 11196
rect 77739 11147 77781 11156
rect 43659 11108 43701 11117
rect 43659 11068 43660 11108
rect 43700 11068 43701 11108
rect 43659 11059 43701 11068
rect 58923 11108 58965 11117
rect 58923 11068 58924 11108
rect 58964 11068 58965 11108
rect 58923 11059 58965 11068
rect 42603 11024 42645 11033
rect 42603 10984 42604 11024
rect 42644 10984 42645 11024
rect 42603 10975 42645 10984
rect 42699 11024 42741 11033
rect 42699 10984 42700 11024
rect 42740 10984 42741 11024
rect 42699 10975 42741 10984
rect 42795 11024 42837 11033
rect 42795 10984 42796 11024
rect 42836 10984 42837 11024
rect 42795 10975 42837 10984
rect 43275 11024 43317 11033
rect 43275 10984 43276 11024
rect 43316 10984 43317 11024
rect 43275 10975 43317 10984
rect 43363 11024 43421 11025
rect 43363 10984 43372 11024
rect 43412 10984 43421 11024
rect 43363 10983 43421 10984
rect 43755 11024 43797 11033
rect 43755 10984 43756 11024
rect 43796 10984 43797 11024
rect 43755 10975 43797 10984
rect 43851 11024 43893 11033
rect 43851 10984 43852 11024
rect 43892 10984 43893 11024
rect 43851 10975 43893 10984
rect 43947 11024 43989 11033
rect 43947 10984 43948 11024
rect 43988 10984 43989 11024
rect 43947 10975 43989 10984
rect 44139 11024 44181 11033
rect 44139 10984 44140 11024
rect 44180 10984 44181 11024
rect 44139 10975 44181 10984
rect 44331 11024 44373 11033
rect 44331 10984 44332 11024
rect 44372 10984 44373 11024
rect 44331 10975 44373 10984
rect 44419 11024 44477 11025
rect 44419 10984 44428 11024
rect 44468 10984 44477 11024
rect 44419 10983 44477 10984
rect 45667 11024 45725 11025
rect 45667 10984 45676 11024
rect 45716 10984 45725 11024
rect 45667 10983 45725 10984
rect 46059 11024 46101 11033
rect 46059 10984 46060 11024
rect 46100 10984 46101 11024
rect 46059 10975 46101 10984
rect 46243 11024 46301 11025
rect 46243 10984 46252 11024
rect 46292 10984 46301 11024
rect 46243 10983 46301 10984
rect 49315 11024 49373 11025
rect 49315 10984 49324 11024
rect 49364 10984 49373 11024
rect 49315 10983 49373 10984
rect 50659 11024 50717 11025
rect 50659 10984 50668 11024
rect 50708 10984 50717 11024
rect 50659 10983 50717 10984
rect 51051 11024 51093 11033
rect 51051 10984 51052 11024
rect 51092 10984 51093 11024
rect 51051 10975 51093 10984
rect 51435 11024 51477 11033
rect 51435 10984 51436 11024
rect 51476 10984 51477 11024
rect 51435 10975 51477 10984
rect 51531 11024 51573 11033
rect 51531 10984 51532 11024
rect 51572 10984 51573 11024
rect 51531 10975 51573 10984
rect 51627 11024 51669 11033
rect 51627 10984 51628 11024
rect 51668 10984 51669 11024
rect 51627 10975 51669 10984
rect 51723 11024 51765 11033
rect 51723 10984 51724 11024
rect 51764 10984 51765 11024
rect 51723 10975 51765 10984
rect 51915 11024 51957 11033
rect 51915 10984 51916 11024
rect 51956 10984 51957 11024
rect 51915 10975 51957 10984
rect 52011 11024 52053 11033
rect 52011 10984 52012 11024
rect 52052 10984 52053 11024
rect 52011 10975 52053 10984
rect 52107 11024 52149 11033
rect 52107 10984 52108 11024
rect 52148 10984 52149 11024
rect 52107 10975 52149 10984
rect 52203 11024 52245 11033
rect 52203 10984 52204 11024
rect 52244 10984 52245 11024
rect 52203 10975 52245 10984
rect 52867 11024 52925 11025
rect 52867 10984 52876 11024
rect 52916 10984 52925 11024
rect 52867 10983 52925 10984
rect 55179 11024 55221 11033
rect 55179 10984 55180 11024
rect 55220 10984 55221 11024
rect 55179 10975 55221 10984
rect 55371 11024 55413 11033
rect 55371 10984 55372 11024
rect 55412 10984 55413 11024
rect 55371 10975 55413 10984
rect 55459 11024 55517 11025
rect 55459 10984 55468 11024
rect 55508 10984 55517 11024
rect 55459 10983 55517 10984
rect 55755 11024 55797 11033
rect 55755 10984 55756 11024
rect 55796 10984 55797 11024
rect 55755 10975 55797 10984
rect 55851 11024 55893 11033
rect 55851 10984 55852 11024
rect 55892 10984 55893 11024
rect 55851 10975 55893 10984
rect 55947 11024 55989 11033
rect 55947 10984 55948 11024
rect 55988 10984 55989 11024
rect 55947 10975 55989 10984
rect 56043 11024 56085 11033
rect 56043 10984 56044 11024
rect 56084 10984 56085 11024
rect 56043 10975 56085 10984
rect 56235 11024 56277 11033
rect 56235 10984 56236 11024
rect 56276 10984 56277 11024
rect 56235 10975 56277 10984
rect 56611 11024 56669 11025
rect 56611 10984 56620 11024
rect 56660 10984 56669 11024
rect 56611 10983 56669 10984
rect 57475 11024 57533 11025
rect 57475 10984 57484 11024
rect 57524 10984 57533 11024
rect 57475 10983 57533 10984
rect 59299 11024 59357 11025
rect 59299 10984 59308 11024
rect 59348 10984 59357 11024
rect 59299 10983 59357 10984
rect 60163 11024 60221 11025
rect 60163 10984 60172 11024
rect 60212 10984 60221 11024
rect 60163 10983 60221 10984
rect 61707 11024 61749 11033
rect 61707 10984 61708 11024
rect 61748 10984 61749 11024
rect 62083 11024 62141 11025
rect 61707 10975 61749 10984
rect 61803 10982 61845 10991
rect 62083 10984 62092 11024
rect 62132 10984 62141 11024
rect 62083 10983 62141 10984
rect 62571 11024 62613 11033
rect 62571 10984 62572 11024
rect 62612 10984 62613 11024
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 45771 10940 45813 10949
rect 45771 10900 45772 10940
rect 45812 10900 45813 10940
rect 45771 10891 45813 10900
rect 45963 10940 46005 10949
rect 45963 10900 45964 10940
rect 46004 10900 46005 10940
rect 45963 10891 46005 10900
rect 50275 10940 50333 10941
rect 50275 10900 50284 10940
rect 50324 10900 50333 10940
rect 50275 10899 50333 10900
rect 50763 10940 50805 10949
rect 50763 10900 50764 10940
rect 50804 10900 50805 10940
rect 50763 10891 50805 10900
rect 50955 10940 50997 10949
rect 61803 10942 61804 10982
rect 61844 10942 61845 10982
rect 62571 10975 62613 10984
rect 62659 11024 62717 11025
rect 62659 10984 62668 11024
rect 62708 10984 62717 11024
rect 62659 10983 62717 10984
rect 63051 11024 63093 11033
rect 63051 10984 63052 11024
rect 63092 10984 63093 11024
rect 63051 10975 63093 10984
rect 63147 11024 63189 11033
rect 63147 10984 63148 11024
rect 63188 10984 63189 11024
rect 63147 10975 63189 10984
rect 63243 11024 63285 11033
rect 63243 10984 63244 11024
rect 63284 10984 63285 11024
rect 63243 10975 63285 10984
rect 63435 11024 63477 11033
rect 63435 10984 63436 11024
rect 63476 10984 63477 11024
rect 63435 10975 63477 10984
rect 63531 11024 63573 11033
rect 63531 10984 63532 11024
rect 63572 10984 63573 11024
rect 63531 10975 63573 10984
rect 63627 11024 63669 11033
rect 63627 10984 63628 11024
rect 63668 10984 63669 11024
rect 63627 10975 63669 10984
rect 63723 11024 63765 11033
rect 63723 10984 63724 11024
rect 63764 10984 63765 11024
rect 63723 10975 63765 10984
rect 65923 11024 65981 11025
rect 65923 10984 65932 11024
rect 65972 10984 65981 11024
rect 65923 10983 65981 10984
rect 66787 11024 66845 11025
rect 66787 10984 66796 11024
rect 66836 10984 66845 11024
rect 66787 10983 66845 10984
rect 67179 11024 67221 11033
rect 67179 10984 67180 11024
rect 67220 10984 67221 11024
rect 67179 10975 67221 10984
rect 67659 11024 67701 11033
rect 67659 10984 67660 11024
rect 67700 10984 67701 11024
rect 67659 10975 67701 10984
rect 67747 11024 67805 11025
rect 67747 10984 67756 11024
rect 67796 10984 67805 11024
rect 67747 10983 67805 10984
rect 69963 11024 70005 11033
rect 69963 10984 69964 11024
rect 70004 10984 70005 11024
rect 69963 10975 70005 10984
rect 70339 11024 70397 11025
rect 70339 10984 70348 11024
rect 70388 10984 70397 11024
rect 70339 10983 70397 10984
rect 71203 11024 71261 11025
rect 71203 10984 71212 11024
rect 71252 10984 71261 11024
rect 71203 10983 71261 10984
rect 72747 11024 72789 11033
rect 72747 10984 72748 11024
rect 72788 10984 72789 11024
rect 72747 10975 72789 10984
rect 72843 11024 72885 11033
rect 72843 10984 72844 11024
rect 72884 10984 72885 11024
rect 72843 10975 72885 10984
rect 72939 11024 72981 11033
rect 72939 10984 72940 11024
rect 72980 10984 72981 11024
rect 72939 10975 72981 10984
rect 73035 11024 73077 11033
rect 73035 10984 73036 11024
rect 73076 10984 73077 11024
rect 73035 10975 73077 10984
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 75043 11024 75101 11025
rect 75043 10984 75052 11024
rect 75092 10984 75101 11024
rect 75043 10983 75101 10984
rect 75907 11024 75965 11025
rect 75907 10984 75916 11024
rect 75956 10984 75965 11024
rect 75907 10983 75965 10984
rect 77547 11024 77589 11033
rect 77547 10984 77548 11024
rect 77588 10984 77589 11024
rect 77547 10975 77589 10984
rect 77635 11024 77693 11025
rect 77635 10984 77644 11024
rect 77684 10984 77693 11024
rect 77635 10983 77693 10984
rect 77923 11024 77981 11025
rect 77923 10984 77932 11024
rect 77972 10984 77981 11024
rect 77923 10983 77981 10984
rect 50955 10900 50956 10940
rect 50996 10900 50997 10940
rect 50955 10891 50997 10900
rect 52387 10940 52445 10941
rect 52387 10900 52396 10940
rect 52436 10900 52445 10940
rect 61803 10933 61845 10942
rect 61995 10940 62037 10949
rect 52387 10899 52445 10900
rect 61995 10900 61996 10940
rect 62036 10900 62037 10940
rect 61995 10891 62037 10900
rect 68899 10940 68957 10941
rect 68899 10900 68908 10940
rect 68948 10900 68957 10940
rect 68899 10899 68957 10900
rect 73507 10940 73565 10941
rect 73507 10900 73516 10940
rect 73556 10900 73565 10940
rect 73507 10899 73565 10900
rect 73891 10940 73949 10941
rect 73891 10900 73900 10940
rect 73940 10900 73949 10940
rect 73891 10899 73949 10900
rect 45867 10856 45909 10865
rect 45867 10816 45868 10856
rect 45908 10816 45909 10856
rect 45867 10807 45909 10816
rect 50859 10856 50901 10865
rect 50859 10816 50860 10856
rect 50900 10816 50901 10856
rect 50859 10807 50901 10816
rect 61899 10856 61941 10865
rect 61899 10816 61900 10856
rect 61940 10816 61941 10856
rect 61899 10807 61941 10816
rect 67371 10856 67413 10865
rect 67371 10816 67372 10856
rect 67412 10816 67413 10856
rect 67371 10807 67413 10816
rect 77259 10856 77301 10865
rect 77259 10816 77260 10856
rect 77300 10816 77301 10856
rect 77259 10807 77301 10816
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 42987 10772 43029 10781
rect 42987 10732 42988 10772
rect 43028 10732 43029 10772
rect 42987 10723 43029 10732
rect 44139 10772 44181 10781
rect 44139 10732 44140 10772
rect 44180 10732 44181 10772
rect 44139 10723 44181 10732
rect 49419 10772 49461 10781
rect 49419 10732 49420 10772
rect 49460 10732 49461 10772
rect 49419 10723 49461 10732
rect 50475 10772 50517 10781
rect 50475 10732 50476 10772
rect 50516 10732 50517 10772
rect 50475 10723 50517 10732
rect 52587 10772 52629 10781
rect 52587 10732 52588 10772
rect 52628 10732 52629 10772
rect 52587 10723 52629 10732
rect 55179 10772 55221 10781
rect 55179 10732 55180 10772
rect 55220 10732 55221 10772
rect 55179 10723 55221 10732
rect 62283 10772 62325 10781
rect 62283 10732 62284 10772
rect 62324 10732 62325 10772
rect 62283 10723 62325 10732
rect 68715 10772 68757 10781
rect 68715 10732 68716 10772
rect 68756 10732 68757 10772
rect 68715 10723 68757 10732
rect 72355 10772 72413 10773
rect 72355 10732 72364 10772
rect 72404 10732 72413 10772
rect 72355 10731 72413 10732
rect 73323 10772 73365 10781
rect 73323 10732 73324 10772
rect 73364 10732 73365 10772
rect 73323 10723 73365 10732
rect 78027 10772 78069 10781
rect 78027 10732 78028 10772
rect 78068 10732 78069 10772
rect 78027 10723 78069 10732
rect 576 10604 79584 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 75112 10604
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75480 10564 79584 10604
rect 576 10540 79584 10564
rect 44715 10436 44757 10445
rect 44715 10396 44716 10436
rect 44756 10396 44757 10436
rect 44715 10387 44757 10396
rect 47779 10436 47837 10437
rect 47779 10396 47788 10436
rect 47828 10396 47837 10436
rect 47779 10395 47837 10396
rect 50371 10436 50429 10437
rect 50371 10396 50380 10436
rect 50420 10396 50429 10436
rect 50371 10395 50429 10396
rect 51147 10436 51189 10445
rect 51147 10396 51148 10436
rect 51188 10396 51189 10436
rect 51147 10387 51189 10396
rect 54115 10436 54173 10437
rect 54115 10396 54124 10436
rect 54164 10396 54173 10436
rect 54115 10395 54173 10396
rect 58443 10436 58485 10445
rect 58443 10396 58444 10436
rect 58484 10396 58485 10436
rect 58443 10387 58485 10396
rect 59595 10436 59637 10445
rect 59595 10396 59596 10436
rect 59636 10396 59637 10436
rect 59595 10387 59637 10396
rect 59979 10436 60021 10445
rect 59979 10396 59980 10436
rect 60020 10396 60021 10436
rect 59979 10387 60021 10396
rect 63339 10436 63381 10445
rect 63339 10396 63340 10436
rect 63380 10396 63381 10436
rect 63339 10387 63381 10396
rect 70059 10436 70101 10445
rect 70059 10396 70060 10436
rect 70100 10396 70101 10436
rect 70059 10387 70101 10396
rect 70347 10436 70389 10445
rect 70347 10396 70348 10436
rect 70388 10396 70389 10436
rect 70347 10387 70389 10396
rect 75235 10436 75293 10437
rect 75235 10396 75244 10436
rect 75284 10396 75293 10436
rect 75235 10395 75293 10396
rect 1515 10352 1557 10361
rect 1515 10312 1516 10352
rect 1556 10312 1557 10352
rect 1515 10303 1557 10312
rect 43275 10352 43317 10361
rect 43275 10312 43276 10352
rect 43316 10312 43317 10352
rect 43275 10303 43317 10312
rect 54987 10352 55029 10361
rect 54987 10312 54988 10352
rect 55028 10312 55029 10352
rect 54987 10303 55029 10312
rect 55851 10352 55893 10361
rect 55851 10312 55852 10352
rect 55892 10312 55893 10352
rect 55851 10303 55893 10312
rect 58923 10352 58965 10361
rect 58923 10312 58924 10352
rect 58964 10312 58965 10352
rect 58923 10303 58965 10312
rect 67179 10352 67221 10361
rect 67179 10312 67180 10352
rect 67220 10312 67221 10352
rect 67179 10303 67221 10312
rect 71883 10352 71925 10361
rect 71883 10312 71884 10352
rect 71924 10312 71925 10352
rect 71883 10303 71925 10312
rect 77163 10352 77205 10361
rect 77163 10312 77164 10352
rect 77204 10312 77205 10352
rect 77163 10303 77205 10312
rect 78123 10352 78165 10361
rect 78123 10312 78124 10352
rect 78164 10312 78165 10352
rect 78123 10303 78165 10312
rect 43172 10278 43230 10279
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 1699 10268 1757 10269
rect 1699 10228 1708 10268
rect 1748 10228 1757 10268
rect 43172 10238 43181 10278
rect 43221 10238 43230 10278
rect 43172 10237 43230 10238
rect 43371 10268 43413 10277
rect 1699 10227 1757 10228
rect 43371 10228 43372 10268
rect 43412 10228 43413 10268
rect 43371 10219 43413 10228
rect 44515 10268 44573 10269
rect 44515 10228 44524 10268
rect 44564 10228 44573 10268
rect 44515 10227 44573 10228
rect 50755 10268 50813 10269
rect 50755 10228 50764 10268
rect 50804 10228 50813 10268
rect 50755 10227 50813 10228
rect 54891 10268 54933 10277
rect 54891 10228 54892 10268
rect 54932 10228 54933 10268
rect 54891 10219 54933 10228
rect 55083 10268 55125 10277
rect 55083 10228 55084 10268
rect 55124 10228 55125 10268
rect 55083 10219 55125 10228
rect 56227 10268 56285 10269
rect 56227 10228 56236 10268
rect 56276 10228 56285 10268
rect 56227 10227 56285 10228
rect 59779 10268 59837 10269
rect 59779 10228 59788 10268
rect 59828 10228 59837 10268
rect 59779 10227 59837 10228
rect 60163 10268 60221 10269
rect 60163 10228 60172 10268
rect 60212 10228 60221 10268
rect 60163 10227 60221 10228
rect 63051 10268 63093 10277
rect 63051 10228 63052 10268
rect 63092 10228 63093 10268
rect 63051 10219 63093 10228
rect 64675 10268 64733 10269
rect 64675 10228 64684 10268
rect 64724 10228 64733 10268
rect 64675 10227 64733 10228
rect 64971 10268 65013 10277
rect 64971 10228 64972 10268
rect 65012 10228 65013 10268
rect 64971 10219 65013 10228
rect 67083 10268 67125 10277
rect 67083 10228 67084 10268
rect 67124 10228 67125 10268
rect 67083 10219 67125 10228
rect 67275 10268 67317 10277
rect 67275 10228 67276 10268
rect 67316 10228 67317 10268
rect 67275 10219 67317 10228
rect 69475 10268 69533 10269
rect 69475 10228 69484 10268
rect 69524 10228 69533 10268
rect 69475 10227 69533 10228
rect 69859 10268 69917 10269
rect 69859 10228 69868 10268
rect 69908 10228 69917 10268
rect 69859 10227 69917 10228
rect 71787 10268 71829 10277
rect 71787 10228 71788 10268
rect 71828 10228 71829 10268
rect 68419 10226 68477 10227
rect 43075 10184 43133 10185
rect 43075 10144 43084 10184
rect 43124 10144 43133 10184
rect 43075 10143 43133 10144
rect 43467 10184 43509 10193
rect 43467 10144 43468 10184
rect 43508 10144 43509 10184
rect 43467 10135 43509 10144
rect 44139 10184 44181 10193
rect 44139 10144 44140 10184
rect 44180 10144 44181 10184
rect 44139 10135 44181 10144
rect 44227 10184 44285 10185
rect 44227 10144 44236 10184
rect 44276 10144 44285 10184
rect 44227 10143 44285 10144
rect 44907 10184 44949 10193
rect 44907 10144 44908 10184
rect 44948 10144 44949 10184
rect 44907 10135 44949 10144
rect 45003 10184 45045 10193
rect 45003 10144 45004 10184
rect 45044 10144 45045 10184
rect 45003 10135 45045 10144
rect 45099 10184 45141 10193
rect 45099 10144 45100 10184
rect 45140 10144 45141 10184
rect 45099 10135 45141 10144
rect 45763 10184 45821 10185
rect 45763 10144 45772 10184
rect 45812 10144 45821 10184
rect 45763 10143 45821 10144
rect 46627 10184 46685 10185
rect 46627 10144 46636 10184
rect 46676 10144 46685 10184
rect 46627 10143 46685 10144
rect 48355 10184 48413 10185
rect 48355 10144 48364 10184
rect 48404 10144 48413 10184
rect 48355 10143 48413 10144
rect 49219 10184 49277 10185
rect 49219 10144 49228 10184
rect 49268 10144 49277 10184
rect 49219 10143 49277 10144
rect 51147 10184 51189 10193
rect 51147 10144 51148 10184
rect 51188 10144 51189 10184
rect 51147 10135 51189 10144
rect 51339 10184 51381 10193
rect 51339 10144 51340 10184
rect 51380 10144 51381 10184
rect 51339 10135 51381 10144
rect 51427 10184 51485 10185
rect 51427 10144 51436 10184
rect 51476 10144 51485 10184
rect 51427 10143 51485 10144
rect 51723 10184 51765 10193
rect 51723 10144 51724 10184
rect 51764 10144 51765 10184
rect 51723 10135 51765 10144
rect 52099 10184 52157 10185
rect 52099 10144 52108 10184
rect 52148 10144 52157 10184
rect 52099 10143 52157 10144
rect 52963 10184 53021 10185
rect 52963 10144 52972 10184
rect 53012 10144 53021 10184
rect 52963 10143 53021 10144
rect 54795 10184 54837 10193
rect 54795 10144 54796 10184
rect 54836 10144 54837 10184
rect 54795 10135 54837 10144
rect 55171 10184 55229 10185
rect 55171 10144 55180 10184
rect 55220 10144 55229 10184
rect 55171 10143 55229 10144
rect 55459 10184 55517 10185
rect 55459 10144 55468 10184
rect 55508 10144 55517 10184
rect 55459 10143 55517 10144
rect 55563 10184 55605 10193
rect 55563 10144 55564 10184
rect 55604 10144 55605 10184
rect 55563 10135 55605 10144
rect 58243 10184 58301 10185
rect 58243 10144 58252 10184
rect 58292 10144 58301 10184
rect 58243 10143 58301 10144
rect 58443 10184 58485 10193
rect 58443 10144 58444 10184
rect 58484 10144 58485 10184
rect 58443 10135 58485 10144
rect 58635 10184 58677 10193
rect 58635 10144 58636 10184
rect 58676 10144 58677 10184
rect 58635 10135 58677 10144
rect 58723 10184 58781 10185
rect 58723 10144 58732 10184
rect 58772 10144 58781 10184
rect 58723 10143 58781 10144
rect 59211 10184 59253 10193
rect 59211 10144 59212 10184
rect 59252 10144 59253 10184
rect 59211 10135 59253 10144
rect 59299 10184 59357 10185
rect 59299 10144 59308 10184
rect 59348 10144 59357 10184
rect 59299 10143 59357 10144
rect 60651 10184 60693 10193
rect 60651 10144 60652 10184
rect 60692 10144 60693 10184
rect 60651 10135 60693 10144
rect 61027 10184 61085 10185
rect 61027 10144 61036 10184
rect 61076 10144 61085 10184
rect 61027 10143 61085 10144
rect 61891 10184 61949 10185
rect 61891 10144 61900 10184
rect 61940 10144 61949 10184
rect 61891 10143 61949 10144
rect 63235 10184 63293 10185
rect 63235 10144 63244 10184
rect 63284 10144 63293 10184
rect 63235 10143 63293 10144
rect 64867 10184 64925 10185
rect 64867 10144 64876 10184
rect 64916 10144 64925 10184
rect 64867 10143 64925 10144
rect 66987 10184 67029 10193
rect 66987 10144 66988 10184
rect 67028 10144 67029 10184
rect 66987 10135 67029 10144
rect 67363 10184 67421 10185
rect 67363 10144 67372 10184
rect 67412 10144 67421 10184
rect 67363 10143 67421 10144
rect 68235 10184 68277 10193
rect 68235 10144 68236 10184
rect 68276 10144 68277 10184
rect 68235 10135 68277 10144
rect 68331 10184 68373 10193
rect 68419 10186 68428 10226
rect 68468 10186 68477 10226
rect 71787 10219 71829 10228
rect 71979 10268 72021 10277
rect 71979 10228 71980 10268
rect 72020 10228 72021 10268
rect 71979 10219 72021 10228
rect 77067 10268 77109 10277
rect 77067 10228 77068 10268
rect 77108 10228 77109 10268
rect 72067 10226 72125 10227
rect 68419 10185 68477 10186
rect 68331 10144 68332 10184
rect 68372 10144 68373 10184
rect 68331 10135 68373 10144
rect 69099 10184 69141 10193
rect 69099 10144 69100 10184
rect 69140 10144 69141 10184
rect 69099 10135 69141 10144
rect 69195 10184 69237 10193
rect 69195 10144 69196 10184
rect 69236 10144 69237 10184
rect 69195 10135 69237 10144
rect 69291 10184 69333 10193
rect 69291 10144 69292 10184
rect 69332 10144 69333 10184
rect 69291 10135 69333 10144
rect 70243 10184 70301 10185
rect 70243 10144 70252 10184
rect 70292 10144 70301 10184
rect 70243 10143 70301 10144
rect 71691 10184 71733 10193
rect 72067 10186 72076 10226
rect 72116 10186 72125 10226
rect 77067 10219 77109 10228
rect 77259 10268 77301 10277
rect 77259 10228 77260 10268
rect 77300 10228 77301 10268
rect 77259 10219 77301 10228
rect 72067 10185 72125 10186
rect 71691 10144 71692 10184
rect 71732 10144 71733 10184
rect 71691 10135 71733 10144
rect 72267 10184 72309 10193
rect 72267 10144 72268 10184
rect 72308 10144 72309 10184
rect 72267 10135 72309 10144
rect 72459 10184 72501 10193
rect 72459 10144 72460 10184
rect 72500 10144 72501 10184
rect 72459 10135 72501 10144
rect 72547 10184 72605 10185
rect 72547 10144 72556 10184
rect 72596 10144 72605 10184
rect 72547 10143 72605 10144
rect 72843 10184 72885 10193
rect 72843 10144 72844 10184
rect 72884 10144 72885 10184
rect 72843 10135 72885 10144
rect 73219 10184 73277 10185
rect 73219 10144 73228 10184
rect 73268 10144 73277 10184
rect 73219 10143 73277 10144
rect 74083 10184 74141 10185
rect 74083 10144 74092 10184
rect 74132 10144 74141 10184
rect 74083 10143 74141 10144
rect 76587 10184 76629 10193
rect 76587 10144 76588 10184
rect 76628 10144 76629 10184
rect 76587 10135 76629 10144
rect 76683 10184 76725 10193
rect 76683 10144 76684 10184
rect 76724 10144 76725 10184
rect 76683 10135 76725 10144
rect 76779 10184 76821 10193
rect 76779 10144 76780 10184
rect 76820 10144 76821 10184
rect 76779 10135 76821 10144
rect 76971 10184 77013 10193
rect 76971 10144 76972 10184
rect 77012 10144 77013 10184
rect 76971 10135 77013 10144
rect 77347 10184 77405 10185
rect 77347 10144 77356 10184
rect 77396 10144 77405 10184
rect 77347 10143 77405 10144
rect 77643 10184 77685 10193
rect 77643 10144 77644 10184
rect 77684 10144 77685 10184
rect 77643 10135 77685 10144
rect 77739 10184 77781 10193
rect 77739 10144 77740 10184
rect 77780 10144 77781 10184
rect 77739 10135 77781 10144
rect 77835 10184 77877 10193
rect 77835 10144 77836 10184
rect 77876 10144 77877 10184
rect 77835 10135 77877 10144
rect 78019 10184 78077 10185
rect 78019 10144 78028 10184
rect 78068 10144 78077 10184
rect 78019 10143 78077 10144
rect 45195 10100 45237 10109
rect 45195 10060 45196 10100
rect 45236 10060 45237 10100
rect 45195 10051 45237 10060
rect 45387 10100 45429 10109
rect 45387 10060 45388 10100
rect 45428 10060 45429 10100
rect 45387 10051 45429 10060
rect 47979 10100 48021 10109
rect 47979 10060 47980 10100
rect 48020 10060 48021 10100
rect 47979 10051 48021 10060
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 47779 10016 47837 10017
rect 47779 9976 47788 10016
rect 47828 9976 47837 10016
rect 47779 9975 47837 9976
rect 50955 10016 50997 10025
rect 50955 9976 50956 10016
rect 50996 9976 50997 10016
rect 50955 9967 50997 9976
rect 56043 10016 56085 10025
rect 56043 9976 56044 10016
rect 56084 9976 56085 10016
rect 56043 9967 56085 9976
rect 58155 10016 58197 10025
rect 58155 9976 58156 10016
rect 58196 9976 58197 10016
rect 58155 9967 58197 9976
rect 59403 10012 59445 10021
rect 59403 9972 59404 10012
rect 59444 9972 59445 10012
rect 55371 9958 55413 9967
rect 59403 9963 59445 9972
rect 59595 10016 59637 10025
rect 59595 9976 59596 10016
rect 59636 9976 59637 10016
rect 59595 9967 59637 9976
rect 64491 10016 64533 10025
rect 64491 9976 64492 10016
rect 64532 9976 64533 10016
rect 64491 9967 64533 9976
rect 68515 10016 68573 10017
rect 68515 9976 68524 10016
rect 68564 9976 68573 10016
rect 68515 9975 68573 9976
rect 68995 10016 69053 10017
rect 68995 9976 69004 10016
rect 69044 9976 69053 10016
rect 68995 9975 69053 9976
rect 69675 10016 69717 10025
rect 69675 9976 69676 10016
rect 69716 9976 69717 10016
rect 69675 9967 69717 9976
rect 72355 10016 72413 10017
rect 72355 9976 72364 10016
rect 72404 9976 72413 10016
rect 72355 9975 72413 9976
rect 76483 10016 76541 10017
rect 76483 9976 76492 10016
rect 76532 9976 76541 10016
rect 76483 9975 76541 9976
rect 77539 10016 77597 10017
rect 77539 9976 77548 10016
rect 77588 9976 77597 10016
rect 77539 9975 77597 9976
rect 55371 9918 55372 9958
rect 55412 9918 55413 9958
rect 55371 9909 55413 9918
rect 576 9848 79584 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 76352 9848
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76720 9808 79584 9848
rect 576 9784 79584 9808
rect 46347 9684 46389 9693
rect 44995 9680 45053 9681
rect 44995 9640 45004 9680
rect 45044 9640 45053 9680
rect 44995 9639 45053 9640
rect 46347 9644 46348 9684
rect 46388 9644 46389 9684
rect 46347 9635 46389 9644
rect 47115 9680 47157 9689
rect 47115 9640 47116 9680
rect 47156 9640 47157 9680
rect 47115 9631 47157 9640
rect 48067 9680 48125 9681
rect 48067 9640 48076 9680
rect 48116 9640 48125 9680
rect 48067 9639 48125 9640
rect 49707 9680 49749 9689
rect 73035 9684 73077 9693
rect 49707 9640 49708 9680
rect 49748 9640 49749 9680
rect 49707 9631 49749 9640
rect 52291 9680 52349 9681
rect 52291 9640 52300 9680
rect 52340 9640 52349 9680
rect 52291 9639 52349 9640
rect 59491 9680 59549 9681
rect 59491 9640 59500 9680
rect 59540 9640 59549 9680
rect 59491 9639 59549 9640
rect 63523 9680 63581 9681
rect 63523 9640 63532 9680
rect 63572 9640 63581 9680
rect 63523 9639 63581 9640
rect 66403 9680 66461 9681
rect 66403 9640 66412 9680
rect 66452 9640 66461 9680
rect 66403 9639 66461 9640
rect 67555 9680 67613 9681
rect 67555 9640 67564 9680
rect 67604 9640 67613 9680
rect 67555 9639 67613 9640
rect 70627 9680 70685 9681
rect 70627 9640 70636 9680
rect 70676 9640 70685 9680
rect 70627 9639 70685 9640
rect 73035 9644 73036 9684
rect 73076 9644 73077 9684
rect 72643 9638 72701 9639
rect 42603 9596 42645 9605
rect 42603 9556 42604 9596
rect 42644 9556 42645 9596
rect 42603 9547 42645 9556
rect 53451 9596 53493 9605
rect 53451 9556 53452 9596
rect 53492 9556 53493 9596
rect 53451 9547 53493 9556
rect 64011 9596 64053 9605
rect 64011 9556 64012 9596
rect 64052 9556 64053 9596
rect 64011 9547 64053 9556
rect 68235 9596 68277 9605
rect 72643 9598 72652 9638
rect 72692 9598 72701 9638
rect 73035 9635 73077 9644
rect 73419 9680 73461 9689
rect 73419 9640 73420 9680
rect 73460 9640 73461 9680
rect 73419 9631 73461 9640
rect 77731 9680 77789 9681
rect 77731 9640 77740 9680
rect 77780 9640 77789 9680
rect 77731 9639 77789 9640
rect 78019 9680 78077 9681
rect 78019 9640 78028 9680
rect 78068 9640 78077 9680
rect 78019 9639 78077 9640
rect 72643 9597 72701 9598
rect 68235 9556 68236 9596
rect 68276 9556 68277 9596
rect 68235 9547 68277 9556
rect 75339 9596 75381 9605
rect 75339 9556 75340 9596
rect 75380 9556 75381 9596
rect 75339 9547 75381 9556
rect 67934 9523 67976 9532
rect 42979 9512 43037 9513
rect 42979 9472 42988 9512
rect 43028 9472 43037 9512
rect 42979 9471 43037 9472
rect 43843 9512 43901 9513
rect 43843 9472 43852 9512
rect 43892 9472 43901 9512
rect 43843 9471 43901 9472
rect 46155 9512 46197 9521
rect 46155 9472 46156 9512
rect 46196 9472 46197 9512
rect 46155 9463 46197 9472
rect 46243 9512 46301 9513
rect 46243 9472 46252 9512
rect 46292 9472 46301 9512
rect 46243 9471 46301 9472
rect 46539 9512 46581 9521
rect 46539 9472 46540 9512
rect 46580 9472 46581 9512
rect 46539 9463 46581 9472
rect 46635 9512 46677 9521
rect 46635 9472 46636 9512
rect 46676 9472 46677 9512
rect 46635 9463 46677 9472
rect 46731 9512 46773 9521
rect 46731 9472 46732 9512
rect 46772 9472 46773 9512
rect 46731 9463 46773 9472
rect 46827 9512 46869 9521
rect 46827 9472 46828 9512
rect 46868 9472 46869 9512
rect 46827 9463 46869 9472
rect 47203 9512 47261 9513
rect 47203 9472 47212 9512
rect 47252 9472 47261 9512
rect 47203 9471 47261 9472
rect 48171 9512 48213 9521
rect 48171 9472 48172 9512
rect 48212 9472 48213 9512
rect 48171 9463 48213 9472
rect 48267 9512 48309 9521
rect 48267 9472 48268 9512
rect 48308 9472 48309 9512
rect 48267 9463 48309 9472
rect 48363 9512 48405 9521
rect 48363 9472 48364 9512
rect 48404 9472 48405 9512
rect 48363 9463 48405 9472
rect 49315 9512 49373 9513
rect 49315 9472 49324 9512
rect 49364 9472 49373 9512
rect 49315 9471 49373 9472
rect 49899 9512 49941 9521
rect 49899 9472 49900 9512
rect 49940 9472 49941 9512
rect 49899 9463 49941 9472
rect 50275 9512 50333 9513
rect 50275 9472 50284 9512
rect 50324 9472 50333 9512
rect 50275 9471 50333 9472
rect 51139 9512 51197 9513
rect 51139 9472 51148 9512
rect 51188 9472 51197 9512
rect 51139 9471 51197 9472
rect 52483 9512 52541 9513
rect 52483 9472 52492 9512
rect 52532 9472 52541 9512
rect 52483 9471 52541 9472
rect 53827 9512 53885 9513
rect 53827 9472 53836 9512
rect 53876 9472 53885 9512
rect 53827 9471 53885 9472
rect 54691 9512 54749 9513
rect 54691 9472 54700 9512
rect 54740 9472 54749 9512
rect 54691 9471 54749 9472
rect 57099 9512 57141 9521
rect 57099 9472 57100 9512
rect 57140 9472 57141 9512
rect 57099 9463 57141 9472
rect 57475 9512 57533 9513
rect 57475 9472 57484 9512
rect 57524 9472 57533 9512
rect 57475 9471 57533 9472
rect 58339 9512 58397 9513
rect 58339 9472 58348 9512
rect 58388 9472 58397 9512
rect 58339 9471 58397 9472
rect 62667 9512 62709 9521
rect 62667 9472 62668 9512
rect 62708 9472 62709 9512
rect 62667 9463 62709 9472
rect 62859 9512 62901 9521
rect 62859 9472 62860 9512
rect 62900 9472 62901 9512
rect 62859 9463 62901 9472
rect 62947 9512 63005 9513
rect 62947 9472 62956 9512
rect 62996 9472 63005 9512
rect 62947 9471 63005 9472
rect 63627 9512 63669 9521
rect 63627 9472 63628 9512
rect 63668 9472 63669 9512
rect 63627 9463 63669 9472
rect 63723 9512 63765 9521
rect 63723 9472 63724 9512
rect 63764 9472 63765 9512
rect 63723 9463 63765 9472
rect 63819 9512 63861 9521
rect 63819 9472 63820 9512
rect 63860 9472 63861 9512
rect 63819 9463 63861 9472
rect 64387 9512 64445 9513
rect 64387 9472 64396 9512
rect 64436 9472 64445 9512
rect 64387 9471 64445 9472
rect 65251 9512 65309 9513
rect 65251 9472 65260 9512
rect 65300 9472 65309 9512
rect 65251 9471 65309 9472
rect 67467 9512 67509 9521
rect 67467 9472 67468 9512
rect 67508 9472 67509 9512
rect 67467 9463 67509 9472
rect 67659 9512 67701 9521
rect 67659 9472 67660 9512
rect 67700 9472 67701 9512
rect 67659 9463 67701 9472
rect 67747 9512 67805 9513
rect 67747 9472 67756 9512
rect 67796 9472 67805 9512
rect 67934 9483 67935 9523
rect 67975 9483 67976 9523
rect 67934 9474 67976 9483
rect 68611 9512 68669 9513
rect 67747 9471 67805 9472
rect 68611 9472 68620 9512
rect 68660 9472 68669 9512
rect 68611 9471 68669 9472
rect 69475 9512 69533 9513
rect 69475 9472 69484 9512
rect 69524 9472 69533 9512
rect 69475 9471 69533 9472
rect 71979 9512 72021 9521
rect 71979 9472 71980 9512
rect 72020 9472 72021 9512
rect 71979 9463 72021 9472
rect 72355 9512 72413 9513
rect 72355 9472 72364 9512
rect 72404 9472 72413 9512
rect 72355 9471 72413 9472
rect 72843 9512 72885 9521
rect 72843 9472 72844 9512
rect 72884 9472 72885 9512
rect 72843 9463 72885 9472
rect 72931 9512 72989 9513
rect 72931 9472 72940 9512
rect 72980 9472 72989 9512
rect 72931 9471 72989 9472
rect 73611 9512 73653 9521
rect 73611 9472 73612 9512
rect 73652 9472 73653 9512
rect 73611 9463 73653 9472
rect 73707 9512 73749 9521
rect 73707 9472 73708 9512
rect 73748 9472 73749 9512
rect 73707 9463 73749 9472
rect 73803 9512 73845 9521
rect 73803 9472 73804 9512
rect 73844 9472 73845 9512
rect 73803 9463 73845 9472
rect 73899 9512 73941 9521
rect 73899 9472 73900 9512
rect 73940 9472 73941 9512
rect 73899 9463 73941 9472
rect 75715 9512 75773 9513
rect 75715 9472 75724 9512
rect 75764 9472 75773 9512
rect 75715 9471 75773 9472
rect 76579 9512 76637 9513
rect 76579 9472 76588 9512
rect 76628 9472 76637 9512
rect 76579 9471 76637 9472
rect 77931 9512 77973 9521
rect 77931 9472 77932 9512
rect 77972 9472 77973 9512
rect 77931 9463 77973 9472
rect 78123 9512 78165 9521
rect 78123 9472 78124 9512
rect 78164 9472 78165 9512
rect 78123 9463 78165 9472
rect 78211 9512 78269 9513
rect 78211 9472 78220 9512
rect 78260 9472 78269 9512
rect 78211 9471 78269 9472
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 45475 9428 45533 9429
rect 45475 9388 45484 9428
rect 45524 9388 45533 9428
rect 45475 9387 45533 9388
rect 49507 9428 49565 9429
rect 49507 9388 49516 9428
rect 49556 9388 49565 9428
rect 49507 9387 49565 9388
rect 56131 9428 56189 9429
rect 56131 9388 56140 9428
rect 56180 9388 56189 9428
rect 56131 9387 56189 9388
rect 60259 9428 60317 9429
rect 60259 9388 60268 9428
rect 60308 9388 60317 9428
rect 60259 9387 60317 9388
rect 61123 9428 61181 9429
rect 61123 9388 61132 9428
rect 61172 9388 61181 9428
rect 61123 9387 61181 9388
rect 63139 9428 63197 9429
rect 63139 9388 63148 9428
rect 63188 9388 63197 9428
rect 63139 9387 63197 9388
rect 72075 9428 72117 9437
rect 72075 9388 72076 9428
rect 72116 9388 72117 9428
rect 72075 9379 72117 9388
rect 72267 9428 72309 9437
rect 72267 9388 72268 9428
rect 72308 9388 72309 9428
rect 72267 9379 72309 9388
rect 73219 9428 73277 9429
rect 73219 9388 73228 9428
rect 73268 9388 73277 9428
rect 73219 9387 73277 9388
rect 78595 9428 78653 9429
rect 78595 9388 78604 9428
rect 78644 9388 78653 9428
rect 78595 9387 78653 9388
rect 45291 9344 45333 9353
rect 45291 9304 45292 9344
rect 45332 9304 45333 9344
rect 45291 9295 45333 9304
rect 45867 9344 45909 9353
rect 45867 9304 45868 9344
rect 45908 9304 45909 9344
rect 45867 9295 45909 9304
rect 63339 9344 63381 9353
rect 63339 9304 63340 9344
rect 63380 9304 63381 9344
rect 63339 9295 63381 9304
rect 72171 9344 72213 9353
rect 72171 9304 72172 9344
rect 72212 9304 72213 9344
rect 72171 9295 72213 9304
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 49227 9260 49269 9269
rect 49227 9220 49228 9260
rect 49268 9220 49269 9260
rect 49227 9211 49269 9220
rect 52587 9260 52629 9269
rect 52587 9220 52588 9260
rect 52628 9220 52629 9260
rect 52587 9211 52629 9220
rect 55843 9260 55901 9261
rect 55843 9220 55852 9260
rect 55892 9220 55901 9260
rect 55843 9219 55901 9220
rect 56331 9260 56373 9269
rect 56331 9220 56332 9260
rect 56372 9220 56373 9260
rect 56331 9211 56373 9220
rect 60075 9260 60117 9269
rect 60075 9220 60076 9260
rect 60116 9220 60117 9260
rect 60075 9211 60117 9220
rect 61323 9260 61365 9269
rect 61323 9220 61324 9260
rect 61364 9220 61365 9260
rect 61323 9211 61365 9220
rect 62667 9260 62709 9269
rect 62667 9220 62668 9260
rect 62708 9220 62709 9260
rect 62667 9211 62709 9220
rect 68043 9260 68085 9269
rect 68043 9220 68044 9260
rect 68084 9220 68085 9260
rect 68043 9211 68085 9220
rect 73419 9260 73461 9269
rect 73419 9220 73420 9260
rect 73460 9220 73461 9260
rect 73419 9211 73461 9220
rect 78411 9260 78453 9269
rect 78411 9220 78412 9260
rect 78452 9220 78453 9260
rect 78411 9211 78453 9220
rect 576 9092 79584 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 75112 9092
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75480 9052 79584 9092
rect 576 9028 79584 9052
rect 45099 8924 45141 8933
rect 45099 8884 45100 8924
rect 45140 8884 45141 8924
rect 45099 8875 45141 8884
rect 50283 8924 50325 8933
rect 50283 8884 50284 8924
rect 50324 8884 50325 8924
rect 50283 8875 50325 8884
rect 51243 8924 51285 8933
rect 51243 8884 51244 8924
rect 51284 8884 51285 8924
rect 51243 8875 51285 8884
rect 55371 8924 55413 8933
rect 55371 8884 55372 8924
rect 55412 8884 55413 8924
rect 55371 8875 55413 8884
rect 58051 8924 58109 8925
rect 58051 8884 58060 8924
rect 58100 8884 58109 8924
rect 58051 8883 58109 8884
rect 62179 8924 62237 8925
rect 62179 8884 62188 8924
rect 62228 8884 62237 8924
rect 62179 8883 62237 8884
rect 65923 8924 65981 8925
rect 65923 8884 65932 8924
rect 65972 8884 65981 8924
rect 65923 8883 65981 8884
rect 68523 8924 68565 8933
rect 68523 8884 68524 8924
rect 68564 8884 68565 8924
rect 68523 8875 68565 8884
rect 72939 8924 72981 8933
rect 72939 8884 72940 8924
rect 72980 8884 72981 8924
rect 72939 8875 72981 8884
rect 74571 8924 74613 8933
rect 74571 8884 74572 8924
rect 74612 8884 74613 8924
rect 74571 8875 74613 8884
rect 44427 8840 44469 8849
rect 44427 8800 44428 8840
rect 44468 8800 44469 8840
rect 44427 8791 44469 8800
rect 45483 8840 45525 8849
rect 45483 8800 45484 8840
rect 45524 8800 45525 8840
rect 45483 8791 45525 8800
rect 48363 8840 48405 8849
rect 48363 8800 48364 8840
rect 48404 8800 48405 8840
rect 48363 8791 48405 8800
rect 50667 8840 50709 8849
rect 50667 8800 50668 8840
rect 50708 8800 50709 8840
rect 50667 8791 50709 8800
rect 52299 8840 52341 8849
rect 52299 8800 52300 8840
rect 52340 8800 52341 8840
rect 52299 8791 52341 8800
rect 58731 8840 58773 8849
rect 58731 8800 58732 8840
rect 58772 8800 58773 8840
rect 58731 8791 58773 8800
rect 59115 8840 59157 8849
rect 59115 8800 59116 8840
rect 59156 8800 59157 8840
rect 59115 8791 59157 8800
rect 63051 8840 63093 8849
rect 63051 8800 63052 8840
rect 63092 8800 63093 8840
rect 63051 8791 63093 8800
rect 63531 8840 63573 8849
rect 63531 8800 63532 8840
rect 63572 8800 63573 8840
rect 63531 8791 63573 8800
rect 74187 8840 74229 8849
rect 74187 8800 74188 8840
rect 74228 8800 74229 8840
rect 74187 8791 74229 8800
rect 76491 8840 76533 8849
rect 76491 8800 76492 8840
rect 76532 8800 76533 8840
rect 76491 8791 76533 8800
rect 73987 8767 74045 8768
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 44611 8756 44669 8757
rect 44611 8716 44620 8756
rect 44660 8716 44669 8756
rect 44611 8715 44669 8716
rect 45387 8756 45429 8765
rect 45387 8716 45388 8756
rect 45428 8716 45429 8756
rect 45387 8707 45429 8716
rect 45579 8756 45621 8765
rect 45579 8716 45580 8756
rect 45620 8716 45621 8756
rect 45579 8707 45621 8716
rect 49699 8756 49757 8757
rect 49699 8716 49708 8756
rect 49748 8716 49757 8756
rect 49699 8715 49757 8716
rect 50083 8756 50141 8757
rect 50083 8716 50092 8756
rect 50132 8716 50141 8756
rect 50083 8715 50141 8716
rect 50571 8756 50613 8765
rect 50571 8716 50572 8756
rect 50612 8716 50613 8756
rect 50571 8707 50613 8716
rect 50763 8756 50805 8765
rect 50763 8716 50764 8756
rect 50804 8716 50805 8756
rect 50763 8707 50805 8716
rect 58635 8756 58677 8765
rect 58635 8716 58636 8756
rect 58676 8716 58677 8756
rect 58635 8707 58677 8716
rect 58827 8756 58869 8765
rect 58827 8716 58828 8756
rect 58868 8716 58869 8756
rect 58827 8707 58869 8716
rect 62955 8756 62997 8765
rect 62955 8716 62956 8756
rect 62996 8716 62997 8756
rect 62955 8707 62997 8716
rect 63147 8756 63189 8765
rect 63147 8716 63148 8756
rect 63188 8716 63189 8756
rect 63147 8707 63189 8716
rect 69379 8756 69437 8757
rect 69379 8716 69388 8756
rect 69428 8716 69437 8756
rect 69379 8715 69437 8716
rect 69675 8756 69717 8765
rect 69675 8716 69676 8756
rect 69716 8716 69717 8756
rect 73987 8727 73996 8767
rect 74036 8727 74045 8767
rect 73987 8726 74045 8727
rect 76395 8756 76437 8765
rect 69675 8707 69717 8716
rect 76395 8716 76396 8756
rect 76436 8716 76437 8756
rect 76395 8707 76437 8716
rect 76587 8756 76629 8765
rect 76587 8716 76588 8756
rect 76628 8716 76629 8756
rect 76587 8707 76629 8716
rect 79275 8756 79317 8765
rect 79275 8716 79276 8756
rect 79316 8716 79317 8756
rect 79275 8707 79317 8716
rect 44803 8672 44861 8673
rect 44803 8632 44812 8672
rect 44852 8632 44861 8672
rect 44803 8631 44861 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 45099 8672 45141 8681
rect 45099 8632 45100 8672
rect 45140 8632 45141 8672
rect 45667 8672 45725 8673
rect 45099 8623 45141 8632
rect 45291 8630 45333 8639
rect 45667 8632 45676 8672
rect 45716 8632 45725 8672
rect 45667 8631 45725 8632
rect 47491 8672 47549 8673
rect 47491 8632 47500 8672
rect 47540 8632 47549 8672
rect 47491 8631 47549 8632
rect 47595 8672 47637 8681
rect 47595 8632 47596 8672
rect 47636 8632 47637 8672
rect 45291 8590 45292 8630
rect 45332 8590 45333 8630
rect 47595 8623 47637 8632
rect 47787 8672 47829 8681
rect 47787 8632 47788 8672
rect 47828 8632 47829 8672
rect 47787 8623 47829 8632
rect 48651 8672 48693 8681
rect 48651 8632 48652 8672
rect 48692 8632 48693 8672
rect 48651 8623 48693 8632
rect 48739 8672 48797 8673
rect 48739 8632 48748 8672
rect 48788 8632 48797 8672
rect 48739 8631 48797 8632
rect 49131 8672 49173 8681
rect 49131 8632 49132 8672
rect 49172 8632 49173 8672
rect 49131 8623 49173 8632
rect 49227 8672 49269 8681
rect 49227 8632 49228 8672
rect 49268 8632 49269 8672
rect 49227 8623 49269 8632
rect 49323 8672 49365 8681
rect 49323 8632 49324 8672
rect 49364 8632 49365 8672
rect 49323 8623 49365 8632
rect 50475 8672 50517 8681
rect 50475 8632 50476 8672
rect 50516 8632 50517 8672
rect 50475 8623 50517 8632
rect 50851 8672 50909 8673
rect 50851 8632 50860 8672
rect 50900 8632 50909 8672
rect 50851 8631 50909 8632
rect 51531 8672 51573 8681
rect 51531 8632 51532 8672
rect 51572 8632 51573 8672
rect 51531 8623 51573 8632
rect 51619 8672 51677 8673
rect 51619 8632 51628 8672
rect 51668 8632 51677 8672
rect 51619 8631 51677 8632
rect 52003 8672 52061 8673
rect 52003 8632 52012 8672
rect 52052 8632 52061 8672
rect 52003 8631 52061 8632
rect 52963 8672 53021 8673
rect 52963 8632 52972 8672
rect 53012 8632 53021 8672
rect 52963 8631 53021 8632
rect 53155 8672 53213 8673
rect 53155 8632 53164 8672
rect 53204 8632 53213 8672
rect 53155 8631 53213 8632
rect 54891 8672 54933 8681
rect 54891 8632 54892 8672
rect 54932 8632 54933 8672
rect 54891 8623 54933 8632
rect 55083 8672 55125 8681
rect 55083 8632 55084 8672
rect 55124 8632 55125 8672
rect 55083 8623 55125 8632
rect 55171 8672 55229 8673
rect 55171 8632 55180 8672
rect 55220 8632 55229 8672
rect 55171 8631 55229 8632
rect 55459 8672 55517 8673
rect 55459 8632 55468 8672
rect 55508 8632 55517 8672
rect 55459 8631 55517 8632
rect 56035 8672 56093 8673
rect 56035 8632 56044 8672
rect 56084 8632 56093 8672
rect 56035 8631 56093 8632
rect 56899 8672 56957 8673
rect 56899 8632 56908 8672
rect 56948 8632 56957 8672
rect 56899 8631 56957 8632
rect 58539 8672 58581 8681
rect 58539 8632 58540 8672
rect 58580 8632 58581 8672
rect 58539 8623 58581 8632
rect 58915 8672 58973 8673
rect 58915 8632 58924 8672
rect 58964 8632 58973 8672
rect 58915 8631 58973 8632
rect 59115 8672 59157 8681
rect 59115 8632 59116 8672
rect 59156 8632 59157 8672
rect 59115 8623 59157 8632
rect 59307 8672 59349 8681
rect 59307 8632 59308 8672
rect 59348 8632 59349 8672
rect 59307 8623 59349 8632
rect 59395 8672 59453 8673
rect 59395 8632 59404 8672
rect 59444 8632 59453 8672
rect 59395 8631 59453 8632
rect 60163 8672 60221 8673
rect 60163 8632 60172 8672
rect 60212 8632 60221 8672
rect 60163 8631 60221 8632
rect 61027 8672 61085 8673
rect 61027 8632 61036 8672
rect 61076 8632 61085 8672
rect 61027 8631 61085 8632
rect 62859 8672 62901 8681
rect 62859 8632 62860 8672
rect 62900 8632 62901 8672
rect 62859 8623 62901 8632
rect 63235 8672 63293 8673
rect 63235 8632 63244 8672
rect 63284 8632 63293 8672
rect 63235 8631 63293 8632
rect 63819 8672 63861 8681
rect 63819 8632 63820 8672
rect 63860 8632 63861 8672
rect 64203 8672 64245 8681
rect 63819 8623 63861 8632
rect 63907 8662 63965 8663
rect 63907 8622 63916 8662
rect 63956 8622 63965 8662
rect 64203 8632 64204 8672
rect 64244 8632 64245 8672
rect 64203 8623 64245 8632
rect 64299 8672 64341 8681
rect 64299 8632 64300 8672
rect 64340 8632 64341 8672
rect 64299 8623 64341 8632
rect 64395 8672 64437 8681
rect 64395 8632 64396 8672
rect 64436 8632 64437 8672
rect 64395 8623 64437 8632
rect 64491 8672 64533 8681
rect 64491 8632 64492 8672
rect 64532 8632 64533 8672
rect 64491 8623 64533 8632
rect 67075 8672 67133 8673
rect 67075 8632 67084 8672
rect 67124 8632 67133 8672
rect 67075 8631 67133 8632
rect 67939 8672 67997 8673
rect 67939 8632 67948 8672
rect 67988 8632 67997 8672
rect 67939 8631 67997 8632
rect 68811 8672 68853 8681
rect 68811 8632 68812 8672
rect 68852 8632 68853 8672
rect 68811 8623 68853 8632
rect 68899 8672 68957 8673
rect 68899 8632 68908 8672
rect 68948 8632 68957 8672
rect 68899 8631 68957 8632
rect 70819 8672 70877 8673
rect 70819 8632 70828 8672
rect 70868 8632 70877 8672
rect 70819 8631 70877 8632
rect 71683 8672 71741 8673
rect 71683 8632 71692 8672
rect 71732 8632 71741 8672
rect 71683 8631 71741 8632
rect 72075 8672 72117 8681
rect 72075 8632 72076 8672
rect 72116 8632 72117 8672
rect 72075 8623 72117 8632
rect 72459 8672 72501 8681
rect 72459 8632 72460 8672
rect 72500 8632 72501 8672
rect 72459 8623 72501 8632
rect 72555 8672 72597 8681
rect 72555 8632 72556 8672
rect 72596 8632 72597 8672
rect 72555 8623 72597 8632
rect 72651 8672 72693 8681
rect 72651 8632 72652 8672
rect 72692 8632 72693 8672
rect 72651 8623 72693 8632
rect 72835 8672 72893 8673
rect 72835 8632 72844 8672
rect 72884 8632 72893 8672
rect 72835 8631 72893 8632
rect 74467 8672 74525 8673
rect 74467 8632 74476 8672
rect 74516 8632 74525 8672
rect 74467 8631 74525 8632
rect 76299 8672 76341 8681
rect 76299 8632 76300 8672
rect 76340 8632 76341 8672
rect 76299 8623 76341 8632
rect 76675 8672 76733 8673
rect 76675 8632 76684 8672
rect 76724 8632 76733 8672
rect 76675 8631 76733 8632
rect 76875 8672 76917 8681
rect 76875 8632 76876 8672
rect 76916 8632 76917 8672
rect 76875 8623 76917 8632
rect 77251 8672 77309 8673
rect 77251 8632 77260 8672
rect 77300 8632 77309 8672
rect 77251 8631 77309 8632
rect 78115 8672 78173 8673
rect 78115 8632 78124 8672
rect 78164 8632 78173 8672
rect 78115 8631 78173 8632
rect 63907 8621 63965 8622
rect 45291 8581 45333 8590
rect 55659 8588 55701 8597
rect 55659 8548 55660 8588
rect 55700 8548 55701 8588
rect 55659 8539 55701 8548
rect 59787 8588 59829 8597
rect 59787 8548 59788 8588
rect 59828 8548 59829 8588
rect 59787 8539 59829 8548
rect 68331 8588 68373 8597
rect 68331 8548 68332 8588
rect 68372 8548 68373 8588
rect 68331 8539 68373 8548
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 47683 8504 47741 8505
rect 47683 8464 47692 8504
rect 47732 8464 47741 8504
rect 47683 8463 47741 8464
rect 48843 8500 48885 8509
rect 48843 8460 48844 8500
rect 48884 8460 48885 8500
rect 49027 8504 49085 8505
rect 49027 8464 49036 8504
rect 49076 8464 49085 8504
rect 49027 8463 49085 8464
rect 49899 8504 49941 8513
rect 49899 8464 49900 8504
rect 49940 8464 49941 8504
rect 48843 8451 48885 8460
rect 49899 8455 49941 8464
rect 54979 8504 55037 8505
rect 54979 8464 54988 8504
rect 55028 8464 55037 8504
rect 54979 8463 55037 8464
rect 69195 8504 69237 8513
rect 69195 8464 69196 8504
rect 69236 8464 69237 8504
rect 69195 8455 69237 8464
rect 72355 8504 72413 8505
rect 72355 8464 72364 8504
rect 72404 8464 72413 8504
rect 72355 8463 72413 8464
rect 51723 8446 51765 8455
rect 51723 8406 51724 8446
rect 51764 8406 51765 8446
rect 51723 8397 51765 8406
rect 64011 8446 64053 8455
rect 64011 8406 64012 8446
rect 64052 8406 64053 8446
rect 64011 8397 64053 8406
rect 69003 8446 69045 8455
rect 69003 8406 69004 8446
rect 69044 8406 69045 8446
rect 69003 8397 69045 8406
rect 576 8336 79584 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 76352 8336
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76720 8296 79584 8336
rect 576 8272 79584 8296
rect 77451 8226 77493 8235
rect 71979 8199 72021 8208
rect 47587 8168 47645 8169
rect 47587 8128 47596 8168
rect 47636 8128 47645 8168
rect 47587 8127 47645 8128
rect 50275 8168 50333 8169
rect 50275 8128 50284 8168
rect 50324 8128 50333 8168
rect 50275 8127 50333 8128
rect 53355 8168 53397 8177
rect 53355 8128 53356 8168
rect 53396 8128 53397 8168
rect 53355 8119 53397 8128
rect 54699 8172 54741 8181
rect 54699 8132 54700 8172
rect 54740 8132 54741 8172
rect 54699 8123 54741 8132
rect 55363 8168 55421 8169
rect 55363 8128 55372 8168
rect 55412 8128 55421 8168
rect 55363 8127 55421 8128
rect 58347 8168 58389 8177
rect 58347 8128 58348 8168
rect 58388 8128 58389 8168
rect 58347 8119 58389 8128
rect 59019 8168 59061 8177
rect 59019 8128 59020 8168
rect 59060 8128 59061 8168
rect 59019 8119 59061 8128
rect 59403 8172 59445 8181
rect 59403 8132 59404 8172
rect 59444 8132 59445 8172
rect 59403 8123 59445 8132
rect 60067 8168 60125 8169
rect 60067 8128 60076 8168
rect 60116 8128 60125 8168
rect 60067 8127 60125 8128
rect 66211 8168 66269 8169
rect 66211 8128 66220 8168
rect 66260 8128 66269 8168
rect 66211 8127 66269 8128
rect 66699 8168 66741 8177
rect 66699 8128 66700 8168
rect 66740 8128 66741 8168
rect 71979 8159 71980 8199
rect 72020 8159 72021 8199
rect 77451 8186 77452 8226
rect 77492 8186 77493 8226
rect 77451 8177 77493 8186
rect 71979 8150 72021 8159
rect 75043 8168 75101 8169
rect 66699 8119 66741 8128
rect 75043 8128 75052 8168
rect 75092 8128 75101 8168
rect 75043 8127 75101 8128
rect 77835 8168 77877 8177
rect 77835 8128 77836 8168
rect 77876 8128 77877 8168
rect 77835 8119 77877 8128
rect 78027 8168 78069 8177
rect 78027 8128 78028 8168
rect 78068 8128 78069 8168
rect 78027 8119 78069 8128
rect 45195 8084 45237 8093
rect 45195 8044 45196 8084
rect 45236 8044 45237 8084
rect 45195 8035 45237 8044
rect 62187 8084 62229 8093
rect 62187 8044 62188 8084
rect 62228 8044 62229 8084
rect 62187 8035 62229 8044
rect 72651 8084 72693 8093
rect 72651 8044 72652 8084
rect 72692 8044 72693 8084
rect 72651 8035 72693 8044
rect 45571 8000 45629 8001
rect 45571 7960 45580 8000
rect 45620 7960 45629 8000
rect 45571 7959 45629 7960
rect 46435 8000 46493 8001
rect 46435 7960 46444 8000
rect 46484 7960 46493 8000
rect 46435 7959 46493 7960
rect 47883 8000 47925 8009
rect 47883 7960 47884 8000
rect 47924 7960 47925 8000
rect 47883 7951 47925 7960
rect 48259 8000 48317 8001
rect 48259 7960 48268 8000
rect 48308 7960 48317 8000
rect 48259 7959 48317 7960
rect 49123 8000 49181 8001
rect 49123 7960 49132 8000
rect 49172 7960 49181 8000
rect 49123 7959 49181 7960
rect 50667 8000 50709 8009
rect 50667 7960 50668 8000
rect 50708 7960 50709 8000
rect 50667 7951 50709 7960
rect 51043 8000 51101 8001
rect 51043 7960 51052 8000
rect 51092 7960 51101 8000
rect 51043 7959 51101 7960
rect 51907 8000 51965 8001
rect 51907 7960 51916 8000
rect 51956 7960 51965 8000
rect 51907 7959 51965 7960
rect 53443 8000 53501 8001
rect 53443 7960 53452 8000
rect 53492 7960 53501 8000
rect 53443 7959 53501 7960
rect 53827 8000 53885 8001
rect 53827 7960 53836 8000
rect 53876 7960 53885 8000
rect 53827 7959 53885 7960
rect 53931 8000 53973 8009
rect 53931 7960 53932 8000
rect 53972 7960 53973 8000
rect 53931 7951 53973 7960
rect 54115 8000 54173 8001
rect 54115 7960 54124 8000
rect 54164 7960 54173 8000
rect 54115 7959 54173 7960
rect 54507 8000 54549 8009
rect 54507 7960 54508 8000
rect 54548 7960 54549 8000
rect 54507 7951 54549 7960
rect 54787 8000 54845 8001
rect 54787 7960 54796 8000
rect 54836 7960 54845 8000
rect 54787 7959 54845 7960
rect 54891 8000 54933 8009
rect 54891 7960 54892 8000
rect 54932 7960 54933 8000
rect 54891 7951 54933 7960
rect 55467 8000 55509 8009
rect 55467 7960 55468 8000
rect 55508 7960 55509 8000
rect 55467 7951 55509 7960
rect 55563 8000 55605 8009
rect 55563 7960 55564 8000
rect 55604 7960 55605 8000
rect 55563 7951 55605 7960
rect 55659 8000 55701 8009
rect 55659 7960 55660 8000
rect 55700 7960 55701 8000
rect 55659 7951 55701 7960
rect 55851 8000 55893 8009
rect 55851 7960 55852 8000
rect 55892 7960 55893 8000
rect 55851 7951 55893 7960
rect 55947 8000 55989 8009
rect 55947 7960 55948 8000
rect 55988 7960 55989 8000
rect 55947 7951 55989 7960
rect 56043 8000 56085 8009
rect 56043 7960 56044 8000
rect 56084 7960 56085 8000
rect 56043 7951 56085 7960
rect 56139 8000 56181 8009
rect 56139 7960 56140 8000
rect 56180 7960 56181 8000
rect 56139 7951 56181 7960
rect 58435 8000 58493 8001
rect 58435 7960 58444 8000
rect 58484 7960 58493 8000
rect 58435 7959 58493 7960
rect 59491 8000 59549 8001
rect 59491 7960 59500 8000
rect 59540 7960 59549 8000
rect 59491 7959 59549 7960
rect 59595 8000 59637 8009
rect 59595 7960 59596 8000
rect 59636 7960 59637 8000
rect 59595 7951 59637 7960
rect 60171 8000 60213 8009
rect 60171 7960 60172 8000
rect 60212 7960 60213 8000
rect 60171 7951 60213 7960
rect 60267 8000 60309 8009
rect 60267 7960 60268 8000
rect 60308 7960 60309 8000
rect 60267 7951 60309 7960
rect 60363 8000 60405 8009
rect 60363 7960 60364 8000
rect 60404 7960 60405 8000
rect 60363 7951 60405 7960
rect 60555 8000 60597 8009
rect 60555 7960 60556 8000
rect 60596 7960 60597 8000
rect 60555 7951 60597 7960
rect 60651 8000 60693 8009
rect 60651 7960 60652 8000
rect 60692 7960 60693 8000
rect 60651 7951 60693 7960
rect 60747 8000 60789 8009
rect 60747 7960 60748 8000
rect 60788 7960 60789 8000
rect 60747 7951 60789 7960
rect 60843 8000 60885 8009
rect 60843 7960 60844 8000
rect 60884 7960 60885 8000
rect 60843 7951 60885 7960
rect 62563 8000 62621 8001
rect 62563 7960 62572 8000
rect 62612 7960 62621 8000
rect 62563 7959 62621 7960
rect 63427 8000 63485 8001
rect 63427 7960 63436 8000
rect 63476 7960 63485 8000
rect 63427 7959 63485 7960
rect 65739 8000 65781 8009
rect 65739 7960 65740 8000
rect 65780 7960 65781 8000
rect 65739 7951 65781 7960
rect 65835 8000 65877 8009
rect 65835 7960 65836 8000
rect 65876 7960 65877 8000
rect 65835 7951 65877 7960
rect 65931 8000 65973 8009
rect 65931 7960 65932 8000
rect 65972 7960 65973 8000
rect 65931 7951 65973 7960
rect 66027 8000 66069 8009
rect 66027 7960 66028 8000
rect 66068 7960 66069 8000
rect 66027 7951 66069 7960
rect 66411 8000 66453 8009
rect 66411 7960 66412 8000
rect 66452 7960 66453 8000
rect 66307 7958 66365 7959
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 53067 7916 53109 7925
rect 53067 7876 53068 7916
rect 53108 7876 53109 7916
rect 53067 7867 53109 7876
rect 54219 7916 54261 7925
rect 54219 7876 54220 7916
rect 54260 7876 54261 7916
rect 54219 7867 54261 7876
rect 54411 7916 54453 7925
rect 66307 7918 66316 7958
rect 66356 7918 66365 7958
rect 66411 7951 66453 7960
rect 66507 8000 66549 8009
rect 66507 7960 66508 8000
rect 66548 7960 66549 8000
rect 66507 7951 66549 7960
rect 66787 8000 66845 8001
rect 66787 7960 66796 8000
rect 66836 7960 66845 8000
rect 66787 7959 66845 7960
rect 67939 8000 67997 8001
rect 67939 7960 67948 8000
rect 67988 7960 67997 8000
rect 67939 7959 67997 7960
rect 68331 8000 68373 8009
rect 68331 7960 68332 8000
rect 68372 7960 68373 8000
rect 68331 7951 68373 7960
rect 71499 8000 71541 8009
rect 71499 7960 71500 8000
rect 71540 7960 71541 8000
rect 71499 7951 71541 7960
rect 71691 8000 71733 8009
rect 71691 7960 71692 8000
rect 71732 7960 71733 8000
rect 71691 7951 71733 7960
rect 71779 8000 71837 8001
rect 71779 7960 71788 8000
rect 71828 7960 71837 8000
rect 71779 7959 71837 7960
rect 72067 8000 72125 8001
rect 72067 7960 72076 8000
rect 72116 7960 72125 8000
rect 72067 7959 72125 7960
rect 72171 8000 72213 8009
rect 72171 7960 72172 8000
rect 72212 7960 72213 8000
rect 72171 7951 72213 7960
rect 73027 8000 73085 8001
rect 73027 7960 73036 8000
rect 73076 7960 73085 8000
rect 73027 7959 73085 7960
rect 73891 8000 73949 8001
rect 73891 7960 73900 8000
rect 73940 7960 73949 8000
rect 73891 7959 73949 7960
rect 76491 8000 76533 8009
rect 76491 7960 76492 8000
rect 76532 7960 76533 8000
rect 76491 7951 76533 7960
rect 76587 8000 76629 8009
rect 76587 7960 76588 8000
rect 76628 7960 76629 8000
rect 76587 7951 76629 7960
rect 76683 8000 76725 8009
rect 76683 7960 76684 8000
rect 76724 7960 76725 8000
rect 76683 7951 76725 7960
rect 76779 8000 76821 8009
rect 76779 7960 76780 8000
rect 76820 7960 76821 8000
rect 76779 7951 76821 7960
rect 77259 8000 77301 8009
rect 77259 7960 77260 8000
rect 77300 7960 77301 8000
rect 77259 7951 77301 7960
rect 77347 8000 77405 8001
rect 77347 7960 77356 8000
rect 77396 7960 77405 8000
rect 77347 7959 77405 7960
rect 78115 8000 78173 8001
rect 78115 7960 78124 8000
rect 78164 7960 78173 8000
rect 78115 7959 78173 7960
rect 66307 7917 66365 7918
rect 54411 7876 54412 7916
rect 54452 7876 54453 7916
rect 54411 7867 54453 7876
rect 58627 7916 58685 7917
rect 58627 7876 58636 7916
rect 58676 7876 58685 7916
rect 58627 7875 58685 7876
rect 59203 7916 59261 7917
rect 59203 7876 59212 7916
rect 59252 7876 59261 7916
rect 59203 7875 59261 7876
rect 64963 7916 65021 7917
rect 64963 7876 64972 7916
rect 65012 7876 65021 7916
rect 64963 7875 65021 7876
rect 68043 7916 68085 7925
rect 68043 7876 68044 7916
rect 68084 7876 68085 7916
rect 68043 7867 68085 7876
rect 68235 7916 68277 7925
rect 68235 7876 68236 7916
rect 68276 7876 68277 7916
rect 68235 7867 68277 7876
rect 68899 7916 68957 7917
rect 68899 7876 68908 7916
rect 68948 7876 68957 7916
rect 68899 7875 68957 7876
rect 69091 7916 69149 7917
rect 69091 7876 69100 7916
rect 69140 7876 69149 7916
rect 69091 7875 69149 7876
rect 77635 7916 77693 7917
rect 77635 7876 77644 7916
rect 77684 7876 77693 7916
rect 77635 7875 77693 7876
rect 54315 7832 54357 7841
rect 54315 7792 54316 7832
rect 54356 7792 54357 7832
rect 54315 7783 54357 7792
rect 68139 7832 68181 7841
rect 68139 7792 68140 7832
rect 68180 7792 68181 7832
rect 68139 7783 68181 7792
rect 76971 7832 77013 7841
rect 76971 7792 76972 7832
rect 77012 7792 77013 7832
rect 76971 7783 77013 7792
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 47587 7748 47645 7749
rect 47587 7708 47596 7748
rect 47636 7708 47645 7748
rect 47587 7707 47645 7708
rect 53355 7748 53397 7757
rect 53355 7708 53356 7748
rect 53396 7708 53397 7748
rect 53355 7699 53397 7708
rect 55179 7748 55221 7757
rect 55179 7708 55180 7748
rect 55220 7708 55221 7748
rect 55179 7699 55221 7708
rect 58827 7748 58869 7757
rect 58827 7708 58828 7748
rect 58868 7708 58869 7748
rect 58827 7699 58869 7708
rect 59883 7748 59925 7757
rect 59883 7708 59884 7748
rect 59924 7708 59925 7748
rect 59883 7699 59925 7708
rect 64579 7748 64637 7749
rect 64579 7708 64588 7748
rect 64628 7708 64637 7748
rect 64579 7707 64637 7708
rect 64779 7748 64821 7757
rect 64779 7708 64780 7748
rect 64820 7708 64821 7748
rect 64779 7699 64821 7708
rect 68715 7748 68757 7757
rect 68715 7708 68716 7748
rect 68756 7708 68757 7748
rect 68715 7699 68757 7708
rect 69291 7748 69333 7757
rect 69291 7708 69292 7748
rect 69332 7708 69333 7748
rect 69291 7699 69333 7708
rect 71499 7748 71541 7757
rect 71499 7708 71500 7748
rect 71540 7708 71541 7748
rect 71499 7699 71541 7708
rect 72459 7748 72501 7757
rect 72459 7708 72460 7748
rect 72500 7708 72501 7748
rect 72459 7699 72501 7708
rect 77835 7748 77877 7757
rect 77835 7708 77836 7748
rect 77876 7708 77877 7748
rect 77835 7699 77877 7708
rect 576 7580 79584 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 79584 7580
rect 576 7516 79584 7540
rect 46827 7412 46869 7421
rect 46827 7372 46828 7412
rect 46868 7372 46869 7412
rect 46827 7363 46869 7372
rect 50379 7412 50421 7421
rect 50379 7372 50380 7412
rect 50420 7372 50421 7412
rect 50379 7363 50421 7372
rect 54595 7412 54653 7413
rect 54595 7372 54604 7412
rect 54644 7372 54653 7412
rect 54595 7371 54653 7372
rect 59491 7412 59549 7413
rect 59491 7372 59500 7412
rect 59540 7372 59549 7412
rect 59491 7371 59549 7372
rect 64011 7412 64053 7421
rect 64011 7372 64012 7412
rect 64052 7372 64053 7412
rect 64011 7363 64053 7372
rect 68515 7412 68573 7413
rect 68515 7372 68524 7412
rect 68564 7372 68573 7412
rect 68515 7371 68573 7372
rect 48075 7328 48117 7337
rect 48075 7288 48076 7328
rect 48116 7288 48117 7328
rect 48075 7279 48117 7288
rect 59883 7328 59925 7337
rect 59883 7288 59884 7328
rect 59924 7288 59925 7328
rect 59883 7279 59925 7288
rect 64587 7328 64629 7337
rect 64587 7288 64588 7328
rect 64628 7288 64629 7328
rect 64587 7279 64629 7288
rect 65643 7328 65685 7337
rect 65643 7288 65644 7328
rect 65684 7288 65685 7328
rect 65643 7279 65685 7288
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 47979 7244 48021 7253
rect 47979 7204 47980 7244
rect 48020 7204 48021 7244
rect 47979 7195 48021 7204
rect 48171 7244 48213 7253
rect 48171 7204 48172 7244
rect 48212 7204 48213 7244
rect 48171 7195 48213 7204
rect 56227 7244 56285 7245
rect 56227 7204 56236 7244
rect 56276 7204 56285 7244
rect 56227 7203 56285 7204
rect 59787 7244 59829 7253
rect 59787 7204 59788 7244
rect 59828 7204 59829 7244
rect 59787 7195 59829 7204
rect 59979 7244 60021 7253
rect 59979 7204 59980 7244
rect 60020 7204 60021 7244
rect 68899 7244 68957 7245
rect 68899 7204 68908 7244
rect 68948 7204 68957 7244
rect 59979 7195 60021 7204
rect 65251 7203 65309 7204
rect 68899 7203 68957 7204
rect 73507 7244 73565 7245
rect 73507 7204 73516 7244
rect 73556 7204 73565 7244
rect 73507 7203 73565 7204
rect 46915 7160 46973 7161
rect 46915 7120 46924 7160
rect 46964 7120 46973 7160
rect 46915 7119 46973 7120
rect 47883 7160 47925 7169
rect 47883 7120 47884 7160
rect 47924 7120 47925 7160
rect 47883 7111 47925 7120
rect 48259 7160 48317 7161
rect 48259 7120 48268 7160
rect 48308 7120 48317 7160
rect 48259 7119 48317 7120
rect 50083 7160 50141 7161
rect 50083 7120 50092 7160
rect 50132 7120 50141 7160
rect 50083 7119 50141 7120
rect 50187 7160 50229 7169
rect 50187 7120 50188 7160
rect 50228 7120 50229 7160
rect 50187 7111 50229 7120
rect 50379 7160 50421 7169
rect 50379 7120 50380 7160
rect 50420 7120 50421 7160
rect 50379 7111 50421 7120
rect 51723 7160 51765 7169
rect 51723 7120 51724 7160
rect 51764 7120 51765 7160
rect 51723 7111 51765 7120
rect 51819 7160 51861 7169
rect 51819 7120 51820 7160
rect 51860 7120 51861 7160
rect 51819 7111 51861 7120
rect 51915 7160 51957 7169
rect 51915 7120 51916 7160
rect 51956 7120 51957 7160
rect 51915 7111 51957 7120
rect 52011 7160 52053 7169
rect 52011 7120 52012 7160
rect 52052 7120 52053 7160
rect 52011 7111 52053 7120
rect 52203 7160 52245 7169
rect 52203 7120 52204 7160
rect 52244 7120 52245 7160
rect 52203 7111 52245 7120
rect 52579 7160 52637 7161
rect 52579 7120 52588 7160
rect 52628 7120 52637 7160
rect 52579 7119 52637 7120
rect 53443 7160 53501 7161
rect 53443 7120 53452 7160
rect 53492 7120 53501 7160
rect 53443 7119 53501 7120
rect 56611 7160 56669 7161
rect 56611 7120 56620 7160
rect 56660 7120 56669 7160
rect 56611 7119 56669 7120
rect 57099 7160 57141 7169
rect 57099 7120 57100 7160
rect 57140 7120 57141 7160
rect 57099 7111 57141 7120
rect 57475 7160 57533 7161
rect 57475 7120 57484 7160
rect 57524 7120 57533 7160
rect 57475 7119 57533 7120
rect 58339 7160 58397 7161
rect 58339 7120 58348 7160
rect 58388 7120 58397 7160
rect 58339 7119 58397 7120
rect 59683 7160 59741 7161
rect 59683 7120 59692 7160
rect 59732 7120 59741 7160
rect 59683 7119 59741 7120
rect 60075 7160 60117 7169
rect 60075 7120 60076 7160
rect 60116 7120 60117 7160
rect 60075 7111 60117 7120
rect 61611 7160 61653 7169
rect 61611 7120 61612 7160
rect 61652 7120 61653 7160
rect 61611 7111 61653 7120
rect 61707 7160 61749 7169
rect 61707 7120 61708 7160
rect 61748 7120 61749 7160
rect 61707 7111 61749 7120
rect 61803 7160 61845 7169
rect 61803 7120 61804 7160
rect 61844 7120 61845 7160
rect 61803 7111 61845 7120
rect 62083 7160 62141 7161
rect 62083 7120 62092 7160
rect 62132 7120 62141 7160
rect 62083 7119 62141 7120
rect 62187 7160 62229 7169
rect 62187 7120 62188 7160
rect 62228 7120 62229 7160
rect 62187 7111 62229 7120
rect 64099 7160 64157 7161
rect 64099 7120 64108 7160
rect 64148 7120 64157 7160
rect 64099 7119 64157 7120
rect 64291 7160 64349 7161
rect 64291 7120 64300 7160
rect 64340 7120 64349 7160
rect 64291 7119 64349 7120
rect 64395 7160 64437 7169
rect 64395 7120 64396 7160
rect 64436 7120 64437 7160
rect 64395 7111 64437 7120
rect 64587 7160 64629 7169
rect 65251 7163 65260 7203
rect 65300 7163 65309 7203
rect 65251 7162 65309 7163
rect 64587 7120 64588 7160
rect 64628 7120 64629 7160
rect 64587 7111 64629 7120
rect 64867 7160 64925 7161
rect 64867 7120 64876 7160
rect 64916 7120 64925 7160
rect 64867 7119 64925 7120
rect 65355 7160 65397 7169
rect 65355 7120 65356 7160
rect 65396 7120 65397 7160
rect 65355 7111 65397 7120
rect 66123 7160 66165 7169
rect 66123 7120 66124 7160
rect 66164 7120 66165 7160
rect 66123 7111 66165 7120
rect 66499 7160 66557 7161
rect 66499 7120 66508 7160
rect 66548 7120 66557 7160
rect 66499 7119 66557 7120
rect 67363 7160 67421 7161
rect 67363 7120 67372 7160
rect 67412 7120 67421 7160
rect 67363 7119 67421 7120
rect 70435 7160 70493 7161
rect 70435 7120 70444 7160
rect 70484 7120 70493 7160
rect 70435 7119 70493 7120
rect 71299 7160 71357 7161
rect 71299 7120 71308 7160
rect 71348 7120 71357 7160
rect 71299 7119 71357 7120
rect 72643 7160 72701 7161
rect 72643 7120 72652 7160
rect 72692 7120 72701 7160
rect 72643 7119 72701 7120
rect 72747 7160 72789 7169
rect 72747 7120 72748 7160
rect 72788 7120 72789 7160
rect 72747 7111 72789 7120
rect 73707 7160 73749 7169
rect 73707 7120 73708 7160
rect 73748 7120 73749 7160
rect 73707 7111 73749 7120
rect 73803 7160 73845 7169
rect 73803 7120 73804 7160
rect 73844 7120 73845 7160
rect 73803 7111 73845 7120
rect 73899 7160 73941 7169
rect 73899 7120 73900 7160
rect 73940 7120 73941 7160
rect 73899 7111 73941 7120
rect 73995 7160 74037 7169
rect 73995 7120 73996 7160
rect 74036 7120 74037 7160
rect 73995 7111 74037 7120
rect 74947 7160 75005 7161
rect 74947 7120 74956 7160
rect 74996 7120 75005 7160
rect 74947 7119 75005 7120
rect 75627 7160 75669 7169
rect 75627 7120 75628 7160
rect 75668 7120 75669 7160
rect 75627 7111 75669 7120
rect 76003 7160 76061 7161
rect 76003 7120 76012 7160
rect 76052 7120 76061 7160
rect 76003 7119 76061 7120
rect 76867 7160 76925 7161
rect 76867 7120 76876 7160
rect 76916 7120 76925 7160
rect 76867 7119 76925 7120
rect 78219 7160 78261 7169
rect 78219 7120 78220 7160
rect 78260 7120 78261 7160
rect 78219 7111 78261 7120
rect 78411 7160 78453 7169
rect 78411 7120 78412 7160
rect 78452 7120 78453 7160
rect 78411 7111 78453 7120
rect 78499 7160 78557 7161
rect 78499 7120 78508 7160
rect 78548 7120 78557 7160
rect 78499 7119 78557 7120
rect 78691 7160 78749 7161
rect 78691 7120 78700 7160
rect 78740 7120 78749 7160
rect 78691 7119 78749 7120
rect 56715 7076 56757 7085
rect 56715 7036 56716 7076
rect 56756 7036 56757 7076
rect 56715 7027 56757 7036
rect 70059 7076 70101 7085
rect 70059 7036 70060 7076
rect 70100 7036 70101 7076
rect 70059 7027 70101 7036
rect 75051 7076 75093 7085
rect 75051 7036 75052 7076
rect 75092 7036 75093 7076
rect 75051 7027 75093 7036
rect 78315 7076 78357 7085
rect 78315 7036 78316 7076
rect 78356 7036 78357 7076
rect 78315 7027 78357 7036
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 56043 6992 56085 7001
rect 56043 6952 56044 6992
rect 56084 6952 56085 6992
rect 56043 6943 56085 6952
rect 61507 6992 61565 6993
rect 61507 6952 61516 6992
rect 61556 6952 61565 6992
rect 61507 6951 61565 6952
rect 64971 6992 65013 7001
rect 64971 6952 64972 6992
rect 65012 6952 65013 6992
rect 64971 6943 65013 6952
rect 68715 6992 68757 7001
rect 68715 6952 68716 6992
rect 68756 6952 68757 6992
rect 68715 6943 68757 6952
rect 72451 6992 72509 6993
rect 72451 6952 72460 6992
rect 72500 6952 72509 6992
rect 72451 6951 72509 6952
rect 73323 6992 73365 7001
rect 73323 6952 73324 6992
rect 73364 6952 73365 6992
rect 73323 6943 73365 6952
rect 78019 6992 78077 6993
rect 78019 6952 78028 6992
rect 78068 6952 78077 6992
rect 78019 6951 78077 6952
rect 78795 6992 78837 7001
rect 78795 6952 78796 6992
rect 78836 6952 78837 6992
rect 78795 6943 78837 6952
rect 65163 6934 65205 6943
rect 65163 6894 65164 6934
rect 65204 6894 65205 6934
rect 65163 6885 65205 6894
rect 576 6824 79584 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 79584 6824
rect 576 6760 79584 6784
rect 52779 6660 52821 6669
rect 52779 6620 52780 6660
rect 52820 6620 52821 6660
rect 52779 6611 52821 6620
rect 57955 6656 58013 6657
rect 57955 6616 57964 6656
rect 58004 6616 58013 6656
rect 57955 6615 58013 6616
rect 59971 6656 60029 6657
rect 59971 6616 59980 6656
rect 60020 6616 60029 6656
rect 59971 6615 60029 6616
rect 63523 6656 63581 6657
rect 63523 6616 63532 6656
rect 63572 6616 63581 6656
rect 63523 6615 63581 6616
rect 63715 6656 63773 6657
rect 63715 6616 63724 6656
rect 63764 6616 63773 6656
rect 63715 6615 63773 6616
rect 70819 6656 70877 6657
rect 70819 6616 70828 6656
rect 70868 6616 70877 6656
rect 70819 6615 70877 6616
rect 72739 6656 72797 6657
rect 72739 6616 72748 6656
rect 72788 6616 72797 6656
rect 72739 6615 72797 6616
rect 75619 6656 75677 6657
rect 75619 6616 75628 6656
rect 75668 6616 75677 6656
rect 75619 6615 75677 6616
rect 79459 6656 79517 6657
rect 79459 6616 79468 6656
rect 79508 6616 79517 6656
rect 79459 6615 79517 6616
rect 55083 6572 55125 6581
rect 55083 6532 55084 6572
rect 55124 6532 55125 6572
rect 55083 6523 55125 6532
rect 55563 6572 55605 6581
rect 55563 6532 55564 6572
rect 55604 6532 55605 6572
rect 55563 6523 55605 6532
rect 73227 6572 73269 6581
rect 73227 6532 73228 6572
rect 73268 6532 73269 6572
rect 73227 6523 73269 6532
rect 68139 6509 68181 6518
rect 52587 6488 52629 6497
rect 52587 6448 52588 6488
rect 52628 6448 52629 6488
rect 52587 6439 52629 6448
rect 52675 6488 52733 6489
rect 52675 6448 52684 6488
rect 52724 6448 52733 6488
rect 52675 6447 52733 6448
rect 52971 6488 53013 6497
rect 52971 6448 52972 6488
rect 53012 6448 53013 6488
rect 52971 6439 53013 6448
rect 53163 6488 53205 6497
rect 53163 6448 53164 6488
rect 53204 6448 53205 6488
rect 53163 6439 53205 6448
rect 53277 6495 53319 6504
rect 53277 6455 53278 6495
rect 53318 6455 53319 6495
rect 53277 6446 53319 6455
rect 53451 6488 53493 6497
rect 53451 6448 53452 6488
rect 53492 6448 53493 6488
rect 53451 6439 53493 6448
rect 53547 6488 53589 6497
rect 53547 6448 53548 6488
rect 53588 6448 53589 6488
rect 53547 6439 53589 6448
rect 53643 6488 53685 6497
rect 53643 6448 53644 6488
rect 53684 6448 53685 6488
rect 53643 6439 53685 6448
rect 53739 6488 53781 6497
rect 53739 6448 53740 6488
rect 53780 6448 53781 6488
rect 53739 6439 53781 6448
rect 55179 6488 55221 6497
rect 55179 6448 55180 6488
rect 55220 6448 55221 6488
rect 55179 6439 55221 6448
rect 55275 6488 55317 6497
rect 55275 6448 55276 6488
rect 55316 6448 55317 6488
rect 55275 6439 55317 6448
rect 55371 6488 55413 6497
rect 55371 6448 55372 6488
rect 55412 6448 55413 6488
rect 55371 6439 55413 6448
rect 55939 6488 55997 6489
rect 55939 6448 55948 6488
rect 55988 6448 55997 6488
rect 55939 6447 55997 6448
rect 56803 6488 56861 6489
rect 56803 6448 56812 6488
rect 56852 6448 56861 6488
rect 56803 6447 56861 6448
rect 59779 6488 59837 6489
rect 59779 6448 59788 6488
rect 59828 6448 59837 6488
rect 59779 6447 59837 6448
rect 59883 6488 59925 6497
rect 59883 6448 59884 6488
rect 59924 6448 59925 6488
rect 59883 6439 59925 6448
rect 60075 6488 60117 6497
rect 60075 6448 60076 6488
rect 60116 6448 60117 6488
rect 60075 6439 60117 6448
rect 60651 6488 60693 6497
rect 60651 6448 60652 6488
rect 60692 6448 60693 6488
rect 60651 6439 60693 6448
rect 60747 6488 60789 6497
rect 60747 6448 60748 6488
rect 60788 6448 60789 6488
rect 60747 6439 60789 6448
rect 60843 6488 60885 6497
rect 60843 6448 60844 6488
rect 60884 6448 60885 6488
rect 60843 6439 60885 6448
rect 60939 6488 60981 6497
rect 60939 6448 60940 6488
rect 60980 6448 60981 6488
rect 60939 6439 60981 6448
rect 61131 6488 61173 6497
rect 61131 6448 61132 6488
rect 61172 6448 61173 6488
rect 61131 6439 61173 6448
rect 61507 6488 61565 6489
rect 61507 6448 61516 6488
rect 61556 6448 61565 6488
rect 61507 6447 61565 6448
rect 62371 6488 62429 6489
rect 62371 6448 62380 6488
rect 62420 6448 62429 6488
rect 62371 6447 62429 6448
rect 64867 6488 64925 6489
rect 64867 6448 64876 6488
rect 64916 6448 64925 6488
rect 64867 6447 64925 6448
rect 65731 6488 65789 6489
rect 65731 6448 65740 6488
rect 65780 6448 65789 6488
rect 65731 6447 65789 6448
rect 66123 6488 66165 6497
rect 66123 6448 66124 6488
rect 66164 6448 66165 6488
rect 66123 6439 66165 6448
rect 67947 6488 67989 6497
rect 67947 6448 67948 6488
rect 67988 6448 67989 6488
rect 67947 6439 67989 6448
rect 68043 6488 68085 6497
rect 68043 6448 68044 6488
rect 68084 6448 68085 6488
rect 68139 6469 68140 6509
rect 68180 6469 68181 6509
rect 68139 6460 68181 6469
rect 68235 6488 68277 6497
rect 68043 6439 68085 6448
rect 68235 6448 68236 6488
rect 68276 6448 68277 6488
rect 68235 6439 68277 6448
rect 68427 6488 68469 6497
rect 68427 6448 68428 6488
rect 68468 6448 68469 6488
rect 68427 6439 68469 6448
rect 68803 6488 68861 6489
rect 68803 6448 68812 6488
rect 68852 6448 68861 6488
rect 68803 6447 68861 6448
rect 69667 6488 69725 6489
rect 69667 6448 69676 6488
rect 69716 6448 69725 6488
rect 69667 6447 69725 6448
rect 71499 6488 71541 6497
rect 71499 6448 71500 6488
rect 71540 6448 71541 6488
rect 71499 6439 71541 6448
rect 71875 6488 71933 6489
rect 71875 6448 71884 6488
rect 71924 6448 71933 6488
rect 71875 6447 71933 6448
rect 72267 6488 72309 6497
rect 72267 6448 72268 6488
rect 72308 6448 72309 6488
rect 72267 6439 72309 6448
rect 72459 6488 72501 6497
rect 72459 6448 72460 6488
rect 72500 6448 72501 6488
rect 72459 6439 72501 6448
rect 72547 6488 72605 6489
rect 72547 6448 72556 6488
rect 72596 6448 72605 6488
rect 72547 6447 72605 6448
rect 72843 6488 72885 6497
rect 72843 6448 72844 6488
rect 72884 6448 72885 6488
rect 72843 6439 72885 6448
rect 72939 6488 72981 6497
rect 72939 6448 72940 6488
rect 72980 6448 72981 6488
rect 72939 6439 72981 6448
rect 73035 6488 73077 6497
rect 73035 6448 73036 6488
rect 73076 6448 73077 6488
rect 73035 6439 73077 6448
rect 73603 6488 73661 6489
rect 73603 6448 73612 6488
rect 73652 6448 73661 6488
rect 73603 6447 73661 6448
rect 74467 6488 74525 6489
rect 74467 6448 74476 6488
rect 74516 6448 74525 6488
rect 74467 6447 74525 6448
rect 76483 6488 76541 6489
rect 76483 6448 76492 6488
rect 76532 6448 76541 6488
rect 76483 6447 76541 6448
rect 76875 6488 76917 6497
rect 76875 6448 76876 6488
rect 76916 6448 76917 6488
rect 76875 6439 76917 6448
rect 77067 6488 77109 6497
rect 77067 6448 77068 6488
rect 77108 6448 77109 6488
rect 77067 6439 77109 6448
rect 77443 6488 77501 6489
rect 77443 6448 77452 6488
rect 77492 6448 77501 6488
rect 77443 6447 77501 6448
rect 78307 6488 78365 6489
rect 78307 6448 78316 6488
rect 78356 6448 78365 6488
rect 78307 6447 78365 6448
rect 71595 6404 71637 6413
rect 71595 6364 71596 6404
rect 71636 6364 71637 6404
rect 71595 6355 71637 6364
rect 71787 6404 71829 6413
rect 71787 6364 71788 6404
rect 71828 6364 71829 6404
rect 71787 6355 71829 6364
rect 76587 6404 76629 6413
rect 76587 6364 76588 6404
rect 76628 6364 76629 6404
rect 76587 6355 76629 6364
rect 76779 6404 76821 6413
rect 76779 6364 76780 6404
rect 76820 6364 76821 6404
rect 76779 6355 76821 6364
rect 52299 6320 52341 6329
rect 52299 6280 52300 6320
rect 52340 6280 52341 6320
rect 52299 6271 52341 6280
rect 71691 6320 71733 6329
rect 71691 6280 71692 6320
rect 71732 6280 71733 6320
rect 71691 6271 71733 6280
rect 76683 6320 76725 6329
rect 76683 6280 76684 6320
rect 76724 6280 76725 6320
rect 76683 6271 76725 6280
rect 52971 6236 53013 6245
rect 52971 6196 52972 6236
rect 53012 6196 53013 6236
rect 52971 6187 53013 6196
rect 72267 6236 72309 6245
rect 72267 6196 72268 6236
rect 72308 6196 72309 6236
rect 72267 6187 72309 6196
rect 576 6068 79584 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 79584 6068
rect 576 6004 79584 6028
rect 77163 5900 77205 5909
rect 77163 5860 77164 5900
rect 77204 5860 77205 5900
rect 77163 5851 77205 5860
rect 55179 5816 55221 5825
rect 55179 5776 55180 5816
rect 55220 5776 55221 5816
rect 55179 5767 55221 5776
rect 60939 5816 60981 5825
rect 60939 5776 60940 5816
rect 60980 5776 60981 5816
rect 60939 5767 60981 5776
rect 64683 5816 64725 5825
rect 64683 5776 64684 5816
rect 64724 5776 64725 5816
rect 64683 5767 64725 5776
rect 68619 5816 68661 5825
rect 68619 5776 68620 5816
rect 68660 5776 68661 5816
rect 68619 5767 68661 5776
rect 72459 5816 72501 5825
rect 72459 5776 72460 5816
rect 72500 5776 72501 5816
rect 72459 5767 72501 5776
rect 72939 5816 72981 5825
rect 72939 5776 72940 5816
rect 72980 5776 72981 5816
rect 72939 5767 72981 5776
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 58059 5732 58101 5741
rect 58059 5692 58060 5732
rect 58100 5692 58101 5732
rect 58059 5683 58101 5692
rect 64587 5732 64629 5741
rect 64587 5692 64588 5732
rect 64628 5692 64629 5732
rect 64587 5683 64629 5692
rect 64779 5732 64821 5741
rect 64779 5692 64780 5732
rect 64820 5692 64821 5732
rect 64779 5683 64821 5692
rect 72363 5732 72405 5741
rect 72363 5692 72364 5732
rect 72404 5692 72405 5732
rect 72363 5683 72405 5692
rect 72555 5732 72597 5741
rect 72555 5692 72556 5732
rect 72596 5692 72597 5732
rect 72555 5683 72597 5692
rect 76875 5732 76917 5741
rect 76875 5692 76876 5732
rect 76916 5692 76917 5732
rect 76875 5683 76917 5692
rect 52099 5648 52157 5649
rect 52099 5608 52108 5648
rect 52148 5608 52157 5648
rect 52099 5607 52157 5608
rect 52963 5648 53021 5649
rect 52963 5608 52972 5648
rect 53012 5608 53021 5648
rect 52963 5607 53021 5608
rect 55467 5648 55509 5657
rect 55467 5608 55468 5648
rect 55508 5608 55509 5648
rect 55467 5599 55509 5608
rect 55555 5648 55613 5649
rect 55555 5608 55564 5648
rect 55604 5608 55613 5648
rect 55555 5607 55613 5608
rect 55947 5648 55989 5657
rect 55947 5608 55948 5648
rect 55988 5608 55989 5648
rect 55947 5599 55989 5608
rect 56043 5648 56085 5657
rect 56043 5608 56044 5648
rect 56084 5608 56085 5648
rect 56043 5599 56085 5608
rect 56139 5648 56181 5657
rect 56139 5608 56140 5648
rect 56180 5608 56181 5648
rect 56139 5599 56181 5608
rect 56235 5648 56277 5657
rect 56235 5608 56236 5648
rect 56276 5608 56277 5648
rect 56235 5599 56277 5608
rect 57955 5648 58013 5649
rect 57955 5608 57964 5648
rect 58004 5608 58013 5648
rect 57955 5607 58013 5608
rect 59395 5648 59453 5649
rect 59395 5608 59404 5648
rect 59444 5608 59453 5648
rect 59395 5607 59453 5608
rect 60259 5648 60317 5649
rect 60259 5608 60268 5648
rect 60308 5608 60317 5648
rect 60259 5607 60317 5608
rect 61227 5648 61269 5657
rect 61227 5608 61228 5648
rect 61268 5608 61269 5648
rect 61227 5599 61269 5608
rect 61315 5648 61373 5649
rect 61315 5608 61324 5648
rect 61364 5608 61373 5648
rect 61315 5607 61373 5608
rect 64491 5648 64533 5657
rect 64491 5608 64492 5648
rect 64532 5608 64533 5648
rect 64491 5599 64533 5608
rect 64867 5648 64925 5649
rect 64867 5608 64876 5648
rect 64916 5608 64925 5648
rect 64867 5607 64925 5608
rect 65163 5648 65205 5657
rect 65163 5608 65164 5648
rect 65204 5608 65205 5648
rect 65163 5599 65205 5608
rect 65259 5648 65301 5657
rect 65259 5608 65260 5648
rect 65300 5608 65301 5648
rect 65259 5599 65301 5608
rect 65355 5648 65397 5657
rect 65355 5608 65356 5648
rect 65396 5608 65397 5648
rect 65355 5599 65397 5608
rect 65643 5648 65685 5657
rect 65643 5608 65644 5648
rect 65684 5608 65685 5648
rect 65643 5599 65685 5608
rect 65739 5648 65781 5657
rect 65739 5608 65740 5648
rect 65780 5608 65781 5648
rect 65739 5599 65781 5608
rect 65835 5648 65877 5657
rect 65835 5608 65836 5648
rect 65876 5608 65877 5648
rect 65835 5599 65877 5608
rect 68139 5648 68181 5657
rect 68139 5608 68140 5648
rect 68180 5608 68181 5648
rect 68139 5599 68181 5608
rect 68331 5648 68373 5657
rect 68331 5608 68332 5648
rect 68372 5608 68373 5648
rect 68331 5599 68373 5608
rect 68419 5648 68477 5649
rect 68419 5608 68428 5648
rect 68468 5608 68477 5648
rect 68419 5607 68477 5608
rect 68907 5648 68949 5657
rect 68907 5608 68908 5648
rect 68948 5608 68949 5648
rect 68907 5599 68949 5608
rect 68995 5648 69053 5649
rect 68995 5608 69004 5648
rect 69044 5608 69053 5648
rect 68995 5607 69053 5608
rect 69387 5648 69429 5657
rect 69387 5608 69388 5648
rect 69428 5608 69429 5648
rect 69387 5599 69429 5608
rect 69483 5648 69525 5657
rect 69483 5608 69484 5648
rect 69524 5608 69525 5648
rect 69483 5599 69525 5608
rect 69579 5648 69621 5657
rect 69579 5608 69580 5648
rect 69620 5608 69621 5648
rect 69579 5599 69621 5608
rect 69675 5648 69717 5657
rect 69675 5608 69676 5648
rect 69716 5608 69717 5648
rect 69675 5599 69717 5608
rect 72267 5648 72309 5657
rect 72267 5608 72268 5648
rect 72308 5608 72309 5648
rect 72267 5599 72309 5608
rect 72643 5648 72701 5649
rect 72643 5608 72652 5648
rect 72692 5608 72701 5648
rect 72643 5607 72701 5608
rect 73227 5648 73269 5657
rect 73227 5608 73228 5648
rect 73268 5608 73269 5648
rect 73227 5599 73269 5608
rect 73315 5648 73373 5649
rect 73315 5608 73324 5648
rect 73364 5608 73373 5648
rect 73315 5607 73373 5608
rect 74283 5648 74325 5657
rect 74283 5608 74284 5648
rect 74324 5608 74325 5648
rect 74283 5599 74325 5608
rect 74379 5648 74421 5657
rect 74379 5608 74380 5648
rect 74420 5608 74421 5648
rect 74379 5599 74421 5608
rect 74475 5648 74517 5657
rect 74475 5608 74476 5648
rect 74516 5608 74517 5648
rect 74475 5599 74517 5608
rect 74571 5648 74613 5657
rect 74571 5608 74572 5648
rect 74612 5608 74613 5648
rect 74571 5599 74613 5608
rect 76963 5648 77021 5649
rect 76963 5608 76972 5648
rect 77012 5608 77021 5648
rect 76963 5607 77021 5608
rect 77451 5648 77493 5657
rect 77451 5608 77452 5648
rect 77492 5608 77493 5648
rect 77451 5599 77493 5608
rect 77539 5648 77597 5649
rect 77539 5608 77548 5648
rect 77588 5608 77597 5648
rect 77539 5607 77597 5608
rect 77835 5648 77877 5657
rect 77835 5608 77836 5648
rect 77876 5608 77877 5648
rect 77835 5599 77877 5608
rect 77931 5648 77973 5657
rect 77931 5608 77932 5648
rect 77972 5608 77973 5648
rect 77931 5599 77973 5608
rect 78027 5648 78069 5657
rect 78027 5608 78028 5648
rect 78068 5608 78069 5648
rect 78027 5599 78069 5608
rect 78123 5648 78165 5657
rect 78123 5608 78124 5648
rect 78164 5608 78165 5648
rect 78123 5599 78165 5608
rect 78403 5648 78461 5649
rect 78403 5608 78412 5648
rect 78452 5608 78461 5648
rect 78403 5607 78461 5608
rect 51723 5564 51765 5573
rect 51723 5524 51724 5564
rect 51764 5524 51765 5564
rect 51723 5515 51765 5524
rect 60651 5564 60693 5573
rect 60651 5524 60652 5564
rect 60692 5524 60693 5564
rect 60651 5515 60693 5524
rect 68235 5564 68277 5573
rect 68235 5524 68236 5564
rect 68276 5524 68277 5564
rect 68235 5515 68277 5524
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 54115 5480 54173 5481
rect 54115 5440 54124 5480
rect 54164 5440 54173 5480
rect 54115 5439 54173 5440
rect 58243 5480 58301 5481
rect 58243 5440 58252 5480
rect 58292 5440 58301 5480
rect 58243 5439 58301 5440
rect 65059 5480 65117 5481
rect 65059 5440 65068 5480
rect 65108 5440 65117 5480
rect 65059 5439 65117 5440
rect 65539 5480 65597 5481
rect 65539 5440 65548 5480
rect 65588 5440 65597 5480
rect 65539 5439 65597 5440
rect 73419 5476 73461 5485
rect 73419 5436 73420 5476
rect 73460 5436 73461 5476
rect 55659 5422 55701 5431
rect 55659 5382 55660 5422
rect 55700 5382 55701 5422
rect 55659 5373 55701 5382
rect 61419 5422 61461 5431
rect 61419 5382 61420 5422
rect 61460 5382 61461 5422
rect 61419 5373 61461 5382
rect 69099 5422 69141 5431
rect 73419 5427 73461 5436
rect 77643 5476 77685 5485
rect 77643 5436 77644 5476
rect 77684 5436 77685 5476
rect 77643 5427 77685 5436
rect 78315 5480 78357 5489
rect 78315 5440 78316 5480
rect 78356 5440 78357 5480
rect 78315 5431 78357 5440
rect 69099 5382 69100 5422
rect 69140 5382 69141 5422
rect 69099 5373 69141 5382
rect 576 5312 79584 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 79584 5312
rect 576 5248 79584 5272
rect 55755 5144 55797 5153
rect 55755 5104 55756 5144
rect 55796 5104 55797 5144
rect 55755 5095 55797 5104
rect 61611 5144 61653 5153
rect 61611 5104 61612 5144
rect 61652 5104 61653 5144
rect 61611 5095 61653 5104
rect 62283 5144 62325 5153
rect 62283 5104 62284 5144
rect 62324 5104 62325 5144
rect 62283 5095 62325 5104
rect 65067 5148 65109 5157
rect 65067 5108 65068 5148
rect 65108 5108 65109 5148
rect 65067 5099 65109 5108
rect 67747 5144 67805 5145
rect 67747 5104 67756 5144
rect 67796 5104 67805 5144
rect 67747 5103 67805 5104
rect 70339 5144 70397 5145
rect 70339 5104 70348 5144
rect 70388 5104 70397 5144
rect 70339 5103 70397 5104
rect 73227 5144 73269 5153
rect 73227 5104 73228 5144
rect 73268 5104 73269 5144
rect 73227 5095 73269 5104
rect 74379 5144 74421 5153
rect 74379 5104 74380 5144
rect 74420 5104 74421 5144
rect 74379 5095 74421 5104
rect 76963 5144 77021 5145
rect 76963 5104 76972 5144
rect 77012 5104 77021 5144
rect 76963 5103 77021 5104
rect 77731 5144 77789 5145
rect 77731 5104 77740 5144
rect 77780 5104 77789 5144
rect 77731 5103 77789 5104
rect 60555 5060 60597 5069
rect 60555 5020 60556 5060
rect 60596 5020 60597 5060
rect 60555 5011 60597 5020
rect 65355 5060 65397 5069
rect 65355 5020 65356 5060
rect 65396 5020 65397 5060
rect 65355 5011 65397 5020
rect 70539 5060 70581 5069
rect 70539 5020 70540 5060
rect 70580 5020 70581 5060
rect 70539 5011 70581 5020
rect 64099 4991 64157 4992
rect 52195 4976 52253 4977
rect 52195 4936 52204 4976
rect 52244 4936 52253 4976
rect 52195 4935 52253 4936
rect 52587 4976 52629 4985
rect 52587 4936 52588 4976
rect 52628 4936 52629 4976
rect 52587 4927 52629 4936
rect 53443 4976 53501 4977
rect 53443 4936 53452 4976
rect 53492 4936 53501 4976
rect 53443 4935 53501 4936
rect 53923 4976 53981 4977
rect 53923 4936 53932 4976
rect 53972 4936 53981 4976
rect 53923 4935 53981 4936
rect 54027 4976 54069 4985
rect 54027 4936 54028 4976
rect 54068 4936 54069 4976
rect 54027 4927 54069 4936
rect 54219 4976 54261 4985
rect 54219 4936 54220 4976
rect 54260 4936 54261 4976
rect 54219 4927 54261 4936
rect 54411 4976 54453 4985
rect 54411 4936 54412 4976
rect 54452 4936 54453 4976
rect 54411 4927 54453 4936
rect 54787 4976 54845 4977
rect 54787 4936 54796 4976
rect 54836 4936 54845 4976
rect 54787 4935 54845 4936
rect 55843 4976 55901 4977
rect 55843 4936 55852 4976
rect 55892 4936 55901 4976
rect 55843 4935 55901 4936
rect 56907 4976 56949 4985
rect 56907 4936 56908 4976
rect 56948 4936 56949 4976
rect 56907 4927 56949 4936
rect 57003 4976 57045 4985
rect 57003 4936 57004 4976
rect 57044 4936 57045 4976
rect 57003 4927 57045 4936
rect 57099 4976 57141 4985
rect 57099 4936 57100 4976
rect 57140 4936 57141 4976
rect 57099 4927 57141 4936
rect 57195 4976 57237 4985
rect 57195 4936 57196 4976
rect 57236 4936 57237 4976
rect 57195 4927 57237 4936
rect 57387 4976 57429 4985
rect 57387 4936 57388 4976
rect 57428 4936 57429 4976
rect 57387 4927 57429 4936
rect 57763 4976 57821 4977
rect 57763 4936 57772 4976
rect 57812 4936 57821 4976
rect 57763 4935 57821 4936
rect 58627 4976 58685 4977
rect 58627 4936 58636 4976
rect 58676 4936 58685 4976
rect 58627 4935 58685 4936
rect 60451 4976 60509 4977
rect 60451 4936 60460 4976
rect 60500 4936 60509 4976
rect 60451 4935 60509 4936
rect 60739 4976 60797 4977
rect 60739 4936 60748 4976
rect 60788 4936 60797 4976
rect 60739 4935 60797 4936
rect 61131 4976 61173 4985
rect 61131 4936 61132 4976
rect 61172 4936 61173 4976
rect 61131 4927 61173 4936
rect 62179 4976 62237 4977
rect 62179 4936 62188 4976
rect 62228 4936 62237 4976
rect 64099 4951 64108 4991
rect 64148 4951 64157 4991
rect 64395 4976 64437 4985
rect 64099 4950 64157 4951
rect 64195 4962 64253 4963
rect 62179 4935 62237 4936
rect 64195 4922 64204 4962
rect 64244 4922 64253 4962
rect 64395 4936 64396 4976
rect 64436 4936 64437 4976
rect 64395 4927 64437 4936
rect 64875 4976 64917 4985
rect 64875 4936 64876 4976
rect 64916 4936 64917 4976
rect 64875 4927 64917 4936
rect 64963 4976 65021 4977
rect 64963 4936 64972 4976
rect 65012 4936 65021 4976
rect 64963 4935 65021 4936
rect 65731 4976 65789 4977
rect 65731 4936 65740 4976
rect 65780 4936 65789 4976
rect 65731 4935 65789 4936
rect 66595 4976 66653 4977
rect 66595 4936 66604 4976
rect 66644 4936 66653 4976
rect 66595 4935 66653 4936
rect 67947 4976 67989 4985
rect 67947 4936 67948 4976
rect 67988 4936 67989 4976
rect 67947 4927 67989 4936
rect 68323 4976 68381 4977
rect 68323 4936 68332 4976
rect 68372 4936 68381 4976
rect 68323 4935 68381 4936
rect 69187 4976 69245 4977
rect 69187 4936 69196 4976
rect 69236 4936 69245 4976
rect 69187 4935 69245 4936
rect 70915 4976 70973 4977
rect 70915 4936 70924 4976
rect 70964 4936 70973 4976
rect 70915 4935 70973 4936
rect 71779 4976 71837 4977
rect 71779 4936 71788 4976
rect 71828 4936 71837 4976
rect 71779 4935 71837 4936
rect 73123 4976 73181 4977
rect 73123 4936 73132 4976
rect 73172 4936 73181 4976
rect 73123 4935 73181 4936
rect 74275 4976 74333 4977
rect 74275 4936 74284 4976
rect 74324 4936 74333 4976
rect 74275 4935 74333 4936
rect 74571 4976 74613 4985
rect 74571 4936 74572 4976
rect 74612 4936 74613 4976
rect 74571 4927 74613 4936
rect 74947 4976 75005 4977
rect 74947 4936 74956 4976
rect 74996 4936 75005 4976
rect 74947 4935 75005 4936
rect 75811 4976 75869 4977
rect 75811 4936 75820 4976
rect 75860 4936 75869 4976
rect 77355 4976 77397 4985
rect 75811 4935 75869 4936
rect 77163 4934 77205 4943
rect 77355 4936 77356 4976
rect 77396 4936 77397 4976
rect 64195 4921 64253 4922
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 52299 4892 52341 4901
rect 52299 4852 52300 4892
rect 52340 4852 52341 4892
rect 52299 4843 52341 4852
rect 52491 4892 52533 4901
rect 52491 4852 52492 4892
rect 52532 4852 52533 4892
rect 52491 4843 52533 4852
rect 53355 4892 53397 4901
rect 53355 4852 53356 4892
rect 53396 4852 53397 4892
rect 53355 4843 53397 4852
rect 54507 4892 54549 4901
rect 54507 4852 54508 4892
rect 54548 4852 54549 4892
rect 54507 4843 54549 4852
rect 54699 4892 54741 4901
rect 54699 4852 54700 4892
rect 54740 4852 54741 4892
rect 54699 4843 54741 4852
rect 60843 4892 60885 4901
rect 60843 4852 60844 4892
rect 60884 4852 60885 4892
rect 60843 4843 60885 4852
rect 61035 4892 61077 4901
rect 77163 4894 77164 4934
rect 77204 4894 77205 4934
rect 61035 4852 61036 4892
rect 61076 4852 61077 4892
rect 61035 4843 61077 4852
rect 61411 4892 61469 4893
rect 61411 4852 61420 4892
rect 61460 4852 61469 4892
rect 61411 4851 61469 4852
rect 61795 4892 61853 4893
rect 61795 4852 61804 4892
rect 61844 4852 61853 4892
rect 77163 4885 77205 4894
rect 77251 4934 77309 4935
rect 77251 4894 77260 4934
rect 77300 4894 77309 4934
rect 77355 4927 77397 4936
rect 77451 4976 77493 4985
rect 77451 4936 77452 4976
rect 77492 4936 77493 4976
rect 77451 4927 77493 4936
rect 77643 4976 77685 4985
rect 77643 4936 77644 4976
rect 77684 4936 77685 4976
rect 77643 4927 77685 4936
rect 77835 4976 77877 4985
rect 77835 4936 77836 4976
rect 77876 4936 77877 4976
rect 77835 4927 77877 4936
rect 77923 4976 77981 4977
rect 77923 4936 77932 4976
rect 77972 4936 77981 4976
rect 77923 4935 77981 4936
rect 77251 4893 77309 4894
rect 61795 4851 61853 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 52395 4808 52437 4817
rect 52395 4768 52396 4808
rect 52436 4768 52437 4808
rect 52395 4759 52437 4768
rect 54603 4808 54645 4817
rect 54603 4768 54604 4808
rect 54644 4768 54645 4808
rect 54603 4759 54645 4768
rect 59779 4808 59837 4809
rect 59779 4768 59788 4808
rect 59828 4768 59837 4808
rect 59779 4767 59837 4768
rect 60939 4808 60981 4817
rect 60939 4768 60940 4808
rect 60980 4768 60981 4808
rect 60939 4759 60981 4768
rect 64587 4808 64629 4817
rect 64587 4768 64588 4808
rect 64628 4768 64629 4808
rect 64587 4759 64629 4768
rect 54219 4724 54261 4733
rect 54219 4684 54220 4724
rect 54260 4684 54261 4724
rect 54219 4675 54261 4684
rect 61611 4724 61653 4733
rect 61611 4684 61612 4724
rect 61652 4684 61653 4724
rect 61611 4675 61653 4684
rect 61995 4724 62037 4733
rect 61995 4684 61996 4724
rect 62036 4684 62037 4724
rect 61995 4675 62037 4684
rect 62283 4724 62325 4733
rect 62283 4684 62284 4724
rect 62324 4684 62325 4724
rect 62283 4675 62325 4684
rect 64395 4724 64437 4733
rect 64395 4684 64396 4724
rect 64436 4684 64437 4724
rect 64395 4675 64437 4684
rect 72931 4724 72989 4725
rect 72931 4684 72940 4724
rect 72980 4684 72989 4724
rect 72931 4683 72989 4684
rect 74379 4724 74421 4733
rect 74379 4684 74380 4724
rect 74420 4684 74421 4724
rect 74379 4675 74421 4684
rect 576 4556 79584 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 79584 4556
rect 576 4492 79584 4516
rect 65835 4388 65877 4397
rect 65835 4348 65836 4388
rect 65876 4348 65877 4388
rect 65835 4339 65877 4348
rect 69291 4388 69333 4397
rect 69291 4348 69292 4388
rect 69332 4348 69333 4388
rect 69291 4339 69333 4348
rect 56227 4304 56285 4305
rect 56227 4264 56236 4304
rect 56276 4264 56285 4304
rect 56227 4263 56285 4264
rect 57003 4304 57045 4313
rect 57003 4264 57004 4304
rect 57044 4264 57045 4304
rect 57003 4255 57045 4264
rect 63043 4304 63101 4305
rect 63043 4264 63052 4304
rect 63092 4264 63101 4304
rect 63043 4263 63101 4264
rect 68523 4304 68565 4313
rect 68523 4264 68524 4304
rect 68564 4264 68565 4304
rect 68523 4255 68565 4264
rect 68907 4304 68949 4313
rect 68907 4264 68908 4304
rect 68948 4264 68949 4304
rect 68907 4255 68949 4264
rect 71691 4304 71733 4313
rect 71691 4264 71692 4304
rect 71732 4264 71733 4304
rect 71691 4255 71733 4264
rect 72555 4304 72597 4313
rect 72555 4264 72556 4304
rect 72596 4264 72597 4304
rect 72555 4255 72597 4264
rect 75139 4304 75197 4305
rect 75139 4264 75148 4304
rect 75188 4264 75197 4304
rect 75139 4263 75197 4264
rect 76299 4304 76341 4313
rect 76299 4264 76300 4304
rect 76340 4264 76341 4304
rect 76299 4255 76341 4264
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 66019 4220 66077 4221
rect 66019 4180 66028 4220
rect 66068 4180 66077 4220
rect 66019 4179 66077 4180
rect 68427 4220 68469 4229
rect 68427 4180 68428 4220
rect 68468 4180 68469 4220
rect 68427 4171 68469 4180
rect 68619 4220 68661 4229
rect 68619 4180 68620 4220
rect 68660 4180 68661 4220
rect 68619 4171 68661 4180
rect 69091 4220 69149 4221
rect 69091 4180 69100 4220
rect 69140 4180 69149 4220
rect 69091 4179 69149 4180
rect 71595 4220 71637 4229
rect 71595 4180 71596 4220
rect 71636 4180 71637 4220
rect 71595 4171 71637 4180
rect 71787 4220 71829 4229
rect 71787 4180 71788 4220
rect 71828 4180 71829 4220
rect 71787 4171 71829 4180
rect 79371 4220 79413 4229
rect 79371 4180 79372 4220
rect 79412 4180 79413 4220
rect 79371 4171 79413 4180
rect 53835 4136 53877 4145
rect 53835 4096 53836 4136
rect 53876 4096 53877 4136
rect 53835 4087 53877 4096
rect 54211 4136 54269 4137
rect 54211 4096 54220 4136
rect 54260 4096 54269 4136
rect 54211 4095 54269 4096
rect 55075 4136 55133 4137
rect 55075 4096 55084 4136
rect 55124 4096 55133 4136
rect 55075 4095 55133 4096
rect 56419 4136 56477 4137
rect 56419 4096 56428 4136
rect 56468 4096 56477 4136
rect 56419 4095 56477 4096
rect 56523 4136 56565 4145
rect 56523 4096 56524 4136
rect 56564 4096 56565 4136
rect 56523 4087 56565 4096
rect 56715 4136 56757 4145
rect 56715 4096 56716 4136
rect 56756 4096 56757 4136
rect 56715 4087 56757 4096
rect 57291 4136 57333 4145
rect 57291 4096 57292 4136
rect 57332 4096 57333 4136
rect 57291 4087 57333 4096
rect 57379 4136 57437 4137
rect 57379 4096 57388 4136
rect 57428 4096 57437 4136
rect 57379 4095 57437 4096
rect 57675 4136 57717 4145
rect 57675 4096 57676 4136
rect 57716 4096 57717 4136
rect 57675 4087 57717 4096
rect 57771 4136 57813 4145
rect 57771 4096 57772 4136
rect 57812 4096 57813 4136
rect 57771 4087 57813 4096
rect 57867 4136 57909 4145
rect 57867 4096 57868 4136
rect 57908 4096 57909 4136
rect 57867 4087 57909 4096
rect 57963 4136 58005 4145
rect 57963 4096 57964 4136
rect 58004 4096 58005 4136
rect 57963 4087 58005 4096
rect 60267 4136 60309 4145
rect 60267 4096 60268 4136
rect 60308 4096 60309 4136
rect 60267 4087 60309 4096
rect 60363 4136 60405 4145
rect 60363 4096 60364 4136
rect 60404 4096 60405 4136
rect 60363 4087 60405 4096
rect 60459 4136 60501 4145
rect 60459 4096 60460 4136
rect 60500 4096 60501 4136
rect 60459 4087 60501 4096
rect 61027 4136 61085 4137
rect 61027 4096 61036 4136
rect 61076 4096 61085 4136
rect 61027 4095 61085 4096
rect 61891 4136 61949 4137
rect 61891 4096 61900 4136
rect 61940 4096 61949 4136
rect 61891 4095 61949 4096
rect 63619 4136 63677 4137
rect 63619 4096 63628 4136
rect 63668 4096 63677 4136
rect 63619 4095 63677 4096
rect 64483 4136 64541 4137
rect 64483 4096 64492 4136
rect 64532 4096 64541 4136
rect 64483 4095 64541 4096
rect 68323 4136 68381 4137
rect 68323 4096 68332 4136
rect 68372 4096 68381 4136
rect 68323 4095 68381 4096
rect 68715 4136 68757 4145
rect 68715 4096 68716 4136
rect 68756 4096 68757 4136
rect 68715 4087 68757 4096
rect 69379 4136 69437 4137
rect 69379 4096 69388 4136
rect 69428 4096 69437 4136
rect 69379 4095 69437 4096
rect 71019 4136 71061 4145
rect 71019 4096 71020 4136
rect 71060 4096 71061 4136
rect 71019 4087 71061 4096
rect 71211 4136 71253 4145
rect 71211 4096 71212 4136
rect 71252 4096 71253 4136
rect 71211 4087 71253 4096
rect 71299 4136 71357 4137
rect 71299 4096 71308 4136
rect 71348 4096 71357 4136
rect 71299 4095 71357 4096
rect 71499 4136 71541 4145
rect 71499 4096 71500 4136
rect 71540 4096 71541 4136
rect 71499 4087 71541 4096
rect 71875 4136 71933 4137
rect 71875 4096 71884 4136
rect 71924 4096 71933 4136
rect 71875 4095 71933 4096
rect 72163 4136 72221 4137
rect 72163 4096 72172 4136
rect 72212 4096 72221 4136
rect 72163 4095 72221 4096
rect 72267 4136 72309 4145
rect 72267 4096 72268 4136
rect 72308 4096 72309 4136
rect 72267 4087 72309 4096
rect 73123 4136 73181 4137
rect 73123 4096 73132 4136
rect 73172 4096 73181 4136
rect 73123 4095 73181 4096
rect 73987 4136 74045 4137
rect 73987 4096 73996 4136
rect 74036 4096 74045 4136
rect 73987 4095 74045 4096
rect 75819 4136 75861 4145
rect 75819 4096 75820 4136
rect 75860 4096 75861 4136
rect 75819 4087 75861 4096
rect 75915 4136 75957 4145
rect 75915 4096 75916 4136
rect 75956 4096 75957 4136
rect 75915 4087 75957 4096
rect 76011 4136 76053 4145
rect 76011 4096 76012 4136
rect 76052 4096 76053 4136
rect 76011 4087 76053 4096
rect 76107 4136 76149 4145
rect 76107 4096 76108 4136
rect 76148 4096 76149 4136
rect 76107 4087 76149 4096
rect 76587 4136 76629 4145
rect 76587 4096 76588 4136
rect 76628 4096 76629 4136
rect 76587 4087 76629 4096
rect 76675 4136 76733 4137
rect 76675 4096 76684 4136
rect 76724 4096 76733 4136
rect 76675 4095 76733 4096
rect 77347 4136 77405 4137
rect 77347 4096 77356 4136
rect 77396 4096 77405 4136
rect 77347 4095 77405 4096
rect 78211 4136 78269 4137
rect 78211 4096 78220 4136
rect 78260 4096 78269 4136
rect 78211 4095 78269 4096
rect 60171 4052 60213 4061
rect 60171 4012 60172 4052
rect 60212 4012 60213 4052
rect 60171 4003 60213 4012
rect 60651 4052 60693 4061
rect 60651 4012 60652 4052
rect 60692 4012 60693 4052
rect 60651 4003 60693 4012
rect 63243 4052 63285 4061
rect 63243 4012 63244 4052
rect 63284 4012 63285 4052
rect 63243 4003 63285 4012
rect 72747 4052 72789 4061
rect 72747 4012 72748 4052
rect 72788 4012 72789 4052
rect 72747 4003 72789 4012
rect 76971 4052 77013 4061
rect 76971 4012 76972 4052
rect 77012 4012 77013 4052
rect 76971 4003 77013 4012
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 56611 3968 56669 3969
rect 56611 3928 56620 3968
rect 56660 3928 56669 3968
rect 56611 3927 56669 3928
rect 65635 3968 65693 3969
rect 65635 3928 65644 3968
rect 65684 3928 65693 3968
rect 65635 3927 65693 3928
rect 71107 3968 71165 3969
rect 71107 3928 71116 3968
rect 71156 3928 71165 3968
rect 71107 3927 71165 3928
rect 72075 3964 72117 3973
rect 72075 3924 72076 3964
rect 72116 3924 72117 3964
rect 57483 3910 57525 3919
rect 72075 3915 72117 3924
rect 57483 3870 57484 3910
rect 57524 3870 57525 3910
rect 57483 3861 57525 3870
rect 76779 3910 76821 3919
rect 76779 3870 76780 3910
rect 76820 3870 76821 3910
rect 76779 3861 76821 3870
rect 576 3800 79584 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 79584 3800
rect 576 3736 79584 3760
rect 5163 3632 5205 3641
rect 5163 3592 5164 3632
rect 5204 3592 5205 3632
rect 5163 3583 5205 3592
rect 60267 3636 60309 3645
rect 60267 3596 60268 3636
rect 60308 3596 60309 3636
rect 60267 3587 60309 3596
rect 61411 3632 61469 3633
rect 61411 3592 61420 3632
rect 61460 3592 61469 3632
rect 61411 3591 61469 3592
rect 61803 3632 61845 3641
rect 61803 3592 61804 3632
rect 61844 3592 61845 3632
rect 61803 3583 61845 3592
rect 64875 3632 64917 3641
rect 64875 3592 64876 3632
rect 64916 3592 64917 3632
rect 64875 3583 64917 3592
rect 68803 3632 68861 3633
rect 68803 3592 68812 3632
rect 68852 3592 68861 3632
rect 68803 3591 68861 3592
rect 69003 3632 69045 3641
rect 69003 3592 69004 3632
rect 69044 3592 69045 3632
rect 69003 3583 69045 3592
rect 72739 3632 72797 3633
rect 72739 3592 72748 3632
rect 72788 3592 72797 3632
rect 72739 3591 72797 3592
rect 73035 3632 73077 3641
rect 73035 3592 73036 3632
rect 73076 3592 73077 3632
rect 73035 3583 73077 3592
rect 73987 3632 74045 3633
rect 73987 3592 73996 3632
rect 74036 3592 74045 3632
rect 73987 3591 74045 3592
rect 77835 3632 77877 3641
rect 77835 3592 77836 3632
rect 77876 3592 77877 3632
rect 77835 3583 77877 3592
rect 69675 3548 69717 3557
rect 69675 3508 69676 3548
rect 69716 3508 69717 3548
rect 69675 3499 69717 3508
rect 5059 3464 5117 3465
rect 5059 3424 5068 3464
rect 5108 3424 5117 3464
rect 5059 3423 5117 3424
rect 56043 3464 56085 3473
rect 56043 3424 56044 3464
rect 56084 3424 56085 3464
rect 56043 3415 56085 3424
rect 56419 3464 56477 3465
rect 56419 3424 56428 3464
rect 56468 3424 56477 3464
rect 56419 3423 56477 3424
rect 57283 3464 57341 3465
rect 57283 3424 57292 3464
rect 57332 3424 57341 3464
rect 57283 3423 57341 3424
rect 60075 3464 60117 3473
rect 60075 3424 60076 3464
rect 60116 3424 60117 3464
rect 60075 3415 60117 3424
rect 60163 3464 60221 3465
rect 60163 3424 60172 3464
rect 60212 3424 60221 3464
rect 60163 3423 60221 3424
rect 60555 3464 60597 3473
rect 60555 3424 60556 3464
rect 60596 3424 60597 3464
rect 60555 3415 60597 3424
rect 60651 3464 60693 3473
rect 60651 3424 60652 3464
rect 60692 3424 60693 3464
rect 60651 3415 60693 3424
rect 60747 3464 60789 3473
rect 60747 3424 60748 3464
rect 60788 3424 60789 3464
rect 60747 3415 60789 3424
rect 60843 3464 60885 3473
rect 60843 3424 60844 3464
rect 60884 3424 60885 3464
rect 60843 3415 60885 3424
rect 61323 3464 61365 3473
rect 61323 3424 61324 3464
rect 61364 3424 61365 3464
rect 61323 3415 61365 3424
rect 61515 3464 61557 3473
rect 61515 3424 61516 3464
rect 61556 3424 61557 3464
rect 64299 3464 64341 3473
rect 61515 3415 61557 3424
rect 61603 3445 61661 3446
rect 61603 3405 61612 3445
rect 61652 3405 61661 3445
rect 64299 3424 64300 3464
rect 64340 3424 64341 3464
rect 64299 3415 64341 3424
rect 64675 3464 64733 3465
rect 64675 3424 64684 3464
rect 64724 3424 64733 3464
rect 64675 3423 64733 3424
rect 64963 3464 65021 3465
rect 64963 3424 64972 3464
rect 65012 3424 65021 3464
rect 64963 3423 65021 3424
rect 65451 3464 65493 3473
rect 65451 3424 65452 3464
rect 65492 3424 65493 3464
rect 65451 3415 65493 3424
rect 65547 3464 65589 3473
rect 65547 3424 65548 3464
rect 65588 3424 65589 3464
rect 65547 3415 65589 3424
rect 65643 3464 65685 3473
rect 65643 3424 65644 3464
rect 65684 3424 65685 3464
rect 65643 3415 65685 3424
rect 65739 3464 65781 3473
rect 65739 3424 65740 3464
rect 65780 3424 65781 3464
rect 65739 3415 65781 3424
rect 65931 3464 65973 3473
rect 65931 3424 65932 3464
rect 65972 3424 65973 3464
rect 65931 3415 65973 3424
rect 66027 3464 66069 3473
rect 66027 3424 66028 3464
rect 66068 3424 66069 3464
rect 66027 3415 66069 3424
rect 66123 3464 66165 3473
rect 66123 3424 66124 3464
rect 66164 3424 66165 3464
rect 66123 3415 66165 3424
rect 66219 3464 66261 3473
rect 66219 3424 66220 3464
rect 66260 3424 66261 3464
rect 66219 3415 66261 3424
rect 66411 3464 66453 3473
rect 66411 3424 66412 3464
rect 66452 3424 66453 3464
rect 66411 3415 66453 3424
rect 66787 3464 66845 3465
rect 66787 3424 66796 3464
rect 66836 3424 66845 3464
rect 66787 3423 66845 3424
rect 67651 3464 67709 3465
rect 67651 3424 67660 3464
rect 67700 3424 67709 3464
rect 67651 3423 67709 3424
rect 70051 3464 70109 3465
rect 70051 3424 70060 3464
rect 70100 3424 70109 3464
rect 70051 3423 70109 3424
rect 70915 3464 70973 3465
rect 70915 3424 70924 3464
rect 70964 3424 70973 3464
rect 70915 3423 70973 3424
rect 72459 3464 72501 3473
rect 72459 3424 72460 3464
rect 72500 3424 72501 3464
rect 72459 3415 72501 3424
rect 72555 3464 72597 3473
rect 72555 3424 72556 3464
rect 72596 3424 72597 3464
rect 72555 3415 72597 3424
rect 72651 3464 72693 3473
rect 72651 3424 72652 3464
rect 72692 3424 72693 3464
rect 72651 3415 72693 3424
rect 72931 3464 72989 3465
rect 72931 3424 72940 3464
rect 72980 3424 72989 3464
rect 72931 3423 72989 3424
rect 73507 3464 73565 3465
rect 73507 3424 73516 3464
rect 73556 3424 73565 3464
rect 73507 3423 73565 3424
rect 74091 3464 74133 3473
rect 74091 3424 74092 3464
rect 74132 3424 74133 3464
rect 74091 3415 74133 3424
rect 74187 3464 74229 3473
rect 74187 3424 74188 3464
rect 74228 3424 74229 3464
rect 74187 3415 74229 3424
rect 74283 3464 74325 3473
rect 74283 3424 74284 3464
rect 74324 3424 74325 3464
rect 74283 3415 74325 3424
rect 76675 3464 76733 3465
rect 76675 3424 76684 3464
rect 76724 3424 76733 3464
rect 76675 3423 76733 3424
rect 76963 3464 77021 3465
rect 76963 3424 76972 3464
rect 77012 3424 77021 3464
rect 76963 3423 77021 3424
rect 77355 3464 77397 3473
rect 77355 3424 77356 3464
rect 77396 3424 77397 3464
rect 77355 3415 77397 3424
rect 78027 3464 78069 3473
rect 78027 3424 78028 3464
rect 78068 3424 78069 3464
rect 78027 3415 78069 3424
rect 78115 3464 78173 3465
rect 78115 3424 78124 3464
rect 78164 3424 78173 3464
rect 78115 3423 78173 3424
rect 61603 3404 61661 3405
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 61987 3380 62045 3381
rect 61987 3340 61996 3380
rect 62036 3340 62045 3380
rect 61987 3339 62045 3340
rect 64395 3380 64437 3389
rect 64395 3340 64396 3380
rect 64436 3340 64437 3380
rect 64395 3331 64437 3340
rect 64587 3380 64629 3389
rect 64587 3340 64588 3380
rect 64628 3340 64629 3380
rect 64587 3331 64629 3340
rect 69187 3380 69245 3381
rect 69187 3340 69196 3380
rect 69236 3340 69245 3380
rect 69187 3339 69245 3340
rect 77067 3380 77109 3389
rect 77067 3340 77068 3380
rect 77108 3340 77109 3380
rect 77067 3331 77109 3340
rect 77259 3380 77301 3389
rect 77259 3340 77260 3380
rect 77300 3340 77301 3380
rect 77259 3331 77301 3340
rect 77635 3380 77693 3381
rect 77635 3340 77644 3380
rect 77684 3340 77693 3380
rect 77635 3339 77693 3340
rect 59787 3296 59829 3305
rect 59787 3256 59788 3296
rect 59828 3256 59829 3296
rect 59787 3247 59829 3256
rect 64491 3296 64533 3305
rect 64491 3256 64492 3296
rect 64532 3256 64533 3296
rect 64491 3247 64533 3256
rect 76779 3296 76821 3305
rect 76779 3256 76780 3296
rect 76820 3256 76821 3296
rect 76779 3247 76821 3256
rect 77163 3296 77205 3305
rect 77163 3256 77164 3296
rect 77204 3256 77205 3296
rect 77163 3247 77205 3256
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 58435 3212 58493 3213
rect 58435 3172 58444 3212
rect 58484 3172 58493 3212
rect 58435 3171 58493 3172
rect 72067 3212 72125 3213
rect 72067 3172 72076 3212
rect 72116 3172 72125 3212
rect 72067 3171 72125 3172
rect 73419 3212 73461 3221
rect 73419 3172 73420 3212
rect 73460 3172 73461 3212
rect 73419 3163 73461 3172
rect 77835 3212 77877 3221
rect 77835 3172 77836 3212
rect 77876 3172 77877 3212
rect 77835 3163 77877 3172
rect 576 3044 79584 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 79584 3044
rect 576 2980 79584 3004
rect 57867 2876 57909 2885
rect 57867 2836 57868 2876
rect 57908 2836 57909 2876
rect 57867 2827 57909 2836
rect 60171 2876 60213 2885
rect 60171 2836 60172 2876
rect 60212 2836 60213 2876
rect 60171 2827 60213 2836
rect 63339 2876 63381 2885
rect 63339 2836 63340 2876
rect 63380 2836 63381 2876
rect 63339 2827 63381 2836
rect 68619 2876 68661 2885
rect 68619 2836 68620 2876
rect 68660 2836 68661 2876
rect 68619 2827 68661 2836
rect 73803 2876 73845 2885
rect 73803 2836 73804 2876
rect 73844 2836 73845 2876
rect 73803 2827 73845 2836
rect 75051 2876 75093 2885
rect 75051 2836 75052 2876
rect 75092 2836 75093 2876
rect 75051 2827 75093 2836
rect 77355 2876 77397 2885
rect 77355 2836 77356 2876
rect 77396 2836 77397 2876
rect 77355 2827 77397 2836
rect 56523 2792 56565 2801
rect 56523 2752 56524 2792
rect 56564 2752 56565 2792
rect 56523 2743 56565 2752
rect 58731 2792 58773 2801
rect 58731 2752 58732 2792
rect 58772 2752 58773 2792
rect 58731 2743 58773 2752
rect 59115 2792 59157 2801
rect 59115 2752 59116 2792
rect 59156 2752 59157 2792
rect 59115 2743 59157 2752
rect 60747 2792 60789 2801
rect 60747 2752 60748 2792
rect 60788 2752 60789 2792
rect 60747 2743 60789 2752
rect 61131 2792 61173 2801
rect 61131 2752 61132 2792
rect 61172 2752 61173 2792
rect 61131 2743 61173 2752
rect 61707 2792 61749 2801
rect 61707 2752 61708 2792
rect 61748 2752 61749 2792
rect 61707 2743 61749 2752
rect 65067 2792 65109 2801
rect 65067 2752 65068 2792
rect 65108 2752 65109 2792
rect 65067 2743 65109 2752
rect 66027 2792 66069 2801
rect 66027 2752 66028 2792
rect 66068 2752 66069 2792
rect 66027 2743 66069 2752
rect 71979 2792 72021 2801
rect 71979 2752 71980 2792
rect 72020 2752 72021 2792
rect 71979 2743 72021 2752
rect 72363 2792 72405 2801
rect 72363 2752 72364 2792
rect 72404 2752 72405 2792
rect 72363 2743 72405 2752
rect 76587 2792 76629 2801
rect 76587 2752 76588 2792
rect 76628 2752 76629 2792
rect 76587 2743 76629 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 56427 2708 56469 2717
rect 56427 2668 56428 2708
rect 56468 2668 56469 2708
rect 56427 2659 56469 2668
rect 56619 2708 56661 2717
rect 56619 2668 56620 2708
rect 56660 2668 56661 2708
rect 56619 2659 56661 2668
rect 59019 2708 59061 2717
rect 59019 2668 59020 2708
rect 59060 2668 59061 2708
rect 59019 2659 59061 2668
rect 59211 2708 59253 2717
rect 59211 2668 59212 2708
rect 59252 2668 59253 2708
rect 59211 2659 59253 2668
rect 61035 2708 61077 2717
rect 61035 2668 61036 2708
rect 61076 2668 61077 2708
rect 61035 2659 61077 2668
rect 61227 2708 61269 2717
rect 61227 2668 61228 2708
rect 61268 2668 61269 2708
rect 61227 2659 61269 2668
rect 64971 2708 65013 2717
rect 64971 2668 64972 2708
rect 65012 2668 65013 2708
rect 64971 2659 65013 2668
rect 65163 2708 65205 2717
rect 65163 2668 65164 2708
rect 65204 2668 65205 2708
rect 65163 2659 65205 2668
rect 71883 2708 71925 2717
rect 71883 2668 71884 2708
rect 71924 2668 71925 2708
rect 71883 2659 71925 2668
rect 72075 2708 72117 2717
rect 72075 2668 72076 2708
rect 72116 2668 72117 2708
rect 72075 2659 72117 2668
rect 56331 2624 56373 2633
rect 56331 2584 56332 2624
rect 56372 2584 56373 2624
rect 56331 2575 56373 2584
rect 56707 2624 56765 2625
rect 56707 2584 56716 2624
rect 56756 2584 56765 2624
rect 56707 2583 56765 2584
rect 57955 2624 58013 2625
rect 57955 2584 57964 2624
rect 58004 2584 58013 2624
rect 57955 2583 58013 2584
rect 58435 2624 58493 2625
rect 58435 2584 58444 2624
rect 58484 2584 58493 2624
rect 58435 2583 58493 2584
rect 58539 2624 58581 2633
rect 58539 2584 58540 2624
rect 58580 2584 58581 2624
rect 58539 2575 58581 2584
rect 58731 2624 58773 2633
rect 58731 2584 58732 2624
rect 58772 2584 58773 2624
rect 58731 2575 58773 2584
rect 58923 2624 58965 2633
rect 58923 2584 58924 2624
rect 58964 2584 58965 2624
rect 58923 2575 58965 2584
rect 59299 2624 59357 2625
rect 59299 2584 59308 2624
rect 59348 2584 59357 2624
rect 59299 2583 59357 2584
rect 60259 2624 60317 2625
rect 60259 2584 60268 2624
rect 60308 2584 60317 2624
rect 60259 2583 60317 2584
rect 60451 2624 60509 2625
rect 60451 2584 60460 2624
rect 60500 2584 60509 2624
rect 60451 2583 60509 2584
rect 60555 2624 60597 2633
rect 60555 2584 60556 2624
rect 60596 2584 60597 2624
rect 60555 2575 60597 2584
rect 60747 2624 60789 2633
rect 60747 2584 60748 2624
rect 60788 2584 60789 2624
rect 60747 2575 60789 2584
rect 60939 2624 60981 2633
rect 60939 2584 60940 2624
rect 60980 2584 60981 2624
rect 60939 2575 60981 2584
rect 61315 2624 61373 2625
rect 61315 2584 61324 2624
rect 61364 2584 61373 2624
rect 61315 2583 61373 2584
rect 61995 2624 62037 2633
rect 61995 2584 61996 2624
rect 62036 2584 62037 2624
rect 61995 2575 62037 2584
rect 62083 2624 62141 2625
rect 62083 2584 62092 2624
rect 62132 2584 62141 2624
rect 62083 2583 62141 2584
rect 62475 2624 62517 2633
rect 62475 2584 62476 2624
rect 62516 2584 62517 2624
rect 62475 2575 62517 2584
rect 62571 2624 62613 2633
rect 62571 2584 62572 2624
rect 62612 2584 62613 2624
rect 62571 2575 62613 2584
rect 62667 2624 62709 2633
rect 62667 2584 62668 2624
rect 62708 2584 62709 2624
rect 62667 2575 62709 2584
rect 62851 2624 62909 2625
rect 62851 2584 62860 2624
rect 62900 2584 62909 2624
rect 62851 2583 62909 2584
rect 63235 2624 63293 2625
rect 63235 2584 63244 2624
rect 63284 2584 63293 2624
rect 63235 2583 63293 2584
rect 64395 2624 64437 2633
rect 64395 2584 64396 2624
rect 64436 2584 64437 2624
rect 64395 2575 64437 2584
rect 64587 2624 64629 2633
rect 64587 2584 64588 2624
rect 64628 2584 64629 2624
rect 64587 2575 64629 2584
rect 64675 2624 64733 2625
rect 64675 2584 64684 2624
rect 64724 2584 64733 2624
rect 64675 2583 64733 2584
rect 64875 2624 64917 2633
rect 64875 2584 64876 2624
rect 64916 2584 64917 2624
rect 64875 2575 64917 2584
rect 65251 2624 65309 2625
rect 65251 2584 65260 2624
rect 65300 2584 65309 2624
rect 65251 2583 65309 2584
rect 65635 2624 65693 2625
rect 65635 2584 65644 2624
rect 65684 2584 65693 2624
rect 65635 2583 65693 2584
rect 65739 2624 65781 2633
rect 65739 2584 65740 2624
rect 65780 2584 65781 2624
rect 65739 2575 65781 2584
rect 66595 2624 66653 2625
rect 66595 2584 66604 2624
rect 66644 2584 66653 2624
rect 66595 2583 66653 2584
rect 66699 2624 66741 2633
rect 66699 2584 66700 2624
rect 66740 2584 66741 2624
rect 66699 2575 66741 2584
rect 66891 2624 66933 2633
rect 66891 2584 66892 2624
rect 66932 2584 66933 2624
rect 66891 2575 66933 2584
rect 68235 2624 68277 2633
rect 68235 2584 68236 2624
rect 68276 2584 68277 2624
rect 68235 2575 68277 2584
rect 68331 2624 68373 2633
rect 68331 2584 68332 2624
rect 68372 2584 68373 2624
rect 68331 2575 68373 2584
rect 68427 2624 68469 2633
rect 68427 2584 68428 2624
rect 68468 2584 68469 2624
rect 68427 2575 68469 2584
rect 68619 2624 68661 2633
rect 68619 2584 68620 2624
rect 68660 2584 68661 2624
rect 68619 2575 68661 2584
rect 68811 2624 68853 2633
rect 68811 2584 68812 2624
rect 68852 2584 68853 2624
rect 68811 2575 68853 2584
rect 68899 2624 68957 2625
rect 68899 2584 68908 2624
rect 68948 2584 68957 2624
rect 68899 2583 68957 2584
rect 69187 2624 69245 2625
rect 69187 2584 69196 2624
rect 69236 2584 69245 2624
rect 69187 2583 69245 2584
rect 71307 2624 71349 2633
rect 71307 2584 71308 2624
rect 71348 2584 71349 2624
rect 71307 2575 71349 2584
rect 71499 2624 71541 2633
rect 71499 2584 71500 2624
rect 71540 2584 71541 2624
rect 71499 2575 71541 2584
rect 71587 2624 71645 2625
rect 71587 2584 71596 2624
rect 71636 2584 71645 2624
rect 71587 2583 71645 2584
rect 71787 2624 71829 2633
rect 71787 2584 71788 2624
rect 71828 2584 71829 2624
rect 71787 2575 71829 2584
rect 72163 2624 72221 2625
rect 72163 2584 72172 2624
rect 72212 2584 72221 2624
rect 72163 2583 72221 2584
rect 72651 2624 72693 2633
rect 72651 2584 72652 2624
rect 72692 2584 72693 2624
rect 72651 2575 72693 2584
rect 72739 2624 72797 2625
rect 72739 2584 72748 2624
rect 72788 2584 72797 2624
rect 72739 2583 72797 2584
rect 73123 2624 73181 2625
rect 73123 2584 73132 2624
rect 73172 2584 73181 2624
rect 73123 2583 73181 2584
rect 74083 2624 74141 2625
rect 74083 2584 74092 2624
rect 74132 2584 74141 2624
rect 74083 2583 74141 2584
rect 74947 2624 75005 2625
rect 74947 2584 74956 2624
rect 74996 2584 75005 2624
rect 74947 2583 75005 2584
rect 76107 2624 76149 2633
rect 76107 2584 76108 2624
rect 76148 2584 76149 2624
rect 76107 2575 76149 2584
rect 76203 2624 76245 2633
rect 76203 2584 76204 2624
rect 76244 2584 76245 2624
rect 76203 2575 76245 2584
rect 76299 2624 76341 2633
rect 76299 2584 76300 2624
rect 76340 2584 76341 2624
rect 76299 2575 76341 2584
rect 76875 2624 76917 2633
rect 76875 2584 76876 2624
rect 76916 2584 76917 2624
rect 76875 2575 76917 2584
rect 76963 2624 77021 2625
rect 76963 2584 76972 2624
rect 77012 2584 77021 2624
rect 76963 2583 77021 2584
rect 77355 2624 77397 2633
rect 77355 2584 77356 2624
rect 77396 2584 77397 2624
rect 77355 2575 77397 2584
rect 77547 2624 77589 2633
rect 77547 2584 77548 2624
rect 77588 2584 77589 2624
rect 77547 2575 77589 2584
rect 77635 2624 77693 2625
rect 77635 2584 77644 2624
rect 77684 2584 77693 2624
rect 77635 2583 77693 2584
rect 77923 2624 77981 2625
rect 77923 2584 77932 2624
rect 77972 2584 77981 2624
rect 77923 2583 77981 2584
rect 64491 2540 64533 2549
rect 64491 2500 64492 2540
rect 64532 2500 64533 2540
rect 64491 2491 64533 2500
rect 77835 2540 77877 2549
rect 77835 2500 77836 2540
rect 77876 2500 77877 2540
rect 77835 2491 77877 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 62187 2452 62229 2461
rect 62187 2412 62188 2452
rect 62228 2412 62229 2452
rect 62371 2456 62429 2457
rect 62371 2416 62380 2456
rect 62420 2416 62429 2456
rect 62371 2415 62429 2416
rect 62955 2456 62997 2465
rect 62955 2416 62956 2456
rect 62996 2416 62997 2456
rect 62187 2403 62229 2412
rect 62955 2407 62997 2416
rect 66787 2456 66845 2457
rect 66787 2416 66796 2456
rect 66836 2416 66845 2456
rect 66787 2415 66845 2416
rect 68131 2456 68189 2457
rect 68131 2416 68140 2456
rect 68180 2416 68189 2456
rect 68131 2415 68189 2416
rect 69099 2456 69141 2465
rect 69099 2416 69100 2456
rect 69140 2416 69141 2456
rect 69099 2407 69141 2416
rect 71395 2456 71453 2457
rect 71395 2416 71404 2456
rect 71444 2416 71453 2456
rect 71395 2415 71453 2416
rect 72843 2452 72885 2461
rect 72843 2412 72844 2452
rect 72884 2412 72885 2452
rect 65547 2398 65589 2407
rect 72843 2403 72885 2412
rect 75051 2456 75093 2465
rect 75051 2416 75052 2456
rect 75092 2416 75093 2456
rect 75051 2407 75093 2416
rect 76387 2456 76445 2457
rect 76387 2416 76396 2456
rect 76436 2416 76445 2456
rect 76387 2415 76445 2416
rect 65547 2358 65548 2398
rect 65588 2358 65589 2398
rect 65547 2349 65589 2358
rect 77067 2398 77109 2407
rect 77067 2358 77068 2398
rect 77108 2358 77109 2398
rect 77067 2349 77109 2358
rect 576 2288 79584 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 79584 2288
rect 576 2224 79584 2248
rect 68619 2178 68661 2187
rect 68619 2138 68620 2178
rect 68660 2138 68661 2178
rect 68619 2129 68661 2138
rect 60739 2120 60797 2121
rect 60739 2080 60748 2120
rect 60788 2080 60797 2120
rect 60739 2079 60797 2080
rect 64771 2120 64829 2121
rect 64771 2080 64780 2120
rect 64820 2080 64829 2120
rect 64771 2079 64829 2080
rect 71203 2120 71261 2121
rect 71203 2080 71212 2120
rect 71252 2080 71261 2120
rect 71203 2079 71261 2080
rect 73795 2120 73853 2121
rect 73795 2080 73804 2120
rect 73844 2080 73853 2120
rect 73795 2079 73853 2080
rect 73987 2120 74045 2121
rect 73987 2080 73996 2120
rect 74036 2080 74045 2120
rect 73987 2079 74045 2080
rect 78403 2120 78461 2121
rect 78403 2080 78412 2120
rect 78452 2080 78461 2120
rect 78403 2079 78461 2080
rect 58347 2036 58389 2045
rect 58347 1996 58348 2036
rect 58388 1996 58389 2036
rect 58347 1987 58389 1996
rect 62379 2036 62421 2045
rect 62379 1996 62380 2036
rect 62420 1996 62421 2036
rect 62379 1987 62421 1996
rect 64971 2036 65013 2045
rect 64971 1996 64972 2036
rect 65012 1996 65013 2036
rect 64971 1987 65013 1996
rect 68811 2036 68853 2045
rect 68811 1996 68812 2036
rect 68852 1996 68853 2036
rect 68811 1987 68853 1996
rect 71403 2036 71445 2045
rect 71403 1996 71404 2036
rect 71444 1996 71445 2036
rect 71403 1987 71445 1996
rect 58723 1952 58781 1953
rect 58723 1912 58732 1952
rect 58772 1912 58781 1952
rect 58723 1911 58781 1912
rect 59587 1952 59645 1953
rect 59587 1912 59596 1952
rect 59636 1912 59645 1952
rect 59587 1911 59645 1912
rect 61323 1952 61365 1961
rect 61323 1912 61324 1952
rect 61364 1912 61365 1952
rect 61323 1903 61365 1912
rect 62755 1952 62813 1953
rect 62755 1912 62764 1952
rect 62804 1912 62813 1952
rect 62755 1911 62813 1912
rect 63619 1952 63677 1953
rect 63619 1912 63628 1952
rect 63668 1912 63677 1952
rect 63619 1911 63677 1912
rect 65347 1952 65405 1953
rect 65347 1912 65356 1952
rect 65396 1912 65405 1952
rect 65347 1911 65405 1912
rect 66211 1952 66269 1953
rect 66211 1912 66220 1952
rect 66260 1912 66269 1952
rect 66211 1911 66269 1912
rect 67563 1952 67605 1961
rect 67563 1912 67564 1952
rect 67604 1912 67605 1952
rect 67939 1952 67997 1953
rect 67563 1903 67605 1912
rect 67659 1910 67701 1919
rect 67939 1912 67948 1952
rect 67988 1912 67997 1952
rect 67939 1911 67997 1912
rect 68427 1952 68469 1961
rect 68427 1912 68428 1952
rect 68468 1912 68469 1952
rect 67659 1870 67660 1910
rect 67700 1870 67701 1910
rect 68427 1903 68469 1912
rect 68515 1952 68573 1953
rect 68515 1912 68524 1952
rect 68564 1912 68573 1952
rect 68515 1911 68573 1912
rect 69187 1952 69245 1953
rect 69187 1912 69196 1952
rect 69236 1912 69245 1952
rect 69187 1911 69245 1912
rect 70051 1952 70109 1953
rect 70051 1912 70060 1952
rect 70100 1912 70109 1952
rect 70051 1911 70109 1912
rect 71779 1952 71837 1953
rect 71779 1912 71788 1952
rect 71828 1912 71837 1952
rect 71779 1911 71837 1912
rect 72643 1952 72701 1953
rect 72643 1912 72652 1952
rect 72692 1912 72701 1952
rect 72643 1911 72701 1912
rect 74091 1952 74133 1961
rect 74091 1912 74092 1952
rect 74132 1912 74133 1952
rect 74091 1903 74133 1912
rect 74187 1952 74229 1961
rect 74187 1912 74188 1952
rect 74228 1912 74229 1952
rect 74187 1903 74229 1912
rect 74283 1952 74325 1961
rect 74283 1912 74284 1952
rect 74324 1912 74325 1952
rect 74283 1903 74325 1912
rect 74467 1952 74525 1953
rect 74467 1912 74476 1952
rect 74516 1912 74525 1952
rect 74467 1911 74525 1912
rect 74571 1952 74613 1961
rect 74571 1912 74572 1952
rect 74612 1912 74613 1952
rect 74571 1903 74613 1912
rect 74763 1952 74805 1961
rect 74763 1912 74764 1952
rect 74804 1912 74805 1952
rect 74763 1903 74805 1912
rect 75435 1952 75477 1961
rect 75435 1912 75436 1952
rect 75476 1912 75477 1952
rect 75435 1903 75477 1912
rect 75811 1952 75869 1953
rect 75811 1912 75820 1952
rect 75860 1912 75869 1952
rect 75811 1911 75869 1912
rect 76011 1952 76053 1961
rect 76011 1912 76012 1952
rect 76052 1912 76053 1952
rect 76011 1903 76053 1912
rect 76387 1952 76445 1953
rect 76387 1912 76396 1952
rect 76436 1912 76445 1952
rect 76387 1911 76445 1912
rect 77251 1952 77309 1953
rect 77251 1912 77260 1952
rect 77300 1912 77309 1952
rect 77251 1911 77309 1912
rect 67659 1861 67701 1870
rect 67851 1868 67893 1877
rect 67851 1828 67852 1868
rect 67892 1828 67893 1868
rect 67851 1819 67893 1828
rect 75531 1868 75573 1877
rect 75531 1828 75532 1868
rect 75572 1828 75573 1868
rect 75531 1819 75573 1828
rect 75723 1868 75765 1877
rect 75723 1828 75724 1868
rect 75764 1828 75765 1868
rect 75723 1819 75765 1828
rect 61899 1784 61941 1793
rect 61899 1744 61900 1784
rect 61940 1744 61941 1784
rect 61899 1735 61941 1744
rect 67755 1784 67797 1793
rect 67755 1744 67756 1784
rect 67796 1744 67797 1784
rect 67755 1735 67797 1744
rect 68139 1784 68181 1793
rect 68139 1744 68140 1784
rect 68180 1744 68181 1784
rect 68139 1735 68181 1744
rect 74763 1784 74805 1793
rect 74763 1744 74764 1784
rect 74804 1744 74805 1784
rect 74763 1735 74805 1744
rect 75627 1784 75669 1793
rect 75627 1744 75628 1784
rect 75668 1744 75669 1784
rect 75627 1735 75669 1744
rect 67363 1700 67421 1701
rect 67363 1660 67372 1700
rect 67412 1660 67421 1700
rect 67363 1659 67421 1660
rect 71203 1700 71261 1701
rect 71203 1660 71212 1700
rect 71252 1660 71261 1700
rect 71203 1659 71261 1660
rect 576 1532 79584 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 79584 1532
rect 576 1468 79584 1492
rect 62275 1364 62333 1365
rect 62275 1324 62284 1364
rect 62324 1324 62333 1364
rect 62275 1323 62333 1324
rect 66123 1364 66165 1373
rect 66123 1324 66124 1364
rect 66164 1324 66165 1364
rect 66123 1315 66165 1324
rect 69187 1364 69245 1365
rect 69187 1324 69196 1364
rect 69236 1324 69245 1364
rect 69187 1323 69245 1324
rect 70731 1364 70773 1373
rect 70731 1324 70732 1364
rect 70772 1324 70773 1364
rect 70731 1315 70773 1324
rect 72267 1364 72309 1373
rect 72267 1324 72268 1364
rect 72308 1324 72309 1364
rect 72267 1315 72309 1324
rect 75619 1364 75677 1365
rect 75619 1324 75628 1364
rect 75668 1324 75677 1364
rect 75619 1323 75677 1324
rect 79371 1196 79413 1205
rect 79371 1156 79372 1196
rect 79412 1156 79413 1196
rect 79371 1147 79413 1156
rect 59587 1112 59645 1113
rect 59587 1072 59596 1112
rect 59636 1072 59645 1112
rect 59587 1071 59645 1072
rect 59883 1112 59925 1121
rect 59883 1072 59884 1112
rect 59924 1072 59925 1112
rect 59883 1063 59925 1072
rect 60259 1112 60317 1113
rect 60259 1072 60268 1112
rect 60308 1072 60317 1112
rect 60259 1071 60317 1072
rect 61123 1112 61181 1113
rect 61123 1072 61132 1112
rect 61172 1072 61181 1112
rect 61123 1071 61181 1072
rect 62571 1112 62613 1121
rect 62571 1072 62572 1112
rect 62612 1072 62613 1112
rect 62571 1063 62613 1072
rect 62667 1112 62709 1121
rect 62667 1072 62668 1112
rect 62708 1072 62709 1112
rect 62667 1063 62709 1072
rect 62763 1112 62805 1121
rect 62763 1072 62764 1112
rect 62804 1072 62805 1112
rect 62763 1063 62805 1072
rect 62859 1112 62901 1121
rect 62859 1072 62860 1112
rect 62900 1072 62901 1112
rect 62859 1063 62901 1072
rect 66211 1112 66269 1113
rect 66211 1072 66220 1112
rect 66260 1072 66269 1112
rect 66211 1071 66269 1072
rect 66795 1112 66837 1121
rect 66795 1072 66796 1112
rect 66836 1072 66837 1112
rect 66795 1063 66837 1072
rect 67171 1112 67229 1113
rect 67171 1072 67180 1112
rect 67220 1072 67229 1112
rect 67171 1071 67229 1072
rect 68035 1112 68093 1113
rect 68035 1072 68044 1112
rect 68084 1072 68093 1112
rect 68035 1071 68093 1072
rect 69483 1112 69525 1121
rect 69483 1072 69484 1112
rect 69524 1072 69525 1112
rect 69483 1063 69525 1072
rect 69579 1112 69621 1121
rect 69579 1072 69580 1112
rect 69620 1072 69621 1112
rect 69579 1063 69621 1072
rect 69675 1112 69717 1121
rect 69675 1072 69676 1112
rect 69716 1072 69717 1112
rect 69675 1063 69717 1072
rect 69771 1112 69813 1121
rect 69771 1072 69772 1112
rect 69812 1072 69813 1112
rect 69771 1063 69813 1072
rect 70051 1112 70109 1113
rect 70051 1072 70060 1112
rect 70100 1072 70109 1112
rect 70051 1071 70109 1072
rect 70243 1112 70301 1113
rect 70243 1072 70252 1112
rect 70292 1072 70301 1112
rect 70243 1071 70301 1072
rect 71115 1112 71157 1121
rect 71115 1072 71116 1112
rect 71156 1072 71157 1112
rect 71115 1063 71157 1072
rect 71499 1112 71541 1121
rect 71499 1072 71500 1112
rect 71540 1072 71541 1112
rect 71499 1063 71541 1072
rect 71595 1112 71637 1121
rect 71595 1072 71596 1112
rect 71636 1072 71637 1112
rect 71595 1063 71637 1072
rect 71691 1112 71733 1121
rect 71691 1072 71692 1112
rect 71732 1072 71733 1112
rect 71691 1063 71733 1072
rect 72843 1112 72885 1121
rect 72843 1072 72844 1112
rect 72884 1072 72885 1112
rect 72843 1063 72885 1072
rect 73603 1112 73661 1113
rect 73603 1072 73612 1112
rect 73652 1072 73661 1112
rect 73603 1071 73661 1072
rect 74467 1112 74525 1113
rect 74467 1072 74476 1112
rect 74516 1072 74525 1112
rect 74467 1071 74525 1072
rect 76491 1112 76533 1121
rect 76491 1072 76492 1112
rect 76532 1072 76533 1112
rect 76491 1063 76533 1072
rect 76587 1112 76629 1121
rect 76587 1072 76588 1112
rect 76628 1072 76629 1112
rect 76587 1063 76629 1072
rect 76683 1112 76725 1121
rect 76683 1072 76684 1112
rect 76724 1072 76725 1112
rect 76683 1063 76725 1072
rect 76779 1112 76821 1121
rect 76779 1072 76780 1112
rect 76820 1072 76821 1112
rect 76779 1063 76821 1072
rect 76971 1112 77013 1121
rect 76971 1072 76972 1112
rect 77012 1072 77013 1112
rect 76971 1063 77013 1072
rect 77347 1112 77405 1113
rect 77347 1072 77356 1112
rect 77396 1072 77405 1112
rect 77347 1071 77405 1072
rect 78211 1112 78269 1113
rect 78211 1072 78220 1112
rect 78260 1072 78269 1112
rect 78211 1071 78269 1072
rect 71787 1028 71829 1037
rect 71787 988 71788 1028
rect 71828 988 71829 1028
rect 71787 979 71829 988
rect 73227 1028 73269 1037
rect 73227 988 73228 1028
rect 73268 988 73269 1028
rect 73227 979 73269 988
rect 576 776 79584 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 79584 776
rect 576 712 79584 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 57676 38200 57716 38240
rect 59884 38200 59924 38240
rect 61228 38200 61268 38240
rect 61420 38200 61460 38240
rect 61516 38200 61556 38240
rect 64684 38200 64724 38240
rect 65260 38200 65300 38240
rect 65452 38200 65492 38240
rect 65548 38200 65588 38240
rect 65740 38200 65780 38240
rect 66892 38200 66932 38240
rect 68332 38200 68372 38240
rect 68716 38200 68756 38240
rect 69580 38200 69620 38240
rect 69964 38200 70004 38240
rect 70060 38200 70100 38240
rect 70156 38200 70196 38240
rect 70252 38200 70292 38240
rect 73996 38200 74036 38240
rect 74188 38200 74228 38240
rect 74284 38200 74324 38240
rect 74476 38200 74516 38240
rect 74572 38200 74612 38240
rect 74668 38200 74708 38240
rect 74764 38200 74804 38240
rect 75628 38200 75668 38240
rect 75916 38200 75956 38240
rect 652 38116 692 38156
rect 64876 38116 64916 38156
rect 70444 38116 70484 38156
rect 71020 38116 71060 38156
rect 77260 38116 77300 38156
rect 67756 38032 67796 38072
rect 844 37948 884 37988
rect 57580 37948 57620 37988
rect 59980 37948 60020 37988
rect 61228 37948 61268 37988
rect 65068 37948 65108 37988
rect 65260 37948 65300 37988
rect 65836 37948 65876 37988
rect 66700 37948 66740 37988
rect 70636 37948 70676 37988
rect 70828 37948 70868 37988
rect 73996 37948 74036 37988
rect 76204 37948 76244 37988
rect 77452 37948 77492 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 73132 37528 73172 37568
rect 56620 37444 56660 37484
rect 56812 37444 56852 37484
rect 57100 37444 57140 37484
rect 60268 37444 60308 37484
rect 64204 37444 64244 37484
rect 56524 37360 56564 37400
rect 64108 37402 64148 37442
rect 64396 37444 64436 37484
rect 67372 37444 67412 37484
rect 56908 37360 56948 37400
rect 58636 37360 58676 37400
rect 59500 37360 59540 37400
rect 60940 37360 60980 37400
rect 61804 37360 61844 37400
rect 64492 37360 64532 37400
rect 65932 37360 65972 37400
rect 66796 37360 66836 37400
rect 68908 37360 68948 37400
rect 69772 37360 69812 37400
rect 70156 37360 70196 37400
rect 71500 37360 71540 37400
rect 72364 37360 72404 37400
rect 73420 37360 73460 37400
rect 73516 37360 73556 37400
rect 74188 37360 74228 37400
rect 75052 37360 75092 37400
rect 76588 37360 76628 37400
rect 77164 37360 77204 37400
rect 78028 37360 78068 37400
rect 56716 37234 56756 37274
rect 59884 37276 59924 37316
rect 60556 37276 60596 37316
rect 57292 37192 57332 37232
rect 57484 37192 57524 37232
rect 64300 37234 64340 37274
rect 67180 37276 67220 37316
rect 72748 37276 72788 37316
rect 73804 37276 73844 37316
rect 76780 37276 76820 37316
rect 60076 37192 60116 37232
rect 62956 37192 62996 37232
rect 64780 37192 64820 37232
rect 67564 37192 67604 37232
rect 67756 37192 67796 37232
rect 70348 37192 70388 37232
rect 76204 37192 76244 37232
rect 76492 37192 76532 37232
rect 79180 37192 79220 37232
rect 73612 37134 73652 37174
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 67660 36914 67700 36954
rect 59404 36856 59444 36896
rect 60172 36860 60212 36900
rect 60844 36856 60884 36896
rect 69388 36856 69428 36896
rect 74092 36856 74132 36896
rect 56236 36772 56276 36812
rect 64108 36772 64148 36812
rect 73324 36772 73364 36812
rect 56620 36688 56660 36728
rect 57484 36688 57524 36728
rect 59596 36688 59636 36728
rect 59980 36688 60020 36728
rect 60268 36688 60308 36728
rect 60364 36688 60404 36728
rect 60940 36688 60980 36728
rect 61036 36688 61076 36728
rect 61132 36688 61172 36728
rect 62860 36688 62900 36728
rect 63724 36688 63764 36728
rect 64300 36688 64340 36728
rect 64684 36688 64724 36728
rect 65548 36688 65588 36728
rect 67084 36688 67124 36728
rect 67468 36688 67508 36728
rect 67756 36688 67796 36728
rect 67852 36688 67892 36728
rect 68332 36688 68372 36728
rect 68524 36688 68564 36728
rect 68620 36688 68660 36728
rect 68812 36688 68852 36728
rect 68908 36688 68948 36728
rect 69004 36688 69044 36728
rect 69100 36688 69140 36728
rect 69292 36688 69332 36728
rect 70732 36688 70772 36728
rect 71596 36688 71636 36728
rect 71980 36688 72020 36728
rect 72172 36688 72212 36728
rect 72556 36688 72596 36728
rect 72748 36688 72788 36728
rect 72940 36688 72980 36728
rect 73036 36688 73076 36728
rect 73228 36688 73268 36728
rect 73516 36688 73556 36728
rect 73900 36688 73940 36728
rect 74188 36688 74228 36728
rect 74284 36688 74324 36728
rect 74380 36688 74420 36728
rect 75340 36688 75380 36728
rect 75628 36688 75668 36728
rect 75724 36688 75764 36728
rect 75820 36688 75860 36728
rect 75916 36688 75956 36728
rect 76108 36688 76148 36728
rect 76492 36688 76532 36728
rect 76684 36688 76724 36728
rect 77068 36688 77108 36728
rect 77932 36688 77972 36728
rect 58828 36604 58868 36644
rect 59212 36604 59252 36644
rect 59692 36604 59732 36644
rect 59884 36604 59924 36644
rect 67180 36604 67220 36644
rect 67372 36604 67412 36644
rect 72268 36604 72308 36644
rect 72460 36604 72500 36644
rect 73612 36604 73652 36644
rect 73804 36604 73844 36644
rect 74572 36604 74612 36644
rect 76204 36604 76244 36644
rect 76396 36604 76436 36644
rect 58636 36520 58676 36560
rect 59788 36520 59828 36560
rect 60652 36520 60692 36560
rect 67276 36520 67316 36560
rect 68140 36520 68180 36560
rect 68332 36520 68372 36560
rect 72364 36520 72404 36560
rect 72748 36520 72788 36560
rect 73708 36520 73748 36560
rect 74764 36520 74804 36560
rect 76300 36520 76340 36560
rect 59020 36436 59060 36476
rect 59404 36436 59444 36476
rect 61708 36436 61748 36476
rect 66700 36436 66740 36476
rect 69580 36436 69620 36476
rect 75436 36436 75476 36476
rect 79084 36436 79124 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 56428 36100 56468 36140
rect 63916 36100 63956 36140
rect 72172 36100 72212 36140
rect 72940 36100 72980 36140
rect 77260 36100 77300 36140
rect 77452 36100 77492 36140
rect 64588 36016 64628 36056
rect 74284 35932 74324 35972
rect 74668 35932 74708 35972
rect 56044 35848 56084 35888
rect 56140 35848 56180 35888
rect 56236 35848 56276 35888
rect 56716 35848 56756 35888
rect 56812 35848 56852 35888
rect 57100 35848 57140 35888
rect 57196 35848 57236 35888
rect 57292 35848 57332 35888
rect 57388 35827 57428 35867
rect 57676 35848 57716 35888
rect 57868 35848 57908 35888
rect 57964 35848 58004 35888
rect 58156 35848 58196 35888
rect 58252 35848 58292 35888
rect 58444 35848 58484 35888
rect 59020 35848 59060 35888
rect 59884 35848 59924 35888
rect 61228 35848 61268 35888
rect 61324 35848 61364 35888
rect 61420 35848 61460 35888
rect 61516 35848 61556 35888
rect 61708 35837 61748 35877
rect 63820 35848 63860 35888
rect 64204 35848 64244 35888
rect 64300 35848 64340 35888
rect 64780 35848 64820 35888
rect 64876 35848 64916 35888
rect 64972 35848 65012 35888
rect 65068 35848 65108 35888
rect 65260 35848 65300 35888
rect 65356 35848 65396 35888
rect 65452 35848 65492 35888
rect 65548 35848 65588 35888
rect 65836 35848 65876 35888
rect 66796 35848 66836 35888
rect 67660 35848 67700 35888
rect 71308 35848 71348 35888
rect 71404 35848 71444 35888
rect 71596 35848 71636 35888
rect 72076 35848 72116 35888
rect 72556 35848 72596 35888
rect 72652 35848 72692 35888
rect 73804 35848 73844 35888
rect 73900 35848 73940 35888
rect 73996 35848 74036 35888
rect 74092 35848 74132 35888
rect 76300 35848 76340 35888
rect 76396 35848 76436 35888
rect 76492 35848 76532 35888
rect 76588 35848 76628 35888
rect 76876 35848 76916 35888
rect 76972 35848 77012 35888
rect 77452 35848 77492 35888
rect 77644 35848 77684 35888
rect 77740 35848 77780 35888
rect 78028 35848 78068 35888
rect 57772 35764 57812 35804
rect 58636 35764 58676 35804
rect 66412 35764 66452 35804
rect 55948 35680 55988 35720
rect 56908 35676 56948 35716
rect 58348 35680 58388 35720
rect 61036 35680 61076 35720
rect 61804 35680 61844 35720
rect 63916 35680 63956 35720
rect 64108 35676 64148 35716
rect 65740 35680 65780 35720
rect 68812 35680 68852 35720
rect 71500 35680 71540 35720
rect 72460 35676 72500 35716
rect 74476 35680 74516 35720
rect 74860 35680 74900 35720
rect 76780 35676 76820 35716
rect 77932 35680 77972 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 57484 35344 57524 35384
rect 59404 35348 59444 35388
rect 60172 35344 60212 35384
rect 75724 35344 75764 35384
rect 79468 35344 79508 35384
rect 55084 35260 55124 35300
rect 72844 35260 72884 35300
rect 73324 35260 73364 35300
rect 55468 35176 55508 35216
rect 56332 35176 56372 35216
rect 58348 35176 58388 35216
rect 58732 35176 58772 35216
rect 59212 35176 59252 35216
rect 59308 35176 59348 35216
rect 60268 35176 60308 35216
rect 61132 35176 61172 35216
rect 61228 35176 61268 35216
rect 61420 35176 61460 35216
rect 61612 35176 61652 35216
rect 61996 35176 62036 35216
rect 62860 35176 62900 35216
rect 68236 35176 68276 35216
rect 70252 35176 70292 35216
rect 71116 35176 71156 35216
rect 71500 35176 71540 35216
rect 71692 35176 71732 35216
rect 72076 35176 72116 35216
rect 72940 35176 72980 35216
rect 73036 35176 73076 35216
rect 73132 35176 73172 35216
rect 73708 35176 73748 35216
rect 74572 35176 74612 35216
rect 76876 35176 76916 35216
rect 77068 35176 77108 35216
rect 77452 35176 77492 35216
rect 78316 35176 78356 35216
rect 58444 35092 58484 35132
rect 58636 35092 58676 35132
rect 71788 35092 71828 35132
rect 71980 35092 72020 35132
rect 58540 35008 58580 35048
rect 58924 35008 58964 35048
rect 71884 35008 71924 35048
rect 57484 34924 57524 34964
rect 61420 34924 61460 34964
rect 64012 34924 64052 34964
rect 68140 34924 68180 34964
rect 69100 34924 69140 34964
rect 76780 34924 76820 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 57292 34588 57332 34628
rect 71020 34588 71060 34628
rect 52108 34504 52148 34544
rect 62476 34504 62516 34544
rect 64012 34504 64052 34544
rect 52012 34420 52052 34460
rect 52204 34420 52244 34460
rect 62380 34420 62420 34460
rect 62572 34420 62612 34460
rect 67180 34462 67220 34502
rect 67276 34504 67316 34544
rect 67660 34504 67700 34544
rect 71692 34504 71732 34544
rect 77548 34504 77588 34544
rect 67372 34420 67412 34460
rect 51916 34336 51956 34376
rect 52300 34336 52340 34376
rect 52972 34336 53012 34376
rect 53836 34336 53876 34376
rect 55180 34336 55220 34376
rect 55948 34336 55988 34376
rect 56044 34336 56084 34376
rect 56140 34336 56180 34376
rect 57196 34336 57236 34376
rect 58540 34336 58580 34376
rect 58636 34336 58676 34376
rect 58732 34336 58772 34376
rect 59308 34336 59348 34376
rect 60172 34336 60212 34376
rect 62284 34336 62324 34376
rect 62668 34336 62708 34376
rect 63052 34336 63092 34376
rect 63244 34336 63284 34376
rect 63350 34355 63390 34395
rect 63628 34336 63668 34376
rect 63724 34336 63764 34376
rect 64684 34336 64724 34376
rect 65548 34336 65588 34376
rect 67084 34336 67124 34376
rect 67468 34336 67508 34376
rect 67948 34336 67988 34376
rect 68044 34336 68084 34376
rect 68620 34336 68660 34376
rect 68716 34336 68756 34376
rect 68812 34336 68852 34376
rect 68908 34336 68948 34376
rect 69676 34336 69716 34376
rect 70924 34336 70964 34376
rect 71308 34336 71348 34376
rect 71404 34336 71444 34376
rect 71980 34336 72020 34376
rect 72076 34336 72116 34376
rect 72172 34336 72212 34376
rect 72748 34336 72788 34376
rect 73612 34336 73652 34376
rect 76108 34336 76148 34376
rect 76972 34336 77012 34376
rect 77836 34336 77876 34376
rect 77932 34336 77972 34376
rect 78220 34336 78260 34376
rect 78316 34336 78356 34376
rect 78412 34336 78452 34376
rect 78508 34336 78548 34376
rect 52588 34252 52628 34292
rect 58924 34252 58964 34292
rect 64300 34252 64340 34292
rect 71884 34252 71924 34292
rect 72364 34252 72404 34292
rect 77356 34252 77396 34292
rect 54988 34168 55028 34208
rect 55276 34168 55316 34208
rect 55852 34168 55892 34208
rect 57292 34168 57332 34208
rect 58444 34168 58484 34208
rect 61324 34168 61364 34208
rect 63148 34168 63188 34208
rect 66700 34168 66740 34208
rect 68140 34164 68180 34204
rect 69580 34168 69620 34208
rect 71212 34164 71252 34204
rect 74764 34168 74804 34208
rect 74956 34168 74996 34208
rect 78028 34164 78068 34204
rect 63532 34110 63572 34150
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 52012 33832 52052 33872
rect 55468 33836 55508 33876
rect 58060 33832 58100 33872
rect 59308 33832 59348 33872
rect 59980 33832 60020 33872
rect 61996 33832 62036 33872
rect 63532 33832 63572 33872
rect 64012 33832 64052 33872
rect 64492 33832 64532 33872
rect 67372 33832 67412 33872
rect 70156 33832 70196 33872
rect 71788 33832 71828 33872
rect 72652 33832 72692 33872
rect 76876 33832 76916 33872
rect 51724 33748 51764 33788
rect 50476 33664 50516 33704
rect 51340 33664 51380 33704
rect 51916 33664 51956 33704
rect 53452 33664 53492 33704
rect 54316 33664 54356 33704
rect 54700 33664 54740 33704
rect 55276 33664 55316 33704
rect 55372 33664 55412 33704
rect 55660 33664 55700 33704
rect 56044 33664 56084 33704
rect 56908 33664 56948 33704
rect 59404 33664 59444 33704
rect 59500 33664 59540 33704
rect 59596 33664 59636 33704
rect 59884 33664 59924 33704
rect 63628 33664 63668 33704
rect 64108 33664 64148 33704
rect 64204 33664 64244 33704
rect 64300 33664 64340 33704
rect 64588 33664 64628 33704
rect 64684 33664 64724 33704
rect 64780 33664 64820 33704
rect 66796 33664 66836 33704
rect 66892 33664 66932 33704
rect 66988 33664 67028 33704
rect 67084 33664 67124 33704
rect 67276 33664 67316 33704
rect 67468 33664 67508 33704
rect 67564 33664 67604 33704
rect 67756 33664 67796 33704
rect 68140 33664 68180 33704
rect 69004 33664 69044 33704
rect 71308 33664 71348 33704
rect 71404 33664 71444 33704
rect 71596 33664 71636 33704
rect 71884 33664 71924 33704
rect 71980 33664 72020 33704
rect 72076 33664 72116 33704
rect 72556 33664 72596 33704
rect 74764 33664 74804 33704
rect 76300 33664 76340 33704
rect 76396 33664 76436 33704
rect 76588 33664 76628 33704
rect 76684 33664 76724 33704
rect 76780 33664 76820 33704
rect 77068 33664 77108 33704
rect 77452 33664 77492 33704
rect 77644 33664 77684 33704
rect 77836 33664 77876 33704
rect 77932 33664 77972 33704
rect 78220 33664 78260 33704
rect 61804 33580 61844 33620
rect 77164 33580 77204 33620
rect 77356 33580 77396 33620
rect 77260 33496 77300 33536
rect 77644 33496 77684 33536
rect 49324 33412 49364 33452
rect 52012 33412 52052 33452
rect 52300 33412 52340 33452
rect 54988 33412 55028 33452
rect 58060 33412 58100 33452
rect 59980 33412 60020 33452
rect 61996 33412 62036 33452
rect 71596 33412 71636 33452
rect 72652 33412 72692 33452
rect 74860 33412 74900 33452
rect 78124 33412 78164 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 50956 33076 50996 33116
rect 52108 33076 52148 33116
rect 53836 33076 53876 33116
rect 67852 33076 67892 33116
rect 78796 33076 78836 33116
rect 51916 32992 51956 33032
rect 55276 32992 55316 33032
rect 55852 32992 55892 33032
rect 63532 32992 63572 33032
rect 72844 32992 72884 33032
rect 49996 32908 50036 32948
rect 55180 32908 55220 32948
rect 55372 32908 55412 32948
rect 63820 32908 63860 32948
rect 50476 32824 50516 32864
rect 50572 32824 50612 32864
rect 50764 32824 50804 32864
rect 51244 32824 51284 32864
rect 51340 32824 51380 32864
rect 52588 32824 52628 32864
rect 52876 32824 52916 32864
rect 52972 32824 53012 32864
rect 53068 32824 53108 32864
rect 53164 32824 53204 32864
rect 53356 32824 53396 32864
rect 53452 32824 53492 32864
rect 53548 32824 53588 32864
rect 53644 32824 53684 32864
rect 53836 32824 53876 32864
rect 54028 32824 54068 32864
rect 54124 32824 54164 32864
rect 54604 32824 54644 32864
rect 54700 32824 54740 32864
rect 54796 32824 54836 32864
rect 54892 32824 54932 32864
rect 55084 32824 55124 32864
rect 55468 32824 55508 32864
rect 55852 32782 55892 32822
rect 56044 32824 56084 32864
rect 56140 32824 56180 32864
rect 61324 32824 61364 32864
rect 62188 32824 62228 32864
rect 62764 32824 62804 32864
rect 63148 32824 63188 32864
rect 63244 32824 63284 32864
rect 65836 32824 65876 32864
rect 66700 32824 66740 32864
rect 68044 32824 68084 32864
rect 70156 32824 70196 32864
rect 71020 32824 71060 32864
rect 72460 32824 72500 32864
rect 72556 32824 72596 32864
rect 76780 32824 76820 32864
rect 77644 32824 77684 32864
rect 62572 32740 62612 32780
rect 65452 32740 65492 32780
rect 69772 32740 69812 32780
rect 76396 32740 76436 32780
rect 49804 32656 49844 32696
rect 50668 32656 50708 32696
rect 51436 32652 51476 32692
rect 60172 32656 60212 32696
rect 62860 32656 62900 32696
rect 63052 32652 63092 32692
rect 64012 32656 64052 32696
rect 68140 32656 68180 32696
rect 72172 32656 72212 32696
rect 72364 32598 72404 32638
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 67660 32378 67700 32418
rect 76780 32378 76820 32418
rect 68428 32320 68468 32360
rect 68812 32320 68852 32360
rect 72652 32320 72692 32360
rect 56908 32236 56948 32276
rect 50572 32152 50612 32192
rect 50956 32152 50996 32192
rect 51820 32152 51860 32192
rect 53356 32152 53396 32192
rect 55660 32152 55700 32192
rect 56524 32152 56564 32192
rect 57196 32152 57236 32192
rect 57580 32152 57620 32192
rect 58924 32152 58964 32192
rect 59788 32152 59828 32192
rect 60172 32152 60212 32192
rect 60364 32152 60404 32192
rect 60748 32152 60788 32192
rect 61132 32152 61172 32192
rect 61516 32152 61556 32192
rect 61708 32152 61748 32192
rect 61804 32152 61844 32192
rect 62764 32152 62804 32192
rect 63148 32152 63188 32192
rect 63340 32152 63380 32192
rect 63724 32152 63764 32192
rect 64588 32152 64628 32192
rect 66412 32152 66452 32192
rect 66796 32152 66836 32192
rect 67468 32152 67508 32192
rect 67564 32152 67604 32192
rect 71500 32152 71540 32192
rect 71884 32152 71924 32192
rect 72076 32152 72116 32192
rect 72268 32152 72308 32192
rect 72364 32152 72404 32192
rect 72556 32152 72596 32192
rect 72844 32152 72884 32192
rect 73228 32152 73268 32192
rect 74092 32152 74132 32192
rect 76588 32152 76628 32192
rect 76684 32152 76724 32192
rect 76972 32152 77012 32192
rect 77356 32152 77396 32192
rect 78220 32152 78260 32192
rect 57292 32068 57332 32108
rect 57484 32068 57524 32108
rect 60844 32068 60884 32108
rect 61036 32068 61076 32108
rect 62860 32068 62900 32108
rect 63052 32068 63092 32108
rect 66508 32068 66548 32108
rect 66700 32068 66740 32108
rect 68620 32068 68660 32108
rect 69004 32068 69044 32108
rect 71596 32068 71636 32108
rect 71788 32068 71828 32108
rect 57388 31984 57428 32024
rect 60940 31984 60980 32024
rect 61516 31984 61556 32024
rect 62956 31984 62996 32024
rect 66604 31984 66644 32024
rect 71692 31984 71732 32024
rect 52972 31900 53012 31940
rect 54508 31900 54548 31940
rect 57772 31900 57812 31940
rect 60460 31900 60500 31940
rect 65740 31900 65780 31940
rect 67180 31900 67220 31940
rect 68428 31900 68468 31940
rect 72076 31900 72116 31940
rect 75244 31900 75284 31940
rect 76300 31900 76340 31940
rect 79372 31900 79412 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 50188 31564 50228 31604
rect 51820 31564 51860 31604
rect 54604 31564 54644 31604
rect 57196 31564 57236 31604
rect 57868 31564 57908 31604
rect 58636 31564 58676 31604
rect 66220 31564 66260 31604
rect 71596 31564 71636 31604
rect 50572 31480 50612 31520
rect 50956 31480 50996 31520
rect 52492 31480 52532 31520
rect 60844 31480 60884 31520
rect 70444 31480 70484 31520
rect 76684 31480 76724 31520
rect 77068 31480 77108 31520
rect 49996 31396 50036 31436
rect 50476 31396 50516 31436
rect 50668 31396 50708 31436
rect 52396 31396 52436 31436
rect 52588 31396 52628 31436
rect 71404 31396 71444 31436
rect 73228 31396 73268 31436
rect 76588 31396 76628 31436
rect 50380 31312 50420 31352
rect 50764 31312 50804 31352
rect 51244 31312 51284 31352
rect 51340 31312 51380 31352
rect 51820 31323 51860 31363
rect 52012 31312 52052 31352
rect 52108 31312 52148 31352
rect 52300 31312 52340 31352
rect 52684 31312 52724 31352
rect 52972 31312 53012 31352
rect 55276 31312 55316 31352
rect 55372 31312 55412 31352
rect 57100 31312 57140 31352
rect 57484 31312 57524 31352
rect 57580 31312 57620 31352
rect 58060 31312 58100 31352
rect 58156 31312 58196 31352
rect 58252 31312 58292 31352
rect 58348 31312 58388 31352
rect 58636 31312 58676 31352
rect 58828 31312 58868 31352
rect 58924 31312 58964 31352
rect 59212 31312 59252 31352
rect 61132 31312 61172 31352
rect 61228 31312 61268 31352
rect 61516 31312 61556 31352
rect 61612 31312 61652 31352
rect 61708 31312 61748 31352
rect 61804 31312 61844 31352
rect 63340 31354 63380 31394
rect 76780 31396 76820 31436
rect 63244 31312 63284 31352
rect 63436 31312 63476 31352
rect 63532 31312 63572 31352
rect 63724 31312 63764 31352
rect 63820 31312 63860 31352
rect 63916 31312 63956 31352
rect 64012 31312 64052 31352
rect 66220 31312 66260 31352
rect 66412 31312 66452 31352
rect 66508 31312 66548 31352
rect 67180 31312 67220 31352
rect 67276 31312 67316 31352
rect 67372 31312 67412 31352
rect 67948 31312 67988 31352
rect 68812 31312 68852 31352
rect 71788 31312 71828 31352
rect 72364 31312 72404 31352
rect 72460 31312 72500 31352
rect 72556 31312 72596 31352
rect 72748 31312 72788 31352
rect 72844 31312 72884 31352
rect 72940 31312 72980 31352
rect 73036 31312 73076 31352
rect 73612 31312 73652 31352
rect 73708 31312 73748 31352
rect 73804 31291 73844 31331
rect 73900 31312 73940 31352
rect 74476 31312 74516 31352
rect 76012 31312 76052 31352
rect 76108 31312 76148 31352
rect 76204 31312 76244 31352
rect 76492 31312 76532 31352
rect 76876 31312 76916 31352
rect 77068 31312 77108 31352
rect 77260 31312 77300 31352
rect 77356 31312 77396 31352
rect 77548 31312 77588 31352
rect 77644 31312 77684 31352
rect 77740 31312 77780 31352
rect 77836 31312 77876 31352
rect 78124 31312 78164 31352
rect 67564 31228 67604 31268
rect 57196 31144 57236 31184
rect 57772 31186 57812 31226
rect 57388 31140 57428 31180
rect 59116 31144 59156 31184
rect 61324 31140 61364 31180
rect 67084 31144 67124 31184
rect 69964 31144 70004 31184
rect 71596 31144 71636 31184
rect 71884 31144 71924 31184
rect 72268 31144 72308 31184
rect 73420 31144 73460 31184
rect 74380 31144 74420 31184
rect 76300 31144 76340 31184
rect 78028 31144 78068 31184
rect 51436 31086 51476 31126
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 56044 30808 56084 30848
rect 56428 30808 56468 30848
rect 57676 30808 57716 30848
rect 60844 30808 60884 30848
rect 66412 30808 66452 30848
rect 68428 30808 68468 30848
rect 69100 30808 69140 30848
rect 74860 30808 74900 30848
rect 77452 30808 77492 30848
rect 53644 30724 53684 30764
rect 57868 30724 57908 30764
rect 61324 30724 61364 30764
rect 72460 30724 72500 30764
rect 48076 30640 48116 30680
rect 48460 30640 48500 30680
rect 50188 30640 50228 30680
rect 50284 30640 50324 30680
rect 50380 30640 50420 30680
rect 50476 30640 50516 30680
rect 50668 30640 50708 30680
rect 51052 30640 51092 30680
rect 51916 30640 51956 30680
rect 54028 30640 54068 30680
rect 54892 30640 54932 30680
rect 57388 30640 57428 30680
rect 57484 30640 57524 30680
rect 57580 30640 57620 30680
rect 58252 30640 58292 30680
rect 59116 30640 59156 30680
rect 60940 30640 60980 30680
rect 61036 30640 61076 30680
rect 61132 30640 61172 30680
rect 61708 30640 61748 30680
rect 62572 30640 62612 30680
rect 64012 30640 64052 30680
rect 64396 30640 64436 30680
rect 65260 30640 65300 30680
rect 66604 30640 66644 30680
rect 66700 30640 66740 30680
rect 66796 30640 66836 30680
rect 66892 30640 66932 30680
rect 67084 30640 67124 30680
rect 68140 30640 68180 30680
rect 68236 30640 68276 30680
rect 68332 30640 68372 30680
rect 69004 30640 69044 30680
rect 70444 30640 70484 30680
rect 71308 30640 71348 30680
rect 71692 30640 71732 30680
rect 71884 30640 71924 30680
rect 72268 30640 72308 30680
rect 72844 30640 72884 30680
rect 73708 30640 73748 30680
rect 75052 30640 75092 30680
rect 75436 30640 75476 30680
rect 76300 30640 76340 30680
rect 77644 30640 77684 30680
rect 48172 30556 48212 30596
rect 48364 30556 48404 30596
rect 56236 30556 56276 30596
rect 71980 30556 72020 30596
rect 72172 30556 72212 30596
rect 48268 30472 48308 30512
rect 72076 30472 72116 30512
rect 53068 30388 53108 30428
rect 56044 30388 56084 30428
rect 56428 30388 56468 30428
rect 60268 30388 60308 30428
rect 63724 30388 63764 30428
rect 67180 30388 67220 30428
rect 69100 30388 69140 30428
rect 69292 30388 69332 30428
rect 77740 30388 77780 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 53932 30052 53972 30092
rect 55468 30052 55508 30092
rect 59212 30052 59252 30092
rect 59596 30052 59636 30092
rect 60940 30052 60980 30092
rect 61324 30052 61364 30092
rect 70924 30052 70964 30092
rect 71788 30052 71828 30092
rect 72460 30052 72500 30092
rect 72652 30052 72692 30092
rect 73612 30052 73652 30092
rect 74092 30052 74132 30092
rect 61900 29968 61940 30008
rect 65068 29968 65108 30008
rect 65452 29968 65492 30008
rect 65932 29968 65972 30008
rect 75628 29968 75668 30008
rect 76012 29968 76052 30008
rect 76396 29968 76436 30008
rect 40396 29884 40436 29924
rect 48076 29884 48116 29924
rect 51148 29884 51188 29924
rect 55084 29884 55124 29924
rect 55660 29884 55700 29924
rect 59404 29884 59444 29924
rect 59788 29884 59828 29924
rect 60748 29884 60788 29924
rect 61132 29884 61172 29924
rect 61708 29884 61748 29924
rect 62092 29884 62132 29924
rect 46540 29800 46580 29840
rect 47404 29800 47444 29840
rect 47788 29800 47828 29840
rect 47980 29800 48020 29840
rect 48748 29800 48788 29840
rect 49612 29800 49652 29840
rect 51436 29800 51476 29840
rect 51532 29800 51572 29840
rect 51628 29800 51668 29840
rect 51724 29800 51764 29840
rect 52204 29800 52244 29840
rect 54220 29800 54260 29840
rect 54316 29800 54356 29840
rect 54604 29800 54644 29840
rect 54700 29800 54740 29840
rect 54796 29800 54836 29840
rect 54892 29800 54932 29840
rect 56044 29800 56084 29840
rect 56140 29800 56180 29840
rect 56332 29800 56372 29840
rect 57004 29800 57044 29840
rect 57868 29800 57908 29840
rect 64780 29800 64820 29840
rect 64876 29800 64916 29840
rect 65068 29800 65108 29840
rect 65260 29842 65300 29882
rect 65356 29884 65396 29924
rect 65548 29884 65588 29924
rect 70732 29884 70772 29924
rect 71596 29884 71636 29924
rect 72844 29884 72884 29924
rect 65644 29800 65684 29840
rect 66220 29800 66260 29840
rect 66316 29800 66356 29840
rect 67084 29800 67124 29840
rect 67948 29800 67988 29840
rect 71116 29800 71156 29840
rect 71308 29800 71348 29840
rect 71404 29800 71444 29840
rect 72076 29800 72116 29840
rect 72172 29800 72212 29840
rect 73132 29800 73172 29840
rect 73228 29800 73268 29840
rect 73324 29800 73364 29840
rect 73420 29845 73460 29885
rect 73804 29884 73844 29924
rect 75436 29884 75476 29924
rect 75916 29884 75956 29924
rect 76108 29884 76148 29924
rect 73996 29800 74036 29840
rect 75820 29800 75860 29840
rect 76204 29800 76244 29840
rect 76684 29800 76724 29840
rect 76780 29800 76820 29840
rect 77452 29800 77492 29840
rect 78316 29800 78356 29840
rect 48364 29716 48404 29756
rect 56620 29716 56660 29756
rect 66700 29716 66740 29756
rect 77068 29716 77108 29756
rect 40588 29632 40628 29672
rect 45388 29632 45428 29672
rect 50764 29632 50804 29672
rect 50956 29632 50996 29672
rect 52108 29632 52148 29672
rect 54412 29628 54452 29668
rect 55276 29632 55316 29672
rect 56236 29632 56276 29672
rect 59020 29632 59060 29672
rect 59212 29632 59252 29672
rect 60940 29632 60980 29672
rect 61324 29632 61364 29672
rect 61516 29632 61556 29672
rect 66412 29628 66452 29668
rect 69100 29632 69140 29672
rect 71212 29632 71252 29672
rect 71788 29632 71828 29672
rect 71980 29628 72020 29668
rect 72652 29632 72692 29672
rect 74092 29632 74132 29672
rect 76876 29628 76916 29668
rect 79468 29632 79508 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 47980 29354 48020 29394
rect 39916 29296 39956 29336
rect 46732 29296 46772 29336
rect 51052 29296 51092 29336
rect 51820 29296 51860 29336
rect 57484 29300 57524 29340
rect 58156 29296 58196 29336
rect 65452 29296 65492 29336
rect 66316 29296 66356 29336
rect 66988 29296 67028 29336
rect 71116 29296 71156 29336
rect 71308 29300 71348 29340
rect 76588 29296 76628 29336
rect 77452 29296 77492 29336
rect 48652 29212 48692 29252
rect 76972 29212 77012 29252
rect 42604 29128 42644 29168
rect 42700 29128 42740 29168
rect 42796 29128 42836 29168
rect 42892 29128 42932 29168
rect 43084 29128 43124 29168
rect 43276 29128 43316 29168
rect 43180 29086 43220 29126
rect 43372 29128 43412 29168
rect 46636 29128 46676 29168
rect 46828 29128 46868 29168
rect 46924 29128 46964 29168
rect 47116 29128 47156 29168
rect 47500 29128 47540 29168
rect 48076 29128 48116 29168
rect 48172 29128 48212 29168
rect 48748 29128 48788 29168
rect 48844 29128 48884 29168
rect 48940 29128 48980 29168
rect 49708 29128 49748 29168
rect 50572 29128 50612 29168
rect 50956 29128 50996 29168
rect 51148 29128 51188 29168
rect 51244 29128 51284 29168
rect 52204 29128 52244 29168
rect 53164 29128 53204 29168
rect 53356 29128 53396 29168
rect 39724 29044 39764 29084
rect 40108 29044 40148 29084
rect 40684 29044 40724 29084
rect 47212 29044 47252 29084
rect 53260 29086 53300 29126
rect 53452 29128 53492 29168
rect 53644 29128 53684 29168
rect 54028 29128 54068 29168
rect 54892 29128 54932 29168
rect 56428 29128 56468 29168
rect 56812 29128 56852 29168
rect 57292 29128 57332 29168
rect 57388 29128 57428 29168
rect 58252 29128 58292 29168
rect 58828 29128 58868 29168
rect 58924 29128 58964 29168
rect 59116 29128 59156 29168
rect 59308 29128 59348 29168
rect 59692 29128 59732 29168
rect 60556 29128 60596 29168
rect 61900 29128 61940 29168
rect 62284 29128 62324 29168
rect 63148 29128 63188 29168
rect 64492 29128 64532 29168
rect 64876 29128 64916 29168
rect 65836 29128 65876 29168
rect 65932 29128 65972 29168
rect 66028 29128 66068 29168
rect 66124 29128 66164 29168
rect 66412 29128 66452 29168
rect 66508 29128 66548 29168
rect 66604 29128 66644 29168
rect 67372 29128 67412 29168
rect 69580 29128 69620 29168
rect 70444 29128 70484 29168
rect 70828 29128 70868 29168
rect 71020 29128 71060 29168
rect 71404 29128 71444 29168
rect 71500 29128 71540 29168
rect 72172 29128 72212 29168
rect 72556 29128 72596 29168
rect 73453 29128 73493 29168
rect 76492 29128 76532 29168
rect 76684 29128 76724 29168
rect 76780 29128 76820 29168
rect 77068 29120 77108 29160
rect 77260 29128 77300 29168
rect 47404 29044 47444 29084
rect 49516 29044 49556 29084
rect 51628 29044 51668 29084
rect 52012 29044 52052 29084
rect 56524 29044 56564 29084
rect 56716 29044 56756 29084
rect 64588 29044 64628 29084
rect 77164 29086 77204 29126
rect 77548 29128 77588 29168
rect 77644 29128 77684 29168
rect 77740 29128 77780 29168
rect 78028 29128 78068 29168
rect 64780 29044 64820 29084
rect 65260 29044 65300 29084
rect 66796 29044 66836 29084
rect 47308 28960 47348 29000
rect 48460 28960 48500 29000
rect 51436 28960 51476 29000
rect 56620 28960 56660 29000
rect 57004 28960 57044 29000
rect 64684 28960 64724 29000
rect 40300 28876 40340 28916
rect 40492 28876 40532 28916
rect 49324 28876 49364 28916
rect 49996 28876 50036 28916
rect 50380 28876 50420 28916
rect 52300 28876 52340 28916
rect 56044 28876 56084 28916
rect 59116 28876 59156 28916
rect 61708 28876 61748 28916
rect 64300 28876 64340 28916
rect 67468 28876 67508 28916
rect 68428 28876 68468 28916
rect 71116 28876 71156 28916
rect 71788 28876 71828 28916
rect 74572 28876 74612 28916
rect 77932 28876 77972 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 45196 28540 45236 28580
rect 49708 28540 49748 28580
rect 55180 28540 55220 28580
rect 65452 28540 65492 28580
rect 65740 28540 65780 28580
rect 72268 28540 72308 28580
rect 76876 28540 76916 28580
rect 42412 28456 42452 28496
rect 52780 28456 52820 28496
rect 59980 28456 60020 28496
rect 61324 28456 61364 28496
rect 70732 28456 70772 28496
rect 71116 28456 71156 28496
rect 77068 28456 77108 28496
rect 42316 28372 42356 28412
rect 42508 28372 42548 28412
rect 59884 28372 59924 28412
rect 40780 28288 40820 28328
rect 41644 28288 41684 28328
rect 42028 28288 42068 28328
rect 42220 28288 42260 28328
rect 42604 28288 42644 28328
rect 42796 28288 42836 28328
rect 43180 28324 43220 28364
rect 44044 28288 44084 28328
rect 45388 28288 45428 28328
rect 45772 28288 45812 28328
rect 46636 28288 46676 28328
rect 48172 28288 48212 28328
rect 48268 28288 48308 28328
rect 48364 28288 48404 28328
rect 52492 28330 52532 28370
rect 60076 28372 60116 28412
rect 69100 28372 69140 28412
rect 71020 28372 71060 28412
rect 71212 28372 71252 28412
rect 72460 28372 72500 28412
rect 48460 28288 48500 28328
rect 50860 28288 50900 28328
rect 51724 28288 51764 28328
rect 52396 28288 52436 28328
rect 53068 28288 53108 28328
rect 53164 28288 53204 28328
rect 53260 28288 53300 28328
rect 55084 28288 55124 28328
rect 56140 28288 56180 28328
rect 56236 28288 56276 28328
rect 56332 28288 56372 28328
rect 57004 28288 57044 28328
rect 57868 28288 57908 28328
rect 59788 28288 59828 28328
rect 60172 28288 60212 28328
rect 60556 28288 60596 28328
rect 60652 28288 60692 28328
rect 60940 28288 60980 28328
rect 61036 28288 61076 28328
rect 61516 28288 61556 28328
rect 61612 28288 61652 28328
rect 61708 28288 61748 28328
rect 61804 28288 61844 28328
rect 61996 28288 62036 28328
rect 62092 28288 62132 28328
rect 62188 28288 62228 28328
rect 62284 28288 62324 28328
rect 62860 28288 62900 28328
rect 63052 28288 63092 28328
rect 63436 28288 63476 28328
rect 64300 28288 64340 28328
rect 65644 28288 65684 28328
rect 66316 28288 66356 28328
rect 67180 28288 67220 28328
rect 70444 28288 70484 28328
rect 70540 28302 70580 28342
rect 70732 28299 70772 28339
rect 70924 28288 70964 28328
rect 71308 28288 71348 28328
rect 71788 28288 71828 28328
rect 71884 28288 71924 28328
rect 71980 28288 72020 28328
rect 72076 28288 72116 28328
rect 72748 28288 72788 28328
rect 72844 28288 72884 28328
rect 72940 28288 72980 28328
rect 73036 28288 73076 28328
rect 73708 28288 73748 28328
rect 74860 28288 74900 28328
rect 75724 28288 75764 28328
rect 77356 28288 77396 28328
rect 77452 28288 77492 28328
rect 77740 28288 77780 28328
rect 52108 28204 52148 28244
rect 56428 28204 56468 28244
rect 56620 28204 56660 28244
rect 65932 28204 65972 28244
rect 74476 28204 74516 28244
rect 39628 28120 39668 28160
rect 45196 28120 45236 28160
rect 47788 28120 47828 28160
rect 52300 28116 52340 28156
rect 52972 28120 53012 28160
rect 55180 28120 55220 28160
rect 59020 28120 59060 28160
rect 60844 28116 60884 28156
rect 62764 28120 62804 28160
rect 65740 28120 65780 28160
rect 68332 28120 68372 28160
rect 68908 28120 68948 28160
rect 73612 28120 73652 28160
rect 77836 28120 77876 28160
rect 77548 28062 77588 28102
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 65548 27842 65588 27882
rect 42220 27784 42260 27824
rect 42508 27788 42548 27828
rect 46060 27784 46100 27824
rect 47308 27784 47348 27824
rect 47596 27788 47636 27828
rect 57484 27784 57524 27824
rect 59404 27784 59444 27824
rect 47980 27742 48020 27782
rect 66028 27784 66068 27824
rect 71116 27784 71156 27824
rect 71500 27788 71540 27828
rect 40588 27616 40628 27656
rect 40780 27616 40820 27656
rect 40876 27616 40916 27656
rect 42124 27616 42164 27656
rect 42604 27616 42644 27656
rect 42700 27616 42740 27656
rect 43180 27658 43220 27698
rect 53164 27700 53204 27740
rect 43372 27616 43412 27656
rect 43468 27616 43508 27656
rect 43660 27616 43700 27656
rect 44044 27616 44084 27656
rect 47404 27616 47444 27656
rect 47692 27616 47732 27656
rect 47788 27616 47828 27656
rect 48268 27616 48308 27656
rect 48364 27616 48404 27656
rect 48460 27616 48500 27656
rect 48556 27616 48596 27656
rect 48748 27616 48788 27656
rect 49132 27616 49172 27656
rect 49996 27616 50036 27656
rect 52012 27616 52052 27656
rect 52396 27616 52436 27656
rect 52588 27605 52628 27645
rect 52780 27616 52820 27656
rect 52876 27616 52916 27656
rect 53548 27616 53588 27656
rect 54412 27616 54452 27656
rect 57580 27616 57620 27656
rect 57676 27616 57716 27656
rect 57772 27616 57812 27656
rect 58060 27616 58100 27656
rect 60652 27616 60692 27656
rect 61036 27616 61076 27656
rect 61228 27616 61268 27656
rect 61420 27616 61460 27656
rect 61516 27616 61556 27656
rect 62380 27616 62420 27656
rect 62764 27616 62804 27656
rect 63628 27616 63668 27656
rect 65356 27616 65396 27656
rect 65452 27616 65492 27656
rect 65740 27616 65780 27656
rect 65836 27616 65876 27656
rect 65932 27616 65972 27656
rect 66508 27616 66548 27656
rect 69580 27616 69620 27656
rect 70444 27616 70484 27656
rect 70828 27616 70868 27656
rect 71212 27616 71252 27656
rect 71596 27616 71636 27656
rect 71692 27616 71732 27656
rect 75724 27616 75764 27656
rect 75916 27616 75956 27656
rect 76012 27616 76052 27656
rect 76204 27616 76244 27656
rect 76588 27616 76628 27656
rect 76876 27616 76916 27656
rect 77068 27616 77108 27656
rect 77452 27616 77492 27656
rect 78316 27616 78356 27656
rect 40396 27532 40436 27572
rect 44236 27532 44276 27572
rect 45868 27532 45908 27572
rect 52108 27532 52148 27572
rect 52300 27532 52340 27572
rect 58828 27532 58868 27572
rect 59212 27532 59252 27572
rect 59596 27532 59636 27572
rect 59980 27532 60020 27572
rect 60748 27532 60788 27572
rect 60940 27532 60980 27572
rect 68428 27532 68468 27572
rect 76300 27532 76340 27572
rect 76492 27532 76532 27572
rect 42988 27448 43028 27488
rect 43180 27448 43220 27488
rect 43756 27448 43796 27488
rect 52204 27448 52244 27488
rect 52588 27448 52628 27488
rect 60844 27448 60884 27488
rect 65068 27448 65108 27488
rect 76396 27448 76436 27488
rect 40204 27364 40244 27404
rect 40588 27364 40628 27404
rect 43948 27364 43988 27404
rect 44428 27364 44468 27404
rect 46060 27364 46100 27404
rect 51148 27364 51188 27404
rect 55564 27364 55604 27404
rect 58156 27364 58196 27404
rect 59020 27364 59060 27404
rect 59788 27364 59828 27404
rect 60172 27364 60212 27404
rect 61228 27364 61268 27404
rect 64780 27364 64820 27404
rect 66604 27364 66644 27404
rect 71116 27364 71156 27404
rect 71980 27364 72020 27404
rect 75724 27364 75764 27404
rect 76780 27364 76820 27404
rect 79468 27364 79508 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 44524 27028 44564 27068
rect 49132 27028 49172 27068
rect 50860 27028 50900 27068
rect 61420 27028 61460 27068
rect 61900 27028 61940 27068
rect 64396 27028 64436 27068
rect 76972 27028 77012 27068
rect 78124 27028 78164 27068
rect 39916 26944 39956 26984
rect 47788 26944 47828 26984
rect 63916 26944 63956 26984
rect 71020 26944 71060 26984
rect 39820 26860 39860 26900
rect 40012 26860 40052 26900
rect 40780 26860 40820 26900
rect 44908 26860 44948 26900
rect 47692 26860 47732 26900
rect 47884 26860 47924 26900
rect 58444 26860 58484 26900
rect 61612 26860 61652 26900
rect 63820 26860 63860 26900
rect 64012 26860 64052 26900
rect 70924 26860 70964 26900
rect 71116 26860 71156 26900
rect 78316 26860 78356 26900
rect 39436 26776 39476 26816
rect 39532 26776 39572 26816
rect 39724 26776 39764 26816
rect 40108 26776 40148 26816
rect 40300 26755 40340 26795
rect 40396 26776 40436 26816
rect 40492 26776 40532 26816
rect 42508 26776 42548 26816
rect 43372 26776 43412 26816
rect 47116 26776 47156 26816
rect 47308 26776 47348 26816
rect 47404 26776 47444 26816
rect 47596 26776 47636 26816
rect 47980 26776 48020 26816
rect 48172 26776 48212 26816
rect 48268 26776 48308 26816
rect 48364 26776 48404 26816
rect 48460 26776 48500 26816
rect 49036 26776 49076 26816
rect 52012 26776 52052 26816
rect 52876 26776 52916 26816
rect 53452 26776 53492 26816
rect 53548 26776 53588 26816
rect 53644 26776 53684 26816
rect 53740 26776 53780 26816
rect 55180 26776 55220 26816
rect 56044 26776 56084 26816
rect 59980 26776 60020 26816
rect 60844 26776 60884 26816
rect 61228 26776 61268 26816
rect 61804 26776 61844 26816
rect 63724 26776 63764 26816
rect 64108 26776 64148 26816
rect 64396 26776 64436 26816
rect 64588 26776 64628 26816
rect 64684 26776 64724 26816
rect 64876 26776 64916 26816
rect 64972 26776 65012 26816
rect 69196 26776 69236 26816
rect 70060 26776 70100 26816
rect 70828 26776 70868 26816
rect 71212 26776 71252 26816
rect 71404 26776 71444 26816
rect 71500 26776 71540 26816
rect 71692 26776 71732 26816
rect 72364 26776 72404 26816
rect 73228 26776 73268 26816
rect 74956 26776 74996 26816
rect 75820 26776 75860 26816
rect 77164 26776 77204 26816
rect 77260 26776 77300 26816
rect 77356 26776 77396 26816
rect 77452 26776 77492 26816
rect 77644 26776 77684 26816
rect 77740 26776 77780 26816
rect 77836 26776 77876 26816
rect 77932 26776 77972 26816
rect 78604 26776 78644 26816
rect 42124 26692 42164 26732
rect 47212 26692 47252 26732
rect 53260 26692 53300 26732
rect 56428 26692 56468 26732
rect 70444 26692 70484 26732
rect 71980 26692 72020 26732
rect 74572 26692 74612 26732
rect 40588 26608 40628 26648
rect 40972 26608 41012 26648
rect 44716 26608 44756 26648
rect 49132 26608 49172 26648
rect 54028 26608 54068 26648
rect 58636 26608 58676 26648
rect 58828 26608 58868 26648
rect 61900 26608 61940 26648
rect 68044 26608 68084 26648
rect 71596 26608 71636 26648
rect 74380 26608 74420 26648
rect 78508 26608 78548 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 61420 26330 61460 26370
rect 844 26272 884 26312
rect 42412 26272 42452 26312
rect 44140 26276 44180 26316
rect 54604 26272 54644 26312
rect 69964 26272 70004 26312
rect 71212 26272 71252 26312
rect 71788 26272 71828 26312
rect 72652 26272 72692 26312
rect 76684 26276 76724 26316
rect 39340 26188 39380 26228
rect 43084 26188 43124 26228
rect 38092 26104 38132 26144
rect 38956 26104 38996 26144
rect 39532 26104 39572 26144
rect 39628 26104 39668 26144
rect 39724 26104 39764 26144
rect 39820 26104 39860 26144
rect 40012 26104 40052 26144
rect 40396 26104 40436 26144
rect 41260 26104 41300 26144
rect 42988 26104 43028 26144
rect 43180 26146 43220 26186
rect 47788 26188 47828 26228
rect 59116 26188 59156 26228
rect 43276 26104 43316 26144
rect 43468 26104 43508 26144
rect 43852 26104 43892 26144
rect 44236 26104 44276 26144
rect 44332 26104 44372 26144
rect 44812 26104 44852 26144
rect 45196 26104 45236 26144
rect 46060 26104 46100 26144
rect 48172 26104 48212 26144
rect 49036 26104 49076 26144
rect 53164 26104 53204 26144
rect 53356 26104 53396 26144
rect 53452 26104 53492 26144
rect 53644 26104 53684 26144
rect 54028 26104 54068 26144
rect 54796 26104 54836 26144
rect 54988 26104 55028 26144
rect 55084 26104 55124 26144
rect 55852 26104 55892 26144
rect 56140 26104 56180 26144
rect 56524 26104 56564 26144
rect 57868 26104 57908 26144
rect 58732 26104 58772 26144
rect 59308 26104 59348 26144
rect 59692 26104 59732 26144
rect 59980 26104 60020 26144
rect 60172 26104 60212 26144
rect 60268 26104 60308 26144
rect 61228 26104 61268 26144
rect 61324 26104 61364 26144
rect 61708 26104 61748 26144
rect 61804 26104 61844 26144
rect 61900 26104 61940 26144
rect 61996 26104 62036 26144
rect 64396 26104 64436 26144
rect 65260 26104 65300 26144
rect 65644 26104 65684 26144
rect 66124 26104 66164 26144
rect 66508 26104 66548 26144
rect 67372 26104 67412 26144
rect 68812 26104 68852 26144
rect 69196 26104 69236 26144
rect 69484 26104 69524 26144
rect 70540 26146 70580 26186
rect 69676 26104 69716 26144
rect 69772 26104 69812 26144
rect 70924 26104 70964 26144
rect 71116 26104 71156 26144
rect 71884 26104 71924 26144
rect 71980 26104 72020 26144
rect 72076 26104 72116 26144
rect 72748 26104 72788 26144
rect 72844 26104 72884 26144
rect 72940 26104 72980 26144
rect 73324 26104 73364 26144
rect 75628 26104 75668 26144
rect 76012 26104 76052 26144
rect 76492 26104 76532 26144
rect 76588 26104 76628 26144
rect 76876 26104 76916 26144
rect 77260 26104 77300 26144
rect 78124 26104 78164 26144
rect 652 26020 692 26060
rect 42796 26020 42836 26060
rect 43564 26020 43604 26060
rect 43756 26020 43796 26060
rect 53740 26020 53780 26060
rect 53932 26020 53972 26060
rect 54412 26020 54452 26060
rect 56236 26020 56276 26060
rect 56428 26020 56468 26060
rect 59404 26020 59444 26060
rect 59596 26020 59636 26060
rect 60460 26020 60500 26060
rect 68908 26020 68948 26060
rect 69100 26020 69140 26060
rect 70156 26020 70196 26060
rect 70636 26020 70676 26060
rect 70828 26020 70868 26060
rect 75244 26020 75284 26060
rect 75724 26020 75764 26060
rect 75916 26020 75956 26060
rect 36940 25936 36980 25976
rect 43660 25936 43700 25976
rect 47212 25936 47252 25976
rect 53836 25936 53876 25976
rect 54796 25936 54836 25976
rect 55948 25936 55988 25976
rect 56332 25936 56372 25976
rect 59500 25936 59540 25976
rect 59980 25936 60020 25976
rect 60652 25936 60692 25976
rect 60940 25936 60980 25976
rect 63244 25936 63284 25976
rect 69004 25936 69044 25976
rect 69484 25936 69524 25976
rect 70732 25936 70772 25976
rect 73420 25936 73460 25976
rect 75436 25936 75476 25976
rect 75820 25936 75860 25976
rect 76204 25936 76244 25976
rect 42604 25852 42644 25892
rect 44620 25852 44660 25892
rect 50188 25852 50228 25892
rect 53068 25852 53108 25892
rect 54604 25852 54644 25892
rect 56716 25852 56756 25892
rect 68524 25852 68564 25892
rect 79276 25852 79316 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 39724 25516 39764 25556
rect 40780 25516 40820 25556
rect 41932 25516 41972 25556
rect 42316 25516 42356 25556
rect 49132 25516 49172 25556
rect 50764 25516 50804 25556
rect 52300 25516 52340 25556
rect 54124 25516 54164 25556
rect 57004 25516 57044 25556
rect 57484 25516 57524 25556
rect 60364 25516 60404 25556
rect 60556 25516 60596 25556
rect 64588 25516 64628 25556
rect 68716 25516 68756 25556
rect 70252 25516 70292 25556
rect 76108 25516 76148 25556
rect 43276 25432 43316 25472
rect 43660 25432 43700 25472
rect 47788 25432 47828 25472
rect 58924 25432 58964 25472
rect 59116 25432 59156 25472
rect 63724 25432 63764 25472
rect 65932 25432 65972 25472
rect 66316 25432 66356 25472
rect 67180 25432 67220 25472
rect 69004 25432 69044 25472
rect 71500 25432 71540 25472
rect 652 25348 692 25388
rect 39532 25348 39572 25388
rect 40588 25348 40628 25388
rect 41740 25348 41780 25388
rect 42124 25348 42164 25388
rect 42508 25348 42548 25388
rect 43084 25348 43124 25388
rect 43468 25348 43508 25388
rect 43852 25348 43892 25388
rect 50572 25348 50612 25388
rect 51244 25348 51284 25388
rect 52108 25348 52148 25388
rect 58732 25348 58772 25388
rect 59980 25348 60020 25388
rect 60172 25348 60212 25388
rect 60748 25348 60788 25388
rect 65836 25348 65876 25388
rect 66028 25348 66068 25388
rect 69868 25348 69908 25388
rect 70060 25348 70100 25388
rect 37708 25264 37748 25304
rect 38380 25264 38420 25304
rect 38572 25264 38612 25304
rect 38668 25264 38708 25304
rect 40012 25264 40052 25304
rect 40108 25264 40148 25304
rect 40972 25264 41012 25304
rect 44428 25264 44468 25304
rect 44524 25264 44564 25304
rect 44620 25264 44660 25304
rect 44716 25264 44756 25304
rect 44908 25264 44948 25304
rect 45004 25264 45044 25304
rect 45100 25264 45140 25304
rect 45196 25264 45236 25304
rect 45676 25264 45716 25304
rect 48076 25264 48116 25304
rect 48172 25264 48212 25304
rect 49228 25264 49268 25304
rect 50092 25264 50132 25304
rect 50188 25264 50228 25304
rect 50380 25264 50420 25304
rect 51052 25264 51092 25304
rect 51724 25264 51764 25304
rect 51820 25264 51860 25304
rect 51916 25264 51956 25304
rect 53740 25264 53780 25304
rect 53836 25264 53876 25304
rect 54316 25264 54356 25304
rect 54412 25264 54452 25304
rect 54508 25264 54548 25304
rect 54604 25264 54644 25304
rect 56620 25264 56660 25304
rect 56716 25264 56756 25304
rect 57484 25264 57524 25304
rect 57676 25264 57716 25304
rect 57772 25264 57812 25304
rect 58444 25264 58484 25304
rect 59404 25264 59444 25304
rect 59500 25264 59540 25304
rect 61324 25264 61364 25304
rect 62188 25264 62228 25304
rect 64012 25264 64052 25304
rect 64108 25264 64148 25304
rect 45580 25180 45620 25220
rect 844 25096 884 25136
rect 37804 25096 37844 25136
rect 38476 25096 38516 25136
rect 39340 25096 39380 25136
rect 40204 25092 40244 25132
rect 41068 25096 41108 25136
rect 42700 25096 42740 25136
rect 44044 25096 44084 25136
rect 48268 25092 48308 25132
rect 50284 25096 50324 25136
rect 50764 25096 50804 25136
rect 50956 25096 50996 25136
rect 51436 25096 51476 25136
rect 51628 25096 51668 25136
rect 53644 25092 53684 25132
rect 54124 25138 54164 25178
rect 60940 25180 60980 25220
rect 64588 25222 64628 25262
rect 64780 25264 64820 25304
rect 64876 25264 64916 25304
rect 65452 25264 65492 25304
rect 65548 25264 65588 25304
rect 65740 25264 65780 25304
rect 66124 25264 66164 25304
rect 66604 25264 66644 25304
rect 66700 25264 66740 25304
rect 67180 25264 67220 25304
rect 67372 25264 67412 25304
rect 67468 25264 67508 25304
rect 68620 25264 68660 25304
rect 69292 25264 69332 25304
rect 69388 25264 69428 25304
rect 71116 25264 71156 25304
rect 71212 25264 71252 25304
rect 71980 25264 72020 25304
rect 72076 25264 72116 25304
rect 72172 25264 72212 25304
rect 72268 25264 72308 25304
rect 73612 25264 73652 25304
rect 74476 25264 74516 25304
rect 75820 25264 75860 25304
rect 75916 25264 75956 25304
rect 76108 25264 76148 25304
rect 76780 25264 76820 25304
rect 76876 25264 76916 25304
rect 76972 25264 77012 25304
rect 77068 25264 77108 25304
rect 77356 25264 77396 25304
rect 77452 25264 77492 25304
rect 77548 25264 77588 25304
rect 77644 25264 77684 25304
rect 78220 25264 78260 25304
rect 73228 25180 73268 25220
rect 56524 25092 56564 25132
rect 58540 25096 58580 25136
rect 59596 25092 59636 25132
rect 59788 25096 59828 25136
rect 63340 25096 63380 25136
rect 64204 25092 64244 25132
rect 66796 25092 66836 25132
rect 69484 25092 69524 25132
rect 69676 25096 69716 25136
rect 71020 25092 71060 25132
rect 75628 25096 75668 25136
rect 78124 25096 78164 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 37804 24818 37844 24858
rect 844 24760 884 24800
rect 2380 24760 2420 24800
rect 40876 24760 40916 24800
rect 43468 24760 43508 24800
rect 75436 24764 75476 24804
rect 38476 24676 38516 24716
rect 41068 24676 41108 24716
rect 36364 24592 36404 24632
rect 37228 24592 37268 24632
rect 37612 24592 37652 24632
rect 37900 24592 37940 24632
rect 37996 24592 38036 24632
rect 38860 24592 38900 24632
rect 39724 24592 39764 24632
rect 41452 24592 41492 24632
rect 42316 24592 42356 24632
rect 43660 24592 43700 24632
rect 44044 24592 44084 24632
rect 44908 24592 44948 24632
rect 46252 24592 46292 24632
rect 46636 24592 46676 24632
rect 47500 24592 47540 24632
rect 48844 24592 48884 24632
rect 49228 24592 49268 24632
rect 50092 24592 50132 24632
rect 51436 24592 51476 24632
rect 51820 24592 51860 24632
rect 52684 24592 52724 24632
rect 54028 24592 54068 24632
rect 54412 24592 54452 24632
rect 55276 24592 55316 24632
rect 56620 24592 56660 24632
rect 57004 24592 57044 24632
rect 57868 24592 57908 24632
rect 59500 24592 59540 24632
rect 59884 24592 59924 24632
rect 60748 24592 60788 24632
rect 62860 24592 62900 24632
rect 62956 24592 62996 24632
rect 63052 24592 63092 24632
rect 63148 24592 63188 24632
rect 63340 24592 63380 24632
rect 63724 24592 63764 24632
rect 64588 24592 64628 24632
rect 66988 24592 67028 24632
rect 67084 24592 67124 24632
rect 67180 24592 67220 24632
rect 67276 24592 67316 24632
rect 69100 24592 69140 24632
rect 69484 24592 69524 24632
rect 70348 24592 70388 24632
rect 71692 24592 71732 24632
rect 72076 24592 72116 24632
rect 72940 24592 72980 24632
rect 74860 24592 74900 24632
rect 75244 24592 75284 24632
rect 75532 24592 75572 24632
rect 75628 24592 75668 24632
rect 76588 24592 76628 24632
rect 76972 24592 77012 24632
rect 77836 24592 77876 24632
rect 652 24508 692 24548
rect 1804 24508 1844 24548
rect 2188 24508 2228 24548
rect 35212 24508 35252 24548
rect 51244 24508 51284 24548
rect 53836 24508 53876 24548
rect 56428 24508 56468 24548
rect 61900 24508 61940 24548
rect 65740 24508 65780 24548
rect 68716 24508 68756 24548
rect 74092 24508 74132 24548
rect 74956 24508 74996 24548
rect 75148 24508 75188 24548
rect 76204 24508 76244 24548
rect 78988 24508 79028 24548
rect 75052 24424 75092 24464
rect 75916 24424 75956 24464
rect 1996 24340 2036 24380
rect 38284 24340 38324 24380
rect 40876 24340 40916 24380
rect 46060 24340 46100 24380
rect 48652 24340 48692 24380
rect 59020 24340 59060 24380
rect 68908 24340 68948 24380
rect 71500 24340 71540 24380
rect 76396 24340 76436 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 41740 24004 41780 24044
rect 37996 23920 38036 23960
rect 42796 23920 42836 23960
rect 43852 23920 43892 23960
rect 50476 23962 50516 24002
rect 51340 24004 51380 24044
rect 52204 24004 52244 24044
rect 53068 24004 53108 24044
rect 54988 24004 55028 24044
rect 55948 24004 55988 24044
rect 56428 24004 56468 24044
rect 62188 24004 62228 24044
rect 64012 24004 64052 24044
rect 65260 24004 65300 24044
rect 68812 24004 68852 24044
rect 74860 24004 74900 24044
rect 75532 24004 75572 24044
rect 57772 23920 57812 23960
rect 65452 23920 65492 23960
rect 71980 23920 72020 23960
rect 652 23836 692 23876
rect 1804 23836 1844 23876
rect 2188 23836 2228 23876
rect 37900 23836 37940 23876
rect 38092 23836 38132 23876
rect 40492 23836 40532 23876
rect 42700 23836 42740 23876
rect 42892 23836 42932 23876
rect 50380 23836 50420 23876
rect 36172 23710 36212 23750
rect 36364 23752 36404 23792
rect 36460 23752 36500 23792
rect 36748 23752 36788 23792
rect 36844 23752 36884 23792
rect 36940 23752 36980 23792
rect 37804 23752 37844 23792
rect 38188 23752 38228 23792
rect 38668 23752 38708 23792
rect 38764 23752 38804 23792
rect 38860 23752 38900 23792
rect 38956 23752 38996 23792
rect 39148 23752 39188 23792
rect 39244 23752 39284 23792
rect 39340 23752 39380 23792
rect 39436 23752 39476 23792
rect 40876 23752 40916 23792
rect 41068 23752 41108 23792
rect 41164 23752 41204 23792
rect 41452 23752 41492 23792
rect 43468 23795 43508 23835
rect 50572 23836 50612 23876
rect 52012 23836 52052 23876
rect 63244 23836 63284 23876
rect 42604 23752 42644 23792
rect 42988 23752 43028 23792
rect 43564 23752 43604 23792
rect 44140 23752 44180 23792
rect 44236 23752 44276 23792
rect 44332 23752 44372 23792
rect 44428 23752 44468 23792
rect 47308 23752 47348 23792
rect 47404 23752 47444 23792
rect 47500 23752 47540 23792
rect 47596 23752 47636 23792
rect 48172 23752 48212 23792
rect 48268 23752 48308 23792
rect 48364 23752 48404 23792
rect 48460 23752 48500 23792
rect 48748 23752 48788 23792
rect 48844 23752 48884 23792
rect 49804 23752 49844 23792
rect 49900 23752 49940 23792
rect 50092 23752 50132 23792
rect 50284 23752 50324 23792
rect 50956 23752 50996 23792
rect 51052 23752 51092 23792
rect 50668 23710 50708 23750
rect 51628 23794 51668 23834
rect 51532 23752 51572 23792
rect 51724 23752 51764 23792
rect 51820 23760 51860 23800
rect 53164 23752 53204 23792
rect 53836 23752 53876 23792
rect 53932 23752 53972 23792
rect 54028 23752 54068 23792
rect 54124 23752 54164 23792
rect 55084 23752 55124 23792
rect 55660 23752 55700 23792
rect 56044 23752 56084 23792
rect 56332 23752 56372 23792
rect 56620 23752 56660 23792
rect 56716 23752 56756 23792
rect 56812 23752 56852 23792
rect 56908 23752 56948 23792
rect 57100 23752 57140 23792
rect 57196 23752 57236 23792
rect 57292 23752 57332 23792
rect 57388 23752 57428 23792
rect 57868 23752 57908 23792
rect 59308 23752 59348 23792
rect 59404 23752 59444 23792
rect 59500 23752 59540 23792
rect 59596 23752 59636 23792
rect 59788 23752 59828 23792
rect 59884 23752 59924 23792
rect 59980 23752 60020 23792
rect 60076 23752 60116 23792
rect 60364 23752 60404 23792
rect 60940 23752 60980 23792
rect 61036 23752 61076 23792
rect 61132 23752 61172 23792
rect 61228 23752 61268 23792
rect 62092 23752 62132 23792
rect 62572 23752 62612 23792
rect 62668 23752 62708 23792
rect 63916 23752 63956 23792
rect 64204 23752 64244 23792
rect 64300 23752 64340 23792
rect 64396 23752 64436 23792
rect 64492 23752 64532 23792
rect 64780 23752 64820 23792
rect 65164 23752 65204 23792
rect 65932 23752 65972 23792
rect 66028 23752 66068 23792
rect 66124 23752 66164 23792
rect 66796 23752 66836 23792
rect 67660 23752 67700 23792
rect 69100 23752 69140 23792
rect 69196 23752 69236 23792
rect 69292 23752 69332 23792
rect 69388 23752 69428 23792
rect 69964 23752 70004 23792
rect 70060 23752 70100 23792
rect 70156 23752 70196 23792
rect 70252 23752 70292 23792
rect 71212 23752 71252 23792
rect 71308 23752 71348 23792
rect 71404 23752 71444 23792
rect 71500 23752 71540 23792
rect 72076 23752 72116 23792
rect 72460 23752 72500 23792
rect 72748 23752 72788 23792
rect 72844 23752 72884 23792
rect 74860 23752 74900 23792
rect 75052 23752 75092 23792
rect 75148 23752 75188 23792
rect 75628 23752 75668 23792
rect 76204 23752 76244 23792
rect 76300 23752 76340 23792
rect 76396 23752 76436 23792
rect 76588 23752 76628 23792
rect 76684 23752 76724 23792
rect 76780 23752 76820 23792
rect 77260 23752 77300 23792
rect 78796 23752 78836 23792
rect 78988 23752 79028 23792
rect 40972 23668 41012 23708
rect 55564 23668 55604 23708
rect 66220 23668 66260 23708
rect 66412 23668 66452 23708
rect 844 23584 884 23624
rect 1612 23584 1652 23624
rect 1996 23584 2036 23624
rect 36268 23584 36308 23624
rect 36652 23584 36692 23624
rect 40684 23584 40724 23624
rect 49996 23584 50036 23624
rect 50860 23580 50900 23620
rect 55948 23584 55988 23624
rect 60268 23584 60308 23624
rect 64876 23584 64916 23624
rect 65260 23584 65300 23624
rect 72364 23584 72404 23624
rect 76108 23584 76148 23624
rect 76876 23584 76916 23624
rect 77164 23584 77204 23624
rect 78700 23584 78740 23624
rect 79084 23584 79124 23624
rect 43372 23526 43412 23566
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 33772 23248 33812 23288
rect 36844 23252 36884 23292
rect 39820 23248 39860 23288
rect 42412 23248 42452 23288
rect 43372 23248 43412 23288
rect 43852 23248 43892 23288
rect 45004 23248 45044 23288
rect 48844 23248 48884 23288
rect 50284 23248 50324 23288
rect 50860 23248 50900 23288
rect 52396 23164 52436 23204
rect 1516 23080 1556 23120
rect 1708 23080 1748 23120
rect 34924 23080 34964 23120
rect 35788 23080 35828 23120
rect 36172 23080 36212 23120
rect 36652 23080 36692 23120
rect 36748 23080 36788 23120
rect 37036 23080 37076 23120
rect 37420 23080 37460 23120
rect 37804 23080 37844 23120
rect 38668 23080 38708 23120
rect 40012 23080 40052 23120
rect 40396 23080 40436 23120
rect 41260 23080 41300 23120
rect 42604 23080 42644 23120
rect 42700 23080 42740 23120
rect 42796 23101 42836 23141
rect 42892 23080 42932 23120
rect 43084 23080 43124 23120
rect 43468 23080 43508 23120
rect 43948 23080 43988 23120
rect 44044 23080 44084 23120
rect 44140 23080 44180 23120
rect 44908 23080 44948 23120
rect 45964 23080 46004 23120
rect 46060 23080 46100 23120
rect 46156 23080 46196 23120
rect 46252 23080 46292 23120
rect 46444 23080 46484 23120
rect 46828 23080 46868 23120
rect 47692 23080 47732 23120
rect 49228 23080 49268 23120
rect 49708 23080 49748 23120
rect 50092 23080 50132 23120
rect 52012 23080 52052 23120
rect 52108 23080 52148 23120
rect 52300 23080 52340 23120
rect 52684 23080 52724 23120
rect 652 22996 692 23036
rect 1612 22996 1652 23036
rect 49324 22996 49364 23036
rect 49804 22996 49844 23036
rect 49996 22996 50036 23036
rect 50476 22996 50516 23036
rect 50668 22996 50708 23036
rect 51532 22996 51572 23036
rect 844 22912 884 22952
rect 49900 22912 49940 22952
rect 36364 22828 36404 22868
rect 37132 22828 37172 22868
rect 43180 22828 43220 22868
rect 48844 22828 48884 22868
rect 51340 22828 51380 22868
rect 52588 22828 52628 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 31084 22492 31124 22532
rect 32044 22492 32084 22532
rect 37804 22492 37844 22532
rect 39436 22492 39476 22532
rect 42028 22534 42068 22574
rect 43468 22492 43508 22532
rect 46444 22492 46484 22532
rect 47116 22492 47156 22532
rect 52396 22492 52436 22532
rect 52684 22492 52724 22532
rect 652 22408 692 22448
rect 36172 22408 36212 22448
rect 41644 22408 41684 22448
rect 42892 22408 42932 22448
rect 49324 22408 49364 22448
rect 31276 22324 31316 22364
rect 32236 22324 32276 22364
rect 33292 22324 33332 22364
rect 36076 22324 36116 22364
rect 36268 22324 36308 22364
rect 41548 22324 41588 22364
rect 41740 22324 41780 22364
rect 7948 22240 7988 22280
rect 31564 22240 31604 22280
rect 31660 22240 31700 22280
rect 31756 22240 31796 22280
rect 35500 22240 35540 22280
rect 35692 22240 35732 22280
rect 35788 22240 35828 22280
rect 35980 22240 36020 22280
rect 36364 22240 36404 22280
rect 36940 22240 36980 22280
rect 37036 22240 37076 22280
rect 37132 22240 37172 22280
rect 37228 22240 37268 22280
rect 37516 22240 37556 22280
rect 37708 22240 37748 22280
rect 39532 22240 39572 22280
rect 41452 22240 41492 22280
rect 41836 22240 41876 22280
rect 42316 22240 42356 22280
rect 42412 22240 42452 22280
rect 42892 22240 42932 22280
rect 43084 22240 43124 22280
rect 43198 22233 43238 22273
rect 43372 22240 43412 22280
rect 45004 22240 45044 22280
rect 45868 22240 45908 22280
rect 46732 22240 46772 22280
rect 46828 22240 46868 22280
rect 47212 22240 47252 22280
rect 47404 22240 47444 22280
rect 47596 22240 47636 22280
rect 47692 22240 47732 22280
rect 49612 22240 49652 22280
rect 49708 22240 49748 22280
rect 50380 22240 50420 22280
rect 51244 22240 51284 22280
rect 52588 22240 52628 22280
rect 46252 22156 46292 22196
rect 49996 22156 50036 22196
rect 31084 22072 31124 22112
rect 31468 22072 31508 22112
rect 32044 22072 32084 22112
rect 33484 22072 33524 22112
rect 35596 22072 35636 22112
rect 37420 22072 37460 22112
rect 37804 22072 37844 22112
rect 39436 22072 39476 22112
rect 42508 22068 42548 22108
rect 43852 22072 43892 22112
rect 47500 22072 47540 22112
rect 52396 22072 52436 22112
rect 46924 22014 46964 22054
rect 49804 22014 49844 22054
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 36076 21740 36116 21780
rect 42124 21736 42164 21776
rect 45004 21736 45044 21776
rect 46732 21736 46772 21776
rect 49996 21736 50036 21776
rect 30892 21652 30932 21692
rect 37228 21652 37268 21692
rect 37420 21652 37460 21692
rect 3724 21568 3764 21608
rect 3820 21568 3860 21608
rect 3916 21568 3956 21608
rect 4012 21568 4052 21608
rect 4492 21568 4532 21608
rect 4588 21568 4628 21608
rect 4684 21568 4724 21608
rect 4780 21568 4820 21608
rect 4972 21568 5012 21608
rect 5356 21568 5396 21608
rect 6220 21568 6260 21608
rect 7756 21568 7796 21608
rect 8140 21568 8180 21608
rect 9004 21568 9044 21608
rect 11212 21568 11252 21608
rect 11596 21568 11636 21608
rect 12460 21568 12500 21608
rect 31276 21568 31316 21608
rect 32140 21568 32180 21608
rect 34636 21568 34676 21608
rect 35500 21568 35540 21608
rect 35884 21568 35924 21608
rect 36172 21568 36212 21608
rect 36268 21568 36308 21608
rect 36940 21568 36980 21608
rect 37036 21568 37076 21608
rect 37132 21568 37172 21608
rect 37804 21568 37844 21608
rect 38668 21568 38708 21608
rect 40012 21568 40052 21608
rect 40108 21568 40148 21608
rect 40300 21610 40340 21650
rect 42604 21652 42644 21692
rect 49804 21652 49844 21692
rect 42220 21568 42260 21608
rect 42316 21568 42356 21608
rect 42412 21568 42452 21608
rect 42988 21568 43028 21608
rect 43852 21568 43892 21608
rect 45868 21568 45908 21608
rect 45964 21568 46004 21608
rect 46156 21568 46196 21608
rect 46540 21568 46580 21608
rect 46828 21568 46868 21608
rect 46924 21568 46964 21608
rect 47020 21568 47060 21608
rect 48556 21568 48596 21608
rect 49420 21568 49460 21608
rect 50092 21568 50132 21608
rect 50188 21568 50228 21608
rect 50284 21568 50324 21608
rect 50476 21568 50516 21608
rect 50572 21568 50612 21608
rect 50668 21568 50708 21608
rect 50764 21568 50804 21608
rect 51244 21568 51284 21608
rect 51532 21568 51572 21608
rect 51820 21568 51860 21608
rect 52204 21568 52244 21608
rect 52492 21568 52532 21608
rect 3340 21484 3380 21524
rect 7372 21484 7412 21524
rect 29740 21484 29780 21524
rect 30124 21484 30164 21524
rect 30508 21484 30548 21524
rect 39820 21484 39860 21524
rect 46252 21484 46292 21524
rect 46444 21484 46484 21524
rect 51148 21484 51188 21524
rect 46348 21400 46388 21440
rect 52588 21400 52628 21440
rect 3532 21316 3572 21356
rect 10156 21316 10196 21356
rect 13612 21316 13652 21356
rect 29932 21316 29972 21356
rect 30316 21316 30356 21356
rect 30700 21316 30740 21356
rect 33292 21316 33332 21356
rect 33484 21316 33524 21356
rect 36556 21316 36596 21356
rect 40300 21316 40340 21356
rect 47404 21316 47444 21356
rect 51628 21316 51668 21356
rect 51916 21316 51956 21356
rect 52300 21316 52340 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 7948 20980 7988 21020
rect 33004 20980 33044 21020
rect 43660 20980 43700 21020
rect 49612 20980 49652 21020
rect 652 20896 692 20936
rect 3820 20896 3860 20936
rect 6796 20896 6836 20936
rect 10252 20896 10292 20936
rect 32620 20896 32660 20936
rect 1324 20812 1364 20852
rect 2764 20812 2804 20852
rect 3628 20812 3668 20852
rect 6412 20812 6452 20852
rect 6700 20812 6740 20852
rect 6892 20812 6932 20852
rect 10156 20812 10196 20852
rect 10348 20812 10388 20852
rect 16300 20812 16340 20852
rect 29644 20812 29684 20852
rect 32524 20812 32564 20852
rect 32716 20854 32756 20894
rect 35692 20896 35732 20936
rect 52492 20896 52532 20936
rect 35596 20812 35636 20852
rect 35788 20812 35828 20852
rect 37420 20812 37460 20852
rect 40012 20812 40052 20852
rect 42604 20812 42644 20852
rect 43852 20812 43892 20852
rect 46828 20812 46868 20852
rect 49996 20812 50036 20852
rect 50380 20812 50420 20852
rect 50572 20812 50612 20852
rect 3148 20728 3188 20768
rect 3244 20728 3284 20768
rect 3340 20728 3380 20768
rect 4396 20728 4436 20768
rect 5260 20728 5300 20768
rect 6604 20728 6644 20768
rect 6988 20728 7028 20768
rect 7468 20728 7508 20768
rect 8428 20728 8468 20768
rect 9772 20728 9812 20768
rect 10060 20728 10100 20768
rect 10444 20728 10484 20768
rect 10828 20728 10868 20768
rect 10924 20728 10964 20768
rect 11020 20728 11060 20768
rect 11116 20728 11156 20768
rect 13516 20728 13556 20768
rect 13612 20728 13652 20768
rect 13708 20728 13748 20768
rect 14284 20728 14324 20768
rect 15148 20728 15188 20768
rect 30988 20728 31028 20768
rect 31852 20728 31892 20768
rect 32236 20728 32276 20768
rect 32428 20728 32468 20768
rect 32812 20728 32852 20768
rect 33004 20728 33044 20768
rect 33196 20728 33236 20768
rect 33292 20728 33332 20768
rect 35212 20728 35252 20768
rect 35500 20728 35540 20768
rect 35884 20728 35924 20768
rect 36748 20728 36788 20768
rect 36844 20728 36884 20768
rect 36940 20728 36980 20768
rect 37036 20728 37076 20768
rect 40588 20728 40628 20768
rect 41452 20728 41492 20768
rect 42892 20728 42932 20768
rect 47212 20728 47252 20768
rect 48844 20728 48884 20768
rect 49132 20728 49172 20768
rect 49516 20728 49556 20768
rect 52204 20728 52244 20768
rect 52588 20728 52628 20768
rect 4012 20644 4052 20684
rect 13900 20644 13940 20684
rect 40204 20644 40244 20684
rect 1516 20560 1556 20600
rect 2956 20560 2996 20600
rect 3436 20560 3476 20600
rect 9868 20560 9908 20600
rect 13420 20560 13460 20600
rect 29452 20560 29492 20600
rect 29836 20560 29876 20600
rect 35308 20560 35348 20600
rect 37612 20560 37652 20600
rect 39820 20560 39860 20600
rect 42796 20560 42836 20600
rect 43660 20560 43700 20600
rect 46636 20560 46676 20600
rect 47116 20560 47156 20600
rect 49804 20560 49844 20600
rect 50188 20560 50228 20600
rect 50764 20560 50804 20600
rect 52300 20560 52340 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 31660 20282 31700 20322
rect 3340 20228 3380 20268
rect 9292 20224 9332 20264
rect 30508 20224 30548 20264
rect 41740 20224 41780 20264
rect 42412 20228 42452 20268
rect 7660 20140 7700 20180
rect 7852 20140 7892 20180
rect 11692 20140 11732 20180
rect 28492 20140 28532 20180
rect 42796 20140 42836 20180
rect 1900 20056 1940 20096
rect 2764 20056 2804 20096
rect 3148 20056 3188 20096
rect 3436 20056 3476 20096
rect 3532 20056 3572 20096
rect 4012 20056 4052 20096
rect 4204 20056 4244 20096
rect 4300 20056 4340 20096
rect 6412 20056 6452 20096
rect 7276 20056 7316 20096
rect 7948 20056 7988 20096
rect 8044 20056 8084 20096
rect 8140 20056 8180 20096
rect 8332 20056 8372 20096
rect 8428 20056 8468 20096
rect 8524 20056 8564 20096
rect 8620 20056 8660 20096
rect 10444 20056 10484 20096
rect 11308 20056 11348 20096
rect 26956 20056 26996 20096
rect 27628 20056 27668 20096
rect 30700 20056 30740 20096
rect 30796 20056 30836 20096
rect 30892 20056 30932 20096
rect 30988 20056 31028 20096
rect 31468 20056 31508 20096
rect 31564 20056 31604 20096
rect 35692 20056 35732 20096
rect 36556 20056 36596 20096
rect 36940 20056 36980 20096
rect 38572 20056 38612 20096
rect 39436 20056 39476 20096
rect 39820 20056 39860 20096
rect 40492 20056 40532 20096
rect 40876 20056 40916 20096
rect 41644 20077 41684 20117
rect 42220 20056 42260 20096
rect 43180 20069 43220 20109
rect 4684 19972 4724 20012
rect 5260 19972 5300 20012
rect 30316 19972 30356 20012
rect 31948 19972 31988 20012
rect 33196 19972 33236 20012
rect 33580 19972 33620 20012
rect 33964 19972 34004 20012
rect 40108 19972 40148 20012
rect 40588 19972 40628 20012
rect 40780 19972 40820 20012
rect 41068 19972 41108 20012
rect 41452 20011 41492 20051
rect 41548 20014 41588 20054
rect 44044 20056 44084 20096
rect 45388 20056 45428 20096
rect 42316 20014 42356 20054
rect 45772 20056 45812 20096
rect 46636 20056 46676 20096
rect 48364 20056 48404 20096
rect 48748 20056 48788 20096
rect 49612 20056 49652 20096
rect 47788 19972 47828 20012
rect 50956 19972 50996 20012
rect 51340 19972 51380 20012
rect 51916 19972 51956 20012
rect 3820 19888 3860 19928
rect 27916 19888 27956 19928
rect 31180 19888 31220 19928
rect 32140 19888 32180 19928
rect 40684 19888 40724 19928
rect 41932 19888 41972 19928
rect 51148 19888 51188 19928
rect 748 19804 788 19844
rect 4012 19804 4052 19844
rect 4492 19804 4532 19844
rect 33004 19804 33044 19844
rect 33388 19804 33428 19844
rect 33772 19804 33812 19844
rect 34540 19804 34580 19844
rect 37420 19804 37460 19844
rect 40300 19804 40340 19844
rect 41260 19804 41300 19844
rect 45196 19804 45236 19844
rect 50764 19804 50804 19844
rect 51532 19804 51572 19844
rect 51724 19804 51764 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 1228 19468 1268 19508
rect 3052 19468 3092 19508
rect 6412 19468 6452 19508
rect 7084 19468 7124 19508
rect 7276 19468 7316 19508
rect 10732 19468 10772 19508
rect 31660 19468 31700 19508
rect 38860 19468 38900 19508
rect 48076 19468 48116 19508
rect 652 19384 692 19424
rect 3436 19384 3476 19424
rect 4588 19384 4628 19424
rect 13420 19384 13460 19424
rect 32812 19384 32852 19424
rect 36460 19384 36500 19424
rect 36844 19384 36884 19424
rect 38092 19384 38132 19424
rect 39244 19384 39284 19424
rect 39628 19384 39668 19424
rect 40012 19384 40052 19424
rect 41164 19384 41204 19424
rect 44332 19384 44372 19424
rect 45676 19384 45716 19424
rect 46156 19384 46196 19424
rect 48460 19384 48500 19424
rect 1420 19300 1460 19340
rect 1804 19300 1844 19340
rect 2188 19300 2228 19340
rect 3340 19300 3380 19340
rect 3532 19300 3572 19340
rect 4108 19300 4148 19340
rect 5932 19300 5972 19340
rect 30700 19300 30740 19340
rect 32428 19300 32468 19340
rect 36364 19300 36404 19340
rect 36556 19300 36596 19340
rect 38668 19300 38708 19340
rect 39052 19300 39092 19340
rect 39532 19300 39572 19340
rect 39724 19300 39764 19340
rect 2956 19216 2996 19256
rect 3244 19216 3284 19256
rect 3628 19216 3668 19256
rect 4290 19201 4330 19241
rect 4396 19216 4436 19256
rect 4588 19216 4628 19256
rect 6316 19216 6356 19256
rect 6700 19216 6740 19256
rect 6796 19216 6836 19256
rect 7276 19216 7316 19256
rect 7468 19216 7508 19256
rect 7564 19216 7604 19256
rect 9772 19216 9812 19256
rect 9868 19216 9908 19256
rect 9964 19216 10004 19256
rect 10060 19216 10100 19256
rect 10348 19216 10388 19256
rect 10444 19216 10484 19256
rect 10924 19216 10964 19256
rect 11116 19216 11156 19256
rect 11212 19216 11252 19256
rect 12460 19216 12500 19256
rect 12556 19216 12596 19256
rect 12652 19216 12692 19256
rect 12748 19216 12788 19256
rect 13036 19216 13076 19256
rect 13132 19216 13172 19256
rect 31564 19216 31604 19256
rect 33100 19214 33140 19254
rect 33196 19216 33236 19256
rect 33580 19216 33620 19256
rect 33964 19216 34004 19256
rect 34828 19216 34868 19256
rect 36268 19216 36308 19256
rect 36652 19216 36692 19256
rect 37132 19216 37172 19256
rect 37228 19216 37268 19256
rect 37516 19216 37556 19256
rect 37612 19216 37652 19256
rect 38092 19216 38132 19256
rect 38284 19216 38324 19256
rect 38380 19216 38420 19256
rect 39436 19216 39476 19256
rect 39820 19216 39860 19256
rect 40300 19216 40340 19256
rect 40396 19216 40436 19256
rect 40684 19216 40724 19256
rect 40780 19216 40820 19256
rect 40876 19216 40916 19256
rect 40972 19261 41012 19301
rect 45100 19300 45140 19340
rect 45580 19300 45620 19340
rect 45772 19300 45812 19340
rect 47500 19300 47540 19340
rect 48364 19300 48404 19340
rect 48556 19300 48596 19340
rect 41164 19216 41204 19256
rect 41356 19216 41396 19256
rect 41452 19216 41492 19256
rect 41740 19216 41780 19256
rect 43180 19216 43220 19256
rect 44044 19216 44084 19256
rect 44140 19216 44180 19256
rect 44332 19216 44372 19256
rect 45484 19216 45524 19256
rect 45868 19216 45908 19256
rect 46444 19216 46484 19256
rect 46540 19216 46580 19256
rect 46924 19216 46964 19256
rect 47020 19216 47060 19256
rect 47116 19216 47156 19256
rect 47788 19216 47828 19256
rect 47884 19216 47924 19256
rect 48076 19202 48116 19242
rect 48268 19216 48308 19256
rect 48652 19216 48692 19256
rect 49036 19216 49076 19256
rect 49900 19216 49940 19256
rect 50668 19216 50708 19256
rect 51532 19216 51572 19256
rect 11020 19132 11060 19172
rect 50284 19132 50324 19172
rect 1612 19048 1652 19088
rect 1996 19048 2036 19088
rect 3916 19048 3956 19088
rect 5740 19048 5780 19088
rect 6604 19044 6644 19084
rect 10252 19044 10292 19084
rect 30892 19048 30932 19088
rect 32620 19048 32660 19088
rect 35980 19048 36020 19088
rect 37324 19044 37364 19084
rect 12940 18990 12980 19030
rect 40492 19044 40532 19084
rect 45292 19048 45332 19088
rect 46828 19048 46868 19088
rect 47308 19048 47348 19088
rect 49420 19048 49460 19088
rect 52684 19048 52724 19088
rect 33292 18990 33332 19030
rect 46636 18990 46676 19030
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 50092 18770 50132 18810
rect 3916 18716 3956 18756
rect 33484 18712 33524 18752
rect 34156 18712 34196 18752
rect 42604 18712 42644 18752
rect 43564 18712 43604 18752
rect 50284 18712 50324 18752
rect 51628 18712 51668 18752
rect 3436 18544 3476 18584
rect 3532 18544 3572 18584
rect 3628 18544 3668 18584
rect 3724 18544 3764 18584
rect 4012 18544 4052 18584
rect 4108 18544 4148 18584
rect 4588 18544 4628 18584
rect 4972 18544 5012 18584
rect 7276 18544 7316 18584
rect 7372 18544 7412 18584
rect 7468 18544 7508 18584
rect 7564 18544 7604 18584
rect 7756 18544 7796 18584
rect 8140 18544 8180 18584
rect 9004 18544 9044 18584
rect 10636 18544 10676 18584
rect 10732 18544 10772 18584
rect 10828 18544 10868 18584
rect 10924 18544 10964 18584
rect 12076 18544 12116 18584
rect 12460 18544 12500 18584
rect 12652 18544 12692 18584
rect 13036 18544 13076 18584
rect 13900 18544 13940 18584
rect 15244 18544 15284 18584
rect 15340 18544 15380 18584
rect 15436 18544 15476 18584
rect 15532 18544 15572 18584
rect 15724 18544 15764 18584
rect 16108 18544 16148 18584
rect 16972 18544 17012 18584
rect 31372 18544 31412 18584
rect 32236 18544 32276 18584
rect 32812 18586 32852 18626
rect 32620 18544 32660 18584
rect 33196 18544 33236 18584
rect 1324 18460 1364 18500
rect 1708 18460 1748 18500
rect 4684 18460 4724 18500
rect 4876 18460 4916 18500
rect 5356 18460 5396 18500
rect 6796 18460 6836 18500
rect 12172 18460 12212 18500
rect 32935 18502 32975 18542
rect 33388 18544 33428 18584
rect 33676 18544 33716 18584
rect 33868 18544 33908 18584
rect 33964 18544 34004 18584
rect 34252 18544 34292 18584
rect 34348 18544 34388 18584
rect 34444 18544 34484 18584
rect 34636 18544 34676 18584
rect 36460 18544 36500 18584
rect 36556 18544 36596 18584
rect 36652 18544 36692 18584
rect 36748 18544 36788 18584
rect 36940 18544 36980 18584
rect 37324 18544 37364 18584
rect 38188 18544 38228 18584
rect 39532 18544 39572 18584
rect 39628 18544 39668 18584
rect 39724 18544 39764 18584
rect 39820 18544 39860 18584
rect 40012 18544 40052 18584
rect 40396 18544 40436 18584
rect 41260 18544 41300 18584
rect 42700 18544 42740 18584
rect 42796 18544 42836 18584
rect 42892 18544 42932 18584
rect 43468 18544 43508 18584
rect 43756 18544 43796 18584
rect 44140 18544 44180 18584
rect 45004 18544 45044 18584
rect 46348 18544 46388 18584
rect 46732 18544 46772 18584
rect 47596 18544 47636 18584
rect 49132 18544 49172 18584
rect 49324 18544 49364 18584
rect 49420 18544 49460 18584
rect 49900 18544 49940 18584
rect 49996 18544 50036 18584
rect 50380 18544 50420 18584
rect 50476 18544 50516 18584
rect 50572 18544 50612 18584
rect 50956 18544 50996 18584
rect 51052 18544 51092 18584
rect 51148 18544 51188 18584
rect 51244 18544 51284 18584
rect 51820 18544 51860 18584
rect 12364 18460 12404 18500
rect 652 18376 692 18416
rect 4780 18376 4820 18416
rect 6604 18376 6644 18416
rect 12268 18376 12308 18416
rect 18124 18376 18164 18416
rect 33004 18376 33044 18416
rect 33100 18418 33140 18458
rect 42412 18460 42452 18500
rect 43084 18460 43124 18500
rect 51436 18460 51476 18500
rect 43276 18376 43316 18416
rect 49612 18376 49652 18416
rect 1132 18292 1172 18332
rect 1516 18292 1556 18332
rect 4396 18292 4436 18332
rect 5164 18292 5204 18332
rect 10156 18292 10196 18332
rect 15052 18292 15092 18332
rect 30220 18292 30260 18332
rect 33676 18292 33716 18332
rect 34732 18292 34772 18332
rect 39340 18292 39380 18332
rect 46156 18292 46196 18332
rect 48748 18292 48788 18332
rect 49132 18292 49172 18332
rect 51628 18292 51668 18332
rect 51916 18292 51956 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 3820 17956 3860 17996
rect 7180 17956 7220 17996
rect 10348 17956 10388 17996
rect 13132 17956 13172 17996
rect 13612 17956 13652 17996
rect 31948 17956 31988 17996
rect 39724 17956 39764 17996
rect 48748 17956 48788 17996
rect 51052 17956 51092 17996
rect 652 17872 692 17912
rect 49900 17872 49940 17912
rect 1324 17788 1364 17828
rect 1708 17788 1748 17828
rect 4012 17788 4052 17828
rect 7372 17788 7412 17828
rect 31756 17788 31796 17828
rect 39916 17788 39956 17828
rect 40300 17788 40340 17828
rect 40492 17788 40532 17828
rect 48556 17788 48596 17828
rect 49132 17788 49172 17828
rect 49324 17788 49364 17828
rect 49804 17788 49844 17828
rect 49996 17788 50036 17828
rect 3724 17704 3764 17744
rect 5164 17704 5204 17744
rect 6028 17704 6068 17744
rect 6412 17704 6452 17744
rect 6796 17704 6836 17744
rect 6892 17704 6932 17744
rect 9964 17704 10004 17744
rect 10060 17704 10100 17744
rect 10924 17704 10964 17744
rect 11788 17704 11828 17744
rect 13132 17704 13172 17744
rect 13324 17704 13364 17744
rect 13420 17704 13460 17744
rect 13708 17704 13748 17744
rect 32140 17704 32180 17744
rect 32236 17704 32276 17744
rect 32428 17704 32468 17744
rect 32716 17704 32756 17744
rect 32812 17704 32852 17744
rect 32908 17704 32948 17744
rect 33100 17704 33140 17744
rect 33196 17704 33236 17744
rect 33388 17704 33428 17744
rect 33484 17683 33524 17723
rect 33580 17704 33620 17744
rect 33676 17704 33716 17744
rect 37420 17704 37460 17744
rect 37516 17704 37556 17744
rect 37612 17704 37652 17744
rect 37708 17704 37748 17744
rect 38188 17704 38228 17744
rect 41644 17704 41684 17744
rect 42508 17704 42548 17744
rect 43084 17704 43124 17744
rect 43468 17704 43508 17744
rect 43564 17704 43604 17744
rect 44044 17704 44084 17744
rect 44140 17704 44180 17744
rect 44236 17704 44276 17744
rect 44524 17704 44564 17744
rect 44620 17704 44660 17744
rect 44716 17704 44756 17744
rect 44812 17704 44852 17744
rect 45100 17704 45140 17744
rect 46156 17704 46196 17744
rect 46252 17704 46292 17744
rect 46348 17704 46388 17744
rect 46444 17704 46484 17744
rect 47500 17704 47540 17744
rect 49708 17704 49748 17744
rect 50092 17704 50132 17744
rect 50572 17704 50612 17744
rect 50668 17704 50708 17744
rect 50764 17704 50804 17744
rect 50956 17704 50996 17744
rect 51340 17704 51380 17744
rect 52396 17704 52436 17744
rect 52684 17704 52724 17744
rect 10540 17620 10580 17660
rect 42892 17620 42932 17660
rect 1132 17536 1172 17576
rect 1516 17536 1556 17576
rect 7564 17536 7604 17576
rect 9868 17532 9908 17572
rect 12940 17536 12980 17576
rect 32332 17536 32372 17576
rect 32620 17536 32660 17576
rect 38284 17536 38324 17576
rect 40108 17536 40148 17576
rect 43180 17536 43220 17576
rect 43756 17578 43796 17618
rect 43372 17532 43412 17572
rect 44332 17536 44372 17576
rect 45004 17536 45044 17576
rect 47404 17536 47444 17576
rect 48940 17536 48980 17576
rect 49516 17536 49556 17576
rect 50476 17536 50516 17576
rect 51244 17536 51284 17576
rect 52300 17536 52340 17576
rect 52588 17536 52628 17576
rect 6700 17478 6740 17518
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 6316 17200 6356 17240
rect 29164 17200 29204 17240
rect 32716 17204 32756 17244
rect 41260 17200 41300 17240
rect 32908 17116 32948 17156
rect 50092 17116 50132 17156
rect 6028 17032 6068 17072
rect 6124 17032 6164 17072
rect 6220 17032 6260 17072
rect 6508 17032 6548 17072
rect 6892 17032 6932 17072
rect 7084 17032 7124 17072
rect 7468 17032 7508 17072
rect 8332 17032 8372 17072
rect 9772 17032 9812 17072
rect 9868 17032 9908 17072
rect 10060 17032 10100 17072
rect 10348 17032 10388 17072
rect 10732 17032 10772 17072
rect 10924 17032 10964 17072
rect 11020 17032 11060 17072
rect 31180 17032 31220 17072
rect 32524 17032 32564 17072
rect 32620 17032 32660 17072
rect 33292 17032 33332 17072
rect 34156 17032 34196 17072
rect 35596 17032 35636 17072
rect 35980 17032 36020 17072
rect 36844 17032 36884 17072
rect 39052 17032 39092 17072
rect 40972 17043 41012 17083
rect 41164 17032 41204 17072
rect 43276 17032 43316 17072
rect 43660 17032 43700 17072
rect 44140 17032 44180 17072
rect 44332 17032 44372 17072
rect 44428 17032 44468 17072
rect 45484 17032 45524 17072
rect 46156 17032 46196 17072
rect 46252 17032 46292 17072
rect 46348 17032 46388 17072
rect 46444 17032 46484 17072
rect 46636 17032 46676 17072
rect 46732 17032 46772 17072
rect 46828 17032 46868 17072
rect 46924 17032 46964 17072
rect 47404 17032 47444 17072
rect 48844 17032 48884 17072
rect 49708 17032 49748 17072
rect 50284 17032 50324 17072
rect 50668 17032 50708 17072
rect 51532 17032 51572 17072
rect 2668 16948 2708 16988
rect 6604 16948 6644 16988
rect 6796 16948 6836 16988
rect 10444 16948 10484 16988
rect 10636 16948 10676 16988
rect 29740 16948 29780 16988
rect 35308 16948 35348 16988
rect 37996 16948 38036 16988
rect 39148 16948 39188 16988
rect 40492 16948 40532 16988
rect 43372 16948 43412 16988
rect 45772 16948 45812 16988
rect 652 16864 692 16904
rect 1036 16864 1076 16904
rect 6700 16864 6740 16904
rect 10060 16864 10100 16904
rect 10540 16864 10580 16904
rect 32236 16864 32276 16904
rect 43564 16906 43604 16946
rect 2476 16780 2516 16820
rect 9484 16780 9524 16820
rect 40684 16780 40724 16820
rect 40876 16780 40916 16820
rect 43468 16822 43508 16862
rect 44140 16864 44180 16904
rect 45580 16780 45620 16820
rect 45964 16780 46004 16820
rect 47308 16780 47348 16820
rect 47692 16780 47732 16820
rect 52684 16780 52724 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 6604 16444 6644 16484
rect 6892 16444 6932 16484
rect 27628 16444 27668 16484
rect 40492 16444 40532 16484
rect 45484 16444 45524 16484
rect 50380 16444 50420 16484
rect 54892 16444 54932 16484
rect 56332 16444 56372 16484
rect 57004 16444 57044 16484
rect 57292 16444 57332 16484
rect 59596 16444 59636 16484
rect 63916 16444 63956 16484
rect 65740 16444 65780 16484
rect 66124 16444 66164 16484
rect 66700 16444 66740 16484
rect 69292 16444 69332 16484
rect 69964 16444 70004 16484
rect 73420 16444 73460 16484
rect 74188 16444 74228 16484
rect 77836 16444 77876 16484
rect 79468 16444 79508 16484
rect 652 16360 692 16400
rect 32236 16360 32276 16400
rect 46348 16360 46388 16400
rect 71788 16360 71828 16400
rect 1708 16276 1748 16316
rect 10540 16276 10580 16316
rect 32140 16276 32180 16316
rect 32332 16276 32372 16316
rect 49708 16276 49748 16316
rect 56044 16276 56084 16316
rect 59116 16276 59156 16316
rect 60748 16287 60788 16327
rect 70348 16276 70388 16316
rect 70732 16276 70772 16316
rect 70924 16276 70964 16316
rect 75628 16276 75668 16316
rect 76012 16276 76052 16316
rect 78604 16276 78644 16316
rect 6316 16192 6356 16232
rect 6412 16192 6452 16232
rect 6604 16192 6644 16232
rect 6988 16192 7028 16232
rect 28300 16192 28340 16232
rect 29932 16192 29972 16232
rect 32044 16192 32084 16232
rect 32428 16192 32468 16232
rect 32812 16192 32852 16232
rect 32908 16192 32948 16232
rect 33004 16192 33044 16232
rect 33100 16192 33140 16232
rect 33388 16192 33428 16232
rect 33484 16192 33524 16232
rect 35500 16192 35540 16232
rect 35596 16192 35636 16232
rect 35692 16192 35732 16232
rect 35788 16192 35828 16232
rect 36172 16192 36212 16232
rect 36268 16192 36308 16232
rect 36364 16192 36404 16232
rect 36844 16192 36884 16232
rect 37708 16192 37748 16232
rect 37804 16192 37844 16232
rect 37900 16192 37940 16232
rect 38476 16192 38516 16232
rect 39340 16192 39380 16232
rect 41068 16192 41108 16232
rect 42892 16192 42932 16232
rect 43468 16192 43508 16232
rect 44332 16192 44372 16232
rect 45964 16192 46004 16232
rect 46060 16192 46100 16232
rect 46540 16192 46580 16232
rect 46924 16192 46964 16232
rect 47788 16192 47828 16232
rect 49612 16192 49652 16232
rect 49996 16192 50036 16232
rect 50092 16192 50132 16232
rect 50572 16192 50612 16232
rect 50668 16192 50708 16232
rect 50764 16192 50804 16232
rect 50860 16192 50900 16232
rect 51052 16192 51092 16232
rect 52204 16192 52244 16232
rect 52876 16192 52916 16232
rect 53740 16192 53780 16232
rect 55180 16192 55220 16232
rect 55276 16192 55316 16232
rect 55372 16192 55412 16232
rect 56236 16192 56276 16232
rect 56620 16192 56660 16232
rect 56908 16192 56948 16232
rect 57196 16192 57236 16232
rect 58060 16192 58100 16232
rect 58156 16192 58196 16232
rect 58252 16192 58292 16232
rect 58636 16192 58676 16232
rect 58732 16192 58772 16232
rect 58828 16192 58868 16232
rect 59500 16192 59540 16232
rect 60076 16192 60116 16232
rect 60460 16192 60500 16232
rect 60556 16192 60596 16232
rect 61516 16192 61556 16232
rect 62380 16192 62420 16232
rect 63820 16192 63860 16232
rect 65644 16192 65684 16232
rect 66028 16192 66068 16232
rect 66316 16192 66356 16232
rect 66604 16192 66644 16232
rect 67276 16192 67316 16232
rect 68140 16192 68180 16232
rect 69580 16192 69620 16232
rect 69676 16192 69716 16232
rect 69868 16192 69908 16232
rect 72172 16192 72212 16232
rect 72460 16192 72500 16232
rect 73324 16192 73364 16232
rect 74092 16192 74132 16232
rect 75340 16192 75380 16232
rect 77740 16192 77780 16232
rect 78508 16192 78548 16232
rect 79372 16192 79412 16232
rect 37612 16108 37652 16148
rect 38092 16108 38132 16148
rect 42796 16108 42836 16148
rect 43084 16108 43124 16148
rect 52492 16108 52532 16148
rect 61132 16108 61172 16148
rect 66892 16108 66932 16148
rect 1516 16024 1556 16064
rect 10348 16024 10388 16064
rect 36076 16024 36116 16064
rect 36748 16024 36788 16064
rect 41164 16024 41204 16064
rect 45868 16020 45908 16060
rect 48940 16024 48980 16064
rect 49900 16020 49940 16060
rect 51148 16024 51188 16064
rect 52300 16024 52340 16064
rect 55084 16024 55124 16064
rect 55852 16024 55892 16064
rect 56716 16024 56756 16064
rect 57292 16024 57332 16064
rect 58348 16024 58388 16064
rect 58924 16024 58964 16064
rect 59308 16024 59348 16064
rect 60172 16024 60212 16064
rect 60940 16024 60980 16064
rect 63532 16024 63572 16064
rect 66124 16024 66164 16064
rect 66700 16024 66740 16064
rect 69292 16024 69332 16064
rect 69964 16024 70004 16064
rect 70156 16024 70196 16064
rect 70540 16024 70580 16064
rect 71116 16024 71156 16064
rect 72268 16024 72308 16064
rect 72556 16024 72596 16064
rect 73420 16024 73460 16064
rect 74188 16024 74228 16064
rect 75436 16024 75476 16064
rect 75820 16024 75860 16064
rect 76204 16024 76244 16064
rect 76396 16024 76436 16064
rect 77836 16024 77876 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 75532 15746 75572 15786
rect 34060 15688 34100 15728
rect 35980 15692 36020 15732
rect 36172 15688 36212 15728
rect 38188 15692 38228 15732
rect 39820 15688 39860 15728
rect 42412 15688 42452 15728
rect 52300 15688 52340 15728
rect 57772 15688 57812 15728
rect 60364 15688 60404 15728
rect 60940 15688 60980 15728
rect 61612 15688 61652 15728
rect 66892 15688 66932 15728
rect 69868 15688 69908 15728
rect 72748 15688 72788 15728
rect 72940 15688 72980 15728
rect 78796 15688 78836 15728
rect 31660 15604 31700 15644
rect 38380 15604 38420 15644
rect 40012 15604 40052 15644
rect 55372 15604 55412 15644
rect 57964 15604 58004 15644
rect 67468 15604 67508 15644
rect 70348 15604 70388 15644
rect 27628 15520 27668 15560
rect 32044 15520 32084 15560
rect 32908 15520 32948 15560
rect 34252 15520 34292 15560
rect 34348 15520 34388 15560
rect 34540 15520 34580 15560
rect 34732 15520 34772 15560
rect 35116 15520 35156 15560
rect 35788 15520 35828 15560
rect 35884 15520 35924 15560
rect 36268 15520 36308 15560
rect 36652 15520 36692 15560
rect 36748 15520 36788 15560
rect 36940 15509 36980 15549
rect 37996 15520 38036 15560
rect 38092 15520 38132 15560
rect 38476 15520 38516 15560
rect 38572 15520 38612 15560
rect 38668 15520 38708 15560
rect 39532 15520 39572 15560
rect 39628 15520 39668 15560
rect 39724 15520 39764 15560
rect 40396 15520 40436 15560
rect 41260 15520 41300 15560
rect 42604 15520 42644 15560
rect 42988 15520 43028 15560
rect 43852 15520 43892 15560
rect 45676 15520 45716 15560
rect 46732 15520 46772 15560
rect 47116 15520 47156 15560
rect 47308 15520 47348 15560
rect 47500 15520 47540 15560
rect 47596 15520 47636 15560
rect 47788 15520 47828 15560
rect 49036 15520 49076 15560
rect 49132 15520 49172 15560
rect 49228 15520 49268 15560
rect 49324 15520 49364 15560
rect 49708 15520 49748 15560
rect 49804 15520 49844 15560
rect 49900 15520 49940 15560
rect 49996 15520 50036 15560
rect 52396 15520 52436 15560
rect 52492 15520 52532 15560
rect 52588 15520 52628 15560
rect 53068 15520 53108 15560
rect 55756 15520 55796 15560
rect 56620 15520 56660 15560
rect 58348 15520 58388 15560
rect 59212 15520 59252 15560
rect 61036 15520 61076 15560
rect 61132 15520 61172 15560
rect 61228 15520 61268 15560
rect 61804 15520 61844 15560
rect 61900 15520 61940 15560
rect 61996 15541 62036 15581
rect 62092 15520 62132 15560
rect 66988 15520 67028 15560
rect 67084 15520 67124 15560
rect 67180 15520 67220 15560
rect 67564 15520 67604 15560
rect 67948 15520 67988 15560
rect 68044 15520 68084 15560
rect 68140 15520 68180 15560
rect 68236 15520 68276 15560
rect 68428 15520 68468 15560
rect 69964 15520 70004 15560
rect 70060 15520 70100 15560
rect 70156 15520 70196 15560
rect 70732 15520 70772 15560
rect 71596 15520 71636 15560
rect 74092 15520 74132 15560
rect 74956 15520 74996 15560
rect 75340 15520 75380 15560
rect 75628 15520 75668 15560
rect 75724 15520 75764 15560
rect 76396 15520 76436 15560
rect 76780 15520 76820 15560
rect 77644 15520 77684 15560
rect 844 15436 884 15476
rect 1708 15436 1748 15476
rect 34828 15436 34868 15476
rect 35020 15436 35060 15476
rect 46828 15436 46868 15476
rect 47020 15436 47060 15476
rect 61420 15436 61460 15476
rect 62284 15436 62324 15476
rect 65068 15436 65108 15476
rect 68524 15436 68564 15476
rect 69484 15436 69524 15476
rect 1516 15352 1556 15392
rect 34540 15352 34580 15392
rect 34924 15352 34964 15392
rect 35500 15352 35540 15392
rect 46924 15352 46964 15392
rect 47884 15352 47924 15392
rect 652 15268 692 15308
rect 36940 15268 36980 15308
rect 37708 15268 37748 15308
rect 42412 15268 42452 15308
rect 45004 15268 45044 15308
rect 47308 15268 47348 15308
rect 54604 15268 54644 15308
rect 61612 15268 61652 15308
rect 62476 15268 62516 15308
rect 65260 15268 65300 15308
rect 69676 15268 69716 15308
rect 76012 15268 76052 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 36844 14932 36884 14972
rect 38380 14932 38420 14972
rect 48268 14932 48308 14972
rect 51148 14932 51188 14972
rect 52300 14932 52340 14972
rect 53452 14932 53492 14972
rect 58252 14932 58292 14972
rect 58924 14932 58964 14972
rect 65260 14932 65300 14972
rect 70924 14932 70964 14972
rect 37228 14848 37268 14888
rect 51916 14848 51956 14888
rect 55084 14848 55124 14888
rect 61036 14848 61076 14888
rect 67180 14848 67220 14888
rect 70060 14848 70100 14888
rect 75436 14848 75476 14888
rect 844 14764 884 14804
rect 37132 14764 37172 14804
rect 37324 14764 37364 14804
rect 51820 14764 51860 14804
rect 52012 14764 52052 14804
rect 59116 14764 59156 14804
rect 60364 14764 60404 14804
rect 61900 14764 61940 14804
rect 68428 14764 68468 14804
rect 69292 14764 69332 14804
rect 70732 14764 70772 14804
rect 73439 14759 73479 14799
rect 75340 14764 75380 14804
rect 34444 14680 34484 14720
rect 34828 14680 34868 14720
rect 35692 14680 35732 14720
rect 37036 14680 37076 14720
rect 37420 14680 37460 14720
rect 38476 14680 38516 14720
rect 38668 14680 38708 14720
rect 38764 14680 38804 14720
rect 38956 14680 38996 14720
rect 39244 14680 39284 14720
rect 42412 14680 42452 14720
rect 42508 14680 42548 14720
rect 42604 14680 42644 14720
rect 42700 14680 42740 14720
rect 43084 14680 43124 14720
rect 43180 14680 43220 14720
rect 43276 14680 43316 14720
rect 45484 14680 45524 14720
rect 45580 14680 45620 14720
rect 45676 14680 45716 14720
rect 46252 14680 46292 14720
rect 47116 14680 47156 14720
rect 48748 14680 48788 14720
rect 49132 14680 49172 14720
rect 49996 14680 50036 14720
rect 51340 14680 51380 14720
rect 51724 14680 51764 14720
rect 52108 14680 52148 14720
rect 52588 14680 52628 14720
rect 52684 14680 52724 14720
rect 52972 14680 53012 14720
rect 53068 14680 53108 14720
rect 53164 14680 53204 14720
rect 53260 14659 53300 14699
rect 53548 14680 53588 14720
rect 53932 14680 53972 14720
rect 54028 14680 54068 14720
rect 54220 14680 54260 14720
rect 54412 14680 54452 14720
rect 55372 14680 55412 14720
rect 55468 14680 55508 14720
rect 55756 14680 55796 14720
rect 55852 14680 55892 14720
rect 55948 14680 55988 14720
rect 56044 14680 56084 14720
rect 58540 14680 58580 14720
rect 58636 14680 58676 14720
rect 61324 14680 61364 14720
rect 61420 14680 61460 14720
rect 62380 14680 62420 14720
rect 62476 14680 62516 14720
rect 62572 14680 62612 14720
rect 63244 14680 63284 14720
rect 64108 14680 64148 14720
rect 65548 14680 65588 14720
rect 65644 14680 65684 14720
rect 65740 14680 65780 14720
rect 67468 14680 67508 14720
rect 67564 14680 67604 14720
rect 68812 14680 68852 14720
rect 68908 14680 68948 14720
rect 69100 14680 69140 14720
rect 70348 14680 70388 14720
rect 70444 14680 70484 14720
rect 71116 14680 71156 14720
rect 71212 14680 71252 14720
rect 71308 14680 71348 14720
rect 71404 14680 71444 14720
rect 71884 14680 71924 14720
rect 71980 14680 72020 14720
rect 72076 14680 72116 14720
rect 75244 14680 75284 14720
rect 75532 14722 75572 14762
rect 75628 14722 75668 14762
rect 75916 14680 75956 14720
rect 76012 14680 76052 14720
rect 76108 14680 76148 14720
rect 76204 14680 76244 14720
rect 76684 14680 76724 14720
rect 76780 14680 76820 14720
rect 76876 14680 76916 14720
rect 76972 14680 77012 14720
rect 45388 14596 45428 14636
rect 45868 14596 45908 14636
rect 62668 14596 62708 14636
rect 62860 14596 62900 14636
rect 652 14512 692 14552
rect 38860 14512 38900 14552
rect 41260 14512 41300 14552
rect 42988 14512 43028 14552
rect 48268 14512 48308 14552
rect 52780 14508 52820 14548
rect 54124 14512 54164 14552
rect 54508 14512 54548 14552
rect 58924 14512 58964 14552
rect 60172 14512 60212 14552
rect 62092 14512 62132 14552
rect 65452 14512 65492 14552
rect 68620 14512 68660 14552
rect 69004 14512 69044 14552
rect 69484 14512 69524 14552
rect 70924 14512 70964 14552
rect 71788 14512 71828 14552
rect 73612 14512 73652 14552
rect 55564 14454 55604 14494
rect 58732 14454 58772 14494
rect 61516 14454 61556 14494
rect 67660 14454 67700 14494
rect 70540 14454 70580 14494
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 39052 14176 39092 14216
rect 40396 14180 40436 14220
rect 41068 14176 41108 14216
rect 42892 14180 42932 14220
rect 45292 14180 45332 14220
rect 53932 14176 53972 14216
rect 66988 14176 67028 14216
rect 70540 14176 70580 14216
rect 74284 14176 74324 14216
rect 75820 14176 75860 14216
rect 79372 14176 79412 14216
rect 36652 14092 36692 14132
rect 46732 14092 46772 14132
rect 51532 14092 51572 14132
rect 64588 14092 64628 14132
rect 71884 14092 71924 14132
rect 37036 14008 37076 14048
rect 37900 14008 37940 14048
rect 39340 14008 39380 14048
rect 39724 14008 39764 14048
rect 40204 14008 40244 14048
rect 40300 14008 40340 14048
rect 40588 14008 40628 14048
rect 40684 14008 40724 14048
rect 40780 14008 40820 14048
rect 40876 14008 40916 14048
rect 41164 14008 41204 14048
rect 41644 14008 41684 14048
rect 42028 14008 42068 14048
rect 42700 13991 42740 14031
rect 42796 14008 42836 14048
rect 45100 14008 45140 14048
rect 45196 14008 45236 14048
rect 45580 14008 45620 14048
rect 46540 14008 46580 14048
rect 46828 14008 46868 14048
rect 46924 14008 46964 14048
rect 47020 14008 47060 14048
rect 48076 14008 48116 14048
rect 48460 14008 48500 14048
rect 48652 14008 48692 14048
rect 49036 14008 49076 14048
rect 49900 14008 49940 14048
rect 51916 14008 51956 14048
rect 52780 14008 52820 14048
rect 54124 14008 54164 14048
rect 54508 14008 54548 14048
rect 55372 14008 55412 14048
rect 58060 14008 58100 14048
rect 58444 14008 58484 14048
rect 59308 14008 59348 14048
rect 59500 14008 59540 14048
rect 59596 14008 59636 14048
rect 59788 14008 59828 14048
rect 59980 14008 60020 14048
rect 60364 14008 60404 14048
rect 61228 14008 61268 14048
rect 62572 14008 62612 14048
rect 63148 14008 63188 14048
rect 63244 14008 63284 14048
rect 63340 14029 63380 14069
rect 63436 14008 63476 14048
rect 64972 14008 65012 14048
rect 65836 14008 65876 14048
rect 67180 14008 67220 14048
rect 67564 14008 67604 14048
rect 68428 14008 68468 14048
rect 69772 14008 69812 14048
rect 70156 14008 70196 14048
rect 70636 14008 70676 14048
rect 70924 14008 70964 14048
rect 71308 14008 71348 14048
rect 72268 14008 72308 14048
rect 73132 14008 73172 14048
rect 75724 14008 75764 14048
rect 75916 14008 75956 14048
rect 76012 14008 76052 14048
rect 76204 14008 76244 14048
rect 76492 14008 76532 14048
rect 76588 14008 76628 14048
rect 76684 14008 76724 14048
rect 76780 14008 76820 14048
rect 76972 14008 77012 14048
rect 77356 14008 77396 14048
rect 78220 14008 78260 14048
rect 1708 13924 1748 13964
rect 39436 13924 39476 13964
rect 39628 13924 39668 13964
rect 41740 13924 41780 13964
rect 41932 13924 41972 13964
rect 48172 13924 48212 13964
rect 48364 13924 48404 13964
rect 58156 13924 58196 13964
rect 58348 13924 58388 13964
rect 69868 13924 69908 13964
rect 70060 13924 70100 13964
rect 71020 13924 71060 13964
rect 71212 13924 71252 13964
rect 39532 13840 39572 13880
rect 39916 13840 39956 13880
rect 41836 13840 41876 13880
rect 42412 13840 42452 13880
rect 44812 13840 44852 13880
rect 48268 13840 48308 13880
rect 58252 13840 58292 13880
rect 59212 13840 59252 13880
rect 62668 13840 62708 13880
rect 69964 13840 70004 13880
rect 71116 13840 71156 13880
rect 1516 13756 1556 13796
rect 45868 13756 45908 13796
rect 51052 13756 51092 13796
rect 56524 13756 56564 13796
rect 59788 13756 59828 13796
rect 62380 13756 62420 13796
rect 69580 13756 69620 13796
rect 76300 13756 76340 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 41164 13420 41204 13460
rect 49324 13420 49364 13460
rect 51436 13420 51476 13460
rect 52012 13420 52052 13460
rect 55180 13420 55220 13460
rect 59116 13420 59156 13460
rect 60172 13420 60212 13460
rect 62572 13420 62612 13460
rect 65260 13420 65300 13460
rect 71020 13420 71060 13460
rect 71500 13420 71540 13460
rect 71692 13420 71732 13460
rect 73996 13420 74036 13460
rect 76588 13420 76628 13460
rect 76780 13420 76820 13460
rect 78220 13420 78260 13460
rect 50284 13336 50324 13376
rect 54508 13336 54548 13376
rect 60556 13336 60596 13376
rect 62188 13336 62228 13376
rect 66892 13336 66932 13376
rect 67276 13336 67316 13376
rect 844 13252 884 13292
rect 1708 13252 1748 13292
rect 47788 13252 47828 13292
rect 54412 13252 54452 13292
rect 54604 13252 54644 13292
rect 59980 13252 60020 13292
rect 60460 13252 60500 13292
rect 60652 13252 60692 13292
rect 62092 13252 62132 13292
rect 62284 13252 62324 13292
rect 66796 13252 66836 13292
rect 66988 13252 67028 13292
rect 38764 13168 38804 13208
rect 39148 13168 39188 13208
rect 40012 13168 40052 13208
rect 41356 13168 41396 13208
rect 41740 13168 41780 13208
rect 42604 13168 42644 13208
rect 44428 13168 44468 13208
rect 45292 13168 45332 13208
rect 46732 13168 46772 13208
rect 46828 13168 46868 13208
rect 46924 13168 46964 13208
rect 47692 13168 47732 13208
rect 49612 13168 49652 13208
rect 49708 13168 49748 13208
rect 50380 13168 50420 13208
rect 51148 13168 51188 13208
rect 51244 13168 51284 13208
rect 51436 13168 51476 13208
rect 51724 13168 51764 13208
rect 52684 13168 52724 13208
rect 54316 13168 54356 13208
rect 54700 13168 54740 13208
rect 55276 13168 55316 13208
rect 55468 13168 55508 13208
rect 55660 13168 55700 13208
rect 55756 13168 55796 13208
rect 56236 13168 56276 13208
rect 56332 13168 56372 13208
rect 56428 13168 56468 13208
rect 56524 13168 56564 13208
rect 56716 13168 56756 13208
rect 57100 13168 57140 13208
rect 57964 13168 58004 13208
rect 60364 13168 60404 13208
rect 60748 13168 60788 13208
rect 61516 13168 61556 13208
rect 61708 13168 61748 13208
rect 61804 13168 61844 13208
rect 61996 13168 62036 13208
rect 62380 13168 62420 13208
rect 62860 13168 62900 13208
rect 62956 13168 62996 13208
rect 65548 13168 65588 13208
rect 65644 13168 65684 13208
rect 66028 13168 66068 13208
rect 66124 13168 66164 13208
rect 66220 13168 66260 13208
rect 66508 13181 66548 13221
rect 66700 13168 66740 13208
rect 67084 13168 67124 13208
rect 67276 13168 67316 13208
rect 67468 13168 67508 13208
rect 67564 13168 67604 13208
rect 68140 13168 68180 13208
rect 68236 13168 68276 13208
rect 68620 13168 68660 13208
rect 69004 13168 69044 13208
rect 69868 13168 69908 13208
rect 71212 13168 71252 13208
rect 71308 13168 71348 13208
rect 71500 13168 71540 13208
rect 71980 13168 72020 13208
rect 72076 13168 72116 13208
rect 72652 13168 72692 13208
rect 72748 13168 72788 13208
rect 72844 13168 72884 13208
rect 72940 13168 72980 13208
rect 73900 13168 73940 13208
rect 74188 13168 74228 13208
rect 74572 13168 74612 13208
rect 75436 13168 75476 13208
rect 77068 13168 77108 13208
rect 77164 13168 77204 13208
rect 77548 13168 77588 13208
rect 77644 13168 77684 13208
rect 77740 13168 77780 13208
rect 77836 13168 77876 13208
rect 78316 13168 78356 13208
rect 44044 13084 44084 13124
rect 61612 13084 61652 13124
rect 66412 13084 66452 13124
rect 652 13000 692 13040
rect 1516 13000 1556 13040
rect 41164 13000 41204 13040
rect 43756 13000 43796 13040
rect 46444 13000 46484 13040
rect 46636 13000 46676 13040
rect 49804 12996 49844 13036
rect 55564 13000 55604 13040
rect 65740 12996 65780 13036
rect 65932 13000 65972 13040
rect 72172 12996 72212 13036
rect 63052 12942 63092 12982
rect 77260 12942 77300 12982
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 43180 12664 43220 12704
rect 45580 12664 45620 12704
rect 49228 12664 49268 12704
rect 49804 12664 49844 12704
rect 50860 12664 50900 12704
rect 53740 12664 53780 12704
rect 56236 12668 56276 12708
rect 60076 12664 60116 12704
rect 62956 12664 62996 12704
rect 63724 12664 63764 12704
rect 66796 12664 66836 12704
rect 72172 12664 72212 12704
rect 75052 12664 75092 12704
rect 41260 12496 41300 12536
rect 41356 12496 41396 12536
rect 41548 12496 41588 12536
rect 43276 12496 43316 12536
rect 43564 12496 43604 12536
rect 43756 12496 43796 12536
rect 43852 12496 43892 12536
rect 44044 12538 44084 12578
rect 46828 12580 46868 12620
rect 51340 12580 51380 12620
rect 56428 12580 56468 12620
rect 57676 12580 57716 12620
rect 60268 12580 60308 12620
rect 69484 12580 69524 12620
rect 44428 12496 44468 12536
rect 44812 12496 44852 12536
rect 45676 12496 45716 12536
rect 45868 12496 45908 12536
rect 45964 12496 46004 12536
rect 46156 12496 46196 12536
rect 46348 12496 46388 12536
rect 46444 12496 46484 12536
rect 46540 12496 46580 12536
rect 46636 12496 46676 12536
rect 47212 12496 47252 12536
rect 48076 12496 48116 12536
rect 49708 12496 49748 12536
rect 49900 12496 49940 12536
rect 49996 12496 50036 12536
rect 50572 12496 50612 12536
rect 50956 12496 50996 12536
rect 51052 12496 51092 12536
rect 51148 12496 51188 12536
rect 51724 12496 51764 12536
rect 52588 12496 52628 12536
rect 55180 12496 55220 12536
rect 55564 12496 55604 12536
rect 56044 12496 56084 12536
rect 56140 12496 56180 12536
rect 56524 12496 56564 12536
rect 56620 12496 56660 12536
rect 56716 12496 56756 12536
rect 58060 12496 58100 12536
rect 58924 12496 58964 12536
rect 60652 12496 60692 12536
rect 61516 12496 61556 12536
rect 62860 12496 62900 12536
rect 63628 12496 63668 12536
rect 64396 12496 64436 12536
rect 64780 12496 64820 12536
rect 65644 12496 65684 12536
rect 67852 12496 67892 12536
rect 67948 12496 67988 12536
rect 68044 12496 68084 12536
rect 68140 12496 68180 12536
rect 69868 12496 69908 12536
rect 70732 12496 70772 12536
rect 72076 12496 72116 12536
rect 72652 12496 72692 12536
rect 73036 12496 73076 12536
rect 73900 12496 73940 12536
rect 76396 12496 76436 12536
rect 76780 12496 76820 12536
rect 77164 12496 77204 12536
rect 77260 12496 77300 12536
rect 77452 12496 77492 12536
rect 844 12412 884 12452
rect 1708 12412 1748 12452
rect 44524 12412 44564 12452
rect 44716 12412 44756 12452
rect 55276 12412 55316 12452
rect 55468 12412 55508 12452
rect 71884 12412 71924 12452
rect 76492 12412 76532 12452
rect 77356 12454 77396 12494
rect 77644 12496 77684 12536
rect 77740 12496 77780 12536
rect 77836 12496 77876 12536
rect 77932 12496 77972 12536
rect 78220 12507 78260 12547
rect 76684 12412 76724 12452
rect 652 12328 692 12368
rect 41548 12328 41588 12368
rect 44044 12328 44084 12368
rect 44620 12328 44660 12368
rect 55372 12328 55412 12368
rect 55756 12328 55796 12368
rect 76588 12328 76628 12368
rect 1516 12244 1556 12284
rect 43468 12244 43508 12284
rect 46156 12244 46196 12284
rect 50668 12244 50708 12284
rect 53740 12244 53780 12284
rect 62668 12244 62708 12284
rect 63724 12244 63764 12284
rect 78124 12244 78164 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 50668 11908 50708 11948
rect 51340 11908 51380 11948
rect 56524 11908 56564 11948
rect 65164 11908 65204 11948
rect 70060 11908 70100 11948
rect 76492 11908 76532 11948
rect 79372 11908 79412 11948
rect 46924 11824 46964 11864
rect 61228 11824 61268 11864
rect 65548 11824 65588 11864
rect 65932 11824 65972 11864
rect 72844 11824 72884 11864
rect 844 11740 884 11780
rect 1708 11740 1748 11780
rect 43660 11740 43700 11780
rect 53356 11740 53396 11780
rect 59980 11740 60020 11780
rect 61420 11740 61460 11780
rect 65452 11740 65492 11780
rect 41644 11656 41684 11696
rect 42508 11656 42548 11696
rect 45004 11656 45044 11696
rect 45868 11656 45908 11696
rect 46540 11656 46580 11696
rect 46636 11656 46676 11696
rect 48652 11656 48692 11696
rect 49516 11656 49556 11696
rect 50956 11656 50996 11696
rect 51052 11656 51092 11696
rect 51628 11656 51668 11696
rect 51724 11656 51764 11696
rect 55756 11698 55796 11738
rect 51820 11656 51860 11696
rect 54508 11656 54548 11696
rect 55372 11656 55412 11696
rect 56140 11698 56180 11738
rect 65644 11740 65684 11780
rect 56044 11656 56084 11696
rect 56236 11635 56276 11675
rect 56428 11656 56468 11696
rect 59020 11656 59060 11696
rect 59116 11656 59156 11696
rect 59212 11656 59252 11696
rect 59596 11656 59636 11696
rect 59692 11656 59732 11696
rect 59788 11656 59828 11696
rect 62188 11656 62228 11696
rect 62380 11656 62420 11696
rect 62476 11656 62516 11696
rect 63148 11656 63188 11696
rect 64012 11656 64052 11696
rect 65356 11656 65396 11696
rect 65740 11656 65780 11696
rect 65932 11656 65972 11696
rect 66124 11656 66164 11696
rect 66220 11656 66260 11696
rect 66892 11656 66932 11696
rect 67180 11656 67220 11696
rect 67276 11656 67316 11696
rect 67372 11656 67412 11696
rect 68044 11656 68084 11696
rect 68908 11656 68948 11696
rect 71596 11656 71636 11696
rect 71788 11656 71828 11696
rect 71884 11656 71924 11696
rect 72172 11656 72212 11696
rect 72460 11656 72500 11696
rect 72556 11656 72596 11696
rect 73036 11656 73076 11696
rect 73132 11656 73172 11696
rect 73228 11656 73268 11696
rect 73324 11656 73364 11696
rect 73516 11656 73556 11696
rect 73612 11656 73652 11696
rect 73708 11656 73748 11696
rect 73804 11656 73844 11696
rect 76492 11656 76532 11696
rect 76684 11656 76724 11696
rect 76780 11656 76820 11696
rect 76972 11656 77012 11696
rect 77356 11656 77396 11696
rect 78220 11656 78260 11696
rect 41260 11572 41300 11612
rect 46252 11572 46292 11612
rect 48268 11572 48308 11612
rect 51532 11572 51572 11612
rect 652 11488 692 11528
rect 1516 11488 1556 11528
rect 43852 11488 43892 11528
rect 51244 11530 51284 11570
rect 62284 11572 62324 11612
rect 62764 11572 62804 11612
rect 67468 11572 67508 11612
rect 67660 11572 67700 11612
rect 50860 11484 50900 11524
rect 55948 11488 55988 11528
rect 58924 11488 58964 11528
rect 59500 11488 59540 11528
rect 60172 11488 60212 11528
rect 66988 11488 67028 11528
rect 71692 11488 71732 11528
rect 72076 11488 72116 11528
rect 72364 11484 72404 11524
rect 46444 11430 46484 11470
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 67852 11210 67892 11250
rect 42508 11152 42548 11192
rect 43468 11156 43508 11196
rect 46348 11152 46388 11192
rect 49420 11152 49460 11192
rect 52780 11152 52820 11192
rect 58636 11152 58676 11192
rect 61324 11152 61364 11192
rect 62764 11156 62804 11196
rect 62956 11152 62996 11192
rect 64780 11152 64820 11192
rect 72364 11152 72404 11192
rect 74092 11152 74132 11192
rect 77068 11152 77108 11192
rect 77740 11156 77780 11196
rect 43660 11068 43700 11108
rect 58924 11068 58964 11108
rect 42604 10984 42644 11024
rect 42700 10984 42740 11024
rect 42796 10984 42836 11024
rect 43276 10984 43316 11024
rect 43372 10984 43412 11024
rect 43756 10984 43796 11024
rect 43852 10984 43892 11024
rect 43948 10984 43988 11024
rect 44140 10984 44180 11024
rect 44332 10984 44372 11024
rect 44428 10984 44468 11024
rect 45676 10984 45716 11024
rect 46060 10984 46100 11024
rect 46252 10984 46292 11024
rect 49324 10984 49364 11024
rect 50668 10984 50708 11024
rect 51052 10984 51092 11024
rect 51436 10984 51476 11024
rect 51532 10984 51572 11024
rect 51628 10984 51668 11024
rect 51724 10984 51764 11024
rect 51916 10984 51956 11024
rect 52012 10984 52052 11024
rect 52108 10984 52148 11024
rect 52204 10984 52244 11024
rect 52876 10984 52916 11024
rect 55180 10984 55220 11024
rect 55372 10984 55412 11024
rect 55468 10984 55508 11024
rect 55756 10984 55796 11024
rect 55852 10984 55892 11024
rect 55948 10984 55988 11024
rect 56044 10984 56084 11024
rect 56236 10984 56276 11024
rect 56620 10984 56660 11024
rect 57484 10984 57524 11024
rect 59308 10984 59348 11024
rect 60172 10984 60212 11024
rect 61708 10984 61748 11024
rect 62092 10984 62132 11024
rect 62572 10984 62612 11024
rect 844 10900 884 10940
rect 45772 10900 45812 10940
rect 45964 10900 46004 10940
rect 50284 10900 50324 10940
rect 50764 10900 50804 10940
rect 61804 10942 61844 10982
rect 62668 10984 62708 11024
rect 63052 10984 63092 11024
rect 63148 10984 63188 11024
rect 63244 10984 63284 11024
rect 63436 10984 63476 11024
rect 63532 10984 63572 11024
rect 63628 10984 63668 11024
rect 63724 10984 63764 11024
rect 65932 10984 65972 11024
rect 66796 10984 66836 11024
rect 67180 10984 67220 11024
rect 67660 10984 67700 11024
rect 67756 10984 67796 11024
rect 69964 10984 70004 11024
rect 70348 10984 70388 11024
rect 71212 10984 71252 11024
rect 72748 10984 72788 11024
rect 72844 10984 72884 11024
rect 72940 10984 72980 11024
rect 73036 10984 73076 11024
rect 74668 10984 74708 11024
rect 75052 10984 75092 11024
rect 75916 10984 75956 11024
rect 77548 10984 77588 11024
rect 77644 10984 77684 11024
rect 77932 10984 77972 11024
rect 50956 10900 50996 10940
rect 52396 10900 52436 10940
rect 61996 10900 62036 10940
rect 68908 10900 68948 10940
rect 73516 10900 73556 10940
rect 73900 10900 73940 10940
rect 45868 10816 45908 10856
rect 50860 10816 50900 10856
rect 61900 10816 61940 10856
rect 67372 10816 67412 10856
rect 77260 10816 77300 10856
rect 652 10732 692 10772
rect 42988 10732 43028 10772
rect 44140 10732 44180 10772
rect 49420 10732 49460 10772
rect 50476 10732 50516 10772
rect 52588 10732 52628 10772
rect 55180 10732 55220 10772
rect 62284 10732 62324 10772
rect 68716 10732 68756 10772
rect 72364 10732 72404 10772
rect 73324 10732 73364 10772
rect 78028 10732 78068 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 44716 10396 44756 10436
rect 47788 10396 47828 10436
rect 50380 10396 50420 10436
rect 51148 10396 51188 10436
rect 54124 10396 54164 10436
rect 58444 10396 58484 10436
rect 59596 10396 59636 10436
rect 59980 10396 60020 10436
rect 63340 10396 63380 10436
rect 70060 10396 70100 10436
rect 70348 10396 70388 10436
rect 75244 10396 75284 10436
rect 1516 10312 1556 10352
rect 43276 10312 43316 10352
rect 54988 10312 55028 10352
rect 55852 10312 55892 10352
rect 58924 10312 58964 10352
rect 67180 10312 67220 10352
rect 71884 10312 71924 10352
rect 77164 10312 77204 10352
rect 78124 10312 78164 10352
rect 844 10228 884 10268
rect 1708 10228 1748 10268
rect 43181 10238 43221 10278
rect 43372 10228 43412 10268
rect 44524 10228 44564 10268
rect 50764 10228 50804 10268
rect 54892 10228 54932 10268
rect 55084 10228 55124 10268
rect 56236 10228 56276 10268
rect 59788 10228 59828 10268
rect 60172 10228 60212 10268
rect 63052 10228 63092 10268
rect 64684 10228 64724 10268
rect 64972 10228 65012 10268
rect 67084 10228 67124 10268
rect 67276 10228 67316 10268
rect 69484 10228 69524 10268
rect 69868 10228 69908 10268
rect 71788 10228 71828 10268
rect 43084 10144 43124 10184
rect 43468 10144 43508 10184
rect 44140 10144 44180 10184
rect 44236 10144 44276 10184
rect 44908 10144 44948 10184
rect 45004 10144 45044 10184
rect 45100 10144 45140 10184
rect 45772 10144 45812 10184
rect 46636 10144 46676 10184
rect 48364 10144 48404 10184
rect 49228 10144 49268 10184
rect 51148 10144 51188 10184
rect 51340 10144 51380 10184
rect 51436 10144 51476 10184
rect 51724 10144 51764 10184
rect 52108 10144 52148 10184
rect 52972 10144 53012 10184
rect 54796 10144 54836 10184
rect 55180 10144 55220 10184
rect 55468 10144 55508 10184
rect 55564 10144 55604 10184
rect 58252 10144 58292 10184
rect 58444 10144 58484 10184
rect 58636 10144 58676 10184
rect 58732 10144 58772 10184
rect 59212 10144 59252 10184
rect 59308 10144 59348 10184
rect 60652 10144 60692 10184
rect 61036 10144 61076 10184
rect 61900 10144 61940 10184
rect 63244 10144 63284 10184
rect 64876 10144 64916 10184
rect 66988 10144 67028 10184
rect 67372 10144 67412 10184
rect 68236 10144 68276 10184
rect 68428 10186 68468 10226
rect 71980 10228 72020 10268
rect 77068 10228 77108 10268
rect 68332 10144 68372 10184
rect 69100 10144 69140 10184
rect 69196 10144 69236 10184
rect 69292 10144 69332 10184
rect 70252 10144 70292 10184
rect 72076 10186 72116 10226
rect 77260 10228 77300 10268
rect 71692 10144 71732 10184
rect 72268 10144 72308 10184
rect 72460 10144 72500 10184
rect 72556 10144 72596 10184
rect 72844 10144 72884 10184
rect 73228 10144 73268 10184
rect 74092 10144 74132 10184
rect 76588 10144 76628 10184
rect 76684 10144 76724 10184
rect 76780 10144 76820 10184
rect 76972 10144 77012 10184
rect 77356 10144 77396 10184
rect 77644 10144 77684 10184
rect 77740 10144 77780 10184
rect 77836 10144 77876 10184
rect 78028 10144 78068 10184
rect 45196 10060 45236 10100
rect 45388 10060 45428 10100
rect 47980 10060 48020 10100
rect 652 9976 692 10016
rect 47788 9976 47828 10016
rect 50956 9976 50996 10016
rect 56044 9976 56084 10016
rect 58156 9976 58196 10016
rect 59404 9972 59444 10012
rect 59596 9976 59636 10016
rect 64492 9976 64532 10016
rect 68524 9976 68564 10016
rect 69004 9976 69044 10016
rect 69676 9976 69716 10016
rect 72364 9976 72404 10016
rect 76492 9976 76532 10016
rect 77548 9976 77588 10016
rect 55372 9918 55412 9958
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 45004 9640 45044 9680
rect 46348 9644 46388 9684
rect 47116 9640 47156 9680
rect 48076 9640 48116 9680
rect 49708 9640 49748 9680
rect 52300 9640 52340 9680
rect 59500 9640 59540 9680
rect 63532 9640 63572 9680
rect 66412 9640 66452 9680
rect 67564 9640 67604 9680
rect 70636 9640 70676 9680
rect 73036 9644 73076 9684
rect 42604 9556 42644 9596
rect 53452 9556 53492 9596
rect 64012 9556 64052 9596
rect 72652 9598 72692 9638
rect 73420 9640 73460 9680
rect 77740 9640 77780 9680
rect 78028 9640 78068 9680
rect 68236 9556 68276 9596
rect 75340 9556 75380 9596
rect 42988 9472 43028 9512
rect 43852 9472 43892 9512
rect 46156 9472 46196 9512
rect 46252 9472 46292 9512
rect 46540 9472 46580 9512
rect 46636 9472 46676 9512
rect 46732 9472 46772 9512
rect 46828 9472 46868 9512
rect 47212 9472 47252 9512
rect 48172 9472 48212 9512
rect 48268 9472 48308 9512
rect 48364 9472 48404 9512
rect 49324 9472 49364 9512
rect 49900 9472 49940 9512
rect 50284 9472 50324 9512
rect 51148 9472 51188 9512
rect 52492 9472 52532 9512
rect 53836 9472 53876 9512
rect 54700 9472 54740 9512
rect 57100 9472 57140 9512
rect 57484 9472 57524 9512
rect 58348 9472 58388 9512
rect 62668 9472 62708 9512
rect 62860 9472 62900 9512
rect 62956 9472 62996 9512
rect 63628 9472 63668 9512
rect 63724 9472 63764 9512
rect 63820 9472 63860 9512
rect 64396 9472 64436 9512
rect 65260 9472 65300 9512
rect 67468 9472 67508 9512
rect 67660 9472 67700 9512
rect 67756 9472 67796 9512
rect 67935 9483 67975 9523
rect 68620 9472 68660 9512
rect 69484 9472 69524 9512
rect 71980 9472 72020 9512
rect 72364 9472 72404 9512
rect 72844 9472 72884 9512
rect 72940 9472 72980 9512
rect 73612 9472 73652 9512
rect 73708 9472 73748 9512
rect 73804 9472 73844 9512
rect 73900 9472 73940 9512
rect 75724 9472 75764 9512
rect 76588 9472 76628 9512
rect 77932 9472 77972 9512
rect 78124 9472 78164 9512
rect 78220 9472 78260 9512
rect 844 9388 884 9428
rect 45484 9388 45524 9428
rect 49516 9388 49556 9428
rect 56140 9388 56180 9428
rect 60268 9388 60308 9428
rect 61132 9388 61172 9428
rect 63148 9388 63188 9428
rect 72076 9388 72116 9428
rect 72268 9388 72308 9428
rect 73228 9388 73268 9428
rect 78604 9388 78644 9428
rect 45292 9304 45332 9344
rect 45868 9304 45908 9344
rect 63340 9304 63380 9344
rect 72172 9304 72212 9344
rect 652 9220 692 9260
rect 49228 9220 49268 9260
rect 52588 9220 52628 9260
rect 55852 9220 55892 9260
rect 56332 9220 56372 9260
rect 60076 9220 60116 9260
rect 61324 9220 61364 9260
rect 62668 9220 62708 9260
rect 68044 9220 68084 9260
rect 73420 9220 73460 9260
rect 78412 9220 78452 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 45100 8884 45140 8924
rect 50284 8884 50324 8924
rect 51244 8884 51284 8924
rect 55372 8884 55412 8924
rect 58060 8884 58100 8924
rect 62188 8884 62228 8924
rect 65932 8884 65972 8924
rect 68524 8884 68564 8924
rect 72940 8884 72980 8924
rect 74572 8884 74612 8924
rect 44428 8800 44468 8840
rect 45484 8800 45524 8840
rect 48364 8800 48404 8840
rect 50668 8800 50708 8840
rect 52300 8800 52340 8840
rect 58732 8800 58772 8840
rect 59116 8800 59156 8840
rect 63052 8800 63092 8840
rect 63532 8800 63572 8840
rect 74188 8800 74228 8840
rect 76492 8800 76532 8840
rect 844 8716 884 8756
rect 44620 8716 44660 8756
rect 45388 8716 45428 8756
rect 45580 8716 45620 8756
rect 49708 8716 49748 8756
rect 50092 8716 50132 8756
rect 50572 8716 50612 8756
rect 50764 8716 50804 8756
rect 58636 8716 58676 8756
rect 58828 8716 58868 8756
rect 62956 8716 62996 8756
rect 63148 8716 63188 8756
rect 69388 8716 69428 8756
rect 69676 8716 69716 8756
rect 73996 8727 74036 8767
rect 76396 8716 76436 8756
rect 76588 8716 76628 8756
rect 79276 8716 79316 8756
rect 44812 8632 44852 8672
rect 44908 8632 44948 8672
rect 45100 8632 45140 8672
rect 45676 8632 45716 8672
rect 47500 8632 47540 8672
rect 47596 8632 47636 8672
rect 45292 8590 45332 8630
rect 47788 8632 47828 8672
rect 48652 8632 48692 8672
rect 48748 8632 48788 8672
rect 49132 8632 49172 8672
rect 49228 8632 49268 8672
rect 49324 8632 49364 8672
rect 50476 8632 50516 8672
rect 50860 8632 50900 8672
rect 51532 8632 51572 8672
rect 51628 8632 51668 8672
rect 52012 8632 52052 8672
rect 52972 8632 53012 8672
rect 53164 8632 53204 8672
rect 54892 8632 54932 8672
rect 55084 8632 55124 8672
rect 55180 8632 55220 8672
rect 55468 8632 55508 8672
rect 56044 8632 56084 8672
rect 56908 8632 56948 8672
rect 58540 8632 58580 8672
rect 58924 8632 58964 8672
rect 59116 8632 59156 8672
rect 59308 8632 59348 8672
rect 59404 8632 59444 8672
rect 60172 8632 60212 8672
rect 61036 8632 61076 8672
rect 62860 8632 62900 8672
rect 63244 8632 63284 8672
rect 63820 8632 63860 8672
rect 63916 8622 63956 8662
rect 64204 8632 64244 8672
rect 64300 8632 64340 8672
rect 64396 8632 64436 8672
rect 64492 8632 64532 8672
rect 67084 8632 67124 8672
rect 67948 8632 67988 8672
rect 68812 8632 68852 8672
rect 68908 8632 68948 8672
rect 70828 8632 70868 8672
rect 71692 8632 71732 8672
rect 72076 8632 72116 8672
rect 72460 8632 72500 8672
rect 72556 8632 72596 8672
rect 72652 8632 72692 8672
rect 72844 8632 72884 8672
rect 74476 8632 74516 8672
rect 76300 8632 76340 8672
rect 76684 8632 76724 8672
rect 76876 8632 76916 8672
rect 77260 8632 77300 8672
rect 78124 8632 78164 8672
rect 55660 8548 55700 8588
rect 59788 8548 59828 8588
rect 68332 8548 68372 8588
rect 652 8464 692 8504
rect 47692 8464 47732 8504
rect 48844 8460 48884 8500
rect 49036 8464 49076 8504
rect 49900 8464 49940 8504
rect 54988 8464 55028 8504
rect 69196 8464 69236 8504
rect 72364 8464 72404 8504
rect 51724 8406 51764 8446
rect 64012 8406 64052 8446
rect 69004 8406 69044 8446
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 47596 8128 47636 8168
rect 50284 8128 50324 8168
rect 53356 8128 53396 8168
rect 54700 8132 54740 8172
rect 55372 8128 55412 8168
rect 58348 8128 58388 8168
rect 59020 8128 59060 8168
rect 59404 8132 59444 8172
rect 60076 8128 60116 8168
rect 66220 8128 66260 8168
rect 66700 8128 66740 8168
rect 71980 8159 72020 8199
rect 77452 8186 77492 8226
rect 75052 8128 75092 8168
rect 77836 8128 77876 8168
rect 78028 8128 78068 8168
rect 45196 8044 45236 8084
rect 62188 8044 62228 8084
rect 72652 8044 72692 8084
rect 45580 7960 45620 8000
rect 46444 7960 46484 8000
rect 47884 7960 47924 8000
rect 48268 7960 48308 8000
rect 49132 7960 49172 8000
rect 50668 7960 50708 8000
rect 51052 7960 51092 8000
rect 51916 7960 51956 8000
rect 53452 7960 53492 8000
rect 53836 7960 53876 8000
rect 53932 7960 53972 8000
rect 54124 7960 54164 8000
rect 54508 7960 54548 8000
rect 54796 7960 54836 8000
rect 54892 7960 54932 8000
rect 55468 7960 55508 8000
rect 55564 7960 55604 8000
rect 55660 7960 55700 8000
rect 55852 7960 55892 8000
rect 55948 7960 55988 8000
rect 56044 7960 56084 8000
rect 56140 7960 56180 8000
rect 58444 7960 58484 8000
rect 59500 7960 59540 8000
rect 59596 7960 59636 8000
rect 60172 7960 60212 8000
rect 60268 7960 60308 8000
rect 60364 7960 60404 8000
rect 60556 7960 60596 8000
rect 60652 7960 60692 8000
rect 60748 7960 60788 8000
rect 60844 7960 60884 8000
rect 62572 7960 62612 8000
rect 63436 7960 63476 8000
rect 65740 7960 65780 8000
rect 65836 7960 65876 8000
rect 65932 7960 65972 8000
rect 66028 7960 66068 8000
rect 66412 7960 66452 8000
rect 844 7876 884 7916
rect 53068 7876 53108 7916
rect 54220 7876 54260 7916
rect 66316 7918 66356 7958
rect 66508 7960 66548 8000
rect 66796 7960 66836 8000
rect 67948 7960 67988 8000
rect 68332 7960 68372 8000
rect 71500 7960 71540 8000
rect 71692 7960 71732 8000
rect 71788 7960 71828 8000
rect 72076 7960 72116 8000
rect 72172 7960 72212 8000
rect 73036 7960 73076 8000
rect 73900 7960 73940 8000
rect 76492 7960 76532 8000
rect 76588 7960 76628 8000
rect 76684 7960 76724 8000
rect 76780 7960 76820 8000
rect 77260 7960 77300 8000
rect 77356 7960 77396 8000
rect 78124 7960 78164 8000
rect 54412 7876 54452 7916
rect 58636 7876 58676 7916
rect 59212 7876 59252 7916
rect 64972 7876 65012 7916
rect 68044 7876 68084 7916
rect 68236 7876 68276 7916
rect 68908 7876 68948 7916
rect 69100 7876 69140 7916
rect 77644 7876 77684 7916
rect 54316 7792 54356 7832
rect 68140 7792 68180 7832
rect 76972 7792 77012 7832
rect 652 7708 692 7748
rect 47596 7708 47636 7748
rect 53356 7708 53396 7748
rect 55180 7708 55220 7748
rect 58828 7708 58868 7748
rect 59884 7708 59924 7748
rect 64588 7708 64628 7748
rect 64780 7708 64820 7748
rect 68716 7708 68756 7748
rect 69292 7708 69332 7748
rect 71500 7708 71540 7748
rect 72460 7708 72500 7748
rect 77836 7708 77876 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 46828 7372 46868 7412
rect 50380 7372 50420 7412
rect 54604 7372 54644 7412
rect 59500 7372 59540 7412
rect 64012 7372 64052 7412
rect 68524 7372 68564 7412
rect 48076 7288 48116 7328
rect 59884 7288 59924 7328
rect 64588 7288 64628 7328
rect 65644 7288 65684 7328
rect 844 7204 884 7244
rect 47980 7204 48020 7244
rect 48172 7204 48212 7244
rect 56236 7204 56276 7244
rect 59788 7204 59828 7244
rect 59980 7204 60020 7244
rect 68908 7204 68948 7244
rect 73516 7204 73556 7244
rect 46924 7120 46964 7160
rect 47884 7120 47924 7160
rect 48268 7120 48308 7160
rect 50092 7120 50132 7160
rect 50188 7120 50228 7160
rect 50380 7120 50420 7160
rect 51724 7120 51764 7160
rect 51820 7120 51860 7160
rect 51916 7120 51956 7160
rect 52012 7120 52052 7160
rect 52204 7120 52244 7160
rect 52588 7120 52628 7160
rect 53452 7120 53492 7160
rect 56620 7120 56660 7160
rect 57100 7120 57140 7160
rect 57484 7120 57524 7160
rect 58348 7120 58388 7160
rect 59692 7120 59732 7160
rect 60076 7120 60116 7160
rect 61612 7120 61652 7160
rect 61708 7120 61748 7160
rect 61804 7120 61844 7160
rect 62092 7120 62132 7160
rect 62188 7120 62228 7160
rect 64108 7120 64148 7160
rect 64300 7120 64340 7160
rect 64396 7120 64436 7160
rect 65260 7163 65300 7203
rect 64588 7120 64628 7160
rect 64876 7120 64916 7160
rect 65356 7120 65396 7160
rect 66124 7120 66164 7160
rect 66508 7120 66548 7160
rect 67372 7120 67412 7160
rect 70444 7120 70484 7160
rect 71308 7120 71348 7160
rect 72652 7120 72692 7160
rect 72748 7120 72788 7160
rect 73708 7120 73748 7160
rect 73804 7120 73844 7160
rect 73900 7120 73940 7160
rect 73996 7120 74036 7160
rect 74956 7120 74996 7160
rect 75628 7120 75668 7160
rect 76012 7120 76052 7160
rect 76876 7120 76916 7160
rect 78220 7120 78260 7160
rect 78412 7120 78452 7160
rect 78508 7120 78548 7160
rect 78700 7120 78740 7160
rect 56716 7036 56756 7076
rect 70060 7036 70100 7076
rect 75052 7036 75092 7076
rect 78316 7036 78356 7076
rect 652 6952 692 6992
rect 56044 6952 56084 6992
rect 61516 6952 61556 6992
rect 64972 6952 65012 6992
rect 68716 6952 68756 6992
rect 72460 6952 72500 6992
rect 73324 6952 73364 6992
rect 78028 6952 78068 6992
rect 78796 6952 78836 6992
rect 65164 6894 65204 6934
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 52780 6620 52820 6660
rect 57964 6616 58004 6656
rect 59980 6616 60020 6656
rect 63532 6616 63572 6656
rect 63724 6616 63764 6656
rect 70828 6616 70868 6656
rect 72748 6616 72788 6656
rect 75628 6616 75668 6656
rect 79468 6616 79508 6656
rect 55084 6532 55124 6572
rect 55564 6532 55604 6572
rect 73228 6532 73268 6572
rect 52588 6448 52628 6488
rect 52684 6448 52724 6488
rect 52972 6448 53012 6488
rect 53164 6448 53204 6488
rect 53278 6455 53318 6495
rect 53452 6448 53492 6488
rect 53548 6448 53588 6488
rect 53644 6448 53684 6488
rect 53740 6448 53780 6488
rect 55180 6448 55220 6488
rect 55276 6448 55316 6488
rect 55372 6448 55412 6488
rect 55948 6448 55988 6488
rect 56812 6448 56852 6488
rect 59788 6448 59828 6488
rect 59884 6448 59924 6488
rect 60076 6448 60116 6488
rect 60652 6448 60692 6488
rect 60748 6448 60788 6488
rect 60844 6448 60884 6488
rect 60940 6448 60980 6488
rect 61132 6448 61172 6488
rect 61516 6448 61556 6488
rect 62380 6448 62420 6488
rect 64876 6448 64916 6488
rect 65740 6448 65780 6488
rect 66124 6448 66164 6488
rect 67948 6448 67988 6488
rect 68044 6448 68084 6488
rect 68140 6469 68180 6509
rect 68236 6448 68276 6488
rect 68428 6448 68468 6488
rect 68812 6448 68852 6488
rect 69676 6448 69716 6488
rect 71500 6448 71540 6488
rect 71884 6448 71924 6488
rect 72268 6448 72308 6488
rect 72460 6448 72500 6488
rect 72556 6448 72596 6488
rect 72844 6448 72884 6488
rect 72940 6448 72980 6488
rect 73036 6448 73076 6488
rect 73612 6448 73652 6488
rect 74476 6448 74516 6488
rect 76492 6448 76532 6488
rect 76876 6448 76916 6488
rect 77068 6448 77108 6488
rect 77452 6448 77492 6488
rect 78316 6448 78356 6488
rect 71596 6364 71636 6404
rect 71788 6364 71828 6404
rect 76588 6364 76628 6404
rect 76780 6364 76820 6404
rect 52300 6280 52340 6320
rect 71692 6280 71732 6320
rect 76684 6280 76724 6320
rect 52972 6196 53012 6236
rect 72268 6196 72308 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 77164 5860 77204 5900
rect 55180 5776 55220 5816
rect 60940 5776 60980 5816
rect 64684 5776 64724 5816
rect 68620 5776 68660 5816
rect 72460 5776 72500 5816
rect 72940 5776 72980 5816
rect 844 5692 884 5732
rect 58060 5692 58100 5732
rect 64588 5692 64628 5732
rect 64780 5692 64820 5732
rect 72364 5692 72404 5732
rect 72556 5692 72596 5732
rect 76876 5692 76916 5732
rect 52108 5608 52148 5648
rect 52972 5608 53012 5648
rect 55468 5608 55508 5648
rect 55564 5608 55604 5648
rect 55948 5608 55988 5648
rect 56044 5608 56084 5648
rect 56140 5608 56180 5648
rect 56236 5608 56276 5648
rect 57964 5608 58004 5648
rect 59404 5608 59444 5648
rect 60268 5608 60308 5648
rect 61228 5608 61268 5648
rect 61324 5608 61364 5648
rect 64492 5608 64532 5648
rect 64876 5608 64916 5648
rect 65164 5608 65204 5648
rect 65260 5608 65300 5648
rect 65356 5608 65396 5648
rect 65644 5608 65684 5648
rect 65740 5608 65780 5648
rect 65836 5608 65876 5648
rect 68140 5608 68180 5648
rect 68332 5608 68372 5648
rect 68428 5608 68468 5648
rect 68908 5608 68948 5648
rect 69004 5608 69044 5648
rect 69388 5608 69428 5648
rect 69484 5608 69524 5648
rect 69580 5608 69620 5648
rect 69676 5608 69716 5648
rect 72268 5608 72308 5648
rect 72652 5608 72692 5648
rect 73228 5608 73268 5648
rect 73324 5608 73364 5648
rect 74284 5608 74324 5648
rect 74380 5608 74420 5648
rect 74476 5608 74516 5648
rect 74572 5608 74612 5648
rect 76972 5608 77012 5648
rect 77452 5608 77492 5648
rect 77548 5608 77588 5648
rect 77836 5608 77876 5648
rect 77932 5608 77972 5648
rect 78028 5608 78068 5648
rect 78124 5608 78164 5648
rect 78412 5608 78452 5648
rect 51724 5524 51764 5564
rect 60652 5524 60692 5564
rect 68236 5524 68276 5564
rect 652 5440 692 5480
rect 54124 5440 54164 5480
rect 58252 5440 58292 5480
rect 65068 5440 65108 5480
rect 65548 5440 65588 5480
rect 73420 5436 73460 5476
rect 55660 5382 55700 5422
rect 61420 5382 61460 5422
rect 77644 5436 77684 5476
rect 78316 5440 78356 5480
rect 69100 5382 69140 5422
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 55756 5104 55796 5144
rect 61612 5104 61652 5144
rect 62284 5104 62324 5144
rect 65068 5108 65108 5148
rect 67756 5104 67796 5144
rect 70348 5104 70388 5144
rect 73228 5104 73268 5144
rect 74380 5104 74420 5144
rect 76972 5104 77012 5144
rect 77740 5104 77780 5144
rect 60556 5020 60596 5060
rect 65356 5020 65396 5060
rect 70540 5020 70580 5060
rect 52204 4936 52244 4976
rect 52588 4936 52628 4976
rect 53452 4936 53492 4976
rect 53932 4936 53972 4976
rect 54028 4936 54068 4976
rect 54220 4936 54260 4976
rect 54412 4936 54452 4976
rect 54796 4936 54836 4976
rect 55852 4936 55892 4976
rect 56908 4936 56948 4976
rect 57004 4936 57044 4976
rect 57100 4936 57140 4976
rect 57196 4936 57236 4976
rect 57388 4936 57428 4976
rect 57772 4936 57812 4976
rect 58636 4936 58676 4976
rect 60460 4936 60500 4976
rect 60748 4936 60788 4976
rect 61132 4936 61172 4976
rect 62188 4936 62228 4976
rect 64108 4951 64148 4991
rect 64204 4922 64244 4962
rect 64396 4936 64436 4976
rect 64876 4936 64916 4976
rect 64972 4936 65012 4976
rect 65740 4936 65780 4976
rect 66604 4936 66644 4976
rect 67948 4936 67988 4976
rect 68332 4936 68372 4976
rect 69196 4936 69236 4976
rect 70924 4936 70964 4976
rect 71788 4936 71828 4976
rect 73132 4936 73172 4976
rect 74284 4936 74324 4976
rect 74572 4936 74612 4976
rect 74956 4936 74996 4976
rect 75820 4936 75860 4976
rect 77356 4936 77396 4976
rect 844 4852 884 4892
rect 52300 4852 52340 4892
rect 52492 4852 52532 4892
rect 53356 4852 53396 4892
rect 54508 4852 54548 4892
rect 54700 4852 54740 4892
rect 60844 4852 60884 4892
rect 77164 4894 77204 4934
rect 61036 4852 61076 4892
rect 61420 4852 61460 4892
rect 61804 4852 61844 4892
rect 77260 4894 77300 4934
rect 77452 4936 77492 4976
rect 77644 4936 77684 4976
rect 77836 4936 77876 4976
rect 77932 4936 77972 4976
rect 652 4768 692 4808
rect 52396 4768 52436 4808
rect 54604 4768 54644 4808
rect 59788 4768 59828 4808
rect 60940 4768 60980 4808
rect 64588 4768 64628 4808
rect 54220 4684 54260 4724
rect 61612 4684 61652 4724
rect 61996 4684 62036 4724
rect 62284 4684 62324 4724
rect 64396 4684 64436 4724
rect 72940 4684 72980 4724
rect 74380 4684 74420 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 65836 4348 65876 4388
rect 69292 4348 69332 4388
rect 56236 4264 56276 4304
rect 57004 4264 57044 4304
rect 63052 4264 63092 4304
rect 68524 4264 68564 4304
rect 68908 4264 68948 4304
rect 71692 4264 71732 4304
rect 72556 4264 72596 4304
rect 75148 4264 75188 4304
rect 76300 4264 76340 4304
rect 844 4180 884 4220
rect 66028 4180 66068 4220
rect 68428 4180 68468 4220
rect 68620 4180 68660 4220
rect 69100 4180 69140 4220
rect 71596 4180 71636 4220
rect 71788 4180 71828 4220
rect 79372 4180 79412 4220
rect 53836 4096 53876 4136
rect 54220 4096 54260 4136
rect 55084 4096 55124 4136
rect 56428 4096 56468 4136
rect 56524 4096 56564 4136
rect 56716 4096 56756 4136
rect 57292 4096 57332 4136
rect 57388 4096 57428 4136
rect 57676 4096 57716 4136
rect 57772 4096 57812 4136
rect 57868 4096 57908 4136
rect 57964 4096 58004 4136
rect 60268 4096 60308 4136
rect 60364 4096 60404 4136
rect 60460 4096 60500 4136
rect 61036 4096 61076 4136
rect 61900 4096 61940 4136
rect 63628 4096 63668 4136
rect 64492 4096 64532 4136
rect 68332 4096 68372 4136
rect 68716 4096 68756 4136
rect 69388 4096 69428 4136
rect 71020 4096 71060 4136
rect 71212 4096 71252 4136
rect 71308 4096 71348 4136
rect 71500 4096 71540 4136
rect 71884 4096 71924 4136
rect 72172 4096 72212 4136
rect 72268 4096 72308 4136
rect 73132 4096 73172 4136
rect 73996 4096 74036 4136
rect 75820 4096 75860 4136
rect 75916 4096 75956 4136
rect 76012 4096 76052 4136
rect 76108 4096 76148 4136
rect 76588 4096 76628 4136
rect 76684 4096 76724 4136
rect 77356 4096 77396 4136
rect 78220 4096 78260 4136
rect 60172 4012 60212 4052
rect 60652 4012 60692 4052
rect 63244 4012 63284 4052
rect 72748 4012 72788 4052
rect 76972 4012 77012 4052
rect 652 3928 692 3968
rect 56620 3928 56660 3968
rect 65644 3928 65684 3968
rect 71116 3928 71156 3968
rect 72076 3924 72116 3964
rect 57484 3870 57524 3910
rect 76780 3870 76820 3910
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 5164 3592 5204 3632
rect 60268 3596 60308 3636
rect 61420 3592 61460 3632
rect 61804 3592 61844 3632
rect 64876 3592 64916 3632
rect 68812 3592 68852 3632
rect 69004 3592 69044 3632
rect 72748 3592 72788 3632
rect 73036 3592 73076 3632
rect 73996 3592 74036 3632
rect 77836 3592 77876 3632
rect 69676 3508 69716 3548
rect 5068 3424 5108 3464
rect 56044 3424 56084 3464
rect 56428 3424 56468 3464
rect 57292 3424 57332 3464
rect 60076 3424 60116 3464
rect 60172 3424 60212 3464
rect 60556 3424 60596 3464
rect 60652 3424 60692 3464
rect 60748 3424 60788 3464
rect 60844 3424 60884 3464
rect 61324 3424 61364 3464
rect 61516 3424 61556 3464
rect 61612 3405 61652 3445
rect 64300 3424 64340 3464
rect 64684 3424 64724 3464
rect 64972 3424 65012 3464
rect 65452 3424 65492 3464
rect 65548 3424 65588 3464
rect 65644 3424 65684 3464
rect 65740 3424 65780 3464
rect 65932 3424 65972 3464
rect 66028 3424 66068 3464
rect 66124 3424 66164 3464
rect 66220 3424 66260 3464
rect 66412 3424 66452 3464
rect 66796 3424 66836 3464
rect 67660 3424 67700 3464
rect 70060 3424 70100 3464
rect 70924 3424 70964 3464
rect 72460 3424 72500 3464
rect 72556 3424 72596 3464
rect 72652 3424 72692 3464
rect 72940 3424 72980 3464
rect 73516 3424 73556 3464
rect 74092 3424 74132 3464
rect 74188 3424 74228 3464
rect 74284 3424 74324 3464
rect 76684 3424 76724 3464
rect 76972 3424 77012 3464
rect 77356 3424 77396 3464
rect 78028 3424 78068 3464
rect 78124 3424 78164 3464
rect 844 3340 884 3380
rect 61996 3340 62036 3380
rect 64396 3340 64436 3380
rect 64588 3340 64628 3380
rect 69196 3340 69236 3380
rect 77068 3340 77108 3380
rect 77260 3340 77300 3380
rect 77644 3340 77684 3380
rect 59788 3256 59828 3296
rect 64492 3256 64532 3296
rect 76780 3256 76820 3296
rect 77164 3256 77204 3296
rect 652 3172 692 3212
rect 58444 3172 58484 3212
rect 72076 3172 72116 3212
rect 73420 3172 73460 3212
rect 77836 3172 77876 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 57868 2836 57908 2876
rect 60172 2836 60212 2876
rect 63340 2836 63380 2876
rect 68620 2836 68660 2876
rect 73804 2836 73844 2876
rect 75052 2836 75092 2876
rect 77356 2836 77396 2876
rect 56524 2752 56564 2792
rect 58732 2752 58772 2792
rect 59116 2752 59156 2792
rect 60748 2752 60788 2792
rect 61132 2752 61172 2792
rect 61708 2752 61748 2792
rect 65068 2752 65108 2792
rect 66028 2752 66068 2792
rect 71980 2752 72020 2792
rect 72364 2752 72404 2792
rect 76588 2752 76628 2792
rect 844 2668 884 2708
rect 56428 2668 56468 2708
rect 56620 2668 56660 2708
rect 59020 2668 59060 2708
rect 59212 2668 59252 2708
rect 61036 2668 61076 2708
rect 61228 2668 61268 2708
rect 64972 2668 65012 2708
rect 65164 2668 65204 2708
rect 71884 2668 71924 2708
rect 72076 2668 72116 2708
rect 56332 2584 56372 2624
rect 56716 2584 56756 2624
rect 57964 2584 58004 2624
rect 58444 2584 58484 2624
rect 58540 2584 58580 2624
rect 58732 2584 58772 2624
rect 58924 2584 58964 2624
rect 59308 2584 59348 2624
rect 60268 2584 60308 2624
rect 60460 2584 60500 2624
rect 60556 2584 60596 2624
rect 60748 2584 60788 2624
rect 60940 2584 60980 2624
rect 61324 2584 61364 2624
rect 61996 2584 62036 2624
rect 62092 2584 62132 2624
rect 62476 2584 62516 2624
rect 62572 2584 62612 2624
rect 62668 2584 62708 2624
rect 62860 2584 62900 2624
rect 63244 2584 63284 2624
rect 64396 2584 64436 2624
rect 64588 2584 64628 2624
rect 64684 2584 64724 2624
rect 64876 2584 64916 2624
rect 65260 2584 65300 2624
rect 65644 2584 65684 2624
rect 65740 2584 65780 2624
rect 66604 2584 66644 2624
rect 66700 2584 66740 2624
rect 66892 2584 66932 2624
rect 68236 2584 68276 2624
rect 68332 2584 68372 2624
rect 68428 2584 68468 2624
rect 68620 2584 68660 2624
rect 68812 2584 68852 2624
rect 68908 2584 68948 2624
rect 69196 2584 69236 2624
rect 71308 2584 71348 2624
rect 71500 2584 71540 2624
rect 71596 2584 71636 2624
rect 71788 2584 71828 2624
rect 72172 2584 72212 2624
rect 72652 2584 72692 2624
rect 72748 2584 72788 2624
rect 73132 2584 73172 2624
rect 74092 2584 74132 2624
rect 74956 2584 74996 2624
rect 76108 2584 76148 2624
rect 76204 2584 76244 2624
rect 76300 2584 76340 2624
rect 76876 2584 76916 2624
rect 76972 2584 77012 2624
rect 77356 2584 77396 2624
rect 77548 2584 77588 2624
rect 77644 2584 77684 2624
rect 77932 2584 77972 2624
rect 64492 2500 64532 2540
rect 77836 2500 77876 2540
rect 652 2416 692 2456
rect 62188 2412 62228 2452
rect 62380 2416 62420 2456
rect 62956 2416 62996 2456
rect 66796 2416 66836 2456
rect 68140 2416 68180 2456
rect 69100 2416 69140 2456
rect 71404 2416 71444 2456
rect 72844 2412 72884 2452
rect 75052 2416 75092 2456
rect 76396 2416 76436 2456
rect 65548 2358 65588 2398
rect 77068 2358 77108 2398
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 68620 2138 68660 2178
rect 60748 2080 60788 2120
rect 64780 2080 64820 2120
rect 71212 2080 71252 2120
rect 73804 2080 73844 2120
rect 73996 2080 74036 2120
rect 78412 2080 78452 2120
rect 58348 1996 58388 2036
rect 62380 1996 62420 2036
rect 64972 1996 65012 2036
rect 68812 1996 68852 2036
rect 71404 1996 71444 2036
rect 58732 1912 58772 1952
rect 59596 1912 59636 1952
rect 61324 1912 61364 1952
rect 62764 1912 62804 1952
rect 63628 1912 63668 1952
rect 65356 1912 65396 1952
rect 66220 1912 66260 1952
rect 67564 1912 67604 1952
rect 67948 1912 67988 1952
rect 68428 1912 68468 1952
rect 67660 1870 67700 1910
rect 68524 1912 68564 1952
rect 69196 1912 69236 1952
rect 70060 1912 70100 1952
rect 71788 1912 71828 1952
rect 72652 1912 72692 1952
rect 74092 1912 74132 1952
rect 74188 1912 74228 1952
rect 74284 1912 74324 1952
rect 74476 1912 74516 1952
rect 74572 1912 74612 1952
rect 74764 1912 74804 1952
rect 75436 1912 75476 1952
rect 75820 1912 75860 1952
rect 76012 1912 76052 1952
rect 76396 1912 76436 1952
rect 77260 1912 77300 1952
rect 67852 1828 67892 1868
rect 75532 1828 75572 1868
rect 75724 1828 75764 1868
rect 61900 1744 61940 1784
rect 67756 1744 67796 1784
rect 68140 1744 68180 1784
rect 74764 1744 74804 1784
rect 75628 1744 75668 1784
rect 67372 1660 67412 1700
rect 71212 1660 71252 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 62284 1324 62324 1364
rect 66124 1324 66164 1364
rect 69196 1324 69236 1364
rect 70732 1324 70772 1364
rect 72268 1324 72308 1364
rect 75628 1324 75668 1364
rect 79372 1156 79412 1196
rect 59596 1072 59636 1112
rect 59884 1072 59924 1112
rect 60268 1072 60308 1112
rect 61132 1072 61172 1112
rect 62572 1072 62612 1112
rect 62668 1072 62708 1112
rect 62764 1072 62804 1112
rect 62860 1072 62900 1112
rect 66220 1072 66260 1112
rect 66796 1072 66836 1112
rect 67180 1072 67220 1112
rect 68044 1072 68084 1112
rect 69484 1072 69524 1112
rect 69580 1072 69620 1112
rect 69676 1072 69716 1112
rect 69772 1072 69812 1112
rect 70060 1072 70100 1112
rect 70252 1072 70292 1112
rect 71116 1072 71156 1112
rect 71500 1072 71540 1112
rect 71596 1072 71636 1112
rect 71692 1072 71732 1112
rect 72844 1072 72884 1112
rect 73612 1072 73652 1112
rect 74476 1072 74516 1112
rect 76492 1072 76532 1112
rect 76588 1072 76628 1112
rect 76684 1072 76724 1112
rect 76780 1072 76820 1112
rect 76972 1072 77012 1112
rect 77356 1072 77396 1112
rect 78220 1072 78260 1112
rect 71788 988 71828 1028
rect 73228 988 73268 1028
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 69579 38408 69621 38417
rect 75915 38408 75957 38417
rect 69579 38368 69580 38408
rect 69620 38368 69621 38408
rect 69579 38359 69621 38368
rect 69868 38368 70196 38408
rect 57676 38240 57716 38249
rect 59884 38240 59924 38249
rect 57716 38200 58580 38240
rect 57676 38191 57716 38200
rect 652 38156 692 38165
rect 652 37577 692 38116
rect 844 37988 884 37997
rect 651 37568 693 37577
rect 651 37528 652 37568
rect 692 37528 693 37568
rect 651 37519 693 37528
rect 844 37460 884 37948
rect 57580 37988 57620 37997
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 56620 37484 56660 37493
rect 844 37420 1364 37460
rect 843 26564 885 26573
rect 843 26524 844 26564
rect 884 26524 885 26564
rect 843 26515 885 26524
rect 844 26312 884 26515
rect 844 26263 884 26272
rect 652 26060 692 26069
rect 652 25817 692 26020
rect 651 25808 693 25817
rect 651 25768 652 25808
rect 692 25768 693 25808
rect 651 25759 693 25768
rect 652 25388 692 25397
rect 652 24977 692 25348
rect 844 25136 884 25145
rect 884 25096 1076 25136
rect 844 25087 884 25096
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 844 24800 884 24809
rect 844 24557 884 24760
rect 652 24548 692 24557
rect 652 24137 692 24508
rect 843 24548 885 24557
rect 843 24508 844 24548
rect 884 24508 885 24548
rect 843 24499 885 24508
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23876 692 23885
rect 652 23297 692 23836
rect 844 23624 884 23633
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 844 23129 884 23584
rect 939 23288 981 23297
rect 939 23248 940 23288
rect 980 23248 981 23288
rect 939 23239 981 23248
rect 843 23120 885 23129
rect 843 23080 844 23120
rect 884 23080 885 23120
rect 843 23071 885 23080
rect 652 23036 692 23045
rect 556 22996 652 23036
rect 556 22457 596 22996
rect 652 22987 692 22996
rect 844 22952 884 22961
rect 940 22952 980 23239
rect 884 22912 980 22952
rect 844 22903 884 22912
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 1036 21533 1076 25096
rect 1035 21524 1077 21533
rect 1035 21484 1036 21524
rect 1076 21484 1077 21524
rect 1035 21475 1077 21484
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 1324 20852 1364 37420
rect 56523 37400 56565 37409
rect 56523 37360 56524 37400
rect 56564 37360 56565 37400
rect 56523 37351 56565 37360
rect 56524 37266 56564 37351
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 56620 36896 56660 37444
rect 56812 37484 56852 37493
rect 56428 36856 56660 36896
rect 56716 37274 56756 37283
rect 56235 36812 56277 36821
rect 56235 36772 56236 36812
rect 56276 36772 56277 36812
rect 56235 36763 56277 36772
rect 36651 36728 36693 36737
rect 36651 36688 36652 36728
rect 36692 36688 36693 36728
rect 36651 36679 36693 36688
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 29739 29924 29781 29933
rect 29739 29884 29740 29924
rect 29780 29884 29781 29924
rect 29739 29875 29781 29884
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 7179 25556 7221 25565
rect 7084 25516 7180 25556
rect 7220 25516 7221 25556
rect 2379 25220 2421 25229
rect 2379 25180 2380 25220
rect 2420 25180 2421 25220
rect 2379 25171 2421 25180
rect 2380 24809 2420 25171
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 1803 24800 1845 24809
rect 1803 24760 1804 24800
rect 1844 24760 1845 24800
rect 1803 24751 1845 24760
rect 2379 24800 2421 24809
rect 2379 24760 2380 24800
rect 2420 24760 2421 24800
rect 2379 24751 2421 24760
rect 1804 24548 1844 24751
rect 2380 24666 2420 24751
rect 1804 24499 1844 24508
rect 2187 24548 2229 24557
rect 2187 24508 2188 24548
rect 2228 24508 2229 24548
rect 2187 24499 2229 24508
rect 2188 24414 2228 24499
rect 1996 24380 2036 24389
rect 1996 23885 2036 24340
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 1804 23876 1844 23885
rect 1612 23624 1652 23633
rect 1804 23624 1844 23836
rect 1995 23876 2037 23885
rect 1995 23836 1996 23876
rect 2036 23836 2037 23876
rect 1995 23827 2037 23836
rect 2187 23876 2229 23885
rect 2187 23836 2188 23876
rect 2228 23836 2229 23876
rect 2187 23827 2229 23836
rect 2188 23742 2228 23827
rect 1996 23624 2036 23633
rect 1652 23584 1748 23624
rect 1804 23584 1996 23624
rect 2036 23584 2132 23624
rect 1612 23575 1652 23584
rect 1516 23129 1556 23214
rect 1515 23120 1557 23129
rect 1515 23080 1516 23120
rect 1556 23080 1557 23120
rect 1515 23071 1557 23080
rect 1708 23120 1748 23584
rect 1996 23575 2036 23584
rect 1611 23036 1653 23045
rect 1611 22996 1612 23036
rect 1652 22996 1653 23036
rect 1611 22987 1653 22996
rect 1612 22902 1652 22987
rect 1708 20945 1748 23080
rect 1707 20936 1749 20945
rect 1707 20896 1708 20936
rect 1748 20896 1749 20936
rect 1707 20887 1749 20896
rect 1324 20803 1364 20812
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 1899 20768 1941 20777
rect 1899 20728 1900 20768
rect 1940 20728 1941 20768
rect 1899 20719 1941 20728
rect 1515 20600 1557 20609
rect 1420 20560 1516 20600
rect 1556 20560 1557 20600
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19424 692 19879
rect 652 19375 692 19384
rect 748 19844 788 19853
rect 748 19349 788 19804
rect 1227 19508 1269 19517
rect 1227 19468 1228 19508
rect 1268 19468 1269 19508
rect 1227 19459 1269 19468
rect 1228 19374 1268 19459
rect 747 19340 789 19349
rect 747 19300 748 19340
rect 788 19300 789 19340
rect 747 19291 789 19300
rect 1420 19340 1460 20560
rect 1515 20551 1557 20560
rect 1516 20466 1556 20551
rect 1707 20096 1749 20105
rect 1707 20056 1708 20096
rect 1748 20056 1749 20096
rect 1707 20047 1749 20056
rect 1900 20096 1940 20719
rect 1900 20047 1940 20056
rect 1420 19291 1460 19300
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 1612 19088 1652 19097
rect 652 18416 692 19039
rect 1323 19004 1365 19013
rect 1323 18964 1324 19004
rect 1364 18964 1365 19004
rect 1323 18955 1365 18964
rect 1227 18752 1269 18761
rect 1227 18712 1228 18752
rect 1268 18712 1269 18752
rect 1227 18703 1269 18712
rect 652 18367 692 18376
rect 1132 18332 1172 18341
rect 748 18292 1132 18332
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 18199
rect 652 17863 692 17872
rect 555 17576 597 17585
rect 555 17536 556 17576
rect 596 17536 597 17576
rect 555 17527 597 17536
rect 459 16064 501 16073
rect 459 16024 460 16064
rect 500 16024 501 16064
rect 459 16015 501 16024
rect 460 7757 500 16015
rect 459 7748 501 7757
rect 459 7708 460 7748
rect 500 7708 501 7748
rect 459 7699 501 7708
rect 556 2708 596 17527
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 16904 692 17359
rect 652 16855 692 16864
rect 652 16400 692 16409
rect 652 15737 692 16360
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 652 12234 692 12319
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 748 7244 788 18292
rect 1132 18283 1172 18292
rect 1228 18164 1268 18703
rect 1324 18500 1364 18955
rect 1612 18761 1652 19048
rect 1611 18752 1653 18761
rect 1611 18712 1612 18752
rect 1652 18712 1653 18752
rect 1611 18703 1653 18712
rect 1324 18451 1364 18460
rect 1708 18500 1748 20047
rect 1803 20012 1845 20021
rect 1803 19972 1804 20012
rect 1844 19972 1845 20012
rect 1803 19963 1845 19972
rect 1804 19340 1844 19963
rect 1804 19291 1844 19300
rect 1708 18451 1748 18460
rect 1996 19088 2036 19097
rect 1516 18332 1556 18341
rect 940 18124 1268 18164
rect 1420 18292 1516 18332
rect 844 15476 884 15487
rect 844 15401 884 15436
rect 843 15392 885 15401
rect 843 15352 844 15392
rect 884 15352 885 15392
rect 843 15343 885 15352
rect 844 14804 884 14813
rect 940 14804 980 18124
rect 1323 17828 1365 17837
rect 1323 17788 1324 17828
rect 1364 17788 1365 17828
rect 1323 17779 1365 17788
rect 1324 17694 1364 17779
rect 1131 17576 1173 17585
rect 1131 17536 1132 17576
rect 1172 17536 1173 17576
rect 1131 17527 1173 17536
rect 1132 17442 1172 17527
rect 1131 17324 1173 17333
rect 1131 17284 1132 17324
rect 1172 17284 1173 17324
rect 1420 17300 1460 18292
rect 1516 18283 1556 18292
rect 1707 17996 1749 18005
rect 1707 17956 1708 17996
rect 1748 17956 1749 17996
rect 1707 17947 1749 17956
rect 1708 17828 1748 17947
rect 1708 17779 1748 17788
rect 1131 17275 1173 17284
rect 1036 16904 1076 16913
rect 1036 16577 1076 16864
rect 1035 16568 1077 16577
rect 1035 16528 1036 16568
rect 1076 16528 1077 16568
rect 1035 16519 1077 16528
rect 884 14764 980 14804
rect 844 14755 884 14764
rect 843 13292 885 13301
rect 843 13252 844 13292
rect 884 13252 885 13292
rect 843 13243 885 13252
rect 844 13158 884 13243
rect 843 13040 885 13049
rect 1132 13040 1172 17275
rect 843 13000 844 13040
rect 884 13000 885 13040
rect 843 12991 885 13000
rect 1036 13000 1172 13040
rect 1324 17260 1460 17300
rect 1516 17576 1556 17585
rect 1516 17300 1556 17536
rect 1996 17333 2036 19048
rect 2092 18677 2132 23584
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 7084 23045 7124 25516
rect 7179 25507 7221 25516
rect 7180 25488 7220 25507
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 13707 23876 13749 23885
rect 13707 23836 13708 23876
rect 13748 23836 13749 23876
rect 13707 23827 13749 23836
rect 3627 23036 3669 23045
rect 3627 22996 3628 23036
rect 3668 22996 3669 23036
rect 3627 22987 3669 22996
rect 7083 23036 7125 23045
rect 7083 22996 7084 23036
rect 7124 22996 7125 23036
rect 7083 22987 7125 22996
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 3339 21524 3381 21533
rect 3339 21484 3340 21524
rect 3380 21484 3381 21524
rect 3339 21475 3381 21484
rect 3340 21390 3380 21475
rect 2763 21356 2805 21365
rect 2763 21316 2764 21356
rect 2804 21316 2805 21356
rect 2763 21307 2805 21316
rect 3531 21356 3573 21365
rect 3531 21316 3532 21356
rect 3572 21316 3573 21356
rect 3531 21307 3573 21316
rect 2764 20852 2804 21307
rect 3532 21222 3572 21307
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 3531 21020 3573 21029
rect 3531 20980 3532 21020
rect 3572 20980 3573 21020
rect 3531 20971 3573 20980
rect 3339 20936 3381 20945
rect 3339 20896 3340 20936
rect 3380 20896 3381 20936
rect 3339 20887 3381 20896
rect 2764 20803 2804 20812
rect 2859 20852 2901 20861
rect 2859 20812 2860 20852
rect 2900 20812 2901 20852
rect 2859 20803 2901 20812
rect 3243 20852 3285 20861
rect 3243 20812 3244 20852
rect 3284 20812 3285 20852
rect 3243 20803 3285 20812
rect 2763 20684 2805 20693
rect 2763 20644 2764 20684
rect 2804 20644 2805 20684
rect 2763 20635 2805 20644
rect 2764 20096 2804 20635
rect 2764 19517 2804 20056
rect 2763 19508 2805 19517
rect 2763 19468 2764 19508
rect 2804 19468 2805 19508
rect 2763 19459 2805 19468
rect 2187 19340 2229 19349
rect 2187 19300 2188 19340
rect 2228 19300 2229 19340
rect 2187 19291 2229 19300
rect 2188 19206 2228 19291
rect 2091 18668 2133 18677
rect 2091 18628 2092 18668
rect 2132 18628 2133 18668
rect 2091 18619 2133 18628
rect 1995 17324 2037 17333
rect 1516 17260 1844 17300
rect 1995 17284 1996 17324
rect 2036 17284 2037 17324
rect 1995 17275 2037 17284
rect 844 12452 884 12991
rect 844 12403 884 12412
rect 843 11780 885 11789
rect 843 11740 844 11780
rect 884 11740 885 11780
rect 843 11731 885 11740
rect 844 11646 884 11731
rect 843 11528 885 11537
rect 843 11488 844 11528
rect 884 11488 885 11528
rect 843 11479 885 11488
rect 844 10940 884 11479
rect 844 10891 884 10900
rect 843 10352 885 10361
rect 843 10312 844 10352
rect 884 10312 885 10352
rect 843 10303 885 10312
rect 844 10268 884 10303
rect 844 10217 884 10228
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 844 8756 884 8765
rect 1036 8756 1076 13000
rect 884 8716 1076 8756
rect 844 8707 884 8716
rect 844 7916 884 7925
rect 1324 7916 1364 17260
rect 1707 16316 1749 16325
rect 1707 16276 1708 16316
rect 1748 16276 1749 16316
rect 1707 16267 1749 16276
rect 1708 16182 1748 16267
rect 1516 16064 1556 16073
rect 1556 16024 1652 16064
rect 1516 16015 1556 16024
rect 1515 15392 1557 15401
rect 1515 15352 1516 15392
rect 1556 15352 1557 15392
rect 1515 15343 1557 15352
rect 1516 15258 1556 15343
rect 1516 13796 1556 13805
rect 1516 13301 1556 13756
rect 1515 13292 1557 13301
rect 1515 13252 1516 13292
rect 1556 13252 1557 13292
rect 1515 13243 1557 13252
rect 1515 13040 1557 13049
rect 1515 13000 1516 13040
rect 1556 13000 1557 13040
rect 1515 12991 1557 13000
rect 1516 12906 1556 12991
rect 1516 12284 1556 12293
rect 1516 11789 1556 12244
rect 1515 11780 1557 11789
rect 1515 11740 1516 11780
rect 1556 11740 1557 11780
rect 1515 11731 1557 11740
rect 1419 11612 1461 11621
rect 1419 11572 1420 11612
rect 1460 11572 1556 11612
rect 1419 11563 1461 11572
rect 1516 11528 1556 11572
rect 1516 11479 1556 11488
rect 1612 11360 1652 16024
rect 1707 15476 1749 15485
rect 1707 15436 1708 15476
rect 1748 15436 1749 15476
rect 1707 15427 1749 15436
rect 1708 15342 1748 15427
rect 1707 13964 1749 13973
rect 1707 13924 1708 13964
rect 1748 13924 1749 13964
rect 1707 13915 1749 13924
rect 1708 13830 1748 13915
rect 1707 13292 1749 13301
rect 1707 13252 1708 13292
rect 1748 13252 1749 13292
rect 1707 13243 1749 13252
rect 1708 13158 1748 13243
rect 1707 12452 1749 12461
rect 1707 12412 1708 12452
rect 1748 12412 1749 12452
rect 1707 12403 1749 12412
rect 1708 12318 1748 12403
rect 1707 11780 1749 11789
rect 1707 11740 1708 11780
rect 1748 11740 1749 11780
rect 1707 11731 1749 11740
rect 1708 11646 1748 11731
rect 884 7876 1364 7916
rect 1420 11320 1652 11360
rect 844 7867 884 7876
rect 939 7748 981 7757
rect 939 7708 940 7748
rect 980 7708 981 7748
rect 939 7699 981 7708
rect 844 7244 884 7253
rect 748 7204 844 7244
rect 844 7195 884 7204
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 843 5732 885 5741
rect 843 5692 844 5732
rect 884 5692 885 5732
rect 843 5683 885 5692
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 844 5598 884 5683
rect 652 5431 692 5440
rect 844 4892 884 4901
rect 940 4892 980 7699
rect 884 4852 980 4892
rect 844 4843 884 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4674 692 4759
rect 1420 4229 1460 11320
rect 1515 10352 1557 10361
rect 1515 10312 1516 10352
rect 1556 10312 1557 10352
rect 1515 10303 1557 10312
rect 1516 10218 1556 10303
rect 1707 10268 1749 10277
rect 1707 10228 1708 10268
rect 1748 10228 1749 10268
rect 1707 10219 1749 10228
rect 1708 10134 1748 10219
rect 1804 7220 1844 17260
rect 2667 16988 2709 16997
rect 2667 16948 2668 16988
rect 2708 16948 2709 16988
rect 2667 16939 2709 16948
rect 2668 16854 2708 16939
rect 1612 7180 1844 7220
rect 2476 16820 2516 16829
rect 1612 5741 1652 7180
rect 1611 5732 1653 5741
rect 1611 5692 1612 5732
rect 1652 5692 1653 5732
rect 1611 5683 1653 5692
rect 843 4220 885 4229
rect 843 4180 844 4220
rect 884 4180 885 4220
rect 843 4171 885 4180
rect 1419 4220 1461 4229
rect 1419 4180 1420 4220
rect 1460 4180 1461 4220
rect 1419 4171 1461 4180
rect 844 4086 884 4171
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 2476 3389 2516 16780
rect 2860 15485 2900 20803
rect 3148 20768 3188 20777
rect 2956 20600 2996 20609
rect 3148 20600 3188 20728
rect 3244 20768 3284 20803
rect 3244 20717 3284 20728
rect 3340 20768 3380 20887
rect 3340 20719 3380 20728
rect 3532 20684 3572 20971
rect 3628 20852 3668 22987
rect 7948 22280 7988 22289
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3628 20803 3668 20812
rect 3724 21608 3764 21617
rect 3532 20644 3668 20684
rect 2996 20560 3188 20600
rect 2956 20551 2996 20560
rect 3148 20432 3188 20560
rect 3436 20600 3476 20609
rect 3476 20560 3572 20600
rect 3436 20551 3476 20560
rect 3148 20392 3476 20432
rect 3340 20268 3380 20277
rect 2956 20228 3340 20264
rect 2956 20224 3380 20228
rect 2956 19508 2996 20224
rect 3340 20219 3380 20224
rect 3148 20096 3188 20105
rect 3148 19844 3188 20056
rect 3436 20096 3476 20392
rect 3436 19928 3476 20056
rect 3532 20096 3572 20560
rect 3532 20047 3572 20056
rect 3628 20012 3668 20644
rect 3724 20525 3764 21568
rect 3820 21608 3860 21617
rect 3820 21197 3860 21568
rect 3915 21608 3957 21617
rect 3915 21568 3916 21608
rect 3956 21568 3957 21608
rect 3915 21559 3957 21568
rect 4012 21608 4052 21619
rect 3916 21474 3956 21559
rect 4012 21533 4052 21568
rect 4492 21608 4532 21619
rect 7948 21617 7988 22240
rect 4492 21533 4532 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 4684 21608 4724 21617
rect 4011 21524 4053 21533
rect 4011 21484 4012 21524
rect 4052 21484 4053 21524
rect 4011 21475 4053 21484
rect 4491 21524 4533 21533
rect 4491 21484 4492 21524
rect 4532 21484 4533 21524
rect 4491 21475 4533 21484
rect 3819 21188 3861 21197
rect 3819 21148 3820 21188
rect 3860 21148 3861 21188
rect 3819 21139 3861 21148
rect 3915 21020 3957 21029
rect 3915 20980 3916 21020
rect 3956 20980 3957 21020
rect 3915 20971 3957 20980
rect 3820 20936 3860 20945
rect 3820 20852 3860 20896
rect 3916 20852 3956 20971
rect 4012 20945 4052 21475
rect 4588 21474 4628 21559
rect 4107 21356 4149 21365
rect 4107 21316 4108 21356
rect 4148 21316 4149 21356
rect 4107 21307 4149 21316
rect 4011 20936 4053 20945
rect 4011 20896 4012 20936
rect 4052 20896 4053 20936
rect 4011 20887 4053 20896
rect 3820 20812 3956 20852
rect 4012 20684 4052 20693
rect 4012 20525 4052 20644
rect 3723 20516 3765 20525
rect 3723 20476 3724 20516
rect 3764 20476 3765 20516
rect 3723 20467 3765 20476
rect 4011 20516 4053 20525
rect 4011 20476 4012 20516
rect 4052 20476 4053 20516
rect 4011 20467 4053 20476
rect 4011 20180 4053 20189
rect 4011 20140 4012 20180
rect 4052 20140 4053 20180
rect 4011 20131 4053 20140
rect 4012 20096 4052 20131
rect 4012 20045 4052 20056
rect 3628 19972 3860 20012
rect 3436 19888 3668 19928
rect 3148 19804 3572 19844
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3052 19508 3092 19517
rect 3339 19508 3381 19517
rect 3532 19508 3572 19804
rect 3628 19685 3668 19888
rect 3627 19676 3669 19685
rect 3627 19636 3628 19676
rect 3668 19636 3669 19676
rect 3627 19627 3669 19636
rect 3724 19601 3764 19972
rect 3820 19928 3860 19972
rect 3820 19879 3860 19888
rect 4012 19844 4052 19853
rect 3916 19804 4012 19844
rect 3723 19592 3765 19601
rect 3723 19552 3724 19592
rect 3764 19552 3765 19592
rect 3723 19543 3765 19552
rect 2956 19468 3052 19508
rect 3092 19468 3284 19508
rect 3052 19459 3092 19468
rect 2955 19340 2997 19349
rect 2955 19300 2956 19340
rect 2996 19300 2997 19340
rect 2955 19291 2997 19300
rect 2956 19256 2996 19291
rect 2956 19205 2996 19216
rect 3244 19256 3284 19468
rect 3339 19468 3340 19508
rect 3380 19468 3381 19508
rect 3339 19459 3381 19468
rect 3436 19468 3572 19508
rect 3340 19340 3380 19459
rect 3436 19424 3476 19468
rect 3916 19424 3956 19804
rect 4012 19795 4052 19804
rect 3436 19375 3476 19384
rect 3532 19384 3956 19424
rect 3340 19291 3380 19300
rect 3532 19340 3572 19384
rect 3532 19291 3572 19300
rect 4108 19340 4148 21307
rect 4203 21020 4245 21029
rect 4203 20980 4204 21020
rect 4244 20980 4245 21020
rect 4203 20971 4245 20980
rect 4204 20273 4244 20971
rect 4396 20768 4436 20779
rect 4396 20693 4436 20728
rect 4395 20684 4437 20693
rect 4395 20644 4396 20684
rect 4436 20644 4437 20684
rect 4395 20635 4437 20644
rect 4684 20600 4724 21568
rect 4780 21608 4820 21617
rect 4972 21608 5012 21617
rect 4820 21568 4972 21608
rect 4780 21559 4820 21568
rect 4972 21559 5012 21568
rect 5356 21608 5396 21617
rect 5067 21524 5109 21533
rect 5067 21484 5068 21524
rect 5108 21484 5109 21524
rect 5067 21475 5109 21484
rect 4684 20560 5012 20600
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4203 20264 4245 20273
rect 4203 20224 4204 20264
rect 4244 20224 4245 20264
rect 4203 20215 4245 20224
rect 4683 20264 4725 20273
rect 4683 20224 4684 20264
rect 4724 20224 4725 20264
rect 4683 20215 4725 20224
rect 4491 20180 4533 20189
rect 4491 20140 4492 20180
rect 4532 20140 4533 20180
rect 4491 20131 4533 20140
rect 4204 20096 4244 20105
rect 4204 19424 4244 20056
rect 4299 20096 4341 20105
rect 4299 20056 4300 20096
rect 4340 20056 4341 20096
rect 4299 20047 4341 20056
rect 4300 19962 4340 20047
rect 4492 19844 4532 20131
rect 4684 20012 4724 20215
rect 4684 19937 4724 19972
rect 4683 19928 4725 19937
rect 4683 19888 4684 19928
rect 4724 19888 4725 19928
rect 4683 19879 4725 19888
rect 4492 19601 4532 19804
rect 4491 19592 4533 19601
rect 4491 19552 4492 19592
rect 4532 19552 4533 19592
rect 4491 19543 4533 19552
rect 4204 19384 4436 19424
rect 4108 19291 4148 19300
rect 3244 19207 3284 19216
rect 3627 19256 3669 19265
rect 3627 19216 3628 19256
rect 3668 19216 3669 19256
rect 4396 19256 4436 19384
rect 4492 19265 4532 19543
rect 4588 19424 4628 19433
rect 4972 19424 5012 20560
rect 5068 19853 5108 21475
rect 5356 21281 5396 21568
rect 6220 21608 6260 21617
rect 5931 21440 5973 21449
rect 5931 21400 5932 21440
rect 5972 21400 5973 21440
rect 5931 21391 5973 21400
rect 5355 21272 5397 21281
rect 5355 21232 5356 21272
rect 5396 21232 5397 21272
rect 5355 21223 5397 21232
rect 5259 20768 5301 20777
rect 5259 20728 5260 20768
rect 5300 20728 5301 20768
rect 5259 20719 5301 20728
rect 5260 20634 5300 20719
rect 5356 20693 5396 21223
rect 5355 20684 5397 20693
rect 5355 20644 5356 20684
rect 5396 20644 5397 20684
rect 5355 20635 5397 20644
rect 5932 20609 5972 21391
rect 6220 20768 6260 21568
rect 7371 21608 7413 21617
rect 7371 21568 7372 21608
rect 7412 21568 7413 21608
rect 7371 21559 7413 21568
rect 7659 21608 7701 21617
rect 7659 21568 7660 21608
rect 7700 21568 7701 21608
rect 7659 21559 7701 21568
rect 7756 21608 7796 21617
rect 7947 21608 7989 21617
rect 7796 21568 7892 21608
rect 7756 21559 7796 21568
rect 7372 21524 7412 21559
rect 7372 21473 7412 21484
rect 7660 21104 7700 21559
rect 7660 21064 7796 21104
rect 6795 20936 6837 20945
rect 6795 20896 6796 20936
rect 6836 20896 6837 20936
rect 6795 20887 6837 20896
rect 7659 20936 7701 20945
rect 7659 20896 7660 20936
rect 7700 20896 7701 20936
rect 7659 20887 7701 20896
rect 6411 20852 6453 20861
rect 6411 20812 6412 20852
rect 6452 20812 6453 20852
rect 6411 20803 6453 20812
rect 6700 20852 6740 20861
rect 6315 20768 6357 20777
rect 6220 20728 6316 20768
rect 6356 20728 6357 20768
rect 6315 20719 6357 20728
rect 5931 20600 5973 20609
rect 5931 20560 5932 20600
rect 5972 20560 5973 20600
rect 5931 20551 5973 20560
rect 5259 20096 5301 20105
rect 5259 20056 5260 20096
rect 5300 20056 5301 20096
rect 5259 20047 5301 20056
rect 5260 20012 5300 20047
rect 5260 19961 5300 19972
rect 5067 19844 5109 19853
rect 5067 19804 5068 19844
rect 5108 19804 5109 19844
rect 5067 19795 5109 19804
rect 5355 19592 5397 19601
rect 5355 19552 5356 19592
rect 5396 19552 5397 19592
rect 5355 19543 5397 19552
rect 4628 19384 4916 19424
rect 4972 19384 5108 19424
rect 4588 19375 4628 19384
rect 3627 19207 3669 19216
rect 4290 19241 4330 19250
rect 3628 19122 3668 19207
rect 4290 19181 4330 19201
rect 4290 19172 4341 19181
rect 4204 19132 4300 19172
rect 4340 19132 4341 19172
rect 3916 19088 3956 19097
rect 3956 19048 4052 19088
rect 3916 19039 3956 19048
rect 3916 18756 3956 18765
rect 3531 18668 3573 18677
rect 3531 18628 3532 18668
rect 3572 18628 3573 18668
rect 3531 18619 3573 18628
rect 3435 18584 3477 18593
rect 3435 18544 3436 18584
rect 3476 18544 3477 18584
rect 3435 18535 3477 18544
rect 3532 18584 3572 18619
rect 3436 18450 3476 18535
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3532 17921 3572 18544
rect 3628 18584 3668 18593
rect 3628 18341 3668 18544
rect 3724 18584 3764 18593
rect 3724 18425 3764 18544
rect 3916 18509 3956 18716
rect 4012 18584 4052 19048
rect 3915 18500 3957 18509
rect 3915 18460 3916 18500
rect 3956 18460 3957 18500
rect 3915 18451 3957 18460
rect 3723 18416 3765 18425
rect 3723 18376 3724 18416
rect 3764 18376 3765 18416
rect 3723 18367 3765 18376
rect 3627 18332 3669 18341
rect 3627 18292 3628 18332
rect 3668 18292 3669 18332
rect 3627 18283 3669 18292
rect 3531 17912 3573 17921
rect 3531 17872 3532 17912
rect 3572 17872 3573 17912
rect 3531 17863 3573 17872
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 2859 15476 2901 15485
rect 2859 15436 2860 15476
rect 2900 15436 2901 15476
rect 2859 15427 2901 15436
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3628 10277 3668 18283
rect 3820 17996 3860 18005
rect 3916 17996 3956 18451
rect 4012 18425 4052 18544
rect 4107 18584 4149 18593
rect 4107 18544 4108 18584
rect 4148 18544 4149 18584
rect 4107 18535 4149 18544
rect 4108 18450 4148 18535
rect 4011 18416 4053 18425
rect 4011 18376 4012 18416
rect 4052 18376 4053 18416
rect 4011 18367 4053 18376
rect 4012 18164 4052 18367
rect 4012 18124 4148 18164
rect 3860 17956 3956 17996
rect 3820 17947 3860 17956
rect 4012 17828 4052 17837
rect 3724 17788 4012 17828
rect 3724 17744 3764 17788
rect 3724 17695 3764 17704
rect 4012 16997 4052 17788
rect 4108 17669 4148 18124
rect 4204 17837 4244 19132
rect 4290 19123 4341 19132
rect 4290 19018 4330 19123
rect 4396 19097 4436 19216
rect 4491 19256 4533 19265
rect 4491 19216 4492 19256
rect 4532 19216 4533 19256
rect 4491 19207 4533 19216
rect 4588 19256 4628 19265
rect 4683 19256 4725 19265
rect 4628 19216 4684 19256
rect 4724 19216 4725 19256
rect 4588 19207 4628 19216
rect 4683 19207 4725 19216
rect 4395 19088 4437 19097
rect 4395 19048 4396 19088
rect 4436 19048 4437 19088
rect 4395 19039 4437 19048
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4588 18584 4628 18595
rect 4588 18509 4628 18544
rect 4683 18584 4725 18593
rect 4683 18544 4684 18584
rect 4724 18544 4725 18584
rect 4683 18535 4725 18544
rect 4587 18500 4629 18509
rect 4587 18460 4588 18500
rect 4628 18460 4629 18500
rect 4587 18451 4629 18460
rect 4684 18500 4724 18535
rect 4396 18332 4436 18341
rect 4684 18332 4724 18460
rect 4876 18500 4916 19384
rect 4971 19256 5013 19265
rect 4971 19216 4972 19256
rect 5012 19216 5013 19256
rect 4971 19207 5013 19216
rect 4876 18451 4916 18460
rect 4972 18584 5012 19207
rect 5068 18593 5108 19384
rect 4779 18416 4821 18425
rect 4779 18376 4780 18416
rect 4820 18376 4821 18416
rect 4779 18367 4821 18376
rect 4436 18292 4724 18332
rect 4396 18283 4436 18292
rect 4780 18282 4820 18367
rect 4972 18332 5012 18544
rect 5067 18584 5109 18593
rect 5067 18544 5068 18584
rect 5108 18544 5109 18584
rect 5067 18535 5109 18544
rect 5356 18500 5396 19543
rect 5932 19340 5972 20551
rect 6219 20096 6261 20105
rect 6219 20056 6220 20096
rect 6260 20056 6261 20096
rect 6316 20096 6356 20719
rect 6412 20357 6452 20803
rect 6604 20768 6644 20777
rect 6508 20728 6604 20768
rect 6411 20348 6453 20357
rect 6411 20308 6412 20348
rect 6452 20308 6453 20348
rect 6411 20299 6453 20308
rect 6412 20096 6452 20105
rect 6316 20056 6412 20096
rect 6219 20047 6261 20056
rect 6412 20047 6452 20056
rect 5932 19291 5972 19300
rect 6220 19256 6260 20047
rect 6412 19508 6452 19517
rect 6508 19508 6548 20728
rect 6604 20719 6644 20728
rect 6700 20105 6740 20812
rect 6796 20802 6836 20887
rect 6891 20852 6933 20861
rect 6891 20812 6892 20852
rect 6932 20812 6933 20852
rect 6891 20803 6933 20812
rect 7371 20852 7413 20861
rect 7371 20812 7372 20852
rect 7412 20812 7413 20852
rect 7371 20803 7413 20812
rect 6892 20718 6932 20803
rect 6988 20768 7028 20777
rect 6988 20264 7028 20728
rect 6796 20224 7028 20264
rect 6699 20096 6741 20105
rect 6699 20056 6700 20096
rect 6740 20056 6741 20096
rect 6699 20047 6741 20056
rect 6699 19676 6741 19685
rect 6699 19636 6700 19676
rect 6740 19636 6741 19676
rect 6699 19627 6741 19636
rect 6452 19468 6644 19508
rect 6412 19459 6452 19468
rect 6316 19256 6356 19265
rect 6220 19216 6316 19256
rect 6316 19207 6356 19216
rect 5356 18451 5396 18460
rect 5740 19088 5780 19097
rect 5164 18332 5204 18341
rect 4972 18292 5164 18332
rect 5204 18292 5300 18332
rect 5164 18283 5204 18292
rect 5067 17912 5109 17921
rect 5067 17872 5068 17912
rect 5108 17872 5109 17912
rect 5067 17863 5109 17872
rect 4203 17828 4245 17837
rect 4203 17788 4204 17828
rect 4244 17788 4245 17828
rect 4203 17779 4245 17788
rect 4107 17660 4149 17669
rect 4107 17620 4108 17660
rect 4148 17620 4149 17660
rect 4107 17611 4149 17620
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 5068 17333 5108 17863
rect 5163 17744 5205 17753
rect 5163 17704 5164 17744
rect 5204 17704 5205 17744
rect 5163 17695 5205 17704
rect 5164 17610 5204 17695
rect 5067 17324 5109 17333
rect 5067 17284 5068 17324
rect 5108 17284 5109 17324
rect 5067 17275 5109 17284
rect 4011 16988 4053 16997
rect 4011 16948 4012 16988
rect 4052 16948 4053 16988
rect 4011 16939 4053 16948
rect 4012 16241 4052 16939
rect 4011 16232 4053 16241
rect 4011 16192 4012 16232
rect 4052 16192 4053 16232
rect 4011 16183 4053 16192
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 3627 10268 3669 10277
rect 3627 10228 3628 10268
rect 3668 10228 3669 10268
rect 3627 10219 3669 10228
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 5068 3464 5108 17275
rect 5260 17081 5300 18292
rect 5740 18080 5780 19048
rect 6507 19088 6549 19097
rect 6507 19048 6508 19088
rect 6548 19048 6549 19088
rect 6507 19039 6549 19048
rect 6604 19084 6644 19468
rect 6700 19256 6740 19627
rect 6796 19601 6836 20224
rect 6891 20096 6933 20105
rect 7276 20096 7316 20105
rect 6891 20056 6892 20096
rect 6932 20056 6933 20096
rect 6891 20047 6933 20056
rect 6988 20056 7276 20096
rect 6795 19592 6837 19601
rect 6795 19552 6796 19592
rect 6836 19552 6837 19592
rect 6795 19543 6837 19552
rect 6892 19517 6932 20047
rect 6891 19508 6933 19517
rect 6891 19468 6892 19508
rect 6932 19468 6933 19508
rect 6891 19459 6933 19468
rect 6700 19207 6740 19216
rect 6795 19256 6837 19265
rect 6795 19216 6796 19256
rect 6836 19216 6837 19256
rect 6795 19207 6837 19216
rect 6796 19122 6836 19207
rect 6219 18500 6261 18509
rect 6219 18460 6220 18500
rect 6260 18460 6261 18500
rect 6219 18451 6261 18460
rect 5740 18040 6068 18080
rect 6028 17744 6068 18040
rect 6028 17417 6068 17704
rect 6123 17660 6165 17669
rect 6123 17620 6124 17660
rect 6164 17620 6165 17660
rect 6123 17611 6165 17620
rect 6027 17408 6069 17417
rect 6027 17368 6028 17408
rect 6068 17368 6069 17408
rect 6027 17359 6069 17368
rect 6124 17300 6164 17611
rect 6220 17333 6260 18451
rect 6411 18416 6453 18425
rect 6411 18376 6412 18416
rect 6452 18376 6453 18416
rect 6411 18367 6453 18376
rect 6508 18416 6548 19039
rect 6604 19035 6644 19044
rect 6796 18500 6836 18509
rect 6604 18416 6644 18425
rect 6508 18376 6604 18416
rect 6412 17744 6452 18367
rect 6412 17695 6452 17704
rect 6028 17260 6164 17300
rect 6219 17324 6261 17333
rect 6219 17284 6220 17324
rect 6260 17284 6261 17324
rect 6508 17300 6548 18376
rect 6604 18367 6644 18376
rect 6796 18257 6836 18460
rect 6988 18425 7028 20056
rect 7276 20047 7316 20056
rect 7083 19508 7125 19517
rect 7083 19468 7084 19508
rect 7124 19468 7125 19508
rect 7083 19459 7125 19468
rect 7276 19508 7316 19517
rect 7372 19508 7412 20803
rect 7467 20768 7509 20777
rect 7467 20728 7468 20768
rect 7508 20728 7509 20768
rect 7467 20719 7509 20728
rect 7468 20634 7508 20719
rect 7563 20180 7605 20189
rect 7563 20140 7564 20180
rect 7604 20140 7605 20180
rect 7563 20131 7605 20140
rect 7660 20180 7700 20887
rect 7660 20131 7700 20140
rect 7316 19468 7412 19508
rect 7276 19459 7316 19468
rect 7084 19374 7124 19459
rect 7275 19340 7317 19349
rect 7275 19300 7276 19340
rect 7316 19300 7317 19340
rect 7275 19291 7317 19300
rect 7276 19256 7316 19291
rect 7276 19205 7316 19216
rect 7468 19256 7508 19265
rect 7468 19097 7508 19216
rect 7564 19256 7604 20131
rect 7467 19088 7509 19097
rect 7467 19048 7468 19088
rect 7508 19048 7509 19088
rect 7467 19039 7509 19048
rect 7468 18761 7508 19039
rect 7564 19013 7604 19216
rect 7563 19004 7605 19013
rect 7563 18964 7564 19004
rect 7604 18964 7605 19004
rect 7563 18955 7605 18964
rect 7467 18752 7509 18761
rect 7467 18712 7468 18752
rect 7508 18712 7509 18752
rect 7756 18752 7796 21064
rect 7852 20180 7892 21568
rect 7947 21568 7948 21608
rect 7988 21568 7989 21608
rect 7947 21559 7989 21568
rect 8140 21608 8180 21617
rect 7948 21020 7988 21559
rect 8140 21449 8180 21568
rect 9003 21608 9045 21617
rect 9003 21568 9004 21608
rect 9044 21568 9045 21608
rect 9003 21559 9045 21568
rect 10539 21608 10581 21617
rect 10539 21568 10540 21608
rect 10580 21568 10581 21608
rect 10539 21559 10581 21568
rect 11212 21608 11252 21617
rect 9004 21474 9044 21559
rect 8139 21440 8181 21449
rect 8139 21400 8140 21440
rect 8180 21400 8181 21440
rect 8139 21391 8181 21400
rect 8140 21281 8180 21391
rect 10156 21356 10196 21365
rect 8139 21272 8181 21281
rect 8139 21232 8140 21272
rect 8180 21232 8181 21272
rect 8139 21223 8181 21232
rect 10156 21113 10196 21316
rect 10155 21104 10197 21113
rect 10155 21064 10156 21104
rect 10196 21064 10197 21104
rect 10155 21055 10197 21064
rect 7948 20971 7988 20980
rect 10251 20936 10293 20945
rect 10251 20896 10252 20936
rect 10292 20896 10293 20936
rect 10251 20887 10293 20896
rect 10155 20852 10197 20861
rect 10155 20812 10156 20852
rect 10196 20812 10197 20852
rect 10155 20803 10197 20812
rect 8427 20768 8469 20777
rect 8427 20728 8428 20768
rect 8468 20728 8469 20768
rect 8427 20719 8469 20728
rect 9772 20768 9812 20777
rect 8428 20634 8468 20719
rect 9292 20264 9332 20275
rect 9292 20189 9332 20224
rect 9772 20189 9812 20728
rect 10060 20768 10100 20777
rect 9868 20600 9908 20609
rect 10060 20600 10100 20728
rect 10156 20718 10196 20803
rect 10252 20802 10292 20887
rect 10348 20852 10388 20861
rect 9908 20560 10100 20600
rect 9868 20551 9908 20560
rect 7852 20131 7892 20140
rect 9291 20180 9333 20189
rect 9291 20140 9292 20180
rect 9332 20140 9333 20180
rect 9291 20131 9333 20140
rect 9771 20180 9813 20189
rect 9771 20140 9772 20180
rect 9812 20140 9813 20180
rect 10060 20180 10100 20560
rect 10251 20180 10293 20189
rect 10060 20140 10196 20180
rect 9771 20131 9813 20140
rect 7947 20096 7989 20105
rect 7947 20056 7948 20096
rect 7988 20056 7989 20096
rect 7947 20047 7989 20056
rect 8044 20096 8084 20105
rect 7948 19962 7988 20047
rect 8044 19013 8084 20056
rect 8140 20096 8180 20105
rect 8140 19853 8180 20056
rect 8332 20096 8372 20105
rect 8139 19844 8181 19853
rect 8139 19804 8140 19844
rect 8180 19804 8181 19844
rect 8139 19795 8181 19804
rect 8332 19265 8372 20056
rect 8428 20096 8468 20105
rect 8428 19853 8468 20056
rect 8523 20096 8565 20105
rect 8523 20056 8524 20096
rect 8564 20056 8565 20096
rect 8523 20047 8565 20056
rect 8620 20096 8660 20105
rect 8524 19962 8564 20047
rect 8427 19844 8469 19853
rect 8427 19804 8428 19844
rect 8468 19804 8469 19844
rect 8427 19795 8469 19804
rect 8620 19685 8660 20056
rect 9963 19844 10005 19853
rect 9963 19804 9964 19844
rect 10004 19804 10005 19844
rect 9963 19795 10005 19804
rect 8619 19676 8661 19685
rect 8619 19636 8620 19676
rect 8660 19636 8661 19676
rect 8619 19627 8661 19636
rect 9867 19676 9909 19685
rect 9867 19636 9868 19676
rect 9908 19636 9909 19676
rect 9867 19627 9909 19636
rect 9387 19508 9429 19517
rect 9387 19468 9388 19508
rect 9428 19468 9429 19508
rect 9387 19459 9429 19468
rect 9771 19508 9813 19517
rect 9771 19468 9772 19508
rect 9812 19468 9813 19508
rect 9771 19459 9813 19468
rect 8331 19256 8373 19265
rect 8331 19216 8332 19256
rect 8372 19216 8373 19256
rect 8331 19207 8373 19216
rect 8043 19004 8085 19013
rect 8043 18964 8044 19004
rect 8084 18964 8085 19004
rect 8043 18955 8085 18964
rect 7756 18712 7892 18752
rect 7467 18703 7509 18712
rect 7083 18668 7125 18677
rect 7083 18628 7084 18668
rect 7124 18628 7125 18668
rect 7083 18619 7125 18628
rect 7563 18668 7605 18677
rect 7563 18628 7564 18668
rect 7604 18628 7605 18668
rect 7563 18619 7605 18628
rect 6987 18416 7029 18425
rect 6987 18376 6988 18416
rect 7028 18376 7029 18416
rect 6987 18367 7029 18376
rect 6795 18248 6837 18257
rect 6795 18208 6796 18248
rect 6836 18208 6837 18248
rect 6795 18199 6837 18208
rect 7084 17996 7124 18619
rect 7276 18584 7316 18593
rect 7276 18332 7316 18544
rect 7371 18584 7413 18593
rect 7371 18544 7372 18584
rect 7412 18544 7413 18584
rect 7371 18535 7413 18544
rect 7468 18584 7508 18593
rect 7372 18450 7412 18535
rect 7468 18416 7508 18544
rect 7564 18584 7604 18619
rect 7564 18533 7604 18544
rect 7659 18584 7701 18593
rect 7659 18544 7660 18584
rect 7700 18544 7701 18584
rect 7659 18535 7701 18544
rect 7756 18584 7796 18593
rect 7660 18416 7700 18535
rect 7468 18376 7700 18416
rect 7756 18332 7796 18544
rect 7852 18341 7892 18712
rect 8140 18584 8180 18593
rect 8140 18425 8180 18544
rect 9004 18584 9044 18595
rect 9004 18509 9044 18544
rect 8331 18500 8373 18509
rect 8331 18460 8332 18500
rect 8372 18460 8373 18500
rect 8331 18451 8373 18460
rect 9003 18500 9045 18509
rect 9003 18460 9004 18500
rect 9044 18460 9045 18500
rect 9003 18451 9045 18460
rect 8139 18416 8181 18425
rect 8139 18376 8140 18416
rect 8180 18376 8181 18416
rect 8139 18367 8181 18376
rect 7276 18292 7796 18332
rect 7851 18332 7893 18341
rect 7851 18292 7852 18332
rect 7892 18292 7893 18332
rect 7851 18283 7893 18292
rect 7180 17996 7220 18005
rect 7084 17956 7180 17996
rect 6604 17788 6836 17828
rect 6604 17669 6644 17788
rect 6796 17744 6836 17788
rect 6796 17695 6836 17704
rect 6892 17744 6932 17753
rect 6932 17704 7028 17744
rect 6892 17695 6932 17704
rect 6603 17660 6645 17669
rect 6603 17620 6604 17660
rect 6644 17620 6645 17660
rect 6603 17611 6645 17620
rect 6700 17518 6740 17527
rect 6740 17478 6932 17492
rect 6700 17452 6932 17478
rect 6219 17275 6261 17284
rect 5259 17072 5301 17081
rect 5259 17032 5260 17072
rect 5300 17032 5301 17072
rect 5259 17023 5301 17032
rect 6028 17072 6068 17260
rect 6028 17023 6068 17032
rect 6124 17072 6164 17081
rect 6124 16997 6164 17032
rect 6220 17072 6260 17275
rect 6412 17260 6548 17300
rect 6795 17324 6837 17333
rect 6795 17284 6796 17324
rect 6836 17284 6837 17324
rect 6795 17275 6837 17284
rect 6315 17240 6357 17249
rect 6315 17200 6316 17240
rect 6356 17200 6357 17240
rect 6315 17191 6357 17200
rect 6316 17106 6356 17191
rect 6220 17023 6260 17032
rect 6123 16988 6165 16997
rect 6123 16948 6124 16988
rect 6164 16948 6165 16988
rect 6123 16939 6165 16948
rect 6124 11789 6164 16939
rect 6315 16232 6357 16241
rect 6315 16192 6316 16232
rect 6356 16192 6357 16232
rect 6315 16183 6357 16192
rect 6412 16232 6452 17260
rect 6507 17072 6549 17081
rect 6507 17032 6508 17072
rect 6548 17032 6549 17072
rect 6507 17023 6549 17032
rect 6699 17072 6741 17081
rect 6699 17032 6700 17072
rect 6740 17032 6741 17072
rect 6699 17023 6741 17032
rect 6508 16232 6548 17023
rect 6604 16988 6644 16997
rect 6604 16484 6644 16948
rect 6700 16904 6740 17023
rect 6796 16988 6836 17275
rect 6796 16939 6836 16948
rect 6892 17072 6932 17452
rect 6988 17249 7028 17704
rect 7084 17333 7124 17956
rect 7180 17928 7220 17956
rect 8140 17837 8180 18367
rect 7372 17828 7412 17837
rect 7083 17324 7125 17333
rect 7083 17284 7084 17324
rect 7124 17284 7125 17324
rect 7083 17275 7125 17284
rect 6987 17240 7029 17249
rect 6987 17200 6988 17240
rect 7028 17200 7029 17240
rect 6987 17191 7029 17200
rect 6700 16855 6740 16864
rect 6604 16435 6644 16444
rect 6892 16484 6932 17032
rect 7083 17072 7125 17081
rect 7083 17032 7084 17072
rect 7124 17032 7125 17072
rect 7083 17023 7125 17032
rect 7084 16938 7124 17023
rect 6892 16435 6932 16444
rect 6987 16316 7029 16325
rect 6987 16276 6988 16316
rect 7028 16276 7029 16316
rect 6987 16267 7029 16276
rect 6604 16232 6644 16241
rect 6508 16192 6604 16232
rect 6412 16183 6452 16192
rect 6604 16183 6644 16192
rect 6988 16232 7028 16267
rect 6316 16098 6356 16183
rect 6988 16181 7028 16192
rect 6123 11780 6165 11789
rect 6123 11740 6124 11780
rect 6164 11740 6165 11780
rect 6123 11731 6165 11740
rect 7372 3641 7412 17788
rect 8139 17828 8181 17837
rect 8139 17788 8140 17828
rect 8180 17788 8181 17828
rect 8139 17779 8181 17788
rect 7563 17576 7605 17585
rect 7563 17536 7564 17576
rect 7604 17536 7605 17576
rect 7563 17527 7605 17536
rect 7564 17442 7604 17527
rect 8140 17417 8180 17779
rect 8332 17753 8372 18451
rect 8331 17744 8373 17753
rect 8331 17704 8332 17744
rect 8372 17704 8373 17744
rect 8331 17695 8373 17704
rect 7467 17408 7509 17417
rect 7467 17368 7468 17408
rect 7508 17368 7509 17408
rect 7467 17359 7509 17368
rect 8139 17408 8181 17417
rect 8139 17368 8140 17408
rect 8180 17368 8181 17408
rect 8139 17359 8181 17368
rect 7468 17072 7508 17359
rect 7468 17023 7508 17032
rect 8332 17072 8372 17695
rect 8332 17023 8372 17032
rect 9388 13973 9428 19459
rect 9772 19256 9812 19459
rect 9772 19207 9812 19216
rect 9868 19256 9908 19627
rect 9868 19097 9908 19216
rect 9964 19256 10004 19795
rect 9964 19207 10004 19216
rect 10059 19256 10101 19265
rect 10059 19216 10060 19256
rect 10100 19216 10101 19256
rect 10156 19256 10196 20140
rect 10251 20140 10252 20180
rect 10292 20140 10293 20180
rect 10251 20131 10293 20140
rect 10252 19433 10292 20131
rect 10348 19592 10388 20812
rect 10444 20768 10484 20777
rect 10444 20273 10484 20728
rect 10443 20264 10485 20273
rect 10443 20224 10444 20264
rect 10484 20224 10485 20264
rect 10443 20215 10485 20224
rect 10444 20096 10484 20105
rect 10540 20096 10580 21559
rect 10635 21104 10677 21113
rect 10635 21064 10636 21104
rect 10676 21064 10677 21104
rect 10635 21055 10677 21064
rect 10636 20105 10676 21055
rect 11020 20861 11060 20892
rect 11019 20852 11061 20861
rect 11019 20812 11020 20852
rect 11060 20812 11061 20852
rect 11019 20803 11061 20812
rect 10828 20768 10868 20777
rect 10484 20056 10580 20096
rect 10635 20096 10677 20105
rect 10635 20056 10636 20096
rect 10676 20056 10677 20096
rect 10444 20047 10484 20056
rect 10635 20047 10677 20056
rect 10828 19853 10868 20728
rect 10924 20768 10964 20777
rect 10924 20609 10964 20728
rect 11020 20768 11060 20803
rect 10923 20600 10965 20609
rect 10923 20560 10924 20600
rect 10964 20560 10965 20600
rect 10923 20551 10965 20560
rect 10827 19844 10869 19853
rect 10827 19804 10828 19844
rect 10868 19804 10869 19844
rect 10827 19795 10869 19804
rect 10348 19552 10676 19592
rect 10251 19424 10293 19433
rect 10251 19384 10252 19424
rect 10292 19384 10293 19424
rect 10251 19375 10293 19384
rect 10636 19340 10676 19552
rect 10732 19508 10772 19517
rect 11020 19508 11060 20728
rect 11116 20768 11156 20777
rect 11212 20768 11252 21568
rect 11596 21608 11636 21617
rect 11596 21449 11636 21568
rect 12459 21608 12501 21617
rect 12459 21568 12460 21608
rect 12500 21568 12501 21608
rect 12459 21559 12501 21568
rect 12460 21474 12500 21559
rect 11595 21440 11637 21449
rect 11595 21400 11596 21440
rect 11636 21400 11637 21440
rect 11595 21391 11637 21400
rect 13612 21356 13652 21367
rect 13612 21281 13652 21316
rect 12939 21272 12981 21281
rect 12939 21232 12940 21272
rect 12980 21232 12981 21272
rect 12939 21223 12981 21232
rect 13611 21272 13653 21281
rect 13611 21232 13612 21272
rect 13652 21232 13653 21272
rect 13611 21223 13653 21232
rect 11691 20936 11733 20945
rect 11691 20896 11692 20936
rect 11732 20896 11733 20936
rect 11691 20887 11733 20896
rect 11156 20728 11252 20768
rect 11116 20719 11156 20728
rect 11692 20180 11732 20887
rect 11692 20131 11732 20140
rect 12075 20180 12117 20189
rect 12075 20140 12076 20180
rect 12116 20140 12117 20180
rect 12075 20131 12117 20140
rect 11308 20096 11348 20105
rect 11115 19592 11157 19601
rect 11115 19552 11116 19592
rect 11156 19552 11157 19592
rect 11115 19543 11157 19552
rect 10772 19468 11060 19508
rect 10732 19459 10772 19468
rect 10828 19384 11060 19424
rect 10828 19340 10868 19384
rect 10636 19300 10868 19340
rect 10348 19256 10388 19265
rect 10156 19216 10348 19256
rect 10059 19207 10101 19216
rect 10348 19207 10388 19216
rect 10443 19256 10485 19265
rect 10443 19216 10444 19256
rect 10484 19216 10485 19256
rect 10443 19207 10485 19216
rect 10924 19256 10964 19265
rect 10060 19122 10100 19207
rect 10444 19122 10484 19207
rect 9867 19088 9909 19097
rect 9867 19048 9868 19088
rect 9908 19048 9909 19088
rect 9867 19039 9909 19048
rect 10251 19088 10293 19097
rect 10251 19044 10252 19088
rect 10292 19044 10293 19088
rect 10251 19039 10293 19044
rect 10252 18953 10292 19039
rect 9771 18752 9813 18761
rect 9771 18712 9772 18752
rect 9812 18712 9813 18752
rect 10924 18752 10964 19216
rect 11020 19172 11060 19384
rect 11020 19123 11060 19132
rect 11116 19256 11156 19543
rect 11116 18761 11156 19216
rect 11212 19256 11252 19265
rect 11115 18752 11157 18761
rect 10924 18712 11060 18752
rect 9771 18703 9813 18712
rect 9772 17300 9812 18703
rect 10732 18677 10772 18708
rect 10731 18668 10773 18677
rect 10731 18628 10732 18668
rect 10772 18628 10773 18668
rect 10731 18619 10773 18628
rect 10636 18584 10676 18593
rect 10060 18544 10636 18584
rect 9963 17744 10005 17753
rect 9963 17704 9964 17744
rect 10004 17704 10005 17744
rect 9963 17695 10005 17704
rect 10060 17744 10100 18544
rect 10636 18535 10676 18544
rect 10732 18584 10772 18619
rect 10732 18425 10772 18544
rect 10828 18584 10868 18593
rect 10731 18416 10773 18425
rect 10731 18376 10732 18416
rect 10772 18376 10773 18416
rect 10731 18367 10773 18376
rect 10060 17695 10100 17704
rect 10156 18332 10196 18341
rect 9867 17660 9909 17669
rect 9867 17620 9868 17660
rect 9908 17620 9909 17660
rect 9867 17611 9909 17620
rect 9868 17572 9908 17611
rect 9964 17610 10004 17695
rect 9868 17523 9908 17532
rect 9772 17260 9908 17300
rect 9772 17072 9812 17081
rect 9484 16820 9524 16829
rect 9772 16820 9812 17032
rect 9868 17072 9908 17260
rect 10059 17156 10101 17165
rect 10059 17116 10060 17156
rect 10100 17116 10101 17156
rect 10059 17107 10101 17116
rect 9868 17023 9908 17032
rect 10060 17072 10100 17107
rect 10060 17021 10100 17032
rect 10156 16997 10196 18292
rect 10347 18332 10389 18341
rect 10347 18292 10348 18332
rect 10388 18292 10389 18332
rect 10347 18283 10389 18292
rect 10635 18332 10677 18341
rect 10635 18292 10636 18332
rect 10676 18292 10677 18332
rect 10635 18283 10677 18292
rect 10251 18080 10293 18089
rect 10251 18040 10252 18080
rect 10292 18040 10293 18080
rect 10251 18031 10293 18040
rect 10155 16988 10197 16997
rect 10155 16948 10156 16988
rect 10196 16948 10197 16988
rect 10155 16939 10197 16948
rect 10059 16904 10101 16913
rect 10059 16864 10060 16904
rect 10100 16864 10101 16904
rect 10059 16855 10101 16864
rect 9524 16780 9812 16820
rect 9484 16325 9524 16780
rect 10060 16770 10100 16855
rect 9483 16316 9525 16325
rect 9483 16276 9484 16316
rect 9524 16276 9525 16316
rect 9483 16267 9525 16276
rect 9387 13964 9429 13973
rect 9387 13924 9388 13964
rect 9428 13924 9429 13964
rect 9387 13915 9429 13924
rect 10252 12461 10292 18031
rect 10348 17996 10388 18283
rect 10348 17947 10388 17956
rect 10540 17660 10580 17669
rect 10347 17576 10389 17585
rect 10347 17536 10348 17576
rect 10388 17536 10389 17576
rect 10347 17527 10389 17536
rect 10348 17165 10388 17527
rect 10347 17156 10389 17165
rect 10347 17116 10348 17156
rect 10388 17116 10389 17156
rect 10347 17107 10389 17116
rect 10348 17072 10388 17107
rect 10348 17021 10388 17032
rect 10444 16988 10484 16999
rect 10444 16913 10484 16948
rect 10443 16904 10485 16913
rect 10443 16864 10444 16904
rect 10484 16864 10485 16904
rect 10443 16855 10485 16864
rect 10540 16904 10580 17620
rect 10636 16988 10676 18283
rect 10828 18089 10868 18544
rect 10923 18584 10965 18593
rect 10923 18544 10924 18584
rect 10964 18544 10965 18584
rect 10923 18535 10965 18544
rect 10827 18080 10869 18089
rect 10827 18040 10828 18080
rect 10868 18040 10869 18080
rect 10827 18031 10869 18040
rect 10924 17912 10964 18535
rect 10828 17872 10964 17912
rect 10731 17744 10773 17753
rect 10731 17704 10732 17744
rect 10772 17704 10773 17744
rect 10731 17695 10773 17704
rect 10732 17072 10772 17695
rect 10828 17669 10868 17872
rect 10923 17744 10965 17753
rect 10923 17704 10924 17744
rect 10964 17704 10965 17744
rect 10923 17695 10965 17704
rect 10827 17660 10869 17669
rect 10827 17620 10828 17660
rect 10868 17620 10869 17660
rect 10827 17611 10869 17620
rect 10924 17610 10964 17695
rect 11020 17585 11060 18712
rect 11115 18712 11116 18752
rect 11156 18712 11157 18752
rect 11115 18703 11157 18712
rect 11212 18005 11252 19216
rect 11211 17996 11253 18005
rect 11211 17956 11212 17996
rect 11252 17956 11253 17996
rect 11211 17947 11253 17956
rect 11308 17753 11348 20056
rect 11979 19256 12021 19265
rect 11979 19216 11980 19256
rect 12020 19216 12021 19256
rect 11979 19207 12021 19216
rect 11787 18584 11829 18593
rect 11787 18544 11788 18584
rect 11828 18544 11829 18584
rect 11787 18535 11829 18544
rect 11307 17744 11349 17753
rect 11307 17704 11308 17744
rect 11348 17704 11349 17744
rect 11307 17695 11349 17704
rect 11788 17744 11828 18535
rect 11788 17695 11828 17704
rect 11499 17660 11541 17669
rect 11499 17620 11500 17660
rect 11540 17620 11541 17660
rect 11499 17611 11541 17620
rect 11019 17576 11061 17585
rect 11019 17536 11020 17576
rect 11060 17536 11061 17576
rect 11019 17527 11061 17536
rect 10924 17072 10964 17081
rect 10772 17032 10924 17072
rect 10732 17023 10772 17032
rect 10924 17023 10964 17032
rect 11019 17072 11061 17081
rect 11019 17032 11020 17072
rect 11060 17032 11061 17072
rect 11019 17023 11061 17032
rect 10636 16939 10676 16948
rect 10540 16855 10580 16864
rect 11020 16325 11060 17023
rect 11500 16997 11540 17611
rect 11499 16988 11541 16997
rect 11499 16948 11500 16988
rect 11540 16948 11541 16988
rect 11499 16939 11541 16948
rect 10539 16316 10581 16325
rect 10539 16276 10540 16316
rect 10580 16276 10581 16316
rect 10539 16267 10581 16276
rect 11019 16316 11061 16325
rect 11019 16276 11020 16316
rect 11060 16276 11061 16316
rect 11019 16267 11061 16276
rect 10540 16182 10580 16267
rect 10347 16064 10389 16073
rect 10347 16024 10348 16064
rect 10388 16024 10389 16064
rect 10347 16015 10389 16024
rect 10348 15930 10388 16015
rect 11980 13301 12020 19207
rect 12076 18584 12116 20131
rect 12940 19517 12980 21223
rect 13611 21020 13653 21029
rect 13611 20980 13612 21020
rect 13652 20980 13653 21020
rect 13611 20971 13653 20980
rect 13516 20768 13556 20777
rect 13324 20728 13516 20768
rect 12939 19508 12981 19517
rect 12939 19468 12940 19508
rect 12980 19468 12981 19508
rect 12939 19459 12981 19468
rect 12363 19424 12405 19433
rect 12363 19384 12364 19424
rect 12404 19384 12405 19424
rect 13324 19424 13364 20728
rect 13516 20719 13556 20728
rect 13612 20768 13652 20971
rect 13708 20945 13748 23827
rect 28779 23792 28821 23801
rect 28779 23752 28780 23792
rect 28820 23752 28821 23792
rect 28779 23743 28821 23752
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 14283 21440 14325 21449
rect 14283 21400 14284 21440
rect 14324 21400 14325 21440
rect 14283 21391 14325 21400
rect 13707 20936 13749 20945
rect 13707 20896 13708 20936
rect 13748 20896 13749 20936
rect 13707 20887 13749 20896
rect 13612 20719 13652 20728
rect 13708 20768 13748 20887
rect 13708 20719 13748 20728
rect 14284 20768 14324 21391
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 16300 20852 16340 20861
rect 16108 20812 16300 20852
rect 15148 20768 15188 20777
rect 14284 20719 14324 20728
rect 14956 20728 15148 20768
rect 13900 20684 13940 20693
rect 13420 20600 13460 20609
rect 13900 20600 13940 20644
rect 13460 20560 13940 20600
rect 13420 20551 13460 20560
rect 13515 19592 13557 19601
rect 13515 19552 13516 19592
rect 13556 19552 13557 19592
rect 13515 19543 13557 19552
rect 13419 19424 13461 19433
rect 13324 19384 13420 19424
rect 13460 19384 13461 19424
rect 12363 19375 12405 19384
rect 13419 19375 13461 19384
rect 12076 18535 12116 18544
rect 12172 18500 12212 18509
rect 12172 18005 12212 18460
rect 12364 18500 12404 19375
rect 13420 19290 13460 19375
rect 12460 19256 12500 19265
rect 12460 18845 12500 19216
rect 12555 19256 12597 19265
rect 12555 19216 12556 19256
rect 12596 19216 12597 19256
rect 12555 19207 12597 19216
rect 12652 19256 12692 19265
rect 12556 19122 12596 19207
rect 12459 18836 12501 18845
rect 12459 18796 12460 18836
rect 12500 18796 12501 18836
rect 12459 18787 12501 18796
rect 12652 18752 12692 19216
rect 12747 19256 12789 19265
rect 12747 19216 12748 19256
rect 12788 19216 12789 19256
rect 12747 19207 12789 19216
rect 13036 19256 13076 19265
rect 12748 19122 12788 19207
rect 12940 19030 12980 19039
rect 12652 18712 12788 18752
rect 12459 18668 12501 18677
rect 12459 18628 12460 18668
rect 12500 18628 12501 18668
rect 12459 18619 12501 18628
rect 12460 18584 12500 18619
rect 12460 18533 12500 18544
rect 12652 18584 12692 18593
rect 12364 18451 12404 18460
rect 12268 18416 12308 18425
rect 12268 18332 12308 18376
rect 12652 18332 12692 18544
rect 12748 18425 12788 18712
rect 12940 18677 12980 18990
rect 13036 18845 13076 19216
rect 13131 19256 13173 19265
rect 13131 19216 13132 19256
rect 13172 19216 13173 19256
rect 13131 19207 13173 19216
rect 13132 19122 13172 19207
rect 13035 18836 13077 18845
rect 13035 18796 13036 18836
rect 13076 18796 13077 18836
rect 13035 18787 13077 18796
rect 12939 18668 12981 18677
rect 12939 18628 12940 18668
rect 12980 18628 12981 18668
rect 12939 18619 12981 18628
rect 13036 18584 13076 18593
rect 12747 18416 12789 18425
rect 12747 18376 12748 18416
rect 12788 18376 12789 18416
rect 12747 18367 12789 18376
rect 12268 18292 12692 18332
rect 13036 18257 13076 18544
rect 13035 18248 13077 18257
rect 13035 18208 13036 18248
rect 13076 18208 13077 18248
rect 13035 18199 13077 18208
rect 12171 17996 12213 18005
rect 12171 17956 12172 17996
rect 12212 17956 12213 17996
rect 12171 17947 12213 17956
rect 13036 17753 13076 18199
rect 13131 17996 13173 18005
rect 13131 17956 13132 17996
rect 13172 17956 13173 17996
rect 13131 17947 13173 17956
rect 13132 17862 13172 17947
rect 13035 17744 13077 17753
rect 13035 17704 13036 17744
rect 13076 17704 13077 17744
rect 13035 17695 13077 17704
rect 13132 17744 13172 17753
rect 13132 17585 13172 17704
rect 13324 17744 13364 17753
rect 12940 17576 12980 17585
rect 12940 17081 12980 17536
rect 13131 17576 13173 17585
rect 13131 17536 13132 17576
rect 13172 17536 13173 17576
rect 13131 17527 13173 17536
rect 13324 17081 13364 17704
rect 13420 17744 13460 17753
rect 13516 17744 13556 19543
rect 13611 18668 13653 18677
rect 13611 18628 13612 18668
rect 13652 18628 13653 18668
rect 13611 18619 13653 18628
rect 13612 17996 13652 18619
rect 14956 18593 14996 20728
rect 15148 20719 15188 20728
rect 16108 20525 16148 20812
rect 16300 20803 16340 20812
rect 28780 20777 28820 23743
rect 29740 21533 29780 29875
rect 31659 27908 31701 27917
rect 31659 27868 31660 27908
rect 31700 27868 31701 27908
rect 31659 27859 31701 27868
rect 31467 27572 31509 27581
rect 31467 27532 31468 27572
rect 31508 27532 31509 27572
rect 31467 27523 31509 27532
rect 31083 22532 31125 22541
rect 31083 22492 31084 22532
rect 31124 22492 31125 22532
rect 31083 22483 31125 22492
rect 31084 22398 31124 22483
rect 31276 22364 31316 22373
rect 31316 22324 31412 22364
rect 31276 22315 31316 22324
rect 30123 22280 30165 22289
rect 30123 22240 30124 22280
rect 30164 22240 30165 22280
rect 30123 22231 30165 22240
rect 29739 21524 29781 21533
rect 29739 21484 29740 21524
rect 29780 21484 29781 21524
rect 29739 21475 29781 21484
rect 30124 21524 30164 22231
rect 31084 22112 31124 22121
rect 30891 21692 30933 21701
rect 30891 21652 30892 21692
rect 30932 21652 30933 21692
rect 30891 21643 30933 21652
rect 30892 21558 30932 21643
rect 29740 21390 29780 21475
rect 30124 21449 30164 21484
rect 30507 21524 30549 21533
rect 30507 21484 30508 21524
rect 30548 21484 30549 21524
rect 30507 21475 30549 21484
rect 30123 21440 30165 21449
rect 30123 21400 30124 21440
rect 30164 21400 30165 21440
rect 30123 21391 30165 21400
rect 29931 21356 29973 21365
rect 29931 21316 29932 21356
rect 29972 21316 29973 21356
rect 29931 21307 29973 21316
rect 30316 21356 30356 21365
rect 29932 21222 29972 21307
rect 29644 20852 29684 20861
rect 27627 20768 27669 20777
rect 27627 20728 27628 20768
rect 27668 20728 27669 20768
rect 27627 20719 27669 20728
rect 28779 20768 28821 20777
rect 28779 20728 28780 20768
rect 28820 20728 28821 20768
rect 28779 20719 28821 20728
rect 16107 20516 16149 20525
rect 16107 20476 16108 20516
rect 16148 20476 16149 20516
rect 16107 20467 16149 20476
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 16108 19349 16148 20467
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 16971 20096 17013 20105
rect 16971 20056 16972 20096
rect 17012 20056 17013 20096
rect 16971 20047 17013 20056
rect 26955 20096 26997 20105
rect 26955 20056 26956 20096
rect 26996 20056 26997 20096
rect 26955 20047 26997 20056
rect 27628 20096 27668 20719
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 28491 20180 28533 20189
rect 28491 20140 28492 20180
rect 28532 20140 28533 20180
rect 28491 20131 28533 20140
rect 27628 20047 27668 20056
rect 27915 20096 27957 20105
rect 27915 20056 27916 20096
rect 27956 20056 27957 20096
rect 27915 20047 27957 20056
rect 16107 19340 16149 19349
rect 16107 19300 16108 19340
rect 16148 19300 16149 19340
rect 16107 19291 16149 19300
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 15339 18752 15381 18761
rect 15339 18712 15340 18752
rect 15380 18712 15381 18752
rect 15339 18703 15381 18712
rect 13899 18584 13941 18593
rect 13899 18544 13900 18584
rect 13940 18544 13941 18584
rect 13899 18535 13941 18544
rect 14955 18584 14997 18593
rect 14955 18544 14956 18584
rect 14996 18544 14997 18584
rect 14955 18535 14997 18544
rect 15244 18584 15284 18593
rect 13900 18450 13940 18535
rect 15244 18425 15284 18544
rect 15340 18584 15380 18703
rect 16972 18593 17012 20047
rect 26956 19962 26996 20047
rect 27916 19928 27956 20047
rect 28492 20046 28532 20131
rect 27916 19879 27956 19888
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 15340 18535 15380 18544
rect 15436 18584 15476 18593
rect 15243 18416 15285 18425
rect 15243 18376 15244 18416
rect 15284 18376 15285 18416
rect 15243 18367 15285 18376
rect 15436 18341 15476 18544
rect 15532 18584 15572 18593
rect 15724 18584 15764 18593
rect 15572 18544 15724 18584
rect 15532 18535 15572 18544
rect 15724 18535 15764 18544
rect 16108 18584 16148 18593
rect 15052 18332 15092 18341
rect 13612 17947 13652 17956
rect 14956 18292 15052 18332
rect 14956 17921 14996 18292
rect 15052 18283 15092 18292
rect 15435 18332 15477 18341
rect 15435 18292 15436 18332
rect 15476 18292 15477 18332
rect 15435 18283 15477 18292
rect 16108 18257 16148 18544
rect 16971 18584 17013 18593
rect 16971 18544 16972 18584
rect 17012 18544 17013 18584
rect 16971 18535 17013 18544
rect 27627 18584 27669 18593
rect 27627 18544 27628 18584
rect 27668 18544 27669 18584
rect 27627 18535 27669 18544
rect 16972 18450 17012 18535
rect 18123 18416 18165 18425
rect 18123 18376 18124 18416
rect 18164 18376 18165 18416
rect 18123 18367 18165 18376
rect 16107 18248 16149 18257
rect 16107 18208 16108 18248
rect 16148 18208 16149 18248
rect 16107 18199 16149 18208
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 18124 18089 18164 18367
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 18123 18080 18165 18089
rect 18123 18040 18124 18080
rect 18164 18040 18165 18080
rect 18123 18031 18165 18040
rect 13707 17912 13749 17921
rect 13707 17872 13708 17912
rect 13748 17872 13749 17912
rect 13707 17863 13749 17872
rect 14955 17912 14997 17921
rect 14955 17872 14956 17912
rect 14996 17872 14997 17912
rect 14955 17863 14997 17872
rect 13460 17704 13556 17744
rect 13708 17744 13748 17863
rect 13420 17695 13460 17704
rect 13708 17695 13748 17704
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 12939 17072 12981 17081
rect 12939 17032 12940 17072
rect 12980 17032 12981 17072
rect 12939 17023 12981 17032
rect 13323 17072 13365 17081
rect 13323 17032 13324 17072
rect 13364 17032 13365 17072
rect 13323 17023 13365 17032
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 27628 16484 27668 18535
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 28780 17249 28820 20719
rect 29452 20600 29492 20609
rect 28299 17240 28341 17249
rect 28299 17200 28300 17240
rect 28340 17200 28341 17240
rect 28299 17191 28341 17200
rect 28779 17240 28821 17249
rect 28779 17200 28780 17240
rect 28820 17200 28821 17240
rect 28779 17191 28821 17200
rect 29163 17240 29205 17249
rect 29163 17200 29164 17240
rect 29204 17200 29205 17240
rect 29163 17191 29205 17200
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 27628 15569 27668 16444
rect 28300 16232 28340 17191
rect 29164 17106 29204 17191
rect 28300 16183 28340 16192
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 27627 15560 27669 15569
rect 27627 15520 27628 15560
rect 27668 15520 27669 15560
rect 27627 15511 27669 15520
rect 27628 15426 27668 15511
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 11979 13292 12021 13301
rect 11979 13252 11980 13292
rect 12020 13252 12021 13292
rect 11979 13243 12021 13252
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 10251 12452 10293 12461
rect 10251 12412 10252 12452
rect 10292 12412 10293 12452
rect 10251 12403 10293 12412
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 29452 9437 29492 20560
rect 29644 20441 29684 20812
rect 30316 20693 30356 21316
rect 30411 21356 30453 21365
rect 30411 21316 30412 21356
rect 30452 21316 30453 21356
rect 30411 21307 30453 21316
rect 30315 20684 30357 20693
rect 30315 20644 30316 20684
rect 30356 20644 30357 20684
rect 30315 20635 30357 20644
rect 29836 20600 29876 20609
rect 29643 20432 29685 20441
rect 29643 20392 29644 20432
rect 29684 20392 29685 20432
rect 29643 20383 29685 20392
rect 29836 19181 29876 20560
rect 30316 20012 30356 20021
rect 30412 20012 30452 21307
rect 30508 20945 30548 21475
rect 30700 21356 30740 21365
rect 30740 21316 30836 21356
rect 30700 21307 30740 21316
rect 30507 20936 30549 20945
rect 30507 20896 30508 20936
rect 30548 20896 30549 20936
rect 30507 20887 30549 20896
rect 30507 20600 30549 20609
rect 30507 20560 30508 20600
rect 30548 20560 30549 20600
rect 30507 20551 30549 20560
rect 30508 20264 30548 20551
rect 30508 20215 30548 20224
rect 30699 20096 30741 20105
rect 30699 20056 30700 20096
rect 30740 20056 30741 20096
rect 30699 20047 30741 20056
rect 30796 20096 30836 21316
rect 30988 20768 31028 20777
rect 30891 20432 30933 20441
rect 30891 20392 30892 20432
rect 30932 20392 30933 20432
rect 30891 20383 30933 20392
rect 30356 19972 30644 20012
rect 30316 19963 30356 19972
rect 30604 19340 30644 19972
rect 30700 19962 30740 20047
rect 30796 19937 30836 20056
rect 30892 20096 30932 20383
rect 30988 20273 31028 20728
rect 31084 20432 31124 22072
rect 31275 21608 31317 21617
rect 31275 21568 31276 21608
rect 31316 21568 31317 21608
rect 31275 21559 31317 21568
rect 31276 21474 31316 21559
rect 31372 20693 31412 22324
rect 31468 22289 31508 27523
rect 31467 22280 31509 22289
rect 31467 22240 31468 22280
rect 31508 22240 31509 22280
rect 31467 22231 31509 22240
rect 31564 22280 31604 22289
rect 31468 22112 31508 22121
rect 31468 21701 31508 22072
rect 31467 21692 31509 21701
rect 31467 21652 31468 21692
rect 31508 21652 31509 21692
rect 31467 21643 31509 21652
rect 31564 21020 31604 22240
rect 31660 22280 31700 27859
rect 33195 27740 33237 27749
rect 33195 27700 33196 27740
rect 33236 27700 33237 27740
rect 33195 27691 33237 27700
rect 32043 23372 32085 23381
rect 32043 23332 32044 23372
rect 32084 23332 32085 23372
rect 32043 23323 32085 23332
rect 32044 22532 32084 23323
rect 32044 22483 32084 22492
rect 32235 22364 32277 22373
rect 32235 22324 32236 22364
rect 32276 22324 32277 22364
rect 32235 22315 32277 22324
rect 31660 22231 31700 22240
rect 31756 22280 31796 22289
rect 31756 21701 31796 22240
rect 32236 22230 32276 22315
rect 33196 22196 33236 27691
rect 36459 25304 36501 25313
rect 36459 25264 36460 25304
rect 36500 25264 36501 25304
rect 36459 25255 36501 25264
rect 34923 24632 34965 24641
rect 34923 24592 34924 24632
rect 34964 24592 34965 24632
rect 34923 24583 34965 24592
rect 36363 24632 36405 24641
rect 36363 24592 36364 24632
rect 36404 24592 36405 24632
rect 36363 24583 36405 24592
rect 33772 23288 33812 23297
rect 33772 23129 33812 23248
rect 33771 23120 33813 23129
rect 33771 23080 33772 23120
rect 33812 23080 33813 23120
rect 33771 23071 33813 23080
rect 34924 23120 34964 24583
rect 35211 24548 35253 24557
rect 35211 24508 35212 24548
rect 35252 24508 35253 24548
rect 35211 24499 35253 24508
rect 35212 24414 35252 24499
rect 36364 24498 36404 24583
rect 36460 24557 36500 25255
rect 36459 24548 36501 24557
rect 36459 24508 36460 24548
rect 36500 24508 36501 24548
rect 36459 24499 36501 24508
rect 36363 24212 36405 24221
rect 36363 24172 36364 24212
rect 36404 24172 36405 24212
rect 36363 24163 36405 24172
rect 36364 23792 36404 24163
rect 36172 23750 36212 23759
rect 35595 23708 35637 23717
rect 36364 23717 36404 23752
rect 36460 23792 36500 24499
rect 36652 24473 36692 36679
rect 56236 36678 56276 36763
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 55467 36224 55509 36233
rect 55467 36184 55468 36224
rect 55508 36184 55509 36224
rect 55467 36175 55509 36184
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 55083 35300 55125 35309
rect 55083 35260 55084 35300
rect 55124 35260 55125 35300
rect 55083 35251 55125 35260
rect 55084 35166 55124 35251
rect 55468 35216 55508 36175
rect 56428 36149 56468 36856
rect 56716 36821 56756 37234
rect 56715 36812 56757 36821
rect 56715 36772 56716 36812
rect 56756 36772 56757 36812
rect 56715 36763 56757 36772
rect 56523 36728 56565 36737
rect 56523 36688 56524 36728
rect 56564 36688 56565 36728
rect 56523 36679 56565 36688
rect 56620 36728 56660 36737
rect 56427 36140 56469 36149
rect 56427 36100 56428 36140
rect 56468 36100 56469 36140
rect 56427 36091 56469 36100
rect 56043 35972 56085 35981
rect 56043 35932 56044 35972
rect 56084 35932 56085 35972
rect 56043 35923 56085 35932
rect 56044 35888 56084 35923
rect 56044 35837 56084 35848
rect 56140 35888 56180 35897
rect 55948 35720 55988 35729
rect 55948 35309 55988 35680
rect 55947 35300 55989 35309
rect 55947 35260 55948 35300
rect 55988 35260 55989 35300
rect 55947 35251 55989 35260
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 51723 34544 51765 34553
rect 51723 34504 51724 34544
rect 51764 34504 51765 34544
rect 51723 34495 51765 34504
rect 52107 34544 52149 34553
rect 52107 34504 52108 34544
rect 52148 34504 52149 34544
rect 52107 34495 52149 34504
rect 50763 34376 50805 34385
rect 50763 34336 50764 34376
rect 50804 34336 50805 34376
rect 50763 34327 50805 34336
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 50475 33704 50517 33713
rect 50475 33664 50476 33704
rect 50516 33664 50517 33704
rect 50475 33655 50517 33664
rect 50476 33570 50516 33655
rect 49323 33452 49365 33461
rect 49323 33412 49324 33452
rect 49364 33412 49365 33452
rect 49323 33403 49365 33412
rect 50475 33452 50517 33461
rect 50475 33412 50476 33452
rect 50516 33412 50517 33452
rect 50475 33403 50517 33412
rect 49324 33318 49364 33403
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 49996 32948 50036 32957
rect 49900 32908 49996 32948
rect 49803 32696 49845 32705
rect 49803 32656 49804 32696
rect 49844 32656 49845 32696
rect 49803 32647 49845 32656
rect 49804 32562 49844 32647
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 48364 30808 48596 30848
rect 48076 30680 48116 30689
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 46635 30260 46677 30269
rect 46635 30220 46636 30260
rect 46676 30220 46677 30260
rect 46635 30211 46677 30220
rect 47979 30260 48021 30269
rect 48076 30260 48116 30640
rect 48172 30596 48212 30605
rect 48172 30269 48212 30556
rect 48364 30596 48404 30808
rect 48364 30547 48404 30556
rect 48460 30680 48500 30689
rect 48268 30512 48308 30521
rect 47979 30220 47980 30260
rect 48020 30220 48116 30260
rect 48171 30260 48213 30269
rect 48171 30220 48172 30260
rect 48212 30220 48213 30260
rect 47979 30211 48021 30220
rect 48171 30211 48213 30220
rect 40587 30008 40629 30017
rect 40587 29968 40588 30008
rect 40628 29968 40629 30008
rect 40587 29959 40629 29968
rect 40395 29924 40437 29933
rect 40395 29884 40396 29924
rect 40436 29884 40437 29924
rect 40395 29875 40437 29884
rect 40396 29790 40436 29875
rect 40588 29681 40628 29959
rect 46540 29840 46580 29849
rect 40587 29672 40629 29681
rect 40587 29632 40588 29672
rect 40628 29632 40629 29672
rect 40587 29623 40629 29632
rect 45388 29672 45428 29681
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 39915 29336 39957 29345
rect 39915 29296 39916 29336
rect 39956 29296 39957 29336
rect 39915 29287 39957 29296
rect 40683 29336 40725 29345
rect 40683 29296 40684 29336
rect 40724 29296 40725 29336
rect 40683 29287 40725 29296
rect 39916 29202 39956 29287
rect 39723 29084 39765 29093
rect 39723 29044 39724 29084
rect 39764 29044 39765 29084
rect 39723 29035 39765 29044
rect 40108 29084 40148 29093
rect 39724 28950 39764 29035
rect 40108 28925 40148 29044
rect 40684 29084 40724 29287
rect 45388 29177 45428 29632
rect 40684 29035 40724 29044
rect 42604 29168 42644 29177
rect 40107 28916 40149 28925
rect 40107 28876 40108 28916
rect 40148 28876 40149 28916
rect 40107 28867 40149 28876
rect 40300 28916 40340 28925
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 40300 28421 40340 28876
rect 40491 28916 40533 28925
rect 40491 28876 40492 28916
rect 40532 28876 40533 28916
rect 40491 28867 40533 28876
rect 41067 28916 41109 28925
rect 41067 28876 41068 28916
rect 41108 28876 41109 28916
rect 41067 28867 41109 28876
rect 40492 28782 40532 28867
rect 40299 28412 40341 28421
rect 40299 28372 40300 28412
rect 40340 28372 40341 28412
rect 40299 28363 40341 28372
rect 40779 28328 40821 28337
rect 40779 28288 40780 28328
rect 40820 28288 40821 28328
rect 40779 28279 40821 28288
rect 40780 28194 40820 28279
rect 39628 28160 39668 28169
rect 39628 27665 39668 28120
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 39627 27656 39669 27665
rect 40588 27656 40628 27665
rect 39627 27616 39628 27656
rect 39668 27616 39669 27656
rect 39627 27607 39669 27616
rect 40492 27616 40588 27656
rect 40396 27572 40436 27581
rect 40204 27404 40244 27413
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 40204 27161 40244 27364
rect 40203 27152 40245 27161
rect 40203 27112 40204 27152
rect 40244 27112 40245 27152
rect 40203 27103 40245 27112
rect 40396 27077 40436 27532
rect 40395 27068 40437 27077
rect 39340 27028 39956 27068
rect 38379 26984 38421 26993
rect 38379 26944 38380 26984
rect 38420 26944 38421 26984
rect 38379 26935 38421 26944
rect 38092 26144 38132 26153
rect 36939 25976 36981 25985
rect 36939 25936 36940 25976
rect 36980 25936 36981 25976
rect 36939 25927 36981 25936
rect 36940 25842 36980 25927
rect 37707 25304 37749 25313
rect 37707 25264 37708 25304
rect 37748 25264 37749 25304
rect 37707 25255 37749 25264
rect 37708 25170 37748 25255
rect 37803 25136 37845 25145
rect 37803 25096 37804 25136
rect 37844 25096 37845 25136
rect 37803 25087 37845 25096
rect 37804 24858 37844 25087
rect 37804 24809 37844 24818
rect 38092 24641 38132 26104
rect 38380 25304 38420 26935
rect 38667 26816 38709 26825
rect 38667 26776 38668 26816
rect 38708 26776 38709 26816
rect 38667 26767 38709 26776
rect 38668 25985 38708 26767
rect 39340 26228 39380 27028
rect 39916 26984 39956 27028
rect 40395 27028 40396 27068
rect 40436 27028 40437 27068
rect 40395 27019 40437 27028
rect 40492 26993 40532 27616
rect 40588 27607 40628 27616
rect 40780 27656 40820 27665
rect 40588 27404 40628 27413
rect 39916 26935 39956 26944
rect 40107 26984 40149 26993
rect 40107 26944 40108 26984
rect 40148 26944 40149 26984
rect 40107 26935 40149 26944
rect 40491 26984 40533 26993
rect 40491 26944 40492 26984
rect 40532 26944 40533 26984
rect 40491 26935 40533 26944
rect 39820 26900 39860 26909
rect 39435 26816 39477 26825
rect 39435 26776 39436 26816
rect 39476 26776 39477 26816
rect 39435 26767 39477 26776
rect 39532 26816 39572 26825
rect 39723 26816 39765 26825
rect 39572 26776 39724 26816
rect 39764 26776 39765 26816
rect 39532 26767 39572 26776
rect 39723 26767 39765 26776
rect 39436 26682 39476 26767
rect 39724 26682 39764 26767
rect 39820 26312 39860 26860
rect 40011 26900 40053 26909
rect 40011 26860 40012 26900
rect 40052 26860 40053 26900
rect 40011 26851 40053 26860
rect 40012 26766 40052 26851
rect 40108 26816 40148 26935
rect 40588 26909 40628 27364
rect 40780 27245 40820 27616
rect 40875 27656 40917 27665
rect 40875 27616 40876 27656
rect 40916 27616 40917 27656
rect 40875 27607 40917 27616
rect 40876 27522 40916 27607
rect 40779 27236 40821 27245
rect 40779 27196 40780 27236
rect 40820 27196 40821 27236
rect 40779 27187 40821 27196
rect 40780 26909 40820 26994
rect 40587 26900 40629 26909
rect 40587 26860 40588 26900
rect 40628 26860 40629 26900
rect 40587 26851 40629 26860
rect 40779 26900 40821 26909
rect 40779 26860 40780 26900
rect 40820 26860 40821 26900
rect 40779 26851 40821 26860
rect 40108 26767 40148 26776
rect 40203 26816 40245 26825
rect 40203 26776 40204 26816
rect 40244 26776 40245 26816
rect 40203 26767 40245 26776
rect 40300 26795 40340 26827
rect 40107 26648 40149 26657
rect 40107 26608 40108 26648
rect 40148 26608 40149 26648
rect 40107 26599 40149 26608
rect 39340 26179 39380 26188
rect 39724 26272 39860 26312
rect 38956 26144 38996 26153
rect 39532 26144 39572 26153
rect 38860 26104 38956 26144
rect 38667 25976 38709 25985
rect 38667 25936 38668 25976
rect 38708 25936 38709 25976
rect 38667 25927 38709 25936
rect 38380 25255 38420 25264
rect 38572 25304 38612 25313
rect 38187 25136 38229 25145
rect 38476 25136 38516 25145
rect 38187 25096 38188 25136
rect 38228 25096 38229 25136
rect 38187 25087 38229 25096
rect 38380 25096 38476 25136
rect 37228 24632 37268 24641
rect 36651 24464 36693 24473
rect 36651 24424 36652 24464
rect 36692 24424 36693 24464
rect 36651 24415 36693 24424
rect 37228 24305 37268 24592
rect 37612 24632 37652 24641
rect 37227 24296 37269 24305
rect 37227 24256 37228 24296
rect 37268 24256 37269 24296
rect 37227 24247 37269 24256
rect 37035 24128 37077 24137
rect 37035 24088 37036 24128
rect 37076 24088 37077 24128
rect 37035 24079 37077 24088
rect 36460 23743 36500 23752
rect 36748 23792 36788 23801
rect 36172 23708 36212 23710
rect 35595 23668 35596 23708
rect 35636 23668 35637 23708
rect 35595 23659 35637 23668
rect 35884 23668 36212 23708
rect 36363 23708 36405 23717
rect 36363 23668 36364 23708
rect 36404 23668 36405 23708
rect 35307 23204 35349 23213
rect 35307 23164 35308 23204
rect 35348 23164 35349 23204
rect 35307 23155 35349 23164
rect 34924 23071 34964 23080
rect 33292 22408 33620 22448
rect 33292 22364 33332 22408
rect 33292 22315 33332 22324
rect 33196 22156 33332 22196
rect 32044 22112 32084 22121
rect 31948 22072 32044 22112
rect 31755 21692 31797 21701
rect 31755 21652 31756 21692
rect 31796 21652 31797 21692
rect 31755 21643 31797 21652
rect 31756 21533 31796 21643
rect 31851 21608 31893 21617
rect 31851 21568 31852 21608
rect 31892 21568 31893 21608
rect 31851 21559 31893 21568
rect 31755 21524 31797 21533
rect 31755 21484 31756 21524
rect 31796 21484 31797 21524
rect 31755 21475 31797 21484
rect 31564 20980 31796 21020
rect 31659 20768 31701 20777
rect 31659 20728 31660 20768
rect 31700 20728 31701 20768
rect 31659 20719 31701 20728
rect 31371 20684 31413 20693
rect 31371 20644 31372 20684
rect 31412 20644 31413 20684
rect 31371 20635 31413 20644
rect 31084 20392 31604 20432
rect 30987 20264 31029 20273
rect 30987 20224 30988 20264
rect 31028 20224 31029 20264
rect 30987 20215 31029 20224
rect 30892 20047 30932 20056
rect 30988 20096 31028 20105
rect 31084 20096 31124 20392
rect 31179 20264 31221 20273
rect 31179 20224 31180 20264
rect 31220 20224 31221 20264
rect 31179 20215 31221 20224
rect 31028 20056 31124 20096
rect 30988 20047 31028 20056
rect 30795 19928 30837 19937
rect 30795 19888 30796 19928
rect 30836 19888 30837 19928
rect 30795 19879 30837 19888
rect 31180 19928 31220 20215
rect 31371 20180 31413 20189
rect 31371 20140 31372 20180
rect 31412 20140 31413 20180
rect 31371 20131 31413 20140
rect 31180 19879 31220 19888
rect 30700 19340 30740 19349
rect 30604 19300 30700 19340
rect 30700 19291 30740 19300
rect 29835 19172 29877 19181
rect 29835 19132 29836 19172
rect 29876 19132 29877 19172
rect 29835 19123 29877 19132
rect 30891 19088 30933 19097
rect 30891 19048 30892 19088
rect 30932 19048 30933 19088
rect 30891 19039 30933 19048
rect 30892 18954 30932 19039
rect 31372 18584 31412 20131
rect 31467 20096 31509 20105
rect 31467 20056 31468 20096
rect 31508 20056 31509 20096
rect 31467 20047 31509 20056
rect 31564 20096 31604 20392
rect 31564 20047 31604 20056
rect 31660 20322 31700 20719
rect 31468 19962 31508 20047
rect 31660 19508 31700 20282
rect 31756 20273 31796 20980
rect 31852 20768 31892 21559
rect 31852 20609 31892 20728
rect 31851 20600 31893 20609
rect 31851 20560 31852 20600
rect 31892 20560 31893 20600
rect 31851 20551 31893 20560
rect 31755 20264 31797 20273
rect 31755 20224 31756 20264
rect 31796 20224 31797 20264
rect 31755 20215 31797 20224
rect 31948 20012 31988 22072
rect 32044 22063 32084 22072
rect 33195 22028 33237 22037
rect 33195 21988 33196 22028
rect 33236 21988 33237 22028
rect 33195 21979 33237 21988
rect 32140 21608 32180 21617
rect 32140 20189 32180 21568
rect 33004 21020 33044 21029
rect 32236 20980 32660 21020
rect 32236 20768 32276 20980
rect 32620 20936 32660 20980
rect 32620 20887 32660 20896
rect 32716 20980 33004 21020
rect 32716 20894 32756 20980
rect 33004 20971 33044 20980
rect 32524 20852 32564 20861
rect 32716 20845 32756 20854
rect 32236 20719 32276 20728
rect 32427 20768 32469 20777
rect 32427 20728 32428 20768
rect 32468 20728 32469 20768
rect 32427 20719 32469 20728
rect 32428 20634 32468 20719
rect 32235 20600 32277 20609
rect 32235 20560 32236 20600
rect 32276 20560 32277 20600
rect 32235 20551 32277 20560
rect 32139 20180 32181 20189
rect 32139 20140 32140 20180
rect 32180 20140 32181 20180
rect 32139 20131 32181 20140
rect 31948 19963 31988 19972
rect 32140 19928 32180 19937
rect 32236 19928 32276 20551
rect 32524 20273 32564 20812
rect 33004 20777 33044 20862
rect 32811 20768 32853 20777
rect 32811 20728 32812 20768
rect 32852 20728 32853 20768
rect 32811 20719 32853 20728
rect 33003 20768 33045 20777
rect 33003 20728 33004 20768
rect 33044 20728 33045 20768
rect 33003 20719 33045 20728
rect 33196 20768 33236 21979
rect 33292 21356 33332 22156
rect 33484 22112 33524 22123
rect 33484 22037 33524 22072
rect 33483 22028 33525 22037
rect 33483 21988 33484 22028
rect 33524 21988 33525 22028
rect 33483 21979 33525 21988
rect 33484 21356 33524 21365
rect 33332 21316 33428 21356
rect 33292 21307 33332 21316
rect 33196 20719 33236 20728
rect 33291 20768 33333 20777
rect 33291 20728 33292 20768
rect 33332 20728 33333 20768
rect 33291 20719 33333 20728
rect 32812 20609 32852 20719
rect 33292 20634 33332 20719
rect 32811 20600 32853 20609
rect 32811 20560 32812 20600
rect 32852 20560 32853 20600
rect 32811 20551 32853 20560
rect 33388 20441 33428 21316
rect 33484 20777 33524 21316
rect 33483 20768 33525 20777
rect 33483 20728 33484 20768
rect 33524 20728 33525 20768
rect 33483 20719 33525 20728
rect 33387 20432 33429 20441
rect 33387 20392 33388 20432
rect 33428 20392 33429 20432
rect 33387 20383 33429 20392
rect 32523 20264 32565 20273
rect 32523 20224 32524 20264
rect 32564 20224 32565 20264
rect 32523 20215 32565 20224
rect 33580 20180 33620 22408
rect 33963 22364 34005 22373
rect 33963 22324 33964 22364
rect 34004 22324 34005 22364
rect 33963 22315 34005 22324
rect 33964 20861 34004 22315
rect 35308 21617 35348 23155
rect 35500 22280 35540 22291
rect 35596 22280 35636 23659
rect 35884 23381 35924 23668
rect 36363 23659 36405 23668
rect 36268 23624 36308 23633
rect 36364 23628 36404 23659
rect 36748 23633 36788 23752
rect 36844 23792 36884 23801
rect 36076 23584 36268 23624
rect 35883 23372 35925 23381
rect 35883 23332 35884 23372
rect 35924 23332 35925 23372
rect 35883 23323 35925 23332
rect 35787 23204 35829 23213
rect 35787 23164 35788 23204
rect 35828 23164 35829 23204
rect 35787 23155 35829 23164
rect 35691 23120 35733 23129
rect 35691 23080 35692 23120
rect 35732 23080 35733 23120
rect 35691 23071 35733 23080
rect 35788 23120 35828 23155
rect 35692 22700 35732 23071
rect 35788 23069 35828 23080
rect 35692 22660 35828 22700
rect 35692 22280 35732 22289
rect 35596 22240 35692 22280
rect 35500 22205 35540 22240
rect 35499 22196 35541 22205
rect 35404 22156 35500 22196
rect 35540 22156 35541 22196
rect 34636 21608 34676 21617
rect 33963 20852 34005 20861
rect 33963 20812 33964 20852
rect 34004 20812 34005 20852
rect 33963 20803 34005 20812
rect 33675 20600 33717 20609
rect 33675 20560 33676 20600
rect 33716 20560 33717 20600
rect 33675 20551 33717 20560
rect 33484 20140 33620 20180
rect 33196 20012 33236 20023
rect 33196 19937 33236 19972
rect 32180 19888 32276 19928
rect 33195 19928 33237 19937
rect 33195 19888 33196 19928
rect 33236 19888 33237 19928
rect 32140 19879 32180 19888
rect 33195 19879 33237 19888
rect 33004 19844 33044 19853
rect 31660 19459 31700 19468
rect 32524 19804 33004 19844
rect 32427 19340 32469 19349
rect 32427 19300 32428 19340
rect 32468 19300 32469 19340
rect 32427 19291 32469 19300
rect 31564 19256 31604 19267
rect 31564 19181 31604 19216
rect 32428 19206 32468 19291
rect 31563 19172 31605 19181
rect 31563 19132 31564 19172
rect 31604 19132 31605 19172
rect 31563 19123 31605 19132
rect 32235 19172 32277 19181
rect 32235 19132 32236 19172
rect 32276 19132 32277 19172
rect 32235 19123 32277 19132
rect 32236 18593 32276 19123
rect 31372 18535 31412 18544
rect 32235 18584 32277 18593
rect 32235 18544 32236 18584
rect 32276 18544 32277 18584
rect 32235 18535 32277 18544
rect 32236 18450 32276 18535
rect 30220 18332 30260 18341
rect 30220 17753 30260 18292
rect 32427 18248 32469 18257
rect 32427 18208 32428 18248
rect 32468 18208 32469 18248
rect 32427 18199 32469 18208
rect 31948 18005 31988 18090
rect 31947 17996 31989 18005
rect 31947 17956 31948 17996
rect 31988 17956 31989 17996
rect 31947 17947 31989 17956
rect 32139 17996 32181 18005
rect 32139 17956 32140 17996
rect 32180 17956 32181 17996
rect 32139 17947 32181 17956
rect 31755 17828 31797 17837
rect 31755 17788 31756 17828
rect 31796 17788 31797 17828
rect 31755 17779 31797 17788
rect 30219 17744 30261 17753
rect 30219 17704 30220 17744
rect 30260 17704 30261 17744
rect 30219 17695 30261 17704
rect 31180 17072 31220 17081
rect 29740 16988 29780 16997
rect 29780 16948 29972 16988
rect 29740 16939 29780 16948
rect 29932 16232 29972 16948
rect 31180 16829 31220 17032
rect 31179 16820 31221 16829
rect 31179 16780 31180 16820
rect 31220 16780 31221 16820
rect 31179 16771 31221 16780
rect 31659 16400 31701 16409
rect 31659 16360 31660 16400
rect 31700 16360 31701 16400
rect 31659 16351 31701 16360
rect 29932 16183 29972 16192
rect 31660 15644 31700 16351
rect 31660 15595 31700 15604
rect 31756 9437 31796 17779
rect 32140 17753 32180 17947
rect 32235 17912 32277 17921
rect 32235 17872 32236 17912
rect 32276 17872 32277 17912
rect 32235 17863 32277 17872
rect 32139 17744 32181 17753
rect 32139 17704 32140 17744
rect 32180 17704 32181 17744
rect 32139 17695 32181 17704
rect 32236 17744 32276 17863
rect 32140 17610 32180 17695
rect 32236 17585 32276 17704
rect 32428 17744 32468 18199
rect 32524 17921 32564 19804
rect 33004 19795 33044 19804
rect 33388 19844 33428 19853
rect 32812 19424 32852 19433
rect 32852 19384 32948 19424
rect 32812 19375 32852 19384
rect 32619 19256 32661 19265
rect 32619 19216 32620 19256
rect 32660 19216 32661 19256
rect 32619 19207 32661 19216
rect 32620 19088 32660 19207
rect 32620 19039 32660 19048
rect 32812 18677 32852 18721
rect 32811 18668 32853 18677
rect 32811 18628 32812 18668
rect 32852 18628 32853 18668
rect 32908 18668 32948 19384
rect 33388 19349 33428 19804
rect 33484 19601 33524 20140
rect 33580 20012 33620 20021
rect 33676 20012 33716 20551
rect 33964 20021 34004 20803
rect 34636 20189 34676 21568
rect 35307 21608 35349 21617
rect 35307 21568 35308 21608
rect 35348 21568 35349 21608
rect 35307 21559 35349 21568
rect 35404 20945 35444 22156
rect 35499 22147 35541 22156
rect 35596 22112 35636 22121
rect 35499 21608 35541 21617
rect 35499 21568 35500 21608
rect 35540 21568 35541 21608
rect 35499 21559 35541 21568
rect 35500 21474 35540 21559
rect 35403 20936 35445 20945
rect 35403 20896 35404 20936
rect 35444 20896 35445 20936
rect 35403 20887 35445 20896
rect 35211 20768 35253 20777
rect 35211 20728 35212 20768
rect 35252 20728 35253 20768
rect 35404 20768 35444 20887
rect 35596 20852 35636 22072
rect 35692 22037 35732 22240
rect 35788 22280 35828 22660
rect 35884 22280 35924 23323
rect 35979 23288 36021 23297
rect 35979 23248 35980 23288
rect 36020 23248 36021 23288
rect 35979 23239 36021 23248
rect 35980 22457 36020 23239
rect 35979 22448 36021 22457
rect 35979 22408 35980 22448
rect 36020 22408 36021 22448
rect 35979 22399 36021 22408
rect 36076 22364 36116 23584
rect 36268 23575 36308 23584
rect 36652 23624 36692 23633
rect 36172 23120 36212 23129
rect 36172 22448 36212 23080
rect 36652 23120 36692 23584
rect 36747 23624 36789 23633
rect 36747 23584 36748 23624
rect 36788 23584 36789 23624
rect 36747 23575 36789 23584
rect 36747 23456 36789 23465
rect 36747 23416 36748 23456
rect 36788 23416 36789 23456
rect 36844 23456 36884 23752
rect 36940 23792 36980 23801
rect 37036 23792 37076 24079
rect 36980 23752 37076 23792
rect 36940 23743 36980 23752
rect 37036 23465 37076 23752
rect 37035 23456 37077 23465
rect 36844 23416 36980 23456
rect 36747 23407 36789 23416
rect 36652 23071 36692 23080
rect 36748 23120 36788 23407
rect 36364 22868 36404 22877
rect 36172 22399 36212 22408
rect 36268 22828 36364 22868
rect 36076 22315 36116 22324
rect 36268 22364 36308 22828
rect 36364 22819 36404 22828
rect 36748 22541 36788 23080
rect 36844 23292 36884 23301
rect 36940 23297 36980 23416
rect 37035 23416 37036 23456
rect 37076 23416 37077 23456
rect 37035 23407 37077 23416
rect 36844 22868 36884 23252
rect 36939 23288 36981 23297
rect 36939 23248 36940 23288
rect 36980 23248 36981 23288
rect 36939 23239 36981 23248
rect 37036 23129 37076 23214
rect 37228 23213 37268 24247
rect 37612 23969 37652 24592
rect 37900 24632 37940 24641
rect 37900 24137 37940 24592
rect 37996 24632 38036 24641
rect 37996 24380 38036 24592
rect 38091 24632 38133 24641
rect 38091 24592 38092 24632
rect 38132 24592 38133 24632
rect 38091 24583 38133 24592
rect 37996 24340 38132 24380
rect 37899 24128 37941 24137
rect 37899 24088 37900 24128
rect 37940 24088 37941 24128
rect 37899 24079 37941 24088
rect 38092 24053 38132 24340
rect 38091 24044 38133 24053
rect 38091 24004 38092 24044
rect 38132 24004 38133 24044
rect 38091 23995 38133 24004
rect 37611 23960 37653 23969
rect 37611 23920 37612 23960
rect 37652 23920 37653 23960
rect 37611 23911 37653 23920
rect 37995 23960 38037 23969
rect 37995 23920 37996 23960
rect 38036 23920 38037 23960
rect 37995 23911 38037 23920
rect 37900 23876 37940 23885
rect 37804 23792 37844 23801
rect 37323 23624 37365 23633
rect 37323 23584 37324 23624
rect 37364 23584 37365 23624
rect 37323 23575 37365 23584
rect 37227 23204 37269 23213
rect 37227 23164 37228 23204
rect 37268 23164 37269 23204
rect 37227 23155 37269 23164
rect 37035 23120 37077 23129
rect 37035 23080 37036 23120
rect 37076 23080 37077 23120
rect 37035 23071 37077 23080
rect 37132 22868 37172 22877
rect 36844 22828 37132 22868
rect 36747 22532 36789 22541
rect 36747 22492 36748 22532
rect 36788 22492 36789 22532
rect 36747 22483 36789 22492
rect 36268 22289 36308 22324
rect 35980 22280 36020 22289
rect 35884 22240 35980 22280
rect 35788 22231 35828 22240
rect 35980 22231 36020 22240
rect 36267 22280 36309 22289
rect 36267 22240 36268 22280
rect 36308 22240 36309 22280
rect 36267 22231 36309 22240
rect 36364 22280 36404 22289
rect 36844 22280 36884 22828
rect 37132 22819 37172 22828
rect 37227 22364 37269 22373
rect 37227 22324 37228 22364
rect 37268 22324 37269 22364
rect 37227 22315 37269 22324
rect 36404 22240 36884 22280
rect 36940 22280 36980 22289
rect 36364 22231 36404 22240
rect 35691 22028 35733 22037
rect 35691 21988 35692 22028
rect 35732 21988 35733 22028
rect 35691 21979 35733 21988
rect 36747 22028 36789 22037
rect 36747 21988 36748 22028
rect 36788 21988 36789 22028
rect 36747 21979 36789 21988
rect 36076 21780 36116 21789
rect 36076 21692 36116 21740
rect 35980 21652 36116 21692
rect 35884 21608 35924 21617
rect 35692 21568 35884 21608
rect 35692 20936 35732 21568
rect 35884 21559 35924 21568
rect 35787 21356 35829 21365
rect 35787 21316 35788 21356
rect 35828 21316 35829 21356
rect 35787 21307 35829 21316
rect 35692 20887 35732 20896
rect 35596 20803 35636 20812
rect 35788 20852 35828 21307
rect 35788 20803 35828 20812
rect 35500 20768 35540 20777
rect 35404 20728 35500 20768
rect 35211 20719 35253 20728
rect 35500 20719 35540 20728
rect 35884 20768 35924 20777
rect 35980 20768 36020 21652
rect 35924 20728 36020 20768
rect 36172 21608 36212 21617
rect 35212 20634 35252 20719
rect 35308 20600 35348 20609
rect 35884 20600 35924 20728
rect 36172 20609 36212 21568
rect 36268 21608 36308 21617
rect 36268 20777 36308 21568
rect 36555 21356 36597 21365
rect 36555 21316 36556 21356
rect 36596 21316 36597 21356
rect 36555 21307 36597 21316
rect 36556 21222 36596 21307
rect 36748 21020 36788 21979
rect 36940 21701 36980 22240
rect 37036 22280 37076 22289
rect 37036 22121 37076 22240
rect 37131 22280 37173 22289
rect 37131 22240 37132 22280
rect 37172 22240 37173 22280
rect 37131 22231 37173 22240
rect 37228 22280 37268 22315
rect 37132 22146 37172 22231
rect 37228 22229 37268 22240
rect 37035 22112 37077 22121
rect 37035 22072 37036 22112
rect 37076 22072 37077 22112
rect 37035 22063 37077 22072
rect 36939 21692 36981 21701
rect 36939 21652 36940 21692
rect 36980 21652 36981 21692
rect 36939 21643 36981 21652
rect 37227 21692 37269 21701
rect 37227 21652 37228 21692
rect 37268 21652 37269 21692
rect 37227 21643 37269 21652
rect 36940 21608 36980 21643
rect 36940 21557 36980 21568
rect 37035 21608 37077 21617
rect 37035 21568 37036 21608
rect 37076 21568 37077 21608
rect 37035 21559 37077 21568
rect 37132 21608 37172 21617
rect 37036 21474 37076 21559
rect 37132 21365 37172 21568
rect 37228 21558 37268 21643
rect 37131 21356 37173 21365
rect 37131 21316 37132 21356
rect 37172 21316 37173 21356
rect 37131 21307 37173 21316
rect 36748 20980 36884 21020
rect 36267 20768 36309 20777
rect 36267 20728 36268 20768
rect 36308 20728 36309 20768
rect 36267 20719 36309 20728
rect 36748 20768 36788 20777
rect 36748 20609 36788 20728
rect 36844 20768 36884 20980
rect 37036 20777 37076 20862
rect 36844 20719 36884 20728
rect 36940 20768 36980 20777
rect 35348 20560 35924 20600
rect 36171 20600 36213 20609
rect 36171 20560 36172 20600
rect 36212 20560 36213 20600
rect 35308 20551 35348 20560
rect 36171 20551 36213 20560
rect 36747 20600 36789 20609
rect 36747 20560 36748 20600
rect 36788 20560 36789 20600
rect 36940 20600 36980 20728
rect 37035 20768 37077 20777
rect 37035 20728 37036 20768
rect 37076 20728 37077 20768
rect 37035 20719 37077 20728
rect 37324 20684 37364 23575
rect 37804 23381 37844 23752
rect 37900 23666 37940 23836
rect 37996 23826 38036 23911
rect 38091 23876 38133 23885
rect 38091 23836 38092 23876
rect 38132 23836 38133 23876
rect 38091 23827 38133 23836
rect 38092 23742 38132 23827
rect 38188 23792 38228 25087
rect 38284 24380 38324 24389
rect 38284 23885 38324 24340
rect 38283 23876 38325 23885
rect 38283 23836 38284 23876
rect 38324 23836 38325 23876
rect 38283 23827 38325 23836
rect 38188 23743 38228 23752
rect 38380 23666 38420 25096
rect 38476 25087 38516 25096
rect 38572 24800 38612 25264
rect 38668 25304 38708 25927
rect 38668 25255 38708 25264
rect 38572 24760 38708 24800
rect 38475 24716 38517 24725
rect 38475 24676 38476 24716
rect 38516 24676 38517 24716
rect 38475 24667 38517 24676
rect 38476 24582 38516 24667
rect 38571 24632 38613 24641
rect 38571 24592 38572 24632
rect 38612 24592 38613 24632
rect 38571 24583 38613 24592
rect 38475 24128 38517 24137
rect 38475 24088 38476 24128
rect 38516 24088 38517 24128
rect 38475 24079 38517 24088
rect 38476 23717 38516 24079
rect 37900 23626 38420 23666
rect 38475 23708 38517 23717
rect 38475 23668 38476 23708
rect 38516 23668 38517 23708
rect 38475 23659 38517 23668
rect 37803 23372 37845 23381
rect 37803 23332 37804 23372
rect 37844 23332 37845 23372
rect 37803 23323 37845 23332
rect 37515 23288 37557 23297
rect 37515 23248 37516 23288
rect 37556 23248 37557 23288
rect 37515 23239 37557 23248
rect 37420 23120 37460 23129
rect 37420 22373 37460 23080
rect 37419 22364 37461 22373
rect 37419 22324 37420 22364
rect 37460 22324 37461 22364
rect 37419 22315 37461 22324
rect 37516 22280 37556 23239
rect 37707 23204 37749 23213
rect 37707 23164 37708 23204
rect 37748 23164 37749 23204
rect 37707 23155 37749 23164
rect 37708 22532 37748 23155
rect 37804 23120 37844 23129
rect 38572 23120 38612 24583
rect 38668 24221 38708 24760
rect 38860 24632 38900 26104
rect 38956 26095 38996 26104
rect 39436 26104 39532 26144
rect 39436 25901 39476 26104
rect 39532 26095 39572 26104
rect 39627 26144 39669 26153
rect 39627 26104 39628 26144
rect 39668 26104 39669 26144
rect 39627 26095 39669 26104
rect 39724 26144 39764 26272
rect 39628 26010 39668 26095
rect 39531 25976 39573 25985
rect 39531 25936 39532 25976
rect 39572 25936 39573 25976
rect 39531 25927 39573 25936
rect 39435 25892 39477 25901
rect 39435 25852 39436 25892
rect 39476 25852 39477 25892
rect 39435 25843 39477 25852
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 39532 25388 39572 25927
rect 39627 25892 39669 25901
rect 39627 25852 39628 25892
rect 39668 25852 39669 25892
rect 39627 25843 39669 25852
rect 39532 25339 39572 25348
rect 39628 25145 39668 25843
rect 39724 25556 39764 26104
rect 39820 26144 39860 26153
rect 40012 26144 40052 26153
rect 39860 26104 40012 26144
rect 39820 26095 39860 26104
rect 40012 26095 40052 26104
rect 40108 25976 40148 26599
rect 40204 26144 40244 26767
rect 40395 26816 40437 26825
rect 40395 26776 40396 26816
rect 40436 26776 40437 26816
rect 40395 26767 40437 26776
rect 40492 26816 40532 26827
rect 40300 26741 40340 26755
rect 40299 26732 40341 26741
rect 40299 26692 40300 26732
rect 40340 26692 40341 26732
rect 40299 26683 40341 26692
rect 40396 26682 40436 26767
rect 40492 26741 40532 26776
rect 40875 26816 40917 26825
rect 40875 26776 40876 26816
rect 40916 26776 40917 26816
rect 40875 26767 40917 26776
rect 40491 26732 40533 26741
rect 40491 26692 40492 26732
rect 40532 26692 40533 26732
rect 40491 26683 40533 26692
rect 40588 26657 40628 26742
rect 40779 26732 40821 26741
rect 40779 26692 40780 26732
rect 40820 26692 40821 26732
rect 40779 26683 40821 26692
rect 40587 26648 40629 26657
rect 40587 26608 40588 26648
rect 40628 26608 40629 26648
rect 40587 26599 40629 26608
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 40395 26228 40437 26237
rect 40395 26188 40396 26228
rect 40436 26188 40437 26228
rect 40395 26179 40437 26188
rect 40396 26144 40436 26179
rect 40204 26104 40340 26144
rect 39724 25507 39764 25516
rect 40012 25936 40148 25976
rect 39819 25304 39861 25313
rect 39819 25264 39820 25304
rect 39860 25264 39861 25304
rect 39819 25255 39861 25264
rect 40012 25304 40052 25936
rect 40107 25808 40149 25817
rect 40107 25768 40108 25808
rect 40148 25768 40149 25808
rect 40107 25759 40149 25768
rect 40012 25255 40052 25264
rect 40108 25304 40148 25759
rect 39339 25136 39381 25145
rect 39339 25096 39340 25136
rect 39380 25096 39381 25136
rect 39339 25087 39381 25096
rect 39627 25136 39669 25145
rect 39627 25096 39628 25136
rect 39668 25096 39669 25136
rect 39627 25087 39669 25096
rect 39340 25002 39380 25087
rect 38955 24716 38997 24725
rect 38955 24676 38956 24716
rect 38996 24676 38997 24716
rect 38955 24667 38997 24676
rect 38860 24305 38900 24592
rect 38859 24296 38901 24305
rect 38859 24256 38860 24296
rect 38900 24256 38901 24296
rect 38859 24247 38901 24256
rect 38667 24212 38709 24221
rect 38667 24172 38668 24212
rect 38708 24172 38709 24212
rect 38667 24163 38709 24172
rect 38667 24044 38709 24053
rect 38667 24004 38668 24044
rect 38708 24004 38709 24044
rect 38956 24044 38996 24667
rect 39723 24632 39765 24641
rect 39723 24592 39724 24632
rect 39764 24592 39765 24632
rect 39723 24583 39765 24592
rect 39724 24498 39764 24583
rect 39820 24380 39860 25255
rect 39915 24800 39957 24809
rect 39915 24760 39916 24800
rect 39956 24760 39957 24800
rect 39915 24751 39957 24760
rect 39724 24340 39860 24380
rect 39627 24296 39669 24305
rect 39627 24256 39628 24296
rect 39668 24256 39669 24296
rect 39627 24247 39669 24256
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 38956 24004 39188 24044
rect 38667 23995 38709 24004
rect 38668 23792 38708 23995
rect 38859 23960 38901 23969
rect 38859 23920 38860 23960
rect 38900 23920 38901 23960
rect 38859 23911 38901 23920
rect 38668 23743 38708 23752
rect 38764 23792 38804 23801
rect 38764 23633 38804 23752
rect 38860 23792 38900 23911
rect 38763 23624 38805 23633
rect 38763 23584 38764 23624
rect 38804 23584 38805 23624
rect 38763 23575 38805 23584
rect 38668 23120 38708 23129
rect 38572 23080 38668 23120
rect 37804 23060 37844 23080
rect 37804 23020 37940 23060
rect 37804 22532 37844 22541
rect 37708 22492 37804 22532
rect 37804 22483 37844 22492
rect 37708 22280 37748 22289
rect 37516 22231 37556 22240
rect 37612 22240 37708 22280
rect 37419 22112 37461 22121
rect 37419 22072 37420 22112
rect 37460 22072 37461 22112
rect 37419 22063 37461 22072
rect 37420 21978 37460 22063
rect 37612 22037 37652 22240
rect 37708 22231 37748 22240
rect 37804 22112 37844 22121
rect 37708 22072 37804 22112
rect 37611 22028 37653 22037
rect 37611 21988 37612 22028
rect 37652 21988 37653 22028
rect 37611 21979 37653 21988
rect 37419 21692 37461 21701
rect 37419 21652 37420 21692
rect 37460 21652 37461 21692
rect 37419 21643 37461 21652
rect 37420 21558 37460 21643
rect 37708 21617 37748 22072
rect 37804 22063 37844 22072
rect 37707 21608 37749 21617
rect 37707 21568 37708 21608
rect 37748 21568 37749 21608
rect 37707 21559 37749 21568
rect 37804 21608 37844 21617
rect 37900 21608 37940 23020
rect 38668 21608 38708 23080
rect 38860 22280 38900 23752
rect 38956 23792 38996 23803
rect 38956 23717 38996 23752
rect 39148 23792 39188 24004
rect 39243 23876 39285 23885
rect 39243 23836 39244 23876
rect 39284 23836 39285 23876
rect 39243 23827 39285 23836
rect 39148 23743 39188 23752
rect 39244 23792 39284 23827
rect 39244 23741 39284 23752
rect 39340 23792 39380 23801
rect 38955 23708 38997 23717
rect 38955 23668 38956 23708
rect 38996 23668 38997 23708
rect 38955 23659 38997 23668
rect 39340 23060 39380 23752
rect 39436 23792 39476 23801
rect 39436 23633 39476 23752
rect 39435 23624 39477 23633
rect 39435 23584 39436 23624
rect 39476 23584 39477 23624
rect 39435 23575 39477 23584
rect 39340 23020 39572 23060
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 39436 22532 39476 22541
rect 39532 22532 39572 23020
rect 39476 22492 39572 22532
rect 39436 22483 39476 22492
rect 39532 22280 39572 22289
rect 38860 22240 39532 22280
rect 39532 22231 39572 22240
rect 39436 22112 39476 22123
rect 39436 22037 39476 22072
rect 39435 22028 39477 22037
rect 39435 21988 39436 22028
rect 39476 21988 39477 22028
rect 39435 21979 39477 21988
rect 39628 21608 39668 24247
rect 37844 21568 37940 21608
rect 37804 21559 37844 21568
rect 37900 21449 37940 21568
rect 38572 21568 38668 21608
rect 37899 21440 37941 21449
rect 37899 21400 37900 21440
rect 37940 21400 37941 21440
rect 37899 21391 37941 21400
rect 38283 21440 38325 21449
rect 38283 21400 38284 21440
rect 38324 21400 38325 21440
rect 38283 21391 38325 21400
rect 37419 20852 37461 20861
rect 37419 20812 37420 20852
rect 37460 20812 37461 20852
rect 37419 20803 37461 20812
rect 37420 20718 37460 20803
rect 37228 20644 37364 20684
rect 37228 20600 37268 20644
rect 36940 20560 37268 20600
rect 37612 20600 37652 20609
rect 36747 20551 36789 20560
rect 34635 20180 34677 20189
rect 34635 20140 34636 20180
rect 34676 20140 34677 20180
rect 34635 20131 34677 20140
rect 33620 19972 33716 20012
rect 33963 20012 34005 20021
rect 33963 19972 33964 20012
rect 34004 19972 34005 20012
rect 33580 19963 33620 19972
rect 33963 19963 34005 19972
rect 33964 19878 34004 19963
rect 33772 19844 33812 19853
rect 33483 19592 33525 19601
rect 33483 19552 33484 19592
rect 33524 19552 33525 19592
rect 33483 19543 33525 19552
rect 33579 19508 33621 19517
rect 33579 19468 33580 19508
rect 33620 19468 33621 19508
rect 33579 19459 33621 19468
rect 33387 19340 33429 19349
rect 33387 19300 33388 19340
rect 33428 19300 33429 19340
rect 33387 19291 33429 19300
rect 33100 19254 33140 19263
rect 33100 18929 33140 19214
rect 33195 19256 33237 19265
rect 33195 19216 33196 19256
rect 33236 19216 33237 19256
rect 33195 19207 33237 19216
rect 33196 19122 33236 19207
rect 33292 19030 33332 19039
rect 33388 19013 33428 19291
rect 33580 19256 33620 19459
rect 33772 19433 33812 19804
rect 34539 19844 34581 19853
rect 34539 19804 34540 19844
rect 34580 19804 34581 19844
rect 34539 19795 34581 19804
rect 34251 19508 34293 19517
rect 34251 19468 34252 19508
rect 34292 19468 34293 19508
rect 34251 19459 34293 19468
rect 33771 19424 33813 19433
rect 33580 19207 33620 19216
rect 33676 19384 33772 19424
rect 33812 19384 33813 19424
rect 33099 18920 33141 18929
rect 33099 18880 33100 18920
rect 33140 18880 33141 18920
rect 33099 18871 33141 18880
rect 33195 18752 33237 18761
rect 33195 18712 33196 18752
rect 33236 18712 33237 18752
rect 33195 18703 33237 18712
rect 33292 18752 33332 18990
rect 33387 19004 33429 19013
rect 33387 18964 33388 19004
rect 33428 18964 33429 19004
rect 33387 18955 33429 18964
rect 33579 18920 33621 18929
rect 33579 18880 33580 18920
rect 33620 18880 33621 18920
rect 33579 18871 33621 18880
rect 33484 18752 33524 18761
rect 33292 18712 33484 18752
rect 32908 18628 32975 18668
rect 32811 18626 32853 18628
rect 32811 18619 32812 18626
rect 32620 18584 32660 18593
rect 32852 18619 32853 18626
rect 32812 18577 32852 18586
rect 32620 18248 32660 18544
rect 32935 18542 32975 18628
rect 32715 18500 32757 18509
rect 32935 18500 32975 18502
rect 32715 18460 32716 18500
rect 32756 18460 32975 18500
rect 33196 18584 33236 18703
rect 33292 18593 33332 18712
rect 33484 18703 33524 18712
rect 32715 18451 32757 18460
rect 33100 18458 33140 18467
rect 33004 18416 33044 18425
rect 33004 18248 33044 18376
rect 32620 18208 33044 18248
rect 33100 18089 33140 18418
rect 33196 18341 33236 18544
rect 33291 18584 33333 18593
rect 33291 18544 33292 18584
rect 33332 18544 33333 18584
rect 33291 18535 33333 18544
rect 33388 18584 33428 18593
rect 33195 18332 33237 18341
rect 33195 18292 33196 18332
rect 33236 18292 33237 18332
rect 33195 18283 33237 18292
rect 33099 18080 33141 18089
rect 33099 18040 33100 18080
rect 33140 18040 33141 18080
rect 33099 18031 33141 18040
rect 33388 18005 33428 18544
rect 33387 17996 33429 18005
rect 33387 17956 33388 17996
rect 33428 17956 33429 17996
rect 33387 17947 33429 17956
rect 32523 17912 32565 17921
rect 32523 17872 32524 17912
rect 32564 17872 32565 17912
rect 32523 17863 32565 17872
rect 32907 17912 32949 17921
rect 33580 17912 33620 18871
rect 33676 18761 33716 19384
rect 33771 19375 33813 19384
rect 33771 19256 33813 19265
rect 33771 19216 33772 19256
rect 33812 19216 33813 19256
rect 33771 19207 33813 19216
rect 33964 19256 34004 19267
rect 33675 18752 33717 18761
rect 33675 18712 33676 18752
rect 33716 18712 33717 18752
rect 33675 18703 33717 18712
rect 33676 18584 33716 18703
rect 33676 18535 33716 18544
rect 33676 18332 33716 18341
rect 33676 18089 33716 18292
rect 33675 18080 33717 18089
rect 33675 18040 33676 18080
rect 33716 18040 33717 18080
rect 33675 18031 33717 18040
rect 32907 17872 32908 17912
rect 32948 17872 32949 17912
rect 32907 17863 32949 17872
rect 33484 17872 33620 17912
rect 32812 17753 32852 17838
rect 32716 17744 32756 17753
rect 32235 17576 32277 17585
rect 32235 17536 32236 17576
rect 32276 17536 32277 17576
rect 32235 17527 32277 17536
rect 32332 17576 32372 17585
rect 32235 17324 32277 17333
rect 32235 17284 32236 17324
rect 32276 17284 32277 17324
rect 32235 17275 32277 17284
rect 32043 17156 32085 17165
rect 32043 17116 32044 17156
rect 32084 17116 32085 17156
rect 32043 17107 32085 17116
rect 32044 16241 32084 17107
rect 32236 16904 32276 17275
rect 32140 16864 32236 16904
rect 32140 16316 32180 16864
rect 32236 16855 32276 16864
rect 32235 16400 32277 16409
rect 32235 16360 32236 16400
rect 32276 16360 32277 16400
rect 32235 16351 32277 16360
rect 32140 16267 32180 16276
rect 32236 16266 32276 16351
rect 32332 16316 32372 17536
rect 32332 16267 32372 16276
rect 32043 16232 32085 16241
rect 32043 16192 32044 16232
rect 32084 16192 32085 16232
rect 32043 16183 32085 16192
rect 32428 16232 32468 17704
rect 32524 17704 32716 17744
rect 32524 17333 32564 17704
rect 32716 17695 32756 17704
rect 32811 17744 32853 17753
rect 32811 17704 32812 17744
rect 32852 17704 32853 17744
rect 32811 17695 32853 17704
rect 32908 17744 32948 17863
rect 33291 17828 33333 17837
rect 33484 17828 33524 17872
rect 33291 17788 33292 17828
rect 33332 17788 33333 17828
rect 33291 17779 33333 17788
rect 33388 17788 33524 17828
rect 32908 17660 32948 17704
rect 33099 17744 33141 17753
rect 33099 17704 33100 17744
rect 33140 17704 33141 17744
rect 33099 17695 33141 17704
rect 33196 17744 33236 17753
rect 32908 17620 33044 17660
rect 32620 17576 32660 17585
rect 32660 17536 32948 17576
rect 32620 17527 32660 17536
rect 32523 17324 32565 17333
rect 32523 17284 32524 17324
rect 32564 17284 32565 17324
rect 32523 17275 32565 17284
rect 32811 17324 32853 17333
rect 32811 17284 32812 17324
rect 32852 17284 32853 17324
rect 32811 17275 32853 17284
rect 32716 17244 32756 17253
rect 32716 17165 32756 17204
rect 32715 17156 32757 17165
rect 32715 17116 32716 17156
rect 32756 17116 32757 17156
rect 32715 17107 32757 17116
rect 32524 17072 32564 17081
rect 32524 16652 32564 17032
rect 32517 16612 32564 16652
rect 32620 17072 32660 17081
rect 32517 16568 32557 16612
rect 32517 16528 32564 16568
rect 32524 16232 32564 16528
rect 32620 16409 32660 17032
rect 32812 16736 32852 17275
rect 32908 17156 32948 17536
rect 33004 17333 33044 17620
rect 33100 17610 33140 17695
rect 33003 17324 33045 17333
rect 33003 17284 33004 17324
rect 33044 17284 33045 17324
rect 33003 17275 33045 17284
rect 32908 17107 32948 17116
rect 33196 16997 33236 17704
rect 33292 17618 33332 17779
rect 33388 17744 33428 17788
rect 33579 17744 33621 17753
rect 33388 17695 33428 17704
rect 33484 17723 33524 17732
rect 33579 17704 33580 17744
rect 33620 17704 33621 17744
rect 33579 17695 33621 17704
rect 33676 17744 33716 17753
rect 33772 17744 33812 19207
rect 33964 19181 34004 19216
rect 34059 19256 34101 19265
rect 34059 19216 34060 19256
rect 34100 19216 34101 19256
rect 34059 19207 34101 19216
rect 33963 19172 34005 19181
rect 33963 19132 33964 19172
rect 34004 19132 34005 19172
rect 33963 19123 34005 19132
rect 33963 18752 34005 18761
rect 33963 18712 33964 18752
rect 34004 18712 34005 18752
rect 33963 18703 34005 18712
rect 33716 17704 33812 17744
rect 33868 18584 33908 18593
rect 33484 17618 33524 17683
rect 33292 17578 33524 17618
rect 33580 17610 33620 17695
rect 33291 17072 33333 17081
rect 33291 17032 33292 17072
rect 33332 17032 33333 17072
rect 33291 17023 33333 17032
rect 33003 16988 33045 16997
rect 33003 16948 33004 16988
rect 33044 16948 33045 16988
rect 33003 16939 33045 16948
rect 33195 16988 33237 16997
rect 33195 16948 33196 16988
rect 33236 16948 33237 16988
rect 33195 16939 33237 16948
rect 32812 16696 32949 16736
rect 32909 16568 32949 16696
rect 32908 16528 32949 16568
rect 32619 16400 32661 16409
rect 32619 16360 32620 16400
rect 32660 16360 32661 16400
rect 32619 16351 32661 16360
rect 32812 16232 32852 16241
rect 32524 16192 32812 16232
rect 32428 16183 32468 16192
rect 32812 16183 32852 16192
rect 32908 16232 32948 16528
rect 32908 16183 32948 16192
rect 33004 16232 33044 16939
rect 33099 16400 33141 16409
rect 33099 16360 33100 16400
rect 33140 16360 33141 16400
rect 33099 16351 33141 16360
rect 33004 16183 33044 16192
rect 33100 16232 33140 16351
rect 33100 16183 33140 16192
rect 32044 16098 32084 16183
rect 32044 15560 32084 15569
rect 32044 15233 32084 15520
rect 32907 15560 32949 15569
rect 32907 15520 32908 15560
rect 32948 15520 32949 15560
rect 32907 15511 32949 15520
rect 32908 15426 32948 15511
rect 33292 15233 33332 17023
rect 33676 16409 33716 17704
rect 33868 17585 33908 18544
rect 33964 18584 34004 18703
rect 33964 18535 34004 18544
rect 33867 17576 33909 17585
rect 33867 17536 33868 17576
rect 33908 17536 33909 17576
rect 33867 17527 33909 17536
rect 33868 17417 33908 17527
rect 33867 17408 33909 17417
rect 33867 17368 33868 17408
rect 33908 17368 33909 17408
rect 33867 17359 33909 17368
rect 34060 17072 34100 19207
rect 34156 18752 34196 18761
rect 34252 18752 34292 19459
rect 34540 18761 34580 19795
rect 34636 19265 34676 20131
rect 35692 20096 35732 20105
rect 35692 19265 35732 20056
rect 36555 20096 36597 20105
rect 36555 20056 36556 20096
rect 36596 20056 36597 20096
rect 36555 20047 36597 20056
rect 36940 20096 36980 20105
rect 36556 19962 36596 20047
rect 35787 19928 35829 19937
rect 35787 19888 35788 19928
rect 35828 19888 35829 19928
rect 35787 19879 35829 19888
rect 34635 19256 34677 19265
rect 34635 19216 34636 19256
rect 34676 19216 34677 19256
rect 34635 19207 34677 19216
rect 34827 19256 34869 19265
rect 34827 19216 34828 19256
rect 34868 19216 34869 19256
rect 34827 19207 34869 19216
rect 35691 19256 35733 19265
rect 35691 19216 35692 19256
rect 35732 19216 35733 19256
rect 35691 19207 35733 19216
rect 34828 19122 34868 19207
rect 35692 18929 35732 19207
rect 35691 18920 35733 18929
rect 35691 18880 35692 18920
rect 35732 18880 35733 18920
rect 35691 18871 35733 18880
rect 34196 18712 34292 18752
rect 34539 18752 34581 18761
rect 34539 18712 34540 18752
rect 34580 18712 34581 18752
rect 34156 18703 34196 18712
rect 34539 18703 34581 18712
rect 34251 18584 34293 18593
rect 34251 18544 34252 18584
rect 34292 18544 34293 18584
rect 34251 18535 34293 18544
rect 34348 18584 34388 18593
rect 34252 18450 34292 18535
rect 34348 18341 34388 18544
rect 34444 18584 34484 18595
rect 34444 18509 34484 18544
rect 34635 18584 34677 18593
rect 34635 18544 34636 18584
rect 34676 18544 34677 18584
rect 34635 18535 34677 18544
rect 34443 18500 34485 18509
rect 34443 18460 34444 18500
rect 34484 18460 34485 18500
rect 34443 18451 34485 18460
rect 34347 18332 34389 18341
rect 34347 18292 34348 18332
rect 34388 18292 34389 18332
rect 34347 18283 34389 18292
rect 34347 18164 34389 18173
rect 34347 18124 34348 18164
rect 34388 18124 34389 18164
rect 34347 18115 34389 18124
rect 34156 17072 34196 17081
rect 34060 17032 34156 17072
rect 34156 17023 34196 17032
rect 33675 16400 33717 16409
rect 33675 16360 33676 16400
rect 33716 16360 33717 16400
rect 33675 16351 33717 16360
rect 33387 16232 33429 16241
rect 33387 16192 33388 16232
rect 33428 16192 33429 16232
rect 33387 16183 33429 16192
rect 33484 16232 33524 16241
rect 33524 16192 34100 16232
rect 33484 16183 33524 16192
rect 33388 16098 33428 16183
rect 34060 15728 34100 16192
rect 34348 15821 34388 18115
rect 34444 17837 34484 18451
rect 34539 18248 34581 18257
rect 34539 18208 34540 18248
rect 34580 18208 34581 18248
rect 34539 18199 34581 18208
rect 34443 17828 34485 17837
rect 34443 17788 34444 17828
rect 34484 17788 34485 17828
rect 34443 17779 34485 17788
rect 34443 17408 34485 17417
rect 34443 17368 34444 17408
rect 34484 17368 34485 17408
rect 34443 17359 34485 17368
rect 34347 15812 34389 15821
rect 34347 15772 34348 15812
rect 34388 15772 34389 15812
rect 34347 15763 34389 15772
rect 34100 15688 34292 15728
rect 34060 15679 34100 15688
rect 34252 15560 34292 15688
rect 34444 15644 34484 17359
rect 34252 15511 34292 15520
rect 34348 15604 34484 15644
rect 34348 15560 34388 15604
rect 34348 15511 34388 15520
rect 34444 15485 34484 15604
rect 34540 15560 34580 18199
rect 34636 17753 34676 18535
rect 34731 18332 34773 18341
rect 34731 18292 34732 18332
rect 34772 18292 34773 18332
rect 34731 18283 34773 18292
rect 34732 18198 34772 18283
rect 34635 17744 34677 17753
rect 34635 17704 34636 17744
rect 34676 17704 34677 17744
rect 34635 17695 34677 17704
rect 35596 17072 35636 17081
rect 35500 17032 35596 17072
rect 35307 16988 35349 16997
rect 35307 16948 35308 16988
rect 35348 16948 35349 16988
rect 35307 16939 35349 16948
rect 35308 16854 35348 16939
rect 35500 16232 35540 17032
rect 35596 17023 35636 17032
rect 35788 16325 35828 19879
rect 36940 19760 36980 20056
rect 37035 20096 37077 20105
rect 37035 20056 37036 20096
rect 37076 20056 37077 20096
rect 37035 20047 37077 20056
rect 36460 19720 36980 19760
rect 36460 19424 36500 19720
rect 36651 19508 36693 19517
rect 36651 19468 36652 19508
rect 36692 19468 36693 19508
rect 36651 19459 36693 19468
rect 36460 19375 36500 19384
rect 36555 19424 36597 19433
rect 36555 19384 36556 19424
rect 36596 19384 36597 19424
rect 36555 19375 36597 19384
rect 36364 19340 36404 19349
rect 36267 19256 36309 19265
rect 36267 19216 36268 19256
rect 36308 19216 36309 19256
rect 36267 19207 36309 19216
rect 36268 19122 36308 19207
rect 35980 19088 36020 19097
rect 36364 19088 36404 19300
rect 36556 19340 36596 19375
rect 36556 19289 36596 19300
rect 36652 19256 36692 19459
rect 36844 19424 36884 19433
rect 36652 19207 36692 19216
rect 36748 19384 36844 19424
rect 36748 19088 36788 19384
rect 36844 19375 36884 19384
rect 36364 19048 36788 19088
rect 35980 18593 36020 19048
rect 35979 18584 36021 18593
rect 35979 18544 35980 18584
rect 36020 18544 36021 18584
rect 35979 18535 36021 18544
rect 36460 18584 36500 18593
rect 35980 17921 36020 18535
rect 36460 18509 36500 18544
rect 36556 18584 36596 18593
rect 36459 18500 36501 18509
rect 36459 18460 36460 18500
rect 36500 18460 36501 18500
rect 36459 18451 36501 18460
rect 35979 17912 36021 17921
rect 35979 17872 35980 17912
rect 36020 17872 36021 17912
rect 35979 17863 36021 17872
rect 36460 17333 36500 18451
rect 36556 17585 36596 18544
rect 36652 18584 36692 19048
rect 36652 18535 36692 18544
rect 36748 18584 36788 18593
rect 36940 18584 36980 18593
rect 36788 18544 36940 18584
rect 37036 18584 37076 20047
rect 37132 19937 37172 20560
rect 37131 19928 37173 19937
rect 37131 19888 37132 19928
rect 37172 19888 37173 19928
rect 37131 19879 37173 19888
rect 37420 19844 37460 19853
rect 37132 19256 37172 19265
rect 37132 18761 37172 19216
rect 37228 19256 37268 19265
rect 37131 18752 37173 18761
rect 37131 18712 37132 18752
rect 37172 18712 37173 18752
rect 37228 18752 37268 19216
rect 37323 19256 37365 19265
rect 37323 19216 37324 19256
rect 37364 19216 37365 19256
rect 37323 19207 37365 19216
rect 37324 19084 37364 19207
rect 37324 19035 37364 19044
rect 37420 19013 37460 19804
rect 37515 19844 37557 19853
rect 37515 19804 37516 19844
rect 37556 19804 37557 19844
rect 37515 19795 37557 19804
rect 37516 19256 37556 19795
rect 37612 19517 37652 20560
rect 37611 19508 37653 19517
rect 37611 19468 37612 19508
rect 37652 19468 37653 19508
rect 37611 19459 37653 19468
rect 37516 19207 37556 19216
rect 37611 19256 37653 19265
rect 37611 19216 37612 19256
rect 37652 19216 37653 19256
rect 37611 19207 37653 19216
rect 37612 19122 37652 19207
rect 37419 19004 37461 19013
rect 37419 18964 37420 19004
rect 37460 18964 37461 19004
rect 37419 18955 37461 18964
rect 37707 18752 37749 18761
rect 37228 18712 37460 18752
rect 37131 18703 37173 18712
rect 37324 18584 37364 18593
rect 37036 18544 37324 18584
rect 36748 18535 36788 18544
rect 36940 18535 36980 18544
rect 36555 17576 36597 17585
rect 36555 17536 36556 17576
rect 36596 17536 36597 17576
rect 36555 17527 36597 17536
rect 36171 17324 36213 17333
rect 36171 17284 36172 17324
rect 36212 17284 36213 17324
rect 36171 17275 36213 17284
rect 36459 17324 36501 17333
rect 36459 17284 36460 17324
rect 36500 17284 36501 17324
rect 36459 17275 36501 17284
rect 35980 17072 36020 17081
rect 35980 16661 36020 17032
rect 35979 16652 36021 16661
rect 35979 16612 35980 16652
rect 36020 16612 36021 16652
rect 35979 16603 36021 16612
rect 35787 16316 35829 16325
rect 35787 16276 35788 16316
rect 35828 16276 35829 16316
rect 35787 16267 35829 16276
rect 35500 16183 35540 16192
rect 35596 16232 35636 16241
rect 35115 15728 35157 15737
rect 35115 15688 35116 15728
rect 35156 15688 35157 15728
rect 35115 15679 35157 15688
rect 34732 15560 34772 15569
rect 34580 15520 34732 15560
rect 34540 15511 34580 15520
rect 34732 15511 34772 15520
rect 35116 15560 35156 15679
rect 35116 15511 35156 15520
rect 34443 15476 34485 15485
rect 34443 15436 34444 15476
rect 34484 15436 34485 15476
rect 34443 15427 34485 15436
rect 34828 15476 34868 15485
rect 34540 15392 34580 15401
rect 34828 15392 34868 15436
rect 35020 15476 35060 15485
rect 34580 15352 34868 15392
rect 34924 15392 34964 15401
rect 35020 15392 35060 15436
rect 35500 15392 35540 15401
rect 35596 15392 35636 16192
rect 35692 16232 35732 16241
rect 35692 16073 35732 16192
rect 35788 16232 35828 16267
rect 35788 16182 35828 16192
rect 36172 16232 36212 17275
rect 37324 17081 37364 18544
rect 37420 17744 37460 18712
rect 37707 18712 37708 18752
rect 37748 18712 37749 18752
rect 37707 18703 37749 18712
rect 36844 17072 36884 17081
rect 36556 17032 36844 17072
rect 36363 16400 36405 16409
rect 36363 16360 36364 16400
rect 36404 16360 36405 16400
rect 36363 16351 36405 16360
rect 36172 16183 36212 16192
rect 36267 16232 36309 16241
rect 36267 16192 36268 16232
rect 36308 16192 36309 16232
rect 36267 16183 36309 16192
rect 36364 16232 36404 16351
rect 36268 16098 36308 16183
rect 35691 16064 35733 16073
rect 36076 16064 36116 16073
rect 35691 16024 35692 16064
rect 35732 16024 35733 16064
rect 35691 16015 35733 16024
rect 35788 16024 36076 16064
rect 35691 15560 35733 15569
rect 35691 15520 35692 15560
rect 35732 15520 35733 15560
rect 35691 15511 35733 15520
rect 35788 15560 35828 16024
rect 36076 16015 36116 16024
rect 35980 15737 36020 15823
rect 35979 15732 36021 15737
rect 35979 15688 35980 15732
rect 36020 15688 36021 15732
rect 35979 15679 36021 15688
rect 36171 15728 36213 15737
rect 36171 15688 36172 15728
rect 36212 15688 36213 15728
rect 36171 15679 36213 15688
rect 35883 15644 35925 15653
rect 35883 15604 35884 15644
rect 35924 15604 35925 15644
rect 35883 15595 35925 15604
rect 35788 15511 35828 15520
rect 35884 15560 35924 15595
rect 36172 15594 36212 15679
rect 36364 15653 36404 16192
rect 36363 15644 36405 15653
rect 36363 15604 36364 15644
rect 36404 15604 36405 15644
rect 36363 15595 36405 15604
rect 36556 15569 36596 17032
rect 36844 17023 36884 17032
rect 37323 17072 37365 17081
rect 37323 17032 37324 17072
rect 37364 17032 37365 17072
rect 37323 17023 37365 17032
rect 36939 16988 36981 16997
rect 36939 16948 36940 16988
rect 36980 16948 36981 16988
rect 36939 16939 36981 16948
rect 36843 16232 36885 16241
rect 36940 16232 36980 16939
rect 37420 16409 37460 17704
rect 37515 17744 37557 17753
rect 37515 17704 37516 17744
rect 37556 17704 37557 17744
rect 37515 17695 37557 17704
rect 37612 17744 37652 17753
rect 37516 17610 37556 17695
rect 37612 17333 37652 17704
rect 37708 17744 37748 18703
rect 37708 17695 37748 17704
rect 37611 17324 37653 17333
rect 37611 17284 37612 17324
rect 37652 17284 37653 17324
rect 37611 17275 37653 17284
rect 37803 17072 37845 17081
rect 37803 17032 37804 17072
rect 37844 17032 37845 17072
rect 37803 17023 37845 17032
rect 37419 16400 37461 16409
rect 37419 16360 37420 16400
rect 37460 16360 37461 16400
rect 37419 16351 37461 16360
rect 36843 16192 36844 16232
rect 36884 16192 36980 16232
rect 37708 16232 37748 16241
rect 36843 16183 36885 16192
rect 36844 16098 36884 16183
rect 37611 16148 37653 16157
rect 37611 16108 37612 16148
rect 37652 16108 37653 16148
rect 37611 16099 37653 16108
rect 36747 16064 36789 16073
rect 36747 16024 36748 16064
rect 36788 16024 36789 16064
rect 36747 16015 36789 16024
rect 36748 15930 36788 16015
rect 37612 16014 37652 16099
rect 37035 15644 37077 15653
rect 37035 15604 37036 15644
rect 37076 15604 37077 15644
rect 37035 15595 37077 15604
rect 35020 15352 35500 15392
rect 35540 15352 35636 15392
rect 34540 15343 34580 15352
rect 32043 15224 32085 15233
rect 32043 15184 32044 15224
rect 32084 15184 32085 15224
rect 32043 15175 32085 15184
rect 33291 15224 33333 15233
rect 33291 15184 33292 15224
rect 33332 15184 33333 15224
rect 33291 15175 33333 15184
rect 34827 15224 34869 15233
rect 34827 15184 34828 15224
rect 34868 15184 34869 15224
rect 34827 15175 34869 15184
rect 34443 14720 34485 14729
rect 34443 14680 34444 14720
rect 34484 14680 34485 14720
rect 34443 14671 34485 14680
rect 34828 14720 34868 15175
rect 34924 14729 34964 15352
rect 35500 15343 35540 15352
rect 34444 14586 34484 14671
rect 34828 14057 34868 14680
rect 34923 14720 34965 14729
rect 34923 14680 34924 14720
rect 34964 14680 34965 14720
rect 34923 14671 34965 14680
rect 35692 14720 35732 15511
rect 35884 15509 35924 15520
rect 36268 15560 36308 15569
rect 36268 15392 36308 15520
rect 36555 15560 36597 15569
rect 36555 15520 36556 15560
rect 36596 15520 36597 15560
rect 36555 15511 36597 15520
rect 36652 15560 36692 15569
rect 36652 15392 36692 15520
rect 36748 15560 36788 15571
rect 36748 15485 36788 15520
rect 36940 15549 36980 15558
rect 36747 15476 36789 15485
rect 36940 15476 36980 15509
rect 37036 15476 37076 15595
rect 36747 15436 36748 15476
rect 36788 15436 36789 15476
rect 36747 15427 36789 15436
rect 36844 15436 37076 15476
rect 36268 15352 36692 15392
rect 36652 14972 36692 15352
rect 36844 15140 36884 15436
rect 36940 15308 36980 15317
rect 37708 15308 37748 16192
rect 37804 16232 37844 17023
rect 37900 16661 37940 21391
rect 38092 19433 38132 19518
rect 38091 19424 38133 19433
rect 38091 19384 38092 19424
rect 38132 19384 38133 19424
rect 38091 19375 38133 19384
rect 38091 19256 38133 19265
rect 38091 19216 38092 19256
rect 38132 19216 38133 19256
rect 38091 19207 38133 19216
rect 38284 19256 38324 21391
rect 38572 20096 38612 21568
rect 38668 21559 38708 21568
rect 39532 21568 39668 21608
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 38572 20047 38612 20056
rect 39436 20096 39476 20105
rect 39532 20096 39572 21568
rect 39724 20852 39764 24340
rect 39819 23288 39861 23297
rect 39819 23248 39820 23288
rect 39860 23248 39861 23288
rect 39819 23239 39861 23248
rect 39820 23154 39860 23239
rect 39916 23060 39956 24751
rect 40108 23717 40148 25264
rect 40300 25220 40340 26104
rect 40396 26093 40436 26104
rect 40780 25901 40820 26683
rect 40876 26321 40916 26767
rect 40972 26648 41012 26657
rect 40972 26405 41012 26608
rect 40971 26396 41013 26405
rect 40971 26356 40972 26396
rect 41012 26356 41013 26396
rect 40971 26347 41013 26356
rect 40875 26312 40917 26321
rect 40875 26272 40876 26312
rect 40916 26272 40917 26312
rect 40875 26263 40917 26272
rect 40779 25892 40821 25901
rect 40779 25852 40780 25892
rect 40820 25852 40821 25892
rect 40779 25843 40821 25852
rect 40780 25556 40820 25843
rect 40780 25507 40820 25516
rect 40204 25180 40340 25220
rect 40588 25388 40628 25397
rect 40204 25132 40244 25180
rect 40588 25145 40628 25348
rect 40876 25304 40916 26263
rect 40972 25985 41012 26347
rect 41068 26237 41108 28867
rect 42507 28748 42549 28757
rect 42507 28708 42508 28748
rect 42548 28708 42549 28748
rect 42507 28699 42549 28708
rect 42028 28540 42452 28580
rect 41643 28412 41685 28421
rect 41643 28372 41644 28412
rect 41684 28372 41685 28412
rect 41643 28363 41685 28372
rect 41644 28328 41684 28363
rect 41547 27236 41589 27245
rect 41547 27196 41548 27236
rect 41588 27196 41589 27236
rect 41547 27187 41589 27196
rect 41451 26816 41493 26825
rect 41451 26776 41452 26816
rect 41492 26776 41493 26816
rect 41451 26767 41493 26776
rect 41067 26228 41109 26237
rect 41067 26188 41068 26228
rect 41108 26188 41109 26228
rect 41067 26179 41109 26188
rect 41260 26144 41300 26153
rect 40971 25976 41013 25985
rect 40971 25936 40972 25976
rect 41012 25936 41013 25976
rect 40971 25927 41013 25936
rect 40972 25304 41012 25313
rect 40876 25264 40972 25304
rect 40972 25255 41012 25264
rect 40779 25220 40821 25229
rect 40779 25180 40780 25220
rect 40820 25180 40821 25220
rect 40779 25171 40821 25180
rect 40204 25083 40244 25092
rect 40587 25136 40629 25145
rect 40587 25096 40588 25136
rect 40628 25096 40629 25136
rect 40587 25087 40629 25096
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 40492 23876 40532 23885
rect 40780 23876 40820 25171
rect 41067 25136 41109 25145
rect 41067 25096 41068 25136
rect 41108 25096 41109 25136
rect 41067 25087 41109 25096
rect 41068 25002 41108 25087
rect 40875 24884 40917 24893
rect 40875 24844 40876 24884
rect 40916 24844 40917 24884
rect 40875 24835 40917 24844
rect 40876 24800 40916 24835
rect 40876 24749 40916 24760
rect 41067 24716 41109 24725
rect 41067 24676 41068 24716
rect 41108 24676 41109 24716
rect 41067 24667 41109 24676
rect 41068 24582 41108 24667
rect 41260 24641 41300 26104
rect 41355 25388 41397 25397
rect 41355 25348 41356 25388
rect 41396 25348 41397 25388
rect 41355 25339 41397 25348
rect 41259 24632 41301 24641
rect 41259 24592 41260 24632
rect 41300 24592 41301 24632
rect 41259 24583 41301 24592
rect 40876 24380 40916 24389
rect 40876 23969 40916 24340
rect 41260 24053 41300 24583
rect 41259 24044 41301 24053
rect 41259 24004 41260 24044
rect 41300 24004 41301 24044
rect 41259 23995 41301 24004
rect 40875 23960 40917 23969
rect 40875 23920 40876 23960
rect 40916 23920 40917 23960
rect 40875 23911 40917 23920
rect 41067 23960 41109 23969
rect 41067 23920 41068 23960
rect 41108 23920 41109 23960
rect 41067 23911 41109 23920
rect 40532 23836 40820 23876
rect 40971 23876 41013 23885
rect 40971 23836 40972 23876
rect 41012 23836 41013 23876
rect 40492 23827 40532 23836
rect 40971 23827 41013 23836
rect 40876 23792 40916 23801
rect 40107 23708 40149 23717
rect 40107 23668 40108 23708
rect 40148 23668 40149 23708
rect 40107 23659 40149 23668
rect 40684 23624 40724 23633
rect 40876 23624 40916 23752
rect 40972 23708 41012 23827
rect 41068 23792 41108 23911
rect 41068 23743 41108 23752
rect 41164 23792 41204 23801
rect 40972 23659 41012 23668
rect 40724 23584 40916 23624
rect 40684 23575 40724 23584
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 40779 23372 40821 23381
rect 40779 23332 40780 23372
rect 40820 23332 40821 23372
rect 40779 23323 40821 23332
rect 40012 23129 40052 23214
rect 40011 23120 40053 23129
rect 40011 23080 40012 23120
rect 40052 23080 40053 23120
rect 40011 23071 40053 23080
rect 40396 23120 40436 23129
rect 40780 23120 40820 23323
rect 40436 23080 40820 23120
rect 40396 23071 40436 23080
rect 39820 23020 39956 23060
rect 39820 21953 39860 23020
rect 40011 22448 40053 22457
rect 40011 22408 40012 22448
rect 40052 22408 40053 22448
rect 40011 22399 40053 22408
rect 39819 21944 39861 21953
rect 39819 21904 39820 21944
rect 39860 21904 39861 21944
rect 39819 21895 39861 21904
rect 39820 21524 39860 21895
rect 40012 21608 40052 22399
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 40299 21692 40341 21701
rect 40299 21652 40300 21692
rect 40340 21652 40341 21692
rect 40299 21650 40341 21652
rect 40299 21643 40300 21650
rect 40012 21559 40052 21568
rect 40108 21608 40148 21617
rect 39820 21475 39860 21484
rect 40108 21449 40148 21568
rect 40340 21643 40341 21650
rect 40780 21617 40820 23080
rect 40876 23060 40916 23584
rect 41067 23624 41109 23633
rect 41067 23584 41068 23624
rect 41108 23584 41109 23624
rect 41067 23575 41109 23584
rect 40876 23045 41012 23060
rect 40876 23036 41013 23045
rect 40876 23020 40972 23036
rect 40876 22289 40916 23020
rect 40971 22996 40972 23020
rect 41012 22996 41013 23036
rect 40971 22987 41013 22996
rect 40972 22956 41012 22987
rect 40875 22280 40917 22289
rect 40875 22240 40876 22280
rect 40916 22240 40917 22280
rect 40875 22231 40917 22240
rect 40300 21557 40340 21610
rect 40779 21608 40821 21617
rect 40779 21568 40780 21608
rect 40820 21568 40821 21608
rect 40779 21559 40821 21568
rect 40107 21440 40149 21449
rect 40107 21400 40108 21440
rect 40148 21400 40149 21440
rect 40107 21391 40149 21400
rect 40300 21356 40340 21365
rect 40340 21316 40820 21356
rect 40300 21307 40340 21316
rect 40012 20852 40052 20861
rect 39724 20812 40012 20852
rect 40012 20803 40052 20812
rect 40587 20768 40629 20777
rect 40587 20728 40588 20768
rect 40628 20728 40629 20768
rect 40587 20719 40629 20728
rect 40204 20684 40244 20693
rect 39820 20600 39860 20609
rect 39860 20560 39956 20600
rect 39820 20551 39860 20560
rect 39820 20096 39860 20105
rect 39476 20056 39572 20096
rect 39628 20056 39820 20096
rect 39436 20047 39476 20056
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 38667 19592 38709 19601
rect 38667 19552 38668 19592
rect 38708 19552 38709 19592
rect 38667 19543 38709 19552
rect 38668 19340 38708 19543
rect 38859 19508 38901 19517
rect 38859 19468 38860 19508
rect 38900 19468 38901 19508
rect 38859 19459 38901 19468
rect 38860 19374 38900 19459
rect 39243 19424 39285 19433
rect 39243 19384 39244 19424
rect 39284 19384 39285 19424
rect 39243 19375 39285 19384
rect 39531 19424 39573 19433
rect 39531 19384 39532 19424
rect 39572 19384 39573 19424
rect 39531 19375 39573 19384
rect 39628 19424 39668 20056
rect 39820 20047 39860 20056
rect 39916 19685 39956 20560
rect 40204 20273 40244 20644
rect 40588 20634 40628 20719
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 40203 20264 40245 20273
rect 40203 20224 40204 20264
rect 40244 20224 40245 20264
rect 40203 20215 40245 20224
rect 40683 20264 40725 20273
rect 40683 20224 40684 20264
rect 40724 20224 40725 20264
rect 40683 20215 40725 20224
rect 40587 20180 40629 20189
rect 40587 20140 40588 20180
rect 40628 20140 40629 20180
rect 40587 20131 40629 20140
rect 40491 20096 40533 20105
rect 40491 20056 40492 20096
rect 40532 20056 40533 20096
rect 40491 20047 40533 20056
rect 40107 20012 40149 20021
rect 40107 19972 40108 20012
rect 40148 19972 40149 20012
rect 40107 19963 40149 19972
rect 40108 19878 40148 19963
rect 40492 19962 40532 20047
rect 40588 20012 40628 20131
rect 40588 19963 40628 19972
rect 40684 19928 40724 20215
rect 40780 20189 40820 21316
rect 40779 20180 40821 20189
rect 40779 20140 40780 20180
rect 40820 20140 40821 20180
rect 40779 20131 40821 20140
rect 40876 20096 40916 22231
rect 40971 21608 41013 21617
rect 40971 21568 40972 21608
rect 41012 21568 41013 21608
rect 40971 21559 41013 21568
rect 40972 20777 41012 21559
rect 40971 20768 41013 20777
rect 40971 20728 40972 20768
rect 41012 20728 41013 20768
rect 40971 20719 41013 20728
rect 40876 20047 40916 20056
rect 40779 20012 40821 20021
rect 40779 19972 40780 20012
rect 40820 19972 40821 20012
rect 40779 19963 40821 19972
rect 41068 20012 41108 23575
rect 41164 23297 41204 23752
rect 41163 23288 41205 23297
rect 41163 23248 41164 23288
rect 41204 23248 41205 23288
rect 41163 23239 41205 23248
rect 41260 23120 41300 23995
rect 41356 23633 41396 25339
rect 41452 24632 41492 26767
rect 41452 24137 41492 24592
rect 41451 24128 41493 24137
rect 41451 24088 41452 24128
rect 41492 24088 41493 24128
rect 41451 24079 41493 24088
rect 41451 23792 41493 23801
rect 41451 23752 41452 23792
rect 41492 23752 41493 23792
rect 41451 23743 41493 23752
rect 41452 23658 41492 23743
rect 41355 23624 41397 23633
rect 41355 23584 41356 23624
rect 41396 23584 41397 23624
rect 41355 23575 41397 23584
rect 41260 23060 41300 23080
rect 41260 23020 41396 23060
rect 41259 22616 41301 22625
rect 41259 22576 41260 22616
rect 41300 22576 41301 22616
rect 41259 22567 41301 22576
rect 41260 21449 41300 22567
rect 41259 21440 41301 21449
rect 41259 21400 41260 21440
rect 41300 21400 41301 21440
rect 41259 21391 41301 21400
rect 41163 21356 41205 21365
rect 41163 21316 41164 21356
rect 41204 21316 41205 21356
rect 41163 21307 41205 21316
rect 41068 19963 41108 19972
rect 40684 19879 40724 19888
rect 40780 19878 40820 19963
rect 40300 19844 40340 19853
rect 39915 19676 39957 19685
rect 39915 19636 39916 19676
rect 39956 19636 39957 19676
rect 39915 19627 39957 19636
rect 40300 19601 40340 19804
rect 41164 19676 41204 21307
rect 41356 20768 41396 23020
rect 41548 22625 41588 27187
rect 41644 26825 41684 28288
rect 42028 28328 42068 28540
rect 42412 28496 42452 28540
rect 42412 28447 42452 28456
rect 42315 28412 42357 28421
rect 42315 28372 42316 28412
rect 42356 28372 42357 28412
rect 42315 28363 42357 28372
rect 42508 28412 42548 28699
rect 42604 28496 42644 29128
rect 42700 29168 42740 29177
rect 42700 28673 42740 29128
rect 42795 29168 42837 29177
rect 42795 29128 42796 29168
rect 42836 29128 42837 29168
rect 42795 29119 42837 29128
rect 42892 29168 42932 29177
rect 42796 29034 42836 29119
rect 42892 28841 42932 29128
rect 43084 29168 43124 29177
rect 43276 29168 43316 29177
rect 42891 28832 42933 28841
rect 42891 28792 42892 28832
rect 42932 28792 42933 28832
rect 42891 28783 42933 28792
rect 42699 28664 42741 28673
rect 42699 28624 42700 28664
rect 42740 28624 42741 28664
rect 42699 28615 42741 28624
rect 43084 28589 43124 29128
rect 43180 29126 43220 29135
rect 43180 28757 43220 29086
rect 43179 28748 43221 28757
rect 43179 28708 43180 28748
rect 43220 28708 43221 28748
rect 43179 28699 43221 28708
rect 43276 28673 43316 29128
rect 43372 29168 43412 29177
rect 43275 28664 43317 28673
rect 43275 28624 43276 28664
rect 43316 28624 43317 28664
rect 43275 28615 43317 28624
rect 42795 28580 42837 28589
rect 42795 28540 42796 28580
rect 42836 28540 42837 28580
rect 42795 28531 42837 28540
rect 43083 28580 43125 28589
rect 43083 28540 43084 28580
rect 43124 28540 43125 28580
rect 43083 28531 43125 28540
rect 42604 28456 42740 28496
rect 42028 28279 42068 28288
rect 42220 28328 42260 28337
rect 42220 28160 42260 28288
rect 42316 28278 42356 28363
rect 42028 28120 42260 28160
rect 41835 26900 41877 26909
rect 41835 26860 41836 26900
rect 41876 26860 41877 26900
rect 41835 26851 41877 26860
rect 41643 26816 41685 26825
rect 41643 26776 41644 26816
rect 41684 26776 41685 26816
rect 41643 26767 41685 26776
rect 41739 25556 41781 25565
rect 41739 25516 41740 25556
rect 41780 25516 41781 25556
rect 41739 25507 41781 25516
rect 41740 25388 41780 25507
rect 41740 25339 41780 25348
rect 41836 24221 41876 26851
rect 41931 26060 41973 26069
rect 41931 26020 41932 26060
rect 41972 26020 41973 26060
rect 41931 26011 41973 26020
rect 41932 25556 41972 26011
rect 41932 25507 41972 25516
rect 42028 25229 42068 28120
rect 42220 28001 42260 28120
rect 42508 28085 42548 28372
rect 42604 28328 42644 28337
rect 42507 28076 42549 28085
rect 42507 28036 42508 28076
rect 42548 28036 42549 28076
rect 42507 28027 42549 28036
rect 42219 27992 42261 28001
rect 42219 27952 42220 27992
rect 42260 27952 42261 27992
rect 42219 27943 42261 27952
rect 42220 27824 42260 27833
rect 42508 27828 42548 27948
rect 42260 27788 42508 27824
rect 42604 27824 42644 28288
rect 42548 27788 42644 27824
rect 42260 27784 42644 27788
rect 42220 27775 42260 27784
rect 42508 27779 42548 27784
rect 42123 27656 42165 27665
rect 42123 27616 42124 27656
rect 42164 27616 42165 27656
rect 42123 27607 42165 27616
rect 42603 27656 42645 27665
rect 42603 27616 42604 27656
rect 42644 27616 42645 27656
rect 42603 27607 42645 27616
rect 42700 27656 42740 28456
rect 42796 28328 42836 28531
rect 43179 28496 43221 28505
rect 43179 28456 43180 28496
rect 43220 28456 43221 28496
rect 43179 28447 43221 28456
rect 43083 28412 43125 28421
rect 43083 28372 43084 28412
rect 43124 28372 43125 28412
rect 43083 28363 43125 28372
rect 43180 28364 43220 28447
rect 42796 28279 42836 28288
rect 42987 28076 43029 28085
rect 42987 28036 42988 28076
rect 43028 28036 43029 28076
rect 42987 28027 43029 28036
rect 42700 27607 42740 27616
rect 42124 27522 42164 27607
rect 42604 27522 42644 27607
rect 42988 27488 43028 28027
rect 43084 27488 43124 28363
rect 43180 28315 43220 28324
rect 43275 28328 43317 28337
rect 43275 28288 43276 28328
rect 43316 28288 43317 28328
rect 43275 28279 43317 28288
rect 43179 27992 43221 28001
rect 43179 27952 43180 27992
rect 43220 27952 43221 27992
rect 43179 27943 43221 27952
rect 43180 27698 43220 27943
rect 43180 27649 43220 27658
rect 43180 27488 43220 27497
rect 43084 27448 43180 27488
rect 42988 27439 43028 27448
rect 43180 27420 43220 27448
rect 42507 26816 42549 26825
rect 42507 26776 42508 26816
rect 42548 26776 42549 26816
rect 42507 26767 42549 26776
rect 43083 26816 43125 26825
rect 43083 26776 43084 26816
rect 43124 26776 43125 26816
rect 43276 26816 43316 28279
rect 43372 27833 43412 29128
rect 44139 29168 44181 29177
rect 44139 29128 44140 29168
rect 44180 29128 44181 29168
rect 44139 29119 44181 29128
rect 45387 29168 45429 29177
rect 45387 29128 45388 29168
rect 45428 29128 45429 29168
rect 45387 29119 45429 29128
rect 44043 28328 44085 28337
rect 44043 28288 44044 28328
rect 44084 28288 44085 28328
rect 44043 28279 44085 28288
rect 44044 28194 44084 28279
rect 43371 27824 43413 27833
rect 43371 27784 43372 27824
rect 43412 27784 43413 27824
rect 43371 27775 43413 27784
rect 43468 27784 43796 27824
rect 43372 27656 43412 27665
rect 43372 27329 43412 27616
rect 43468 27656 43508 27784
rect 43468 27607 43508 27616
rect 43659 27656 43701 27665
rect 43659 27616 43660 27656
rect 43700 27616 43701 27656
rect 43756 27656 43796 27784
rect 44140 27665 44180 29119
rect 46443 29084 46485 29093
rect 46443 29044 46444 29084
rect 46484 29044 46485 29084
rect 46443 29035 46485 29044
rect 45387 29000 45429 29009
rect 45387 28960 45388 29000
rect 45428 28960 45429 29000
rect 45387 28951 45429 28960
rect 44331 28664 44373 28673
rect 44331 28624 44332 28664
rect 44372 28624 44373 28664
rect 44331 28615 44373 28624
rect 44044 27656 44084 27665
rect 43756 27616 44044 27656
rect 43659 27607 43701 27616
rect 43660 27522 43700 27607
rect 43755 27488 43797 27497
rect 43755 27448 43756 27488
rect 43796 27448 43797 27488
rect 43755 27439 43797 27448
rect 43756 27354 43796 27439
rect 43948 27404 43988 27413
rect 43371 27320 43413 27329
rect 43371 27280 43372 27320
rect 43412 27280 43413 27320
rect 43371 27271 43413 27280
rect 43372 26993 43412 27271
rect 43371 26984 43413 26993
rect 43371 26944 43372 26984
rect 43412 26944 43413 26984
rect 43371 26935 43413 26944
rect 43372 26816 43412 26825
rect 43276 26776 43372 26816
rect 43083 26767 43125 26776
rect 43372 26767 43412 26776
rect 42124 26732 42164 26741
rect 42124 25985 42164 26692
rect 42508 26682 42548 26767
rect 43084 26564 43124 26767
rect 43084 26524 43220 26564
rect 42795 26480 42837 26489
rect 42795 26440 42796 26480
rect 42836 26440 42837 26480
rect 42795 26431 42837 26440
rect 42411 26312 42453 26321
rect 42411 26272 42412 26312
rect 42452 26272 42453 26312
rect 42411 26263 42453 26272
rect 42412 26178 42452 26263
rect 42796 26069 42836 26431
rect 42987 26312 43029 26321
rect 42987 26272 42988 26312
rect 43028 26272 43029 26312
rect 42987 26263 43029 26272
rect 42988 26144 43028 26263
rect 42892 26104 42988 26144
rect 42795 26060 42837 26069
rect 42795 26020 42796 26060
rect 42836 26020 42837 26060
rect 42795 26011 42837 26020
rect 42123 25976 42165 25985
rect 42123 25936 42124 25976
rect 42164 25936 42165 25976
rect 42123 25927 42165 25936
rect 42796 25926 42836 26011
rect 42604 25892 42644 25901
rect 42315 25556 42357 25565
rect 42315 25516 42316 25556
rect 42356 25516 42357 25556
rect 42315 25507 42357 25516
rect 42507 25556 42549 25565
rect 42507 25516 42508 25556
rect 42548 25516 42549 25556
rect 42507 25507 42549 25516
rect 42316 25422 42356 25507
rect 42123 25388 42165 25397
rect 42123 25348 42124 25388
rect 42164 25348 42165 25388
rect 42123 25339 42165 25348
rect 42508 25388 42548 25507
rect 42604 25397 42644 25852
rect 42795 25808 42837 25817
rect 42795 25768 42796 25808
rect 42836 25768 42837 25808
rect 42795 25759 42837 25768
rect 42508 25339 42548 25348
rect 42603 25388 42645 25397
rect 42603 25348 42604 25388
rect 42644 25348 42645 25388
rect 42603 25339 42645 25348
rect 42124 25254 42164 25339
rect 42796 25313 42836 25759
rect 42795 25304 42837 25313
rect 42795 25264 42796 25304
rect 42836 25264 42837 25304
rect 42795 25255 42837 25264
rect 42027 25220 42069 25229
rect 42027 25180 42028 25220
rect 42068 25180 42069 25220
rect 42027 25171 42069 25180
rect 42699 25220 42741 25229
rect 42699 25180 42700 25220
rect 42740 25180 42741 25220
rect 42699 25171 42741 25180
rect 42700 25136 42740 25171
rect 42700 25085 42740 25096
rect 42892 24884 42932 26104
rect 42988 26095 43028 26104
rect 43084 26228 43124 26237
rect 43084 26069 43124 26188
rect 43180 26186 43220 26524
rect 43467 26312 43509 26321
rect 43467 26272 43468 26312
rect 43508 26272 43509 26312
rect 43467 26263 43509 26272
rect 43659 26312 43701 26321
rect 43659 26272 43660 26312
rect 43700 26272 43701 26312
rect 43659 26263 43701 26272
rect 43948 26312 43988 27364
rect 44044 27068 44084 27616
rect 44139 27656 44181 27665
rect 44139 27616 44140 27656
rect 44180 27616 44181 27656
rect 44139 27607 44181 27616
rect 44235 27572 44277 27581
rect 44235 27532 44236 27572
rect 44276 27532 44277 27572
rect 44235 27523 44277 27532
rect 44236 27438 44276 27523
rect 44332 27497 44372 28615
rect 45195 28580 45237 28589
rect 45195 28540 45196 28580
rect 45236 28540 45237 28580
rect 45195 28531 45237 28540
rect 45196 28446 45236 28531
rect 45388 28328 45428 28951
rect 45388 28279 45428 28288
rect 45772 28328 45812 28337
rect 46155 28328 46197 28337
rect 45812 28288 46100 28328
rect 45772 28279 45812 28288
rect 44907 28244 44949 28253
rect 44907 28204 44908 28244
rect 44948 28204 44949 28244
rect 44907 28195 44949 28204
rect 44331 27488 44373 27497
rect 44331 27448 44332 27488
rect 44372 27448 44373 27488
rect 44331 27439 44373 27448
rect 44908 27413 44948 28195
rect 45196 28160 45236 28169
rect 45196 27665 45236 28120
rect 46060 27824 46100 28288
rect 46155 28288 46156 28328
rect 46196 28288 46197 28328
rect 46155 28279 46197 28288
rect 46060 27775 46100 27784
rect 45195 27656 45237 27665
rect 45195 27616 45196 27656
rect 45236 27616 45237 27656
rect 45195 27607 45237 27616
rect 45868 27572 45908 27581
rect 44427 27404 44469 27413
rect 44427 27364 44428 27404
rect 44468 27364 44469 27404
rect 44427 27355 44469 27364
rect 44907 27404 44949 27413
rect 44907 27364 44908 27404
rect 44948 27364 44949 27404
rect 44907 27355 44949 27364
rect 44428 27270 44468 27355
rect 44524 27068 44564 27077
rect 44044 27028 44524 27068
rect 44524 27019 44564 27028
rect 44908 26900 44948 27355
rect 44908 26851 44948 26860
rect 44716 26648 44756 26657
rect 44716 26564 44756 26608
rect 44716 26524 44948 26564
rect 44715 26396 44757 26405
rect 44715 26356 44716 26396
rect 44756 26356 44757 26396
rect 44715 26347 44757 26356
rect 44140 26316 44180 26325
rect 43948 26276 44140 26312
rect 43948 26272 44180 26276
rect 43083 26060 43125 26069
rect 43083 26020 43084 26060
rect 43124 26020 43125 26060
rect 43083 26011 43125 26020
rect 43180 25724 43220 26146
rect 43276 26144 43316 26153
rect 43468 26144 43508 26263
rect 43660 26153 43700 26263
rect 43316 26104 43412 26144
rect 43276 26095 43316 26104
rect 42604 24844 42932 24884
rect 42988 25684 43220 25724
rect 42316 24641 42356 24726
rect 42315 24632 42357 24641
rect 42315 24592 42316 24632
rect 42356 24592 42357 24632
rect 42315 24583 42357 24592
rect 41835 24212 41877 24221
rect 41835 24172 41836 24212
rect 41876 24172 41877 24212
rect 41835 24163 41877 24172
rect 41643 24128 41685 24137
rect 41643 24088 41644 24128
rect 41684 24088 41685 24128
rect 41643 24079 41685 24088
rect 41644 23381 41684 24079
rect 41739 24044 41781 24053
rect 41739 24004 41740 24044
rect 41780 24004 41781 24044
rect 41739 23995 41781 24004
rect 41740 23910 41780 23995
rect 42604 23792 42644 24844
rect 42795 24716 42837 24725
rect 42795 24676 42796 24716
rect 42836 24676 42837 24716
rect 42795 24667 42837 24676
rect 42796 23960 42836 24667
rect 42988 23960 43028 25684
rect 43275 25472 43317 25481
rect 43275 25432 43276 25472
rect 43316 25432 43317 25472
rect 43275 25423 43317 25432
rect 43084 25388 43124 25399
rect 43084 25313 43124 25348
rect 43276 25338 43316 25423
rect 43083 25304 43125 25313
rect 43083 25264 43084 25304
rect 43124 25264 43125 25304
rect 43083 25255 43125 25264
rect 43372 24800 43412 26104
rect 43468 26095 43508 26104
rect 43659 26144 43701 26153
rect 43659 26104 43660 26144
rect 43700 26104 43701 26144
rect 43659 26095 43701 26104
rect 43852 26144 43892 26153
rect 43948 26144 43988 26272
rect 44140 26267 44180 26272
rect 43892 26104 43988 26144
rect 44043 26144 44085 26153
rect 44236 26144 44276 26153
rect 44043 26104 44044 26144
rect 44084 26104 44085 26144
rect 43852 26095 43892 26104
rect 44043 26095 44085 26104
rect 44140 26104 44236 26144
rect 43563 26060 43605 26069
rect 43563 26020 43564 26060
rect 43604 26020 43605 26060
rect 43563 26011 43605 26020
rect 43755 26060 43797 26069
rect 43755 26020 43756 26060
rect 43796 26020 43797 26060
rect 43755 26011 43797 26020
rect 43564 25926 43604 26011
rect 43659 25976 43701 25985
rect 43659 25936 43660 25976
rect 43700 25936 43701 25976
rect 43659 25927 43701 25936
rect 43660 25842 43700 25927
rect 43756 25926 43796 26011
rect 43563 25640 43605 25649
rect 43563 25600 43564 25640
rect 43604 25600 43605 25640
rect 43563 25591 43605 25600
rect 43467 25472 43509 25481
rect 43467 25432 43468 25472
rect 43508 25432 43509 25472
rect 43564 25472 43604 25591
rect 43660 25472 43700 25481
rect 43564 25432 43660 25472
rect 43700 25432 43892 25472
rect 43467 25423 43509 25432
rect 43660 25423 43700 25432
rect 43468 25388 43508 25423
rect 43468 25337 43508 25348
rect 43852 25388 43892 25432
rect 43852 25339 43892 25348
rect 44044 25304 44084 26095
rect 43948 25264 44084 25304
rect 43468 24800 43508 24809
rect 43372 24760 43468 24800
rect 43083 23960 43125 23969
rect 42988 23920 43084 23960
rect 43124 23920 43125 23960
rect 42796 23911 42836 23920
rect 43083 23911 43125 23920
rect 42699 23876 42741 23885
rect 42699 23836 42700 23876
rect 42740 23836 42741 23876
rect 42699 23827 42741 23836
rect 42892 23876 42932 23885
rect 42508 23752 42604 23792
rect 41643 23372 41685 23381
rect 41643 23332 41644 23372
rect 41684 23332 41685 23372
rect 41643 23323 41685 23332
rect 42411 23288 42453 23297
rect 42411 23248 42412 23288
rect 42452 23248 42453 23288
rect 42411 23239 42453 23248
rect 42412 23154 42452 23239
rect 41643 23120 41685 23129
rect 41643 23080 41644 23120
rect 41684 23080 41685 23120
rect 41643 23071 41685 23080
rect 41547 22616 41589 22625
rect 41547 22576 41548 22616
rect 41588 22576 41589 22616
rect 41547 22567 41589 22576
rect 41547 22448 41589 22457
rect 41547 22408 41548 22448
rect 41588 22408 41589 22448
rect 41547 22399 41589 22408
rect 41644 22448 41684 23071
rect 42508 23045 42548 23752
rect 42604 23743 42644 23752
rect 42700 23742 42740 23827
rect 42795 23792 42837 23801
rect 42795 23752 42796 23792
rect 42836 23752 42837 23792
rect 42795 23743 42837 23752
rect 42699 23540 42741 23549
rect 42699 23500 42700 23540
rect 42740 23500 42741 23540
rect 42699 23491 42741 23500
rect 42604 23120 42644 23129
rect 42507 23036 42549 23045
rect 42507 22996 42508 23036
rect 42548 22996 42549 23036
rect 42507 22987 42549 22996
rect 42411 22952 42453 22961
rect 42411 22912 42412 22952
rect 42452 22912 42453 22952
rect 42411 22903 42453 22912
rect 41644 22399 41684 22408
rect 41740 22576 42068 22616
rect 41548 22364 41588 22399
rect 41548 22313 41588 22324
rect 41740 22364 41780 22576
rect 42028 22574 42068 22576
rect 42028 22525 42068 22534
rect 41451 22280 41493 22289
rect 41451 22240 41452 22280
rect 41492 22240 41493 22280
rect 41451 22231 41493 22240
rect 41452 22146 41492 22231
rect 41740 21701 41780 22324
rect 41836 22289 41876 22374
rect 41835 22280 41877 22289
rect 41835 22240 41836 22280
rect 41876 22240 41877 22280
rect 41835 22231 41877 22240
rect 42316 22280 42356 22289
rect 42316 22121 42356 22240
rect 42412 22280 42452 22903
rect 42507 22868 42549 22877
rect 42507 22828 42508 22868
rect 42548 22828 42549 22868
rect 42507 22819 42549 22828
rect 42508 22289 42548 22819
rect 42412 22205 42452 22240
rect 42507 22280 42549 22289
rect 42507 22240 42508 22280
rect 42548 22240 42549 22280
rect 42507 22231 42549 22240
rect 42411 22196 42453 22205
rect 42411 22156 42412 22196
rect 42452 22156 42453 22196
rect 42411 22147 42453 22156
rect 42315 22112 42357 22121
rect 42315 22072 42316 22112
rect 42356 22072 42357 22112
rect 42315 22063 42357 22072
rect 42508 22108 42548 22231
rect 42604 22121 42644 23080
rect 42700 23120 42740 23491
rect 42796 23456 42836 23743
rect 42892 23633 42932 23836
rect 42987 23792 43029 23801
rect 42987 23752 42988 23792
rect 43028 23752 43029 23792
rect 42987 23743 43029 23752
rect 42988 23658 43028 23743
rect 42891 23624 42933 23633
rect 42891 23584 42892 23624
rect 42932 23584 42933 23624
rect 42891 23575 42933 23584
rect 43084 23540 43124 23911
rect 43275 23792 43317 23801
rect 43275 23752 43276 23792
rect 43316 23752 43317 23792
rect 43275 23743 43317 23752
rect 43084 23500 43220 23540
rect 42796 23416 42932 23456
rect 42795 23288 42837 23297
rect 42795 23248 42796 23288
rect 42836 23248 42837 23288
rect 42795 23239 42837 23248
rect 42796 23141 42836 23239
rect 42796 23092 42836 23101
rect 42892 23120 42932 23416
rect 43083 23372 43125 23381
rect 43083 23332 43084 23372
rect 43124 23332 43125 23372
rect 43083 23323 43125 23332
rect 42987 23288 43029 23297
rect 42987 23248 42988 23288
rect 43028 23248 43029 23288
rect 42987 23239 43029 23248
rect 42988 23129 43028 23239
rect 42508 22059 42548 22068
rect 42603 22112 42645 22121
rect 42603 22072 42604 22112
rect 42644 22072 42645 22112
rect 42700 22112 42740 23080
rect 42795 23036 42837 23045
rect 42795 22996 42796 23036
rect 42836 22996 42837 23036
rect 42795 22987 42837 22996
rect 42796 22280 42836 22987
rect 42892 22961 42932 23080
rect 42987 23120 43029 23129
rect 42987 23080 42988 23120
rect 43028 23080 43029 23120
rect 42987 23071 43029 23080
rect 43084 23120 43124 23323
rect 43180 23129 43220 23500
rect 43276 23288 43316 23743
rect 43372 23708 43412 24760
rect 43468 24751 43508 24760
rect 43660 24632 43700 24641
rect 43948 24632 43988 25264
rect 44140 25145 44180 26104
rect 44236 26095 44276 26104
rect 44332 26144 44372 26153
rect 44332 25985 44372 26104
rect 44427 26144 44469 26153
rect 44427 26104 44428 26144
rect 44468 26104 44469 26144
rect 44427 26095 44469 26104
rect 44331 25976 44373 25985
rect 44331 25936 44332 25976
rect 44372 25936 44373 25976
rect 44331 25927 44373 25936
rect 44428 25304 44468 26095
rect 44523 26060 44565 26069
rect 44523 26020 44524 26060
rect 44564 26020 44565 26060
rect 44523 26011 44565 26020
rect 44428 25255 44468 25264
rect 44524 25892 44564 26011
rect 44620 25892 44660 25901
rect 44524 25852 44620 25892
rect 44524 25304 44564 25852
rect 44620 25843 44660 25852
rect 44524 25255 44564 25264
rect 44620 25304 44660 25315
rect 44620 25229 44660 25264
rect 44716 25304 44756 26347
rect 44811 26144 44853 26153
rect 44811 26104 44812 26144
rect 44852 26104 44853 26144
rect 44811 26095 44853 26104
rect 44812 26010 44852 26095
rect 44908 25901 44948 26524
rect 45771 26396 45813 26405
rect 45771 26356 45772 26396
rect 45812 26356 45813 26396
rect 45771 26347 45813 26356
rect 45195 26312 45237 26321
rect 45387 26312 45429 26321
rect 45195 26272 45196 26312
rect 45236 26272 45237 26312
rect 45195 26263 45237 26272
rect 45292 26272 45388 26312
rect 45428 26272 45429 26312
rect 45196 26153 45236 26263
rect 45195 26144 45237 26153
rect 45195 26104 45196 26144
rect 45236 26104 45237 26144
rect 45195 26095 45237 26104
rect 45195 25976 45237 25985
rect 45195 25936 45196 25976
rect 45236 25936 45237 25976
rect 45195 25927 45237 25936
rect 44907 25892 44949 25901
rect 44907 25852 44908 25892
rect 44948 25852 44949 25892
rect 44907 25843 44949 25852
rect 44908 25649 44948 25843
rect 44907 25640 44949 25649
rect 44907 25600 44908 25640
rect 44948 25600 44949 25640
rect 44907 25591 44949 25600
rect 44716 25255 44756 25264
rect 44908 25304 44948 25313
rect 44619 25220 44661 25229
rect 44619 25180 44620 25220
rect 44660 25180 44661 25220
rect 44619 25171 44661 25180
rect 44908 25145 44948 25264
rect 45003 25304 45045 25313
rect 45003 25264 45004 25304
rect 45044 25264 45045 25304
rect 45003 25255 45045 25264
rect 45100 25304 45140 25313
rect 45004 25170 45044 25255
rect 44044 25136 44084 25145
rect 44139 25136 44181 25145
rect 44084 25096 44140 25136
rect 44180 25096 44181 25136
rect 44044 25087 44084 25096
rect 44139 25087 44181 25096
rect 44907 25136 44949 25145
rect 44907 25096 44908 25136
rect 44948 25096 44949 25136
rect 44907 25087 44949 25096
rect 45100 25132 45140 25264
rect 45196 25304 45236 25927
rect 45196 25255 45236 25264
rect 45100 25092 45236 25132
rect 44044 24632 44084 24641
rect 43948 24592 44044 24632
rect 43468 23885 43508 23930
rect 43467 23876 43509 23885
rect 43467 23836 43468 23876
rect 43508 23836 43509 23876
rect 43467 23835 43509 23836
rect 43467 23827 43468 23835
rect 43508 23827 43509 23835
rect 43468 23786 43508 23795
rect 43563 23792 43605 23801
rect 43563 23752 43564 23792
rect 43604 23752 43605 23792
rect 43563 23743 43605 23752
rect 43372 23668 43508 23708
rect 43372 23566 43412 23575
rect 43372 23288 43412 23526
rect 43276 23248 43372 23288
rect 43372 23239 43412 23248
rect 43084 23071 43124 23080
rect 43179 23120 43221 23129
rect 43179 23080 43180 23120
rect 43220 23080 43221 23120
rect 43179 23071 43221 23080
rect 43468 23120 43508 23668
rect 43564 23658 43604 23743
rect 43660 23288 43700 24592
rect 44044 24583 44084 24592
rect 44140 23969 44180 25087
rect 45196 24977 45236 25092
rect 45195 24968 45237 24977
rect 45195 24928 45196 24968
rect 45236 24928 45237 24968
rect 45195 24919 45237 24928
rect 44907 24632 44949 24641
rect 44907 24592 44908 24632
rect 44948 24592 44949 24632
rect 44907 24583 44949 24592
rect 45099 24632 45141 24641
rect 45099 24592 45100 24632
rect 45140 24592 45141 24632
rect 45099 24583 45141 24592
rect 44908 24498 44948 24583
rect 44331 24380 44373 24389
rect 44331 24340 44332 24380
rect 44372 24340 44373 24380
rect 44331 24331 44373 24340
rect 44907 24380 44949 24389
rect 44907 24340 44908 24380
rect 44948 24340 44949 24380
rect 44907 24331 44949 24340
rect 43852 23960 43892 23969
rect 44139 23960 44181 23969
rect 43892 23920 43988 23960
rect 43852 23911 43892 23920
rect 43852 23633 43892 23652
rect 43851 23624 43893 23633
rect 43948 23624 43988 23920
rect 44139 23920 44140 23960
rect 44180 23920 44181 23960
rect 44139 23911 44181 23920
rect 44139 23792 44181 23801
rect 44139 23752 44140 23792
rect 44180 23752 44181 23792
rect 44139 23743 44181 23752
rect 44236 23792 44276 23801
rect 44140 23658 44180 23743
rect 43851 23584 43852 23624
rect 43892 23584 43988 23624
rect 43851 23575 43893 23584
rect 43852 23288 43892 23297
rect 43660 23248 43852 23288
rect 43852 23239 43892 23248
rect 43468 23071 43508 23080
rect 43948 23120 43988 23584
rect 44043 23624 44085 23633
rect 44043 23584 44044 23624
rect 44084 23584 44085 23624
rect 44043 23575 44085 23584
rect 43948 23071 43988 23080
rect 44044 23120 44084 23575
rect 44236 23549 44276 23752
rect 44332 23792 44372 24331
rect 44427 23876 44469 23885
rect 44427 23836 44428 23876
rect 44468 23836 44469 23876
rect 44427 23827 44469 23836
rect 44332 23743 44372 23752
rect 44428 23792 44468 23827
rect 44428 23741 44468 23752
rect 44235 23540 44277 23549
rect 44044 23071 44084 23080
rect 44140 23500 44236 23540
rect 44276 23500 44277 23540
rect 44140 23120 44180 23500
rect 44235 23491 44277 23500
rect 44140 23071 44180 23080
rect 44908 23120 44948 24331
rect 45003 23624 45045 23633
rect 45003 23584 45004 23624
rect 45044 23584 45045 23624
rect 45003 23575 45045 23584
rect 45004 23288 45044 23575
rect 45004 23239 45044 23248
rect 44908 23071 44948 23080
rect 45100 23060 45140 24583
rect 45196 24557 45236 24919
rect 45195 24548 45237 24557
rect 45195 24508 45196 24548
rect 45236 24508 45237 24548
rect 45195 24499 45237 24508
rect 45004 23020 45140 23060
rect 42891 22952 42933 22961
rect 42891 22912 42892 22952
rect 42932 22912 42933 22952
rect 42891 22903 42933 22912
rect 43083 22952 43125 22961
rect 43083 22912 43084 22952
rect 43124 22912 43125 22952
rect 43083 22903 43125 22912
rect 43371 22952 43413 22961
rect 43371 22912 43372 22952
rect 43412 22912 43413 22952
rect 43371 22903 43413 22912
rect 42892 22457 42932 22542
rect 42891 22448 42933 22457
rect 42891 22408 42892 22448
rect 42932 22408 42933 22448
rect 42891 22399 42933 22408
rect 42892 22280 42932 22289
rect 42796 22240 42892 22280
rect 42700 22072 42836 22112
rect 42603 22063 42645 22072
rect 42123 21776 42165 21785
rect 42123 21736 42124 21776
rect 42164 21736 42165 21776
rect 42123 21727 42165 21736
rect 42603 21776 42645 21785
rect 42603 21736 42604 21776
rect 42644 21736 42645 21776
rect 42603 21727 42645 21736
rect 41739 21692 41781 21701
rect 41739 21652 41740 21692
rect 41780 21652 41781 21692
rect 41739 21643 41781 21652
rect 42124 21642 42164 21727
rect 42604 21692 42644 21727
rect 42604 21641 42644 21652
rect 42796 21617 42836 22072
rect 42892 21785 42932 22240
rect 43084 22280 43124 22903
rect 43179 22868 43221 22877
rect 43179 22828 43180 22868
rect 43220 22828 43221 22868
rect 43179 22819 43221 22828
rect 43180 22734 43220 22819
rect 43372 22289 43412 22903
rect 43467 22532 43509 22541
rect 43467 22492 43468 22532
rect 43508 22492 43509 22532
rect 43467 22483 43509 22492
rect 43468 22398 43508 22483
rect 42891 21776 42933 21785
rect 42891 21736 42892 21776
rect 42932 21736 42933 21776
rect 42891 21727 42933 21736
rect 43084 21617 43124 22240
rect 43198 22273 43238 22282
rect 43198 22121 43238 22233
rect 43371 22280 43413 22289
rect 43371 22240 43372 22280
rect 43412 22240 43413 22280
rect 43371 22231 43413 22240
rect 45004 22280 45044 23020
rect 45292 22289 45332 26272
rect 45387 26263 45429 26272
rect 45387 25892 45429 25901
rect 45387 25852 45388 25892
rect 45428 25852 45429 25892
rect 45387 25843 45429 25852
rect 45388 25061 45428 25843
rect 45772 25808 45812 26347
rect 45868 26153 45908 27532
rect 46060 27404 46100 27413
rect 45964 27364 46060 27404
rect 45867 26144 45909 26153
rect 45867 26104 45868 26144
rect 45908 26104 45909 26144
rect 45867 26095 45909 26104
rect 45964 25985 46004 27364
rect 46060 27355 46100 27364
rect 46060 26144 46100 26153
rect 46156 26144 46196 28279
rect 46100 26104 46196 26144
rect 46060 26095 46100 26104
rect 45963 25976 46005 25985
rect 45963 25936 45964 25976
rect 46004 25936 46005 25976
rect 45963 25927 46005 25936
rect 45772 25768 46004 25808
rect 45483 25640 45525 25649
rect 45483 25600 45484 25640
rect 45524 25600 45525 25640
rect 45483 25591 45525 25600
rect 45675 25640 45717 25649
rect 45675 25600 45676 25640
rect 45716 25600 45717 25640
rect 45675 25591 45717 25600
rect 45484 25145 45524 25591
rect 45676 25313 45716 25591
rect 45675 25304 45717 25313
rect 45675 25264 45676 25304
rect 45716 25264 45717 25304
rect 45675 25255 45717 25264
rect 45579 25220 45621 25229
rect 45579 25180 45580 25220
rect 45620 25180 45621 25220
rect 45579 25171 45621 25180
rect 45483 25136 45525 25145
rect 45483 25096 45484 25136
rect 45524 25096 45525 25136
rect 45483 25087 45525 25096
rect 45580 25086 45620 25171
rect 45676 25170 45716 25255
rect 45387 25052 45429 25061
rect 45387 25012 45388 25052
rect 45428 25012 45429 25052
rect 45387 25003 45429 25012
rect 43372 22146 43412 22231
rect 43852 22121 43892 22206
rect 43197 22112 43239 22121
rect 43197 22072 43198 22112
rect 43238 22072 43239 22112
rect 43197 22063 43239 22072
rect 43851 22112 43893 22121
rect 43851 22072 43852 22112
rect 43892 22072 43893 22112
rect 43851 22063 43893 22072
rect 45004 21953 45044 22240
rect 45291 22280 45333 22289
rect 45291 22240 45292 22280
rect 45332 22240 45333 22280
rect 45291 22231 45333 22240
rect 43851 21944 43893 21953
rect 43851 21904 43852 21944
rect 43892 21904 43893 21944
rect 43851 21895 43893 21904
rect 45003 21944 45045 21953
rect 45003 21904 45004 21944
rect 45044 21904 45045 21944
rect 45003 21895 45045 21904
rect 42219 21608 42261 21617
rect 42219 21568 42220 21608
rect 42260 21568 42261 21608
rect 42219 21559 42261 21568
rect 42316 21608 42356 21617
rect 42220 21474 42260 21559
rect 42316 21449 42356 21568
rect 42411 21608 42453 21617
rect 42411 21568 42412 21608
rect 42452 21568 42453 21608
rect 42411 21559 42453 21568
rect 42795 21608 42837 21617
rect 42795 21568 42796 21608
rect 42836 21568 42837 21608
rect 42795 21559 42837 21568
rect 42988 21608 43028 21617
rect 42315 21440 42357 21449
rect 42315 21400 42316 21440
rect 42356 21400 42357 21440
rect 42315 21391 42357 21400
rect 42412 21104 42452 21559
rect 42220 21064 42452 21104
rect 41452 20768 41492 20777
rect 41356 20728 41452 20768
rect 41452 20719 41492 20728
rect 41739 20432 41781 20441
rect 41739 20392 41740 20432
rect 41780 20392 41781 20432
rect 41739 20383 41781 20392
rect 41740 20264 41780 20383
rect 42220 20273 42260 21064
rect 42604 20852 42644 20861
rect 42644 20812 42932 20852
rect 42604 20803 42644 20812
rect 42892 20768 42932 20812
rect 42988 20777 43028 21568
rect 43083 21608 43125 21617
rect 43083 21568 43084 21608
rect 43124 21568 43125 21608
rect 43083 21559 43125 21568
rect 43659 21608 43701 21617
rect 43659 21568 43660 21608
rect 43700 21568 43701 21608
rect 43659 21559 43701 21568
rect 43852 21608 43892 21895
rect 44235 21776 44277 21785
rect 44235 21736 44236 21776
rect 44276 21736 44277 21776
rect 44235 21727 44277 21736
rect 45004 21776 45044 21785
rect 45292 21776 45332 22231
rect 45044 21736 45332 21776
rect 45004 21727 45044 21736
rect 43852 21559 43892 21568
rect 43660 21020 43700 21559
rect 43660 20971 43700 20980
rect 43851 20852 43893 20861
rect 43851 20812 43852 20852
rect 43892 20812 43893 20852
rect 43851 20803 43893 20812
rect 42796 20600 42836 20609
rect 42700 20560 42796 20600
rect 42412 20273 42452 20359
rect 42700 20273 42740 20560
rect 42796 20551 42836 20560
rect 41740 20215 41780 20224
rect 42219 20264 42261 20273
rect 42219 20224 42220 20264
rect 42260 20224 42261 20264
rect 42219 20215 42261 20224
rect 42411 20268 42453 20273
rect 42411 20224 42412 20268
rect 42452 20224 42453 20268
rect 42411 20215 42453 20224
rect 42699 20264 42741 20273
rect 42699 20224 42700 20264
rect 42740 20224 42741 20264
rect 42699 20215 42741 20224
rect 41355 20180 41397 20189
rect 41355 20140 41356 20180
rect 41396 20140 41397 20180
rect 41355 20131 41397 20140
rect 42795 20180 42837 20189
rect 42795 20140 42796 20180
rect 42836 20140 42837 20180
rect 42795 20131 42837 20140
rect 41356 20012 41396 20131
rect 41644 20117 41684 20126
rect 41684 20096 41876 20117
rect 42220 20096 42260 20105
rect 41684 20077 41972 20096
rect 41644 20068 41684 20077
rect 41452 20051 41492 20060
rect 41356 20011 41452 20012
rect 41356 19972 41492 20011
rect 41068 19636 41204 19676
rect 41260 19844 41300 19853
rect 40299 19592 40341 19601
rect 40299 19552 40300 19592
rect 40340 19552 40341 19592
rect 40299 19543 40341 19552
rect 40012 19424 40052 19433
rect 40300 19424 40340 19543
rect 40395 19508 40437 19517
rect 40395 19468 40396 19508
rect 40436 19468 40437 19508
rect 40395 19459 40437 19468
rect 40971 19508 41013 19517
rect 40971 19468 40972 19508
rect 41012 19468 41013 19508
rect 40971 19459 41013 19468
rect 39628 19375 39668 19384
rect 39724 19384 40012 19424
rect 38668 19291 38708 19300
rect 39052 19340 39092 19349
rect 38092 19122 38132 19207
rect 38284 19181 38324 19216
rect 38380 19256 38420 19265
rect 38283 19172 38325 19181
rect 38283 19132 38284 19172
rect 38324 19132 38325 19172
rect 38283 19123 38325 19132
rect 38380 19013 38420 19216
rect 39052 19181 39092 19300
rect 39244 19290 39284 19375
rect 39532 19340 39572 19375
rect 39532 19289 39572 19300
rect 39724 19340 39764 19384
rect 40012 19375 40052 19384
rect 40204 19384 40340 19424
rect 39435 19256 39477 19265
rect 39435 19216 39436 19256
rect 39476 19216 39477 19256
rect 39435 19207 39477 19216
rect 38763 19172 38805 19181
rect 38763 19132 38764 19172
rect 38804 19132 38805 19172
rect 38763 19123 38805 19132
rect 39051 19172 39093 19181
rect 39051 19132 39052 19172
rect 39092 19132 39093 19172
rect 39051 19123 39093 19132
rect 38379 19004 38421 19013
rect 38379 18964 38380 19004
rect 38420 18964 38421 19004
rect 38379 18955 38421 18964
rect 38187 18920 38229 18929
rect 38187 18880 38188 18920
rect 38228 18880 38229 18920
rect 38187 18871 38229 18880
rect 38188 18584 38228 18871
rect 38188 18535 38228 18544
rect 38187 18248 38229 18257
rect 38187 18208 38188 18248
rect 38228 18208 38229 18248
rect 38187 18199 38229 18208
rect 38188 17753 38228 18199
rect 38187 17744 38229 17753
rect 38187 17704 38188 17744
rect 38228 17704 38229 17744
rect 38187 17695 38229 17704
rect 38188 17610 38228 17695
rect 38283 17576 38325 17585
rect 38283 17536 38284 17576
rect 38324 17536 38325 17576
rect 38283 17527 38325 17536
rect 38284 17442 38324 17527
rect 38379 17324 38421 17333
rect 38379 17284 38380 17324
rect 38420 17284 38421 17324
rect 38379 17275 38421 17284
rect 37995 16988 38037 16997
rect 37995 16948 37996 16988
rect 38036 16948 38037 16988
rect 37995 16939 38037 16948
rect 37996 16854 38036 16939
rect 37899 16652 37941 16661
rect 37899 16612 37900 16652
rect 37940 16612 37941 16652
rect 37899 16603 37941 16612
rect 37899 16316 37941 16325
rect 37899 16276 37900 16316
rect 37940 16276 37941 16316
rect 37899 16267 37941 16276
rect 37804 16183 37844 16192
rect 37900 16232 37940 16267
rect 37900 16181 37940 16192
rect 38091 16148 38133 16157
rect 38091 16108 38092 16148
rect 38132 16108 38133 16148
rect 38091 16099 38133 16108
rect 38092 16014 38132 16099
rect 38380 16064 38420 17275
rect 38571 17072 38613 17081
rect 38571 17032 38572 17072
rect 38612 17032 38613 17072
rect 38571 17023 38613 17032
rect 38475 16652 38517 16661
rect 38475 16612 38476 16652
rect 38516 16612 38517 16652
rect 38475 16603 38517 16612
rect 38476 16232 38516 16603
rect 38476 16183 38516 16192
rect 38380 16024 38516 16064
rect 38091 15812 38133 15821
rect 38091 15772 38092 15812
rect 38132 15772 38133 15812
rect 38091 15763 38133 15772
rect 37995 15644 38037 15653
rect 37995 15604 37996 15644
rect 38036 15604 38037 15644
rect 37995 15595 38037 15604
rect 37899 15560 37941 15569
rect 37899 15520 37900 15560
rect 37940 15520 37941 15560
rect 37899 15511 37941 15520
rect 37996 15560 38036 15595
rect 36980 15268 37172 15308
rect 36940 15259 36980 15268
rect 36844 15100 37076 15140
rect 36844 14972 36884 14981
rect 36652 14932 36844 14972
rect 36844 14923 36884 14932
rect 35692 14671 35732 14680
rect 37036 14720 37076 15100
rect 37132 14804 37172 15268
rect 37132 14755 37172 14764
rect 37228 14888 37268 14897
rect 37036 14645 37076 14680
rect 37035 14636 37077 14645
rect 37035 14596 37036 14636
rect 37076 14596 37077 14636
rect 37035 14587 37077 14596
rect 37036 14556 37076 14587
rect 37228 14468 37268 14848
rect 37708 14813 37748 15268
rect 37323 14804 37365 14813
rect 37323 14764 37324 14804
rect 37364 14764 37365 14804
rect 37323 14755 37365 14764
rect 37707 14804 37749 14813
rect 37707 14764 37708 14804
rect 37748 14764 37749 14804
rect 37707 14755 37749 14764
rect 37324 14670 37364 14755
rect 37419 14720 37461 14729
rect 37419 14680 37420 14720
rect 37460 14680 37461 14720
rect 37419 14671 37461 14680
rect 37420 14586 37460 14671
rect 36940 14428 37268 14468
rect 36652 14132 36692 14141
rect 36940 14132 36980 14428
rect 36692 14092 36980 14132
rect 36652 14083 36692 14092
rect 34827 14048 34869 14057
rect 34827 14008 34828 14048
rect 34868 14008 34869 14048
rect 34827 13999 34869 14008
rect 37035 14048 37077 14057
rect 37035 14008 37036 14048
rect 37076 14008 37077 14048
rect 37035 13999 37077 14008
rect 37900 14048 37940 15511
rect 37996 15509 38036 15520
rect 38092 15560 38132 15763
rect 38188 15732 38228 15741
rect 38228 15692 38324 15728
rect 38188 15688 38324 15692
rect 38188 15683 38228 15688
rect 38092 15511 38132 15520
rect 38284 14972 38324 15688
rect 38379 15644 38421 15653
rect 38379 15604 38380 15644
rect 38420 15604 38421 15644
rect 38379 15595 38421 15604
rect 38380 15510 38420 15595
rect 38476 15560 38516 16024
rect 38476 15511 38516 15520
rect 38572 15560 38612 17023
rect 38667 15812 38709 15821
rect 38667 15772 38668 15812
rect 38708 15772 38709 15812
rect 38667 15763 38709 15772
rect 38572 15511 38612 15520
rect 38668 15560 38708 15763
rect 38380 14972 38420 14981
rect 38284 14932 38380 14972
rect 38284 14729 38324 14932
rect 38380 14923 38420 14932
rect 38668 14897 38708 15520
rect 38764 15485 38804 19123
rect 39436 19122 39476 19207
rect 39531 19172 39573 19181
rect 39531 19132 39532 19172
rect 39572 19132 39573 19172
rect 39531 19123 39573 19132
rect 39532 18584 39572 19123
rect 39340 18341 39380 18426
rect 39339 18332 39381 18341
rect 39339 18292 39340 18332
rect 39380 18292 39381 18332
rect 39339 18283 39381 18292
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 39532 17996 39572 18544
rect 39627 18584 39669 18593
rect 39627 18544 39628 18584
rect 39668 18544 39669 18584
rect 39627 18535 39669 18544
rect 39724 18584 39764 19300
rect 40107 19340 40149 19349
rect 40107 19300 40108 19340
rect 40148 19300 40149 19340
rect 40107 19291 40149 19300
rect 39820 19256 39860 19265
rect 39820 19097 39860 19216
rect 39819 19088 39861 19097
rect 39819 19048 39820 19088
rect 39860 19048 39861 19088
rect 39819 19039 39861 19048
rect 40108 18761 40148 19291
rect 40107 18752 40149 18761
rect 40107 18712 40108 18752
rect 40148 18712 40149 18752
rect 40107 18703 40149 18712
rect 39724 18535 39764 18544
rect 39820 18584 39860 18593
rect 40012 18584 40052 18593
rect 39860 18544 40012 18584
rect 39820 18535 39860 18544
rect 40012 18535 40052 18544
rect 39628 18450 39668 18535
rect 39724 17996 39764 18005
rect 39532 17956 39724 17996
rect 39052 17081 39092 17166
rect 39051 17072 39093 17081
rect 39051 17032 39052 17072
rect 39092 17032 39093 17072
rect 39051 17023 39093 17032
rect 39147 16988 39189 16997
rect 39147 16948 39148 16988
rect 39188 16948 39189 16988
rect 39147 16939 39189 16948
rect 39148 16854 39188 16939
rect 38955 16820 38997 16829
rect 38955 16780 38956 16820
rect 38996 16780 38997 16820
rect 38955 16771 38997 16780
rect 38763 15476 38805 15485
rect 38763 15436 38764 15476
rect 38804 15436 38805 15476
rect 38763 15427 38805 15436
rect 38667 14888 38709 14897
rect 38667 14848 38668 14888
rect 38708 14848 38709 14888
rect 38667 14839 38709 14848
rect 38283 14720 38325 14729
rect 38283 14680 38284 14720
rect 38324 14680 38325 14720
rect 38283 14671 38325 14680
rect 38476 14720 38516 14729
rect 38668 14720 38708 14729
rect 38516 14680 38668 14720
rect 38476 14671 38516 14680
rect 38668 14468 38708 14680
rect 38764 14720 38804 15427
rect 38956 14972 38996 16771
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 39340 16232 39380 16241
rect 39340 15569 39380 16192
rect 39339 15560 39381 15569
rect 39339 15520 39340 15560
rect 39380 15520 39381 15560
rect 39339 15511 39381 15520
rect 39532 15560 39572 17956
rect 39724 17947 39764 17956
rect 39916 17828 39956 17837
rect 39956 17788 40148 17828
rect 39916 17779 39956 17788
rect 40108 17576 40148 17788
rect 40108 17501 40148 17536
rect 40107 17492 40149 17501
rect 40107 17452 40108 17492
rect 40148 17452 40149 17492
rect 40107 17443 40149 17452
rect 40204 17300 40244 19384
rect 40299 19256 40341 19265
rect 40299 19216 40300 19256
rect 40340 19216 40341 19256
rect 40299 19207 40341 19216
rect 40396 19256 40436 19459
rect 40779 19340 40821 19349
rect 40779 19300 40780 19340
rect 40820 19300 40821 19340
rect 40779 19291 40821 19300
rect 40972 19301 41012 19459
rect 40396 19207 40436 19216
rect 40683 19256 40725 19265
rect 40683 19216 40684 19256
rect 40724 19216 40725 19256
rect 40683 19207 40725 19216
rect 40780 19256 40820 19291
rect 40300 19122 40340 19207
rect 40492 19097 40532 19179
rect 40684 19122 40724 19207
rect 40780 19205 40820 19216
rect 40876 19256 40916 19265
rect 40972 19252 41012 19261
rect 40491 19088 40533 19097
rect 40491 19044 40492 19088
rect 40532 19044 40533 19088
rect 40491 19039 40533 19044
rect 40492 19035 40532 19039
rect 40779 19004 40821 19013
rect 40779 18964 40780 19004
rect 40820 18964 40821 19004
rect 40779 18955 40821 18964
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 40683 18752 40725 18761
rect 40683 18712 40684 18752
rect 40724 18712 40725 18752
rect 40683 18703 40725 18712
rect 40396 18584 40436 18593
rect 40396 18425 40436 18544
rect 40395 18416 40437 18425
rect 40395 18376 40396 18416
rect 40436 18376 40437 18416
rect 40395 18367 40437 18376
rect 40299 17828 40341 17837
rect 40299 17788 40300 17828
rect 40340 17788 40341 17828
rect 40299 17779 40341 17788
rect 40492 17828 40532 17839
rect 40684 17837 40724 18703
rect 40300 17694 40340 17779
rect 40492 17753 40532 17788
rect 40683 17828 40725 17837
rect 40683 17788 40684 17828
rect 40724 17788 40725 17828
rect 40683 17779 40725 17788
rect 40491 17744 40533 17753
rect 40491 17704 40492 17744
rect 40532 17704 40533 17744
rect 40491 17695 40533 17704
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 40204 17260 40532 17300
rect 39723 17240 39765 17249
rect 39723 17200 39724 17240
rect 39764 17200 39765 17240
rect 39723 17191 39765 17200
rect 39724 16829 39764 17191
rect 40395 17072 40437 17081
rect 40395 17032 40396 17072
rect 40436 17032 40437 17072
rect 40395 17023 40437 17032
rect 39723 16820 39765 16829
rect 39723 16780 39724 16820
rect 39764 16780 39765 16820
rect 39723 16771 39765 16780
rect 40396 16568 40436 17023
rect 40492 16988 40532 17260
rect 40780 16988 40820 18955
rect 40876 18509 40916 19216
rect 41068 19172 41108 19636
rect 41164 19433 41204 19518
rect 41163 19424 41205 19433
rect 41163 19384 41164 19424
rect 41204 19384 41205 19424
rect 41163 19375 41205 19384
rect 40972 19132 41108 19172
rect 41164 19256 41204 19265
rect 40972 18845 41012 19132
rect 41067 19004 41109 19013
rect 41067 18964 41068 19004
rect 41108 18964 41109 19004
rect 41067 18955 41109 18964
rect 40971 18836 41013 18845
rect 40971 18796 40972 18836
rect 41012 18796 41013 18836
rect 40971 18787 41013 18796
rect 40875 18500 40917 18509
rect 40875 18460 40876 18500
rect 40916 18460 41012 18500
rect 40875 18451 40917 18460
rect 40972 17083 41012 18460
rect 41068 17240 41108 18955
rect 41164 18425 41204 19216
rect 41260 19013 41300 19804
rect 41452 19433 41492 19972
rect 41548 20054 41588 20063
rect 41740 20021 41780 20077
rect 41836 20056 41972 20077
rect 41451 19424 41493 19433
rect 41451 19384 41452 19424
rect 41492 19384 41493 19424
rect 41451 19375 41493 19384
rect 41356 19256 41396 19265
rect 41259 19004 41301 19013
rect 41259 18964 41260 19004
rect 41300 18964 41301 19004
rect 41259 18955 41301 18964
rect 41356 18845 41396 19216
rect 41452 19256 41492 19265
rect 41355 18836 41397 18845
rect 41355 18796 41356 18836
rect 41396 18796 41397 18836
rect 41355 18787 41397 18796
rect 41452 18668 41492 19216
rect 41548 18929 41588 20014
rect 41739 20012 41781 20021
rect 41739 19972 41740 20012
rect 41780 19972 41781 20012
rect 41739 19963 41781 19972
rect 41740 19953 41780 19963
rect 41932 19928 41972 20056
rect 42135 20056 42220 20096
rect 42135 19928 42175 20056
rect 42220 20047 42260 20056
rect 42316 20054 42356 20063
rect 42796 20046 42836 20131
rect 42316 19937 42356 20014
rect 41932 19879 41972 19888
rect 42124 19888 42175 19928
rect 42315 19928 42357 19937
rect 42315 19888 42316 19928
rect 42356 19888 42357 19928
rect 41739 19256 41781 19265
rect 41739 19216 41740 19256
rect 41780 19216 41781 19256
rect 41739 19207 41781 19216
rect 41740 19122 41780 19207
rect 42124 19181 42164 19888
rect 42315 19879 42357 19888
rect 42795 19928 42837 19937
rect 42795 19888 42796 19928
rect 42836 19888 42837 19928
rect 42795 19879 42837 19888
rect 42699 19424 42741 19433
rect 42699 19384 42700 19424
rect 42740 19384 42741 19424
rect 42699 19375 42741 19384
rect 42123 19172 42165 19181
rect 42123 19132 42124 19172
rect 42164 19132 42165 19172
rect 42123 19123 42165 19132
rect 42603 19172 42645 19181
rect 42603 19132 42604 19172
rect 42644 19132 42645 19172
rect 42603 19123 42645 19132
rect 41547 18920 41589 18929
rect 41547 18880 41548 18920
rect 41588 18880 41589 18920
rect 41547 18871 41589 18880
rect 42315 18836 42357 18845
rect 42315 18796 42316 18836
rect 42356 18796 42357 18836
rect 42315 18787 42357 18796
rect 42027 18668 42069 18677
rect 41452 18628 41780 18668
rect 41260 18584 41300 18593
rect 41300 18544 41684 18584
rect 41260 18535 41300 18544
rect 41163 18416 41205 18425
rect 41163 18376 41164 18416
rect 41204 18376 41205 18416
rect 41163 18367 41205 18376
rect 41260 17240 41300 17249
rect 41068 17200 41260 17240
rect 41260 17191 41300 17200
rect 40972 17034 41012 17043
rect 41164 17072 41204 17081
rect 40780 16948 41012 16988
rect 40492 16939 40532 16948
rect 40972 16904 41012 16948
rect 41164 16904 41204 17032
rect 40972 16864 41204 16904
rect 40683 16820 40725 16829
rect 40875 16820 40917 16829
rect 40683 16780 40684 16820
rect 40724 16780 40820 16820
rect 40683 16771 40725 16780
rect 40684 16686 40724 16771
rect 40491 16568 40533 16577
rect 40396 16528 40492 16568
rect 40532 16528 40533 16568
rect 40491 16519 40533 16528
rect 40492 16484 40532 16519
rect 40492 16433 40532 16444
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 39820 15728 39860 15737
rect 39860 15688 40052 15728
rect 39820 15679 39860 15688
rect 39627 15644 39669 15653
rect 39627 15604 39628 15644
rect 39668 15604 39669 15644
rect 39627 15595 39669 15604
rect 40012 15644 40052 15688
rect 40012 15595 40052 15604
rect 39532 15511 39572 15520
rect 39628 15560 39668 15595
rect 40780 15569 40820 16780
rect 40875 16780 40876 16820
rect 40916 16780 40917 16820
rect 40875 16771 40917 16780
rect 40876 16686 40916 16771
rect 41067 16232 41109 16241
rect 41067 16192 41068 16232
rect 41108 16192 41109 16232
rect 41067 16183 41109 16192
rect 41068 16098 41108 16183
rect 41163 16064 41205 16073
rect 41163 16024 41164 16064
rect 41204 16024 41205 16064
rect 41163 16015 41205 16024
rect 41164 15930 41204 16015
rect 39628 15509 39668 15520
rect 39724 15560 39764 15569
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 38956 14932 39284 14972
rect 38764 14671 38804 14680
rect 38956 14720 38996 14731
rect 38956 14645 38996 14680
rect 39244 14720 39284 14932
rect 39244 14671 39284 14680
rect 38955 14636 38997 14645
rect 38955 14596 38956 14636
rect 38996 14596 38997 14636
rect 38955 14587 38997 14596
rect 38860 14552 38900 14561
rect 38860 14468 38900 14512
rect 39244 14512 39476 14552
rect 39244 14468 39284 14512
rect 38668 14428 38804 14468
rect 38860 14428 39284 14468
rect 38764 14384 38804 14428
rect 39339 14384 39381 14393
rect 38764 14344 38996 14384
rect 38956 14216 38996 14344
rect 39339 14344 39340 14384
rect 39380 14344 39381 14384
rect 39339 14335 39381 14344
rect 39052 14216 39092 14225
rect 38956 14176 39052 14216
rect 39052 14167 39092 14176
rect 37900 13999 37940 14008
rect 39340 14048 39380 14335
rect 39340 13999 39380 14008
rect 37036 13914 37076 13999
rect 39436 13964 39476 14512
rect 39724 14468 39764 15520
rect 39915 15560 39957 15569
rect 39915 15520 39916 15560
rect 39956 15520 39957 15560
rect 39915 15511 39957 15520
rect 40395 15560 40437 15569
rect 40395 15520 40396 15560
rect 40436 15520 40437 15560
rect 40395 15511 40437 15520
rect 40779 15560 40821 15569
rect 40779 15520 40780 15560
rect 40820 15520 40821 15560
rect 40779 15511 40821 15520
rect 41260 15560 41300 15569
rect 41356 15560 41396 18544
rect 41547 18416 41589 18425
rect 41547 18376 41548 18416
rect 41588 18376 41589 18416
rect 41547 18367 41589 18376
rect 41451 16652 41493 16661
rect 41451 16612 41452 16652
rect 41492 16612 41493 16652
rect 41451 16603 41493 16612
rect 41300 15520 41396 15560
rect 41260 15511 41300 15520
rect 39916 15140 39956 15511
rect 39916 15100 40052 15140
rect 39915 14888 39957 14897
rect 39915 14848 39916 14888
rect 39956 14848 39957 14888
rect 39915 14839 39957 14848
rect 39436 13915 39476 13924
rect 39628 14428 39764 14468
rect 39628 13964 39668 14428
rect 39723 14216 39765 14225
rect 39723 14176 39724 14216
rect 39764 14176 39765 14216
rect 39723 14167 39765 14176
rect 39724 14048 39764 14167
rect 39916 14141 39956 14839
rect 39915 14132 39957 14141
rect 39915 14092 39916 14132
rect 39956 14092 39957 14132
rect 39915 14083 39957 14092
rect 39724 13999 39764 14008
rect 39532 13880 39572 13889
rect 39628 13880 39668 13924
rect 39916 13880 39956 13889
rect 39628 13840 39916 13880
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 39243 13292 39285 13301
rect 39148 13252 39244 13292
rect 39284 13252 39285 13292
rect 38763 13208 38805 13217
rect 38763 13168 38764 13208
rect 38804 13168 38805 13208
rect 38763 13159 38805 13168
rect 39148 13208 39188 13252
rect 39243 13243 39285 13252
rect 39532 13217 39572 13840
rect 39916 13831 39956 13840
rect 39148 13159 39188 13168
rect 39531 13208 39573 13217
rect 39531 13168 39532 13208
rect 39572 13168 39573 13208
rect 39531 13159 39573 13168
rect 40012 13208 40052 15100
rect 40396 14552 40436 15511
rect 40204 14512 40436 14552
rect 41260 14552 41300 14561
rect 40204 14300 40244 14512
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 40108 14260 40244 14300
rect 40779 14300 40821 14309
rect 40779 14260 40780 14300
rect 40820 14260 40821 14300
rect 40108 13301 40148 14260
rect 40779 14251 40821 14260
rect 40396 14225 40436 14229
rect 40395 14220 40437 14225
rect 40395 14176 40396 14220
rect 40436 14176 40437 14220
rect 40395 14167 40437 14176
rect 40299 14132 40341 14141
rect 40299 14092 40300 14132
rect 40340 14092 40341 14132
rect 40299 14083 40341 14092
rect 40396 14085 40436 14167
rect 40683 14132 40725 14141
rect 40683 14092 40684 14132
rect 40724 14092 40725 14132
rect 40683 14083 40725 14092
rect 40203 14048 40245 14057
rect 40203 14008 40204 14048
rect 40244 14008 40245 14048
rect 40203 13999 40245 14008
rect 40300 14048 40340 14083
rect 40204 13914 40244 13999
rect 40300 13997 40340 14008
rect 40587 14048 40629 14057
rect 40587 14008 40588 14048
rect 40628 14008 40629 14048
rect 40587 13999 40629 14008
rect 40684 14048 40724 14083
rect 40588 13914 40628 13999
rect 40684 13997 40724 14008
rect 40780 14048 40820 14251
rect 41067 14216 41109 14225
rect 41067 14176 41068 14216
rect 41108 14176 41109 14216
rect 41067 14167 41109 14176
rect 41068 14082 41108 14167
rect 40780 13999 40820 14008
rect 40876 14048 40916 14059
rect 41260 14057 41300 14512
rect 41356 14393 41396 15520
rect 41355 14384 41397 14393
rect 41355 14344 41356 14384
rect 41396 14344 41397 14384
rect 41355 14335 41397 14344
rect 40876 13973 40916 14008
rect 41164 14048 41204 14057
rect 40875 13964 40917 13973
rect 40875 13924 40876 13964
rect 40916 13924 40917 13964
rect 40875 13915 40917 13924
rect 41164 13460 41204 14008
rect 41259 14048 41301 14057
rect 41259 14008 41260 14048
rect 41300 14008 41301 14048
rect 41259 13999 41301 14008
rect 41164 13411 41204 13420
rect 40107 13292 40149 13301
rect 40107 13252 40108 13292
rect 40148 13252 40149 13292
rect 40107 13243 40149 13252
rect 40012 13159 40052 13168
rect 41355 13208 41397 13217
rect 41355 13168 41356 13208
rect 41396 13168 41397 13208
rect 41355 13159 41397 13168
rect 38764 13074 38804 13159
rect 41356 13074 41396 13159
rect 41164 13040 41204 13049
rect 41164 12980 41204 13000
rect 41164 12940 41300 12980
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 41260 12536 41300 12940
rect 41260 12487 41300 12496
rect 41356 12536 41396 12545
rect 41452 12536 41492 16603
rect 41548 14048 41588 18367
rect 41644 17744 41684 18544
rect 41740 17753 41780 18628
rect 42027 18628 42028 18668
rect 42068 18628 42069 18668
rect 42027 18619 42069 18628
rect 41644 17695 41684 17704
rect 41739 17744 41781 17753
rect 41739 17704 41740 17744
rect 41780 17704 41781 17744
rect 41739 17695 41781 17704
rect 42028 17249 42068 18619
rect 42219 17828 42261 17837
rect 42219 17788 42220 17828
rect 42260 17788 42261 17828
rect 42219 17779 42261 17788
rect 42027 17240 42069 17249
rect 42027 17200 42028 17240
rect 42068 17200 42069 17240
rect 42027 17191 42069 17200
rect 42220 14729 42260 17779
rect 42316 16661 42356 18787
rect 42604 18752 42644 19123
rect 42604 18703 42644 18712
rect 42700 18584 42740 19375
rect 42796 18740 42836 19879
rect 42892 19265 42932 20728
rect 42987 20768 43029 20777
rect 42987 20728 42988 20768
rect 43028 20728 43029 20768
rect 42987 20719 43029 20728
rect 42988 20516 43028 20719
rect 43852 20718 43892 20803
rect 43660 20600 43700 20609
rect 42988 20476 43220 20516
rect 43180 20109 43220 20476
rect 43660 20189 43700 20560
rect 43659 20180 43701 20189
rect 43659 20140 43660 20180
rect 43700 20140 43701 20180
rect 43659 20131 43701 20140
rect 44139 20180 44181 20189
rect 44139 20140 44140 20180
rect 44180 20140 44181 20180
rect 44139 20131 44181 20140
rect 43180 20060 43220 20069
rect 44043 20096 44085 20105
rect 44043 20056 44044 20096
rect 44084 20056 44085 20096
rect 44043 20047 44085 20056
rect 44044 19962 44084 20047
rect 43947 19592 43989 19601
rect 43947 19552 43948 19592
rect 43988 19552 43989 19592
rect 43947 19543 43989 19552
rect 43371 19508 43413 19517
rect 43371 19468 43372 19508
rect 43412 19468 43413 19508
rect 43371 19459 43413 19468
rect 42891 19256 42933 19265
rect 43180 19256 43220 19265
rect 42891 19216 42892 19256
rect 42932 19216 42933 19256
rect 42891 19207 42933 19216
rect 43084 19216 43180 19256
rect 42796 18700 42932 18740
rect 42796 18584 42836 18593
rect 42700 18535 42740 18544
rect 42795 18544 42796 18551
rect 42892 18584 42932 18700
rect 43084 18677 43124 19216
rect 43180 19188 43220 19216
rect 43083 18668 43125 18677
rect 43083 18628 43084 18668
rect 43124 18628 43125 18668
rect 43083 18619 43125 18628
rect 42836 18544 42837 18551
rect 42795 18542 42837 18544
rect 42411 18500 42453 18509
rect 42411 18460 42412 18500
rect 42452 18460 42453 18500
rect 42795 18502 42796 18542
rect 42836 18502 42837 18542
rect 42892 18535 42932 18544
rect 42795 18493 42837 18502
rect 43084 18500 43124 18509
rect 42411 18451 42453 18460
rect 42412 18005 42452 18451
rect 42796 18449 42836 18493
rect 42987 18332 43029 18341
rect 43084 18332 43124 18460
rect 43275 18416 43317 18425
rect 43275 18376 43276 18416
rect 43316 18376 43317 18416
rect 43275 18367 43317 18376
rect 42987 18292 42988 18332
rect 43028 18292 43124 18332
rect 42987 18283 43029 18292
rect 43276 18282 43316 18367
rect 43178 18164 43220 18173
rect 42988 18124 43179 18164
rect 43219 18124 43220 18164
rect 42988 18005 43028 18124
rect 43178 18115 43220 18124
rect 42411 17996 42453 18005
rect 42411 17956 42412 17996
rect 42452 17956 42453 17996
rect 42411 17947 42453 17956
rect 42987 17996 43029 18005
rect 42987 17956 42988 17996
rect 43028 17956 43029 17996
rect 42987 17947 43029 17956
rect 43372 17912 43412 19459
rect 43563 18836 43605 18845
rect 43563 18796 43564 18836
rect 43604 18796 43605 18836
rect 43563 18787 43605 18796
rect 43564 18752 43604 18787
rect 43948 18761 43988 19543
rect 44043 19256 44085 19265
rect 44043 19216 44044 19256
rect 44084 19216 44085 19256
rect 44043 19207 44085 19216
rect 44140 19256 44180 20131
rect 44236 19256 44276 21727
rect 44619 20936 44661 20945
rect 44619 20896 44620 20936
rect 44660 20896 44661 20936
rect 44619 20887 44661 20896
rect 44523 20852 44565 20861
rect 44523 20812 44524 20852
rect 44564 20812 44565 20852
rect 44523 20803 44565 20812
rect 44332 19433 44372 19518
rect 44331 19424 44373 19433
rect 44331 19384 44332 19424
rect 44372 19384 44373 19424
rect 44331 19375 44373 19384
rect 44332 19256 44372 19265
rect 44236 19216 44332 19256
rect 44140 19207 44180 19216
rect 44332 19207 44372 19216
rect 44044 19122 44084 19207
rect 43564 18701 43604 18712
rect 43947 18752 43989 18761
rect 43947 18712 43948 18752
rect 43988 18712 43989 18752
rect 43947 18703 43989 18712
rect 44139 18752 44181 18761
rect 44139 18712 44140 18752
rect 44180 18712 44181 18752
rect 44139 18703 44181 18712
rect 43468 18584 43508 18595
rect 43468 18509 43508 18544
rect 43756 18584 43796 18593
rect 44140 18584 44180 18703
rect 43796 18544 44084 18584
rect 43756 18535 43796 18544
rect 43467 18500 43509 18509
rect 43467 18460 43468 18500
rect 43508 18460 43509 18500
rect 43467 18451 43509 18460
rect 44044 18080 44084 18544
rect 44140 18535 44180 18544
rect 44524 18341 44564 20803
rect 44523 18332 44565 18341
rect 44523 18292 44524 18332
rect 44564 18292 44565 18332
rect 44523 18283 44565 18292
rect 44620 18089 44660 20887
rect 45388 20264 45428 25003
rect 45867 23120 45909 23129
rect 45867 23080 45868 23120
rect 45908 23080 45909 23120
rect 45867 23071 45909 23080
rect 45964 23120 46004 25768
rect 46444 25733 46484 29035
rect 46540 28328 46580 29800
rect 46636 29168 46676 30211
rect 48268 30092 48308 30472
rect 47788 30052 48308 30092
rect 47403 29840 47445 29849
rect 47403 29800 47404 29840
rect 47444 29800 47445 29840
rect 47403 29791 47445 29800
rect 47788 29840 47828 30052
rect 48460 30008 48500 30640
rect 48076 29968 48500 30008
rect 48076 29924 48116 29968
rect 47980 29840 48020 29849
rect 47788 29791 47828 29800
rect 47884 29800 47980 29840
rect 47404 29345 47444 29791
rect 46732 29336 46772 29345
rect 47403 29336 47445 29345
rect 46772 29296 47252 29336
rect 46732 29287 46772 29296
rect 46828 29168 46868 29177
rect 46636 29093 46676 29128
rect 46732 29128 46828 29168
rect 46635 29084 46677 29093
rect 46635 29044 46636 29084
rect 46676 29044 46677 29084
rect 46635 29035 46677 29044
rect 46635 28328 46677 28337
rect 46540 28288 46636 28328
rect 46676 28288 46677 28328
rect 46635 28279 46677 28288
rect 46636 28194 46676 28279
rect 46732 26144 46772 29128
rect 46828 29119 46868 29128
rect 46923 29168 46965 29177
rect 46923 29128 46924 29168
rect 46964 29128 46965 29168
rect 46923 29119 46965 29128
rect 47116 29168 47156 29177
rect 46924 29034 46964 29119
rect 46540 26104 46772 26144
rect 47116 26816 47156 29128
rect 47212 29084 47252 29296
rect 47403 29296 47404 29336
rect 47444 29296 47445 29336
rect 47403 29287 47445 29296
rect 47884 29177 47924 29800
rect 47980 29791 48020 29800
rect 48076 29672 48116 29884
rect 48364 29756 48404 29765
rect 47980 29632 48116 29672
rect 48268 29716 48364 29756
rect 47980 29394 48020 29632
rect 47980 29345 48020 29354
rect 48171 29252 48213 29261
rect 48171 29212 48172 29252
rect 48212 29212 48213 29252
rect 48171 29203 48213 29212
rect 47500 29168 47540 29177
rect 47212 29035 47252 29044
rect 47403 29084 47445 29093
rect 47403 29044 47404 29084
rect 47444 29044 47445 29084
rect 47403 29035 47445 29044
rect 47307 29000 47349 29009
rect 47307 28960 47308 29000
rect 47348 28960 47349 29000
rect 47307 28951 47349 28960
rect 47308 28866 47348 28951
rect 47404 28950 47444 29035
rect 47308 27824 47348 27833
rect 47500 27828 47540 29128
rect 47883 29168 47925 29177
rect 47883 29128 47884 29168
rect 47924 29128 47925 29168
rect 47883 29119 47925 29128
rect 48075 29168 48117 29177
rect 48075 29128 48076 29168
rect 48116 29128 48117 29168
rect 48075 29119 48117 29128
rect 48172 29168 48212 29203
rect 47979 29084 48021 29093
rect 47979 29044 47980 29084
rect 48020 29044 48021 29084
rect 47979 29035 48021 29044
rect 47788 28160 47828 28169
rect 47596 27828 47636 27856
rect 47788 27833 47828 28120
rect 47500 27824 47596 27828
rect 47348 27788 47596 27824
rect 47348 27784 47540 27788
rect 47308 27775 47348 27784
rect 47596 27779 47636 27788
rect 47787 27824 47829 27833
rect 47787 27784 47788 27824
rect 47828 27784 47829 27824
rect 47787 27775 47829 27784
rect 47980 27824 48020 29035
rect 48076 29034 48116 29119
rect 48172 29117 48212 29128
rect 48268 28916 48308 29716
rect 48364 29707 48404 29716
rect 48460 29000 48500 29009
rect 48556 29000 48596 30808
rect 49900 29849 49940 32908
rect 49996 32899 50036 32908
rect 50476 32864 50516 33403
rect 50476 32815 50516 32824
rect 50572 32864 50612 32873
rect 50572 32621 50612 32824
rect 50764 32864 50804 34327
rect 50859 33872 50901 33881
rect 50859 33832 50860 33872
rect 50900 33832 50901 33872
rect 50859 33823 50901 33832
rect 51339 33872 51381 33881
rect 51339 33832 51340 33872
rect 51380 33832 51381 33872
rect 51339 33823 51381 33832
rect 50668 32696 50708 32705
rect 50571 32612 50613 32621
rect 50571 32572 50572 32612
rect 50612 32572 50613 32612
rect 50571 32563 50613 32572
rect 50572 32192 50612 32201
rect 50187 31604 50229 31613
rect 50187 31564 50188 31604
rect 50228 31564 50229 31604
rect 50187 31555 50229 31564
rect 50188 31470 50228 31555
rect 50476 31529 50516 31560
rect 50475 31520 50517 31529
rect 50475 31480 50476 31520
rect 50516 31480 50517 31520
rect 50475 31471 50517 31480
rect 50572 31520 50612 32152
rect 50572 31471 50612 31480
rect 49996 31436 50036 31445
rect 48747 29840 48789 29849
rect 48747 29800 48748 29840
rect 48788 29800 48789 29840
rect 48747 29791 48789 29800
rect 49515 29840 49557 29849
rect 49515 29800 49516 29840
rect 49556 29800 49557 29840
rect 49515 29791 49557 29800
rect 49612 29840 49652 29849
rect 49899 29840 49941 29849
rect 49652 29800 49748 29840
rect 49612 29791 49652 29800
rect 48748 29706 48788 29791
rect 48651 29252 48693 29261
rect 48651 29212 48652 29252
rect 48692 29212 48693 29252
rect 48651 29203 48693 29212
rect 48652 29118 48692 29203
rect 48748 29168 48788 29177
rect 48172 28876 48308 28916
rect 48364 28960 48460 29000
rect 48500 28960 48596 29000
rect 48172 28328 48212 28876
rect 48364 28832 48404 28960
rect 48460 28951 48500 28960
rect 48172 28279 48212 28288
rect 48268 28792 48404 28832
rect 48268 28328 48308 28792
rect 48268 28279 48308 28288
rect 48364 28328 48404 28337
rect 48364 28001 48404 28288
rect 48460 28328 48500 28337
rect 48748 28328 48788 29128
rect 48844 29168 48884 29179
rect 48844 29093 48884 29128
rect 48939 29168 48981 29177
rect 48939 29128 48940 29168
rect 48980 29128 48981 29168
rect 48939 29119 48981 29128
rect 48843 29084 48885 29093
rect 48843 29044 48844 29084
rect 48884 29044 48885 29084
rect 48843 29035 48885 29044
rect 48500 28288 48788 28328
rect 48460 28279 48500 28288
rect 48363 27992 48405 28001
rect 48363 27952 48364 27992
rect 48404 27952 48405 27992
rect 48363 27943 48405 27952
rect 47980 27784 48500 27824
rect 47980 27782 48020 27784
rect 47980 27733 48020 27742
rect 47403 27656 47445 27665
rect 47403 27616 47404 27656
rect 47444 27616 47445 27656
rect 47403 27607 47445 27616
rect 47692 27656 47732 27665
rect 47307 27320 47349 27329
rect 47307 27280 47308 27320
rect 47348 27280 47349 27320
rect 47307 27271 47349 27280
rect 47211 26900 47253 26909
rect 47211 26860 47212 26900
rect 47252 26860 47253 26900
rect 47211 26851 47253 26860
rect 46443 25724 46485 25733
rect 46443 25684 46444 25724
rect 46484 25684 46485 25724
rect 46443 25675 46485 25684
rect 46252 24632 46292 24641
rect 46059 24380 46101 24389
rect 46059 24340 46060 24380
rect 46100 24340 46101 24380
rect 46059 24331 46101 24340
rect 46060 24246 46100 24331
rect 46252 23801 46292 24592
rect 46251 23792 46293 23801
rect 46251 23752 46252 23792
rect 46292 23752 46293 23792
rect 46251 23743 46293 23752
rect 46059 23204 46101 23213
rect 46059 23164 46060 23204
rect 46100 23164 46101 23204
rect 46059 23155 46101 23164
rect 45964 23071 46004 23080
rect 46060 23120 46100 23155
rect 45868 22280 45908 23071
rect 46060 23069 46100 23080
rect 46156 23120 46196 23129
rect 46156 22532 46196 23080
rect 46252 23120 46292 23129
rect 46444 23120 46484 23129
rect 46292 23080 46444 23120
rect 46252 23071 46292 23080
rect 46444 23071 46484 23080
rect 46540 23045 46580 26104
rect 46635 25976 46677 25985
rect 46635 25936 46636 25976
rect 46676 25936 46677 25976
rect 46635 25927 46677 25936
rect 46636 24632 46676 25927
rect 47116 25901 47156 26776
rect 47212 26732 47252 26851
rect 47308 26816 47348 27271
rect 47308 26767 47348 26776
rect 47404 26816 47444 27607
rect 47692 27245 47732 27616
rect 47788 27656 47828 27665
rect 48268 27656 48308 27665
rect 47828 27616 48212 27656
rect 47788 27607 47828 27616
rect 47691 27236 47733 27245
rect 47691 27196 47692 27236
rect 47732 27196 47733 27236
rect 47691 27187 47733 27196
rect 48075 27236 48117 27245
rect 48075 27196 48076 27236
rect 48116 27196 48117 27236
rect 48075 27187 48117 27196
rect 47788 26984 47828 26993
rect 47691 26900 47733 26909
rect 47691 26860 47692 26900
rect 47732 26860 47733 26900
rect 47691 26851 47733 26860
rect 47404 26767 47444 26776
rect 47596 26816 47636 26825
rect 47212 26683 47252 26692
rect 47212 25976 47252 25985
rect 47115 25892 47157 25901
rect 47115 25852 47116 25892
rect 47156 25852 47157 25892
rect 47115 25843 47157 25852
rect 46923 25808 46965 25817
rect 46923 25768 46924 25808
rect 46964 25768 46965 25808
rect 46923 25759 46965 25768
rect 46924 25481 46964 25759
rect 47212 25649 47252 25936
rect 47596 25733 47636 26776
rect 47692 26766 47732 26851
rect 47788 26228 47828 26944
rect 47788 26179 47828 26188
rect 47884 26900 47924 26909
rect 47307 25724 47349 25733
rect 47307 25684 47308 25724
rect 47348 25684 47349 25724
rect 47307 25675 47349 25684
rect 47595 25724 47637 25733
rect 47595 25684 47596 25724
rect 47636 25684 47637 25724
rect 47595 25675 47637 25684
rect 47211 25640 47253 25649
rect 47211 25600 47212 25640
rect 47252 25600 47253 25640
rect 47211 25591 47253 25600
rect 46923 25472 46965 25481
rect 46923 25432 46924 25472
rect 46964 25432 46965 25472
rect 46923 25423 46965 25432
rect 46676 24592 46868 24632
rect 46636 24583 46676 24592
rect 46635 24464 46677 24473
rect 46635 24424 46636 24464
rect 46676 24424 46677 24464
rect 46635 24415 46677 24424
rect 46539 23036 46581 23045
rect 46539 22996 46540 23036
rect 46580 22996 46581 23036
rect 46539 22987 46581 22996
rect 46444 22532 46484 22541
rect 46156 22492 46444 22532
rect 46059 22364 46101 22373
rect 46059 22324 46060 22364
rect 46100 22324 46101 22364
rect 46059 22315 46101 22324
rect 45292 20224 45428 20264
rect 45772 22240 45868 22280
rect 45003 20096 45045 20105
rect 45003 20056 45004 20096
rect 45044 20056 45045 20096
rect 45003 20047 45045 20056
rect 45004 19097 45044 20047
rect 45196 19844 45236 19853
rect 45100 19340 45140 19349
rect 45100 19181 45140 19300
rect 45099 19172 45141 19181
rect 45099 19132 45100 19172
rect 45140 19132 45141 19172
rect 45099 19123 45141 19132
rect 45003 19088 45045 19097
rect 45003 19048 45004 19088
rect 45044 19048 45045 19088
rect 45003 19039 45045 19048
rect 44907 18752 44949 18761
rect 44907 18712 44908 18752
rect 44948 18712 44949 18752
rect 44907 18703 44949 18712
rect 44619 18080 44661 18089
rect 44044 18040 44564 18080
rect 43467 17912 43509 17921
rect 43372 17872 43468 17912
rect 43508 17872 43509 17912
rect 43467 17863 43509 17872
rect 44043 17912 44085 17921
rect 44043 17872 44044 17912
rect 44084 17872 44085 17912
rect 44043 17863 44085 17872
rect 43468 17753 43508 17863
rect 42508 17744 42548 17753
rect 42508 17585 42548 17704
rect 43083 17744 43125 17753
rect 43083 17704 43084 17744
rect 43124 17704 43125 17744
rect 43083 17695 43125 17704
rect 43467 17744 43509 17753
rect 43467 17704 43468 17744
rect 43508 17704 43509 17744
rect 43467 17695 43509 17704
rect 43564 17744 43604 17753
rect 44044 17744 44084 17863
rect 44140 17753 44180 17838
rect 44235 17828 44277 17837
rect 44235 17788 44236 17828
rect 44276 17788 44277 17828
rect 44235 17779 44277 17788
rect 43604 17704 43988 17744
rect 43564 17695 43604 17704
rect 42892 17660 42932 17669
rect 42507 17576 42549 17585
rect 42507 17536 42508 17576
rect 42548 17536 42549 17576
rect 42507 17527 42549 17536
rect 42411 17072 42453 17081
rect 42411 17032 42412 17072
rect 42452 17032 42453 17072
rect 42411 17023 42453 17032
rect 42315 16652 42357 16661
rect 42315 16612 42316 16652
rect 42356 16612 42357 16652
rect 42315 16603 42357 16612
rect 42412 16241 42452 17023
rect 42892 16913 42932 17620
rect 43084 17610 43124 17695
rect 43468 17610 43508 17695
rect 43756 17618 43796 17627
rect 43179 17576 43221 17585
rect 43179 17536 43180 17576
rect 43220 17536 43221 17576
rect 43179 17527 43221 17536
rect 43371 17576 43413 17585
rect 43755 17578 43756 17585
rect 43796 17578 43797 17585
rect 43755 17576 43797 17578
rect 43371 17532 43372 17576
rect 43412 17532 43413 17576
rect 43371 17527 43413 17532
rect 43564 17536 43756 17576
rect 43796 17536 43797 17576
rect 43948 17576 43988 17704
rect 44044 17695 44084 17704
rect 44139 17744 44181 17753
rect 44139 17704 44140 17744
rect 44180 17704 44181 17744
rect 44139 17695 44181 17704
rect 44236 17744 44276 17779
rect 44236 17693 44276 17704
rect 44524 17744 44564 18040
rect 44619 18040 44620 18080
rect 44660 18040 44661 18080
rect 44619 18031 44661 18040
rect 44811 17828 44853 17837
rect 44811 17788 44812 17828
rect 44852 17788 44853 17828
rect 44811 17779 44853 17788
rect 44524 17695 44564 17704
rect 44620 17744 44660 17753
rect 44620 17585 44660 17704
rect 44716 17744 44756 17753
rect 44332 17576 44372 17585
rect 43948 17536 44332 17576
rect 43180 17072 43220 17527
rect 43372 17441 43412 17527
rect 43276 17072 43316 17081
rect 43564 17072 43604 17536
rect 43755 17527 43797 17536
rect 44332 17527 44372 17536
rect 44619 17576 44661 17585
rect 44619 17536 44620 17576
rect 44660 17536 44661 17576
rect 44619 17527 44661 17536
rect 43756 17442 43796 17527
rect 44619 17408 44661 17417
rect 44619 17368 44620 17408
rect 44660 17368 44661 17408
rect 44619 17359 44661 17368
rect 44140 17081 44180 17166
rect 43180 17032 43276 17072
rect 43276 17023 43316 17032
rect 43372 17032 43604 17072
rect 43659 17072 43701 17081
rect 43659 17032 43660 17072
rect 43700 17032 43701 17072
rect 43372 16988 43412 17032
rect 43659 17023 43701 17032
rect 44139 17072 44181 17081
rect 44139 17032 44140 17072
rect 44180 17032 44181 17072
rect 44139 17023 44181 17032
rect 44332 17072 44372 17081
rect 43372 16939 43412 16948
rect 43564 16946 43604 16955
rect 42891 16904 42933 16913
rect 42891 16864 42892 16904
rect 42932 16864 42933 16904
rect 43563 16906 43564 16913
rect 43660 16938 43700 17023
rect 43604 16906 43605 16913
rect 43563 16904 43605 16906
rect 42891 16855 42933 16864
rect 43468 16862 43508 16871
rect 43563 16864 43564 16904
rect 43604 16864 43605 16904
rect 43563 16855 43605 16864
rect 44139 16904 44181 16913
rect 44139 16864 44140 16904
rect 44180 16864 44181 16904
rect 44139 16855 44181 16864
rect 43468 16745 43508 16822
rect 43564 16811 43604 16855
rect 44140 16770 44180 16855
rect 43467 16736 43509 16745
rect 43467 16696 43468 16736
rect 43508 16696 43509 16736
rect 43467 16687 43509 16696
rect 44332 16661 44372 17032
rect 44427 17072 44469 17081
rect 44427 17032 44428 17072
rect 44468 17032 44469 17072
rect 44427 17023 44469 17032
rect 44428 16938 44468 17023
rect 44331 16652 44373 16661
rect 44331 16612 44332 16652
rect 44372 16612 44373 16652
rect 44331 16603 44373 16612
rect 42411 16232 42453 16241
rect 42411 16192 42412 16232
rect 42452 16192 42453 16232
rect 42411 16183 42453 16192
rect 42892 16232 42932 16241
rect 42412 15728 42452 16183
rect 42795 16148 42837 16157
rect 42412 15679 42452 15688
rect 42700 16108 42796 16148
rect 42836 16108 42837 16148
rect 42604 15560 42644 15569
rect 42508 15520 42604 15560
rect 42412 15308 42452 15317
rect 42316 15268 42412 15308
rect 42219 14720 42261 14729
rect 42219 14680 42220 14720
rect 42260 14680 42261 14720
rect 42219 14671 42261 14680
rect 42220 14225 42260 14671
rect 42316 14309 42356 15268
rect 42412 15259 42452 15268
rect 42508 15056 42548 15520
rect 42604 15511 42644 15520
rect 42700 15224 42740 16108
rect 42795 16099 42837 16108
rect 42796 16014 42836 16099
rect 42892 15317 42932 16192
rect 43468 16232 43508 16241
rect 43084 16148 43124 16157
rect 42987 15560 43029 15569
rect 42987 15520 42988 15560
rect 43028 15520 43029 15560
rect 42987 15511 43029 15520
rect 42988 15426 43028 15511
rect 43084 15401 43124 16108
rect 43468 15569 43508 16192
rect 44332 16232 44372 16241
rect 43467 15560 43509 15569
rect 43467 15520 43468 15560
rect 43508 15520 43509 15560
rect 43467 15511 43509 15520
rect 43852 15560 43892 15569
rect 44332 15560 44372 16192
rect 43892 15520 44372 15560
rect 43083 15392 43125 15401
rect 43083 15352 43084 15392
rect 43124 15352 43125 15392
rect 43083 15343 43125 15352
rect 42891 15308 42933 15317
rect 42891 15268 42892 15308
rect 42932 15268 42933 15308
rect 42891 15259 42933 15268
rect 43179 15308 43221 15317
rect 43179 15268 43180 15308
rect 43220 15268 43221 15308
rect 43179 15259 43221 15268
rect 42412 15016 42548 15056
rect 42604 15184 42740 15224
rect 42412 14720 42452 15016
rect 42412 14671 42452 14680
rect 42508 14720 42548 14729
rect 42315 14300 42357 14309
rect 42315 14260 42316 14300
rect 42356 14260 42357 14300
rect 42315 14251 42357 14260
rect 42219 14216 42261 14225
rect 42219 14176 42220 14216
rect 42260 14176 42261 14216
rect 42219 14167 42261 14176
rect 42027 14132 42069 14141
rect 42027 14092 42028 14132
rect 42068 14092 42069 14132
rect 42027 14083 42069 14092
rect 41644 14048 41684 14057
rect 41548 14008 41644 14048
rect 41548 12629 41588 14008
rect 41644 13999 41684 14008
rect 42028 14048 42068 14083
rect 42028 13997 42068 14008
rect 41740 13964 41780 13973
rect 41740 13460 41780 13924
rect 41932 13964 41972 13973
rect 41644 13420 41780 13460
rect 41836 13880 41876 13889
rect 41932 13880 41972 13924
rect 42412 13880 42452 13889
rect 42508 13880 42548 14680
rect 42604 14720 42644 15184
rect 42700 14729 42740 14814
rect 42604 14671 42644 14680
rect 42699 14720 42741 14729
rect 42699 14680 42700 14720
rect 42740 14680 42741 14720
rect 42699 14671 42741 14680
rect 43083 14720 43125 14729
rect 43083 14680 43084 14720
rect 43124 14680 43125 14720
rect 43083 14671 43125 14680
rect 43180 14720 43220 15259
rect 43180 14671 43220 14680
rect 43275 14720 43317 14729
rect 43275 14680 43276 14720
rect 43316 14680 43317 14720
rect 43275 14671 43317 14680
rect 42988 14552 43028 14561
rect 42700 14512 42988 14552
rect 42603 14384 42645 14393
rect 42603 14344 42604 14384
rect 42644 14344 42645 14384
rect 42603 14335 42645 14344
rect 41932 13840 42412 13880
rect 42452 13840 42548 13880
rect 41547 12620 41589 12629
rect 41547 12580 41548 12620
rect 41588 12580 41589 12620
rect 41547 12571 41589 12580
rect 41396 12496 41492 12536
rect 41356 12487 41396 12496
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 41259 11612 41301 11621
rect 41259 11572 41260 11612
rect 41300 11572 41301 11612
rect 41259 11563 41301 11572
rect 41260 11478 41300 11563
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 41452 11285 41492 12496
rect 41548 12536 41588 12571
rect 41548 12486 41588 12496
rect 41548 12368 41588 12377
rect 41644 12368 41684 13420
rect 41739 13292 41781 13301
rect 41739 13252 41740 13292
rect 41780 13252 41781 13292
rect 41739 13243 41781 13252
rect 41588 12328 41684 12368
rect 41740 13208 41780 13243
rect 41836 13217 41876 13840
rect 42412 13831 42452 13840
rect 41548 12319 41588 12328
rect 41644 11696 41684 11705
rect 41740 11696 41780 13168
rect 41835 13208 41877 13217
rect 41835 13168 41836 13208
rect 41876 13168 41877 13208
rect 41835 13159 41877 13168
rect 42604 13208 42644 14335
rect 42700 14031 42740 14512
rect 42988 14503 43028 14512
rect 42892 14220 42932 14229
rect 42892 14141 42932 14180
rect 42891 14132 42933 14141
rect 42891 14092 42892 14132
rect 42932 14092 42933 14132
rect 42891 14083 42933 14092
rect 42700 13982 42740 13991
rect 42796 14048 42836 14059
rect 42796 13973 42836 14008
rect 42795 13964 42837 13973
rect 42795 13924 42796 13964
rect 42836 13924 42837 13964
rect 42795 13915 42837 13924
rect 42795 13796 42837 13805
rect 42795 13756 42796 13796
rect 42836 13756 42837 13796
rect 42795 13747 42837 13756
rect 42604 12980 42644 13168
rect 41684 11656 41780 11696
rect 42508 12940 42644 12980
rect 42508 11696 42548 12940
rect 41644 11647 41684 11656
rect 42508 11647 42548 11656
rect 42411 11612 42453 11621
rect 42411 11572 42412 11612
rect 42452 11572 42453 11612
rect 42411 11563 42453 11572
rect 41451 11276 41493 11285
rect 41451 11236 41452 11276
rect 41492 11236 41493 11276
rect 41451 11227 41493 11236
rect 42412 11192 42452 11563
rect 42699 11360 42741 11369
rect 42699 11320 42700 11360
rect 42740 11320 42741 11360
rect 42699 11311 42741 11320
rect 42508 11192 42548 11201
rect 42412 11152 42508 11192
rect 42508 11143 42548 11152
rect 42603 11024 42645 11033
rect 42603 10984 42604 11024
rect 42644 10984 42645 11024
rect 42603 10975 42645 10984
rect 42700 11024 42740 11311
rect 42796 11117 42836 13747
rect 42892 12704 42932 14083
rect 43084 13805 43124 14671
rect 43276 13973 43316 14671
rect 43852 14393 43892 15520
rect 43851 14384 43893 14393
rect 43851 14344 43852 14384
rect 43892 14344 43893 14384
rect 43851 14335 43893 14344
rect 44427 14300 44469 14309
rect 44427 14260 44428 14300
rect 44468 14260 44469 14300
rect 44427 14251 44469 14260
rect 43275 13964 43317 13973
rect 43275 13924 43276 13964
rect 43316 13924 43317 13964
rect 43275 13915 43317 13924
rect 43659 13964 43701 13973
rect 43659 13924 43660 13964
rect 43700 13924 43701 13964
rect 43659 13915 43701 13924
rect 43083 13796 43125 13805
rect 43083 13756 43084 13796
rect 43124 13756 43125 13796
rect 43083 13747 43125 13756
rect 43180 12704 43220 12713
rect 42892 12664 43180 12704
rect 43180 12655 43220 12664
rect 43275 12536 43317 12545
rect 43275 12496 43276 12536
rect 43316 12496 43317 12536
rect 43275 12487 43317 12496
rect 43564 12536 43604 12545
rect 43276 12402 43316 12487
rect 43468 12284 43508 12295
rect 43468 12209 43508 12244
rect 43275 12200 43317 12209
rect 43275 12160 43276 12200
rect 43316 12160 43317 12200
rect 43275 12151 43317 12160
rect 43467 12200 43509 12209
rect 43467 12160 43468 12200
rect 43508 12160 43509 12200
rect 43467 12151 43509 12160
rect 43276 11369 43316 12151
rect 43564 12125 43604 12496
rect 43563 12116 43605 12125
rect 43563 12076 43564 12116
rect 43604 12076 43605 12116
rect 43660 12116 43700 13915
rect 44428 13208 44468 14251
rect 44428 13159 44468 13168
rect 44620 13133 44660 17359
rect 44716 16997 44756 17704
rect 44812 17744 44852 17779
rect 44812 17693 44852 17704
rect 44715 16988 44757 16997
rect 44715 16948 44716 16988
rect 44756 16948 44757 16988
rect 44715 16939 44757 16948
rect 44811 14468 44853 14477
rect 44811 14428 44812 14468
rect 44852 14428 44853 14468
rect 44811 14419 44853 14428
rect 44812 13880 44852 14419
rect 44716 13840 44812 13880
rect 44908 13880 44948 18703
rect 45004 18584 45044 19039
rect 45100 18761 45140 19123
rect 45099 18752 45141 18761
rect 45099 18712 45100 18752
rect 45140 18712 45141 18752
rect 45099 18703 45141 18712
rect 45004 18535 45044 18544
rect 45196 18509 45236 19804
rect 45292 19508 45332 20224
rect 45772 20105 45812 22240
rect 45868 22231 45908 22240
rect 45867 22112 45909 22121
rect 45867 22072 45868 22112
rect 45908 22072 45909 22112
rect 45867 22063 45909 22072
rect 45868 21608 45908 22063
rect 45963 21776 46005 21785
rect 45963 21736 45964 21776
rect 46004 21736 46005 21776
rect 45963 21727 46005 21736
rect 45868 21559 45908 21568
rect 45964 21608 46004 21727
rect 45964 21559 46004 21568
rect 46060 20861 46100 22315
rect 46156 22028 46196 22492
rect 46444 22483 46484 22492
rect 46540 22373 46580 22987
rect 46539 22364 46581 22373
rect 46539 22324 46540 22364
rect 46580 22324 46581 22364
rect 46539 22315 46581 22324
rect 46252 22196 46292 22205
rect 46539 22196 46581 22205
rect 46292 22156 46388 22196
rect 46252 22147 46292 22156
rect 46156 21988 46292 22028
rect 46155 21776 46197 21785
rect 46155 21736 46156 21776
rect 46196 21736 46197 21776
rect 46155 21727 46197 21736
rect 46156 21608 46196 21727
rect 46156 21559 46196 21568
rect 46252 21524 46292 21988
rect 46252 21475 46292 21484
rect 46348 21440 46388 22156
rect 46539 22156 46540 22196
rect 46580 22156 46581 22196
rect 46539 22147 46581 22156
rect 46540 21608 46580 22147
rect 46636 21608 46676 24415
rect 46828 23129 46868 24592
rect 46827 23120 46869 23129
rect 46827 23080 46828 23120
rect 46868 23080 46869 23120
rect 46827 23071 46869 23080
rect 46732 22280 46772 22289
rect 46732 21776 46772 22240
rect 46828 22280 46868 22289
rect 46924 22280 46964 25423
rect 47308 23960 47348 25675
rect 47403 25472 47445 25481
rect 47403 25432 47404 25472
rect 47444 25432 47445 25472
rect 47403 25423 47445 25432
rect 47787 25472 47829 25481
rect 47884 25472 47924 26860
rect 48076 26825 48116 27187
rect 47787 25432 47788 25472
rect 47828 25432 47924 25472
rect 47980 26816 48020 26825
rect 47787 25423 47829 25432
rect 47212 23920 47348 23960
rect 47115 23876 47157 23885
rect 47115 23836 47116 23876
rect 47156 23836 47157 23876
rect 47115 23827 47157 23836
rect 47116 23213 47156 23827
rect 47115 23204 47157 23213
rect 47115 23164 47116 23204
rect 47156 23164 47157 23204
rect 47115 23155 47157 23164
rect 47116 22532 47156 23155
rect 47212 23060 47252 23920
rect 47307 23792 47349 23801
rect 47307 23752 47308 23792
rect 47348 23752 47349 23792
rect 47307 23743 47349 23752
rect 47404 23792 47444 25423
rect 47788 25338 47828 25423
rect 47980 25229 48020 26776
rect 48075 26816 48117 26825
rect 48075 26776 48076 26816
rect 48116 26776 48117 26816
rect 48075 26767 48117 26776
rect 48172 26816 48212 27616
rect 48172 26767 48212 26776
rect 48268 26816 48308 27616
rect 48364 27656 48404 27665
rect 48364 27413 48404 27616
rect 48460 27656 48500 27784
rect 48460 27607 48500 27616
rect 48555 27656 48597 27665
rect 48555 27616 48556 27656
rect 48596 27616 48597 27656
rect 48555 27607 48597 27616
rect 48556 27522 48596 27607
rect 48363 27404 48405 27413
rect 48363 27364 48364 27404
rect 48404 27364 48405 27404
rect 48363 27355 48405 27364
rect 48555 27320 48597 27329
rect 48555 27280 48556 27320
rect 48596 27280 48597 27320
rect 48555 27271 48597 27280
rect 48076 25808 48116 26767
rect 48172 26144 48212 26153
rect 48172 25985 48212 26104
rect 48171 25976 48213 25985
rect 48171 25936 48172 25976
rect 48212 25936 48213 25976
rect 48171 25927 48213 25936
rect 48076 25768 48212 25808
rect 48172 25313 48212 25768
rect 48268 25724 48308 26776
rect 48364 26816 48404 26827
rect 48364 26741 48404 26776
rect 48459 26816 48501 26825
rect 48459 26776 48460 26816
rect 48500 26776 48501 26816
rect 48459 26767 48501 26776
rect 48363 26732 48405 26741
rect 48363 26692 48364 26732
rect 48404 26692 48405 26732
rect 48363 26683 48405 26692
rect 48460 26682 48500 26767
rect 48268 25684 48404 25724
rect 48267 25556 48309 25565
rect 48267 25516 48268 25556
rect 48308 25516 48309 25556
rect 48267 25507 48309 25516
rect 48076 25304 48116 25313
rect 47979 25220 48021 25229
rect 47979 25180 47980 25220
rect 48020 25180 48021 25220
rect 47979 25171 48021 25180
rect 47499 24632 47541 24641
rect 47499 24592 47500 24632
rect 47540 24592 47541 24632
rect 47499 24583 47541 24592
rect 47691 24632 47733 24641
rect 47691 24592 47692 24632
rect 47732 24592 47733 24632
rect 47691 24583 47733 24592
rect 47500 24498 47540 24583
rect 47595 24548 47637 24557
rect 47595 24508 47596 24548
rect 47636 24508 47637 24548
rect 47595 24499 47637 24508
rect 47404 23743 47444 23752
rect 47499 23792 47541 23801
rect 47499 23752 47500 23792
rect 47540 23752 47541 23792
rect 47499 23743 47541 23752
rect 47596 23792 47636 24499
rect 47596 23743 47636 23752
rect 47308 23658 47348 23743
rect 47500 23658 47540 23743
rect 47692 23120 47732 24583
rect 48076 23792 48116 25264
rect 48171 25304 48213 25313
rect 48171 25264 48172 25304
rect 48212 25264 48213 25304
rect 48171 25255 48213 25264
rect 48172 25170 48212 25255
rect 48268 25229 48308 25507
rect 48267 25220 48309 25229
rect 48267 25180 48268 25220
rect 48308 25180 48309 25220
rect 48267 25171 48309 25180
rect 48268 25132 48308 25171
rect 48268 25083 48308 25092
rect 48364 24968 48404 25684
rect 48459 25304 48501 25313
rect 48459 25264 48460 25304
rect 48500 25264 48501 25304
rect 48459 25255 48501 25264
rect 48268 24928 48404 24968
rect 48268 24557 48308 24928
rect 48267 24548 48309 24557
rect 48267 24508 48268 24548
rect 48308 24508 48309 24548
rect 48267 24499 48309 24508
rect 48172 23792 48212 23801
rect 48076 23752 48172 23792
rect 48172 23743 48212 23752
rect 48268 23792 48308 24499
rect 48268 23743 48308 23752
rect 48364 23792 48404 23801
rect 48364 23465 48404 23752
rect 48460 23792 48500 25255
rect 48556 24137 48596 27271
rect 48652 26405 48692 28288
rect 48843 27740 48885 27749
rect 48843 27700 48844 27740
rect 48884 27700 48885 27740
rect 48843 27691 48885 27700
rect 48747 27656 48789 27665
rect 48747 27616 48748 27656
rect 48788 27616 48789 27656
rect 48747 27607 48789 27616
rect 48748 27522 48788 27607
rect 48844 27497 48884 27691
rect 48843 27488 48885 27497
rect 48843 27448 48844 27488
rect 48884 27448 48885 27488
rect 48843 27439 48885 27448
rect 48651 26396 48693 26405
rect 48651 26356 48652 26396
rect 48692 26356 48693 26396
rect 48651 26347 48693 26356
rect 48940 25817 48980 29119
rect 49516 29084 49556 29791
rect 49708 29168 49748 29800
rect 49899 29800 49900 29840
rect 49940 29800 49941 29840
rect 49899 29791 49941 29800
rect 49708 29119 49748 29128
rect 49996 29084 50036 31396
rect 50380 31361 50420 31446
rect 50476 31436 50516 31471
rect 50379 31352 50421 31361
rect 50379 31312 50380 31352
rect 50420 31312 50421 31352
rect 50379 31303 50421 31312
rect 50476 31184 50516 31396
rect 50668 31436 50708 32656
rect 50668 31387 50708 31396
rect 50764 31352 50804 32824
rect 50860 32705 50900 33823
rect 51340 33704 51380 33823
rect 51724 33788 51764 34495
rect 52012 34460 52052 34469
rect 51916 34376 51956 34385
rect 51916 33872 51956 34336
rect 52012 34040 52052 34420
rect 52108 34410 52148 34495
rect 52203 34460 52245 34469
rect 52203 34420 52204 34460
rect 52244 34420 52245 34460
rect 52203 34411 52245 34420
rect 53067 34460 53109 34469
rect 53067 34420 53068 34460
rect 53108 34420 53109 34460
rect 53067 34411 53109 34420
rect 52204 34326 52244 34411
rect 52299 34376 52341 34385
rect 52299 34336 52300 34376
rect 52340 34336 52341 34376
rect 52299 34327 52341 34336
rect 52972 34376 53012 34385
rect 52300 34242 52340 34327
rect 52588 34292 52628 34301
rect 52628 34252 52916 34292
rect 52588 34243 52628 34252
rect 52352 34040 52720 34049
rect 52012 34000 52244 34040
rect 52012 33872 52052 33881
rect 51916 33832 52012 33872
rect 52012 33823 52052 33832
rect 51724 33739 51764 33748
rect 51340 33655 51380 33664
rect 51916 33704 51956 33713
rect 51916 33545 51956 33664
rect 52107 33704 52149 33713
rect 52107 33664 52108 33704
rect 52148 33664 52149 33704
rect 52107 33655 52149 33664
rect 51915 33536 51957 33545
rect 51915 33496 51916 33536
rect 51956 33496 51957 33536
rect 51915 33487 51957 33496
rect 51531 33452 51573 33461
rect 51531 33412 51532 33452
rect 51572 33412 51573 33452
rect 51531 33403 51573 33412
rect 52011 33452 52053 33461
rect 52011 33412 52012 33452
rect 52052 33412 52053 33452
rect 52011 33403 52053 33412
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 51532 33140 51572 33403
rect 52012 33318 52052 33403
rect 50955 33116 50997 33125
rect 50955 33076 50956 33116
rect 50996 33076 50997 33116
rect 50955 33067 50997 33076
rect 51436 33100 51572 33140
rect 52108 33116 52148 33655
rect 52204 33125 52244 34000
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 52299 33452 52341 33461
rect 52299 33412 52300 33452
rect 52340 33412 52341 33452
rect 52299 33403 52341 33412
rect 52300 33318 52340 33403
rect 50956 32982 50996 33067
rect 51339 32948 51381 32957
rect 51339 32908 51340 32948
rect 51380 32908 51381 32948
rect 51339 32899 51381 32908
rect 51243 32864 51285 32873
rect 51243 32824 51244 32864
rect 51284 32824 51285 32864
rect 51243 32815 51285 32824
rect 51340 32864 51380 32899
rect 51244 32730 51284 32815
rect 51340 32813 51380 32824
rect 50859 32696 50901 32705
rect 50859 32656 50860 32696
rect 50900 32656 50901 32696
rect 50859 32647 50901 32656
rect 51436 32692 51476 33100
rect 52108 33067 52148 33076
rect 52203 33116 52245 33125
rect 52203 33076 52204 33116
rect 52244 33076 52245 33116
rect 52203 33067 52245 33076
rect 51916 33032 51956 33041
rect 51820 32992 51916 33032
rect 51531 32948 51573 32957
rect 51531 32908 51532 32948
rect 51572 32908 51573 32948
rect 51531 32899 51573 32908
rect 50860 32192 50900 32647
rect 51436 32643 51476 32652
rect 50956 32192 50996 32201
rect 50860 32152 50956 32192
rect 50956 31688 50996 32152
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 50956 31648 51084 31688
rect 51044 31604 51084 31648
rect 51339 31604 51381 31613
rect 51532 31604 51572 32899
rect 51820 32192 51860 32992
rect 51916 32983 51956 32992
rect 52588 32864 52628 32873
rect 52588 32696 52628 32824
rect 52876 32864 52916 34252
rect 52972 33881 53012 34336
rect 52971 33872 53013 33881
rect 52971 33832 52972 33872
rect 53012 33832 53013 33872
rect 52971 33823 53013 33832
rect 53068 33125 53108 34411
rect 55180 34385 55220 34470
rect 55468 34385 55508 35176
rect 56140 34637 56180 35848
rect 56236 35888 56276 35897
rect 56139 34628 56181 34637
rect 56139 34588 56140 34628
rect 56180 34588 56181 34628
rect 56236 34628 56276 35848
rect 56524 35720 56564 36679
rect 56620 36317 56660 36688
rect 56619 36308 56661 36317
rect 56619 36268 56620 36308
rect 56660 36268 56661 36308
rect 56619 36259 56661 36268
rect 56812 36140 56852 37444
rect 57100 37484 57140 37493
rect 56908 37400 56948 37409
rect 56908 36989 56948 37360
rect 57003 37400 57045 37409
rect 57003 37360 57004 37400
rect 57044 37360 57045 37400
rect 57003 37351 57045 37360
rect 56907 36980 56949 36989
rect 56907 36940 56908 36980
rect 56948 36940 56949 36980
rect 56907 36931 56949 36940
rect 56620 36100 56852 36140
rect 56620 35813 56660 36100
rect 56715 35888 56757 35897
rect 56715 35848 56716 35888
rect 56756 35848 56757 35888
rect 56715 35839 56757 35848
rect 56812 35888 56852 35897
rect 56619 35804 56661 35813
rect 56619 35764 56620 35804
rect 56660 35764 56661 35804
rect 56619 35755 56661 35764
rect 56716 35754 56756 35839
rect 56428 35680 56564 35720
rect 56332 35216 56372 35225
rect 56428 35216 56468 35680
rect 56812 35645 56852 35848
rect 56908 35716 56948 35725
rect 57004 35716 57044 37351
rect 57100 36233 57140 37444
rect 57580 37409 57620 37948
rect 57579 37400 57621 37409
rect 57579 37360 57580 37400
rect 57620 37360 57621 37400
rect 57292 37325 57332 37356
rect 57579 37351 57621 37360
rect 57291 37316 57333 37325
rect 57291 37276 57292 37316
rect 57332 37276 57333 37316
rect 57291 37267 57333 37276
rect 57292 37232 57332 37267
rect 57292 36317 57332 37192
rect 57483 37232 57525 37241
rect 57483 37192 57484 37232
rect 57524 37192 57525 37232
rect 57483 37183 57525 37192
rect 57963 37232 58005 37241
rect 57963 37192 57964 37232
rect 58004 37192 58005 37232
rect 57963 37183 58005 37192
rect 57484 37098 57524 37183
rect 57579 36980 57621 36989
rect 57579 36940 57580 36980
rect 57620 36940 57621 36980
rect 57579 36931 57621 36940
rect 57483 36728 57525 36737
rect 57483 36688 57484 36728
rect 57524 36688 57525 36728
rect 57483 36679 57525 36688
rect 57484 36594 57524 36679
rect 57291 36308 57333 36317
rect 57291 36268 57292 36308
rect 57332 36268 57333 36308
rect 57291 36259 57333 36268
rect 57099 36224 57141 36233
rect 57099 36184 57100 36224
rect 57140 36184 57141 36224
rect 57099 36175 57141 36184
rect 57292 35932 57524 35972
rect 57099 35888 57141 35897
rect 57099 35848 57100 35888
rect 57140 35848 57141 35888
rect 57099 35839 57141 35848
rect 57196 35888 57236 35897
rect 57100 35754 57140 35839
rect 56948 35676 57044 35716
rect 56908 35667 56948 35676
rect 56619 35636 56661 35645
rect 56619 35596 56620 35636
rect 56660 35596 56661 35636
rect 56619 35587 56661 35596
rect 56811 35636 56853 35645
rect 56811 35596 56812 35636
rect 56852 35596 56853 35636
rect 56811 35587 56853 35596
rect 56372 35176 56468 35216
rect 56332 35167 56372 35176
rect 56236 34588 56372 34628
rect 56139 34579 56181 34588
rect 55947 34544 55989 34553
rect 55947 34504 55948 34544
rect 55988 34504 55989 34544
rect 55947 34495 55989 34504
rect 53836 34376 53876 34385
rect 53836 33713 53876 34336
rect 54123 34376 54165 34385
rect 54123 34336 54124 34376
rect 54164 34336 54165 34376
rect 54123 34327 54165 34336
rect 55179 34376 55221 34385
rect 55179 34336 55180 34376
rect 55220 34336 55221 34376
rect 55179 34327 55221 34336
rect 55467 34376 55509 34385
rect 55467 34336 55468 34376
rect 55508 34336 55509 34376
rect 55467 34327 55509 34336
rect 55948 34376 55988 34495
rect 55948 34327 55988 34336
rect 56043 34376 56085 34385
rect 56043 34336 56044 34376
rect 56084 34336 56085 34376
rect 56043 34327 56085 34336
rect 56140 34376 56180 34387
rect 53451 33704 53493 33713
rect 53451 33664 53452 33704
rect 53492 33664 53493 33704
rect 53451 33655 53493 33664
rect 53835 33704 53877 33713
rect 53835 33664 53836 33704
rect 53876 33664 53877 33704
rect 53835 33655 53877 33664
rect 53452 33570 53492 33655
rect 54124 33461 54164 34327
rect 56044 34242 56084 34327
rect 56140 34301 56180 34336
rect 56139 34292 56181 34301
rect 56139 34252 56140 34292
rect 56180 34252 56181 34292
rect 56139 34243 56181 34252
rect 54988 34208 55028 34217
rect 55276 34208 55316 34217
rect 55852 34208 55892 34217
rect 54700 34168 54988 34208
rect 54315 34124 54357 34133
rect 54315 34084 54316 34124
rect 54356 34084 54357 34124
rect 54315 34075 54357 34084
rect 54316 33881 54356 34075
rect 54315 33872 54357 33881
rect 54700 33872 54740 34168
rect 54988 34159 55028 34168
rect 55084 34168 55276 34208
rect 55084 33881 55124 34168
rect 55276 34159 55316 34168
rect 55372 34168 55852 34208
rect 55372 33956 55412 34168
rect 55852 34159 55892 34168
rect 56043 34124 56085 34133
rect 56043 34084 56044 34124
rect 56084 34084 56085 34124
rect 56043 34075 56085 34084
rect 55276 33916 55412 33956
rect 54315 33832 54316 33872
rect 54356 33832 54357 33872
rect 54315 33823 54357 33832
rect 54604 33832 54740 33872
rect 55083 33872 55125 33881
rect 55083 33832 55084 33872
rect 55124 33832 55125 33872
rect 54316 33704 54356 33823
rect 54316 33655 54356 33664
rect 54604 33536 54644 33832
rect 55083 33823 55125 33832
rect 54700 33704 54740 33713
rect 54740 33664 54836 33704
rect 54700 33655 54740 33664
rect 54604 33496 54740 33536
rect 54123 33452 54165 33461
rect 54123 33412 54124 33452
rect 54164 33412 54165 33452
rect 54123 33403 54165 33412
rect 53067 33116 53109 33125
rect 53067 33076 53068 33116
rect 53108 33076 53109 33116
rect 53067 33067 53109 33076
rect 53835 33116 53877 33125
rect 53835 33076 53836 33116
rect 53876 33076 53877 33116
rect 53835 33067 53877 33076
rect 52971 33032 53013 33041
rect 52971 32992 52972 33032
rect 53012 32992 53013 33032
rect 52971 32983 53013 32992
rect 52876 32815 52916 32824
rect 52972 32864 53012 32983
rect 53644 32957 53684 32988
rect 53836 32982 53876 33067
rect 53643 32948 53685 32957
rect 53643 32908 53644 32948
rect 53684 32908 53685 32948
rect 53643 32899 53685 32908
rect 54027 32948 54069 32957
rect 54027 32908 54028 32948
rect 54068 32908 54069 32948
rect 54027 32899 54069 32908
rect 52972 32815 53012 32824
rect 53068 32864 53108 32873
rect 52588 32656 52820 32696
rect 52011 32612 52053 32621
rect 52011 32572 52012 32612
rect 52052 32572 52053 32612
rect 52011 32563 52053 32572
rect 51820 32143 51860 32152
rect 51820 31604 51860 31613
rect 51915 31604 51957 31613
rect 51044 31564 51092 31604
rect 50955 31520 50997 31529
rect 50955 31480 50956 31520
rect 50996 31480 50997 31520
rect 50955 31471 50997 31480
rect 50956 31386 50996 31471
rect 50764 31277 50804 31312
rect 50763 31268 50805 31277
rect 50763 31228 50764 31268
rect 50804 31228 50805 31268
rect 50763 31219 50805 31228
rect 50955 31268 50997 31277
rect 50955 31228 50956 31268
rect 50996 31228 50997 31268
rect 50955 31219 50997 31228
rect 50284 31144 50516 31184
rect 50187 30680 50229 30689
rect 50187 30640 50188 30680
rect 50228 30640 50229 30680
rect 50187 30631 50229 30640
rect 50284 30680 50324 31144
rect 50956 31126 50996 31219
rect 50860 31086 50996 31126
rect 50284 30631 50324 30640
rect 50380 30680 50420 30689
rect 50188 30546 50228 30631
rect 50380 30353 50420 30640
rect 50476 30680 50516 30689
rect 50379 30344 50421 30353
rect 50379 30304 50380 30344
rect 50420 30304 50421 30344
rect 50379 30295 50421 30304
rect 50476 29681 50516 30640
rect 50667 30680 50709 30689
rect 50667 30640 50668 30680
rect 50708 30640 50709 30680
rect 50667 30631 50709 30640
rect 50668 30546 50708 30631
rect 50475 29672 50517 29681
rect 50475 29632 50476 29672
rect 50516 29632 50517 29672
rect 50475 29623 50517 29632
rect 50764 29672 50804 29681
rect 49516 28925 49556 29044
rect 49900 29044 50036 29084
rect 50572 29168 50612 29177
rect 49707 29000 49749 29009
rect 49707 28960 49708 29000
rect 49748 28960 49749 29000
rect 49707 28951 49749 28960
rect 49324 28916 49364 28925
rect 49132 28876 49324 28916
rect 49132 27656 49172 28876
rect 49324 28867 49364 28876
rect 49515 28916 49557 28925
rect 49515 28876 49516 28916
rect 49556 28876 49557 28916
rect 49515 28867 49557 28876
rect 49708 28580 49748 28951
rect 49708 28531 49748 28540
rect 49132 27572 49172 27616
rect 49132 27532 49268 27572
rect 49131 27404 49173 27413
rect 49131 27364 49132 27404
rect 49172 27364 49173 27404
rect 49131 27355 49173 27364
rect 49132 27068 49172 27355
rect 49228 27161 49268 27532
rect 49227 27152 49269 27161
rect 49227 27112 49228 27152
rect 49268 27112 49269 27152
rect 49227 27103 49269 27112
rect 49419 27152 49461 27161
rect 49419 27112 49420 27152
rect 49460 27112 49461 27152
rect 49419 27103 49461 27112
rect 49132 27019 49172 27028
rect 49036 26816 49076 26827
rect 49036 26741 49076 26776
rect 49035 26732 49077 26741
rect 49035 26692 49036 26732
rect 49076 26692 49077 26732
rect 49035 26683 49077 26692
rect 49131 26648 49173 26657
rect 49131 26608 49132 26648
rect 49172 26608 49173 26648
rect 49131 26599 49173 26608
rect 49132 26514 49172 26599
rect 49035 26144 49077 26153
rect 49035 26104 49036 26144
rect 49076 26104 49077 26144
rect 49035 26095 49077 26104
rect 49036 26010 49076 26095
rect 49035 25892 49077 25901
rect 49035 25852 49036 25892
rect 49076 25852 49077 25892
rect 49035 25843 49077 25852
rect 48939 25808 48981 25817
rect 48939 25768 48940 25808
rect 48980 25768 48981 25808
rect 48939 25759 48981 25768
rect 48844 24632 48884 24641
rect 48844 24473 48884 24592
rect 48939 24632 48981 24641
rect 48939 24592 48940 24632
rect 48980 24592 48981 24632
rect 48939 24583 48981 24592
rect 48843 24464 48885 24473
rect 48843 24424 48844 24464
rect 48884 24424 48885 24464
rect 48843 24415 48885 24424
rect 48652 24380 48692 24389
rect 48555 24128 48597 24137
rect 48555 24088 48556 24128
rect 48596 24088 48597 24128
rect 48555 24079 48597 24088
rect 48363 23456 48405 23465
rect 48363 23416 48364 23456
rect 48404 23416 48405 23456
rect 48363 23407 48405 23416
rect 47692 23071 47732 23080
rect 47212 23020 47444 23060
rect 47116 22483 47156 22492
rect 46868 22240 46964 22280
rect 47211 22280 47253 22289
rect 47211 22240 47212 22280
rect 47252 22240 47253 22280
rect 46828 22231 46868 22240
rect 47211 22231 47253 22240
rect 47404 22280 47444 23020
rect 46924 22054 46964 22063
rect 46924 21785 46964 22014
rect 47019 21860 47061 21869
rect 47019 21820 47020 21860
rect 47060 21820 47061 21860
rect 47019 21811 47061 21820
rect 46732 21727 46772 21736
rect 46923 21776 46965 21785
rect 46923 21736 46924 21776
rect 46964 21736 46965 21776
rect 46923 21727 46965 21736
rect 46828 21608 46868 21617
rect 46636 21568 46828 21608
rect 46540 21559 46580 21568
rect 46828 21559 46868 21568
rect 46923 21608 46965 21617
rect 46923 21568 46924 21608
rect 46964 21568 46965 21608
rect 46923 21559 46965 21568
rect 47020 21608 47060 21811
rect 47212 21701 47252 22231
rect 47404 22205 47444 22240
rect 47596 22280 47636 22289
rect 47403 22196 47445 22205
rect 47403 22156 47404 22196
rect 47444 22156 47445 22196
rect 47403 22147 47445 22156
rect 47500 22112 47540 22121
rect 47211 21692 47253 21701
rect 47211 21652 47212 21692
rect 47252 21652 47253 21692
rect 47211 21643 47253 21652
rect 47020 21559 47060 21568
rect 46443 21524 46485 21533
rect 46443 21484 46444 21524
rect 46484 21484 46485 21524
rect 46443 21475 46485 21484
rect 46348 21391 46388 21400
rect 46444 21390 46484 21475
rect 46924 21474 46964 21559
rect 47500 21533 47540 22072
rect 47499 21524 47541 21533
rect 47499 21484 47500 21524
rect 47540 21484 47541 21524
rect 47499 21475 47541 21484
rect 47403 21356 47445 21365
rect 47403 21316 47404 21356
rect 47444 21316 47445 21356
rect 47403 21307 47445 21316
rect 47404 21222 47444 21307
rect 47596 20936 47636 22240
rect 47692 22280 47732 22289
rect 47692 21365 47732 22240
rect 48460 21869 48500 23752
rect 48652 23465 48692 24340
rect 48747 23792 48789 23801
rect 48747 23752 48748 23792
rect 48788 23752 48789 23792
rect 48747 23743 48789 23752
rect 48844 23792 48884 23801
rect 48748 23658 48788 23743
rect 48844 23465 48884 23752
rect 48651 23456 48693 23465
rect 48651 23416 48652 23456
rect 48692 23416 48693 23456
rect 48651 23407 48693 23416
rect 48843 23456 48885 23465
rect 48843 23416 48844 23456
rect 48884 23416 48885 23456
rect 48843 23407 48885 23416
rect 48844 23288 48884 23297
rect 48940 23288 48980 24583
rect 48884 23248 48980 23288
rect 48844 23239 48884 23248
rect 48939 23120 48981 23129
rect 48939 23080 48940 23120
rect 48980 23080 48981 23120
rect 48939 23071 48981 23080
rect 48844 22868 48884 22877
rect 48844 22289 48884 22828
rect 48843 22280 48885 22289
rect 48843 22240 48844 22280
rect 48884 22240 48885 22280
rect 48843 22231 48885 22240
rect 48459 21860 48501 21869
rect 48459 21820 48460 21860
rect 48500 21820 48501 21860
rect 48459 21811 48501 21820
rect 48556 21608 48596 21617
rect 47691 21356 47733 21365
rect 47691 21316 47692 21356
rect 47732 21316 47733 21356
rect 47691 21307 47733 21316
rect 47596 20896 47924 20936
rect 46059 20852 46101 20861
rect 46059 20812 46060 20852
rect 46100 20812 46101 20852
rect 46059 20803 46101 20812
rect 46828 20852 46868 20861
rect 46636 20600 46676 20609
rect 46540 20560 46636 20600
rect 45388 20096 45428 20105
rect 45388 19760 45428 20056
rect 45771 20096 45813 20105
rect 45771 20056 45772 20096
rect 45812 20056 45813 20096
rect 45771 20047 45813 20056
rect 45772 19962 45812 20047
rect 45388 19720 45716 19760
rect 45292 19468 45524 19508
rect 45484 19349 45524 19468
rect 45579 19424 45621 19433
rect 45579 19384 45580 19424
rect 45620 19384 45621 19424
rect 45579 19375 45621 19384
rect 45676 19424 45716 19720
rect 46540 19517 46580 20560
rect 46636 20551 46676 20560
rect 46636 20096 46676 20105
rect 46539 19508 46581 19517
rect 46539 19468 46540 19508
rect 46580 19468 46581 19508
rect 46539 19459 46581 19468
rect 46156 19424 46196 19433
rect 45676 19375 45716 19384
rect 45772 19384 46156 19424
rect 45483 19340 45525 19349
rect 45483 19300 45484 19340
rect 45524 19300 45525 19340
rect 45483 19291 45525 19300
rect 45580 19340 45620 19375
rect 45484 19256 45524 19291
rect 45580 19289 45620 19300
rect 45772 19340 45812 19384
rect 45772 19291 45812 19300
rect 45484 19206 45524 19216
rect 45867 19256 45909 19265
rect 45867 19216 45868 19256
rect 45908 19216 45909 19256
rect 45867 19207 45909 19216
rect 45868 19122 45908 19207
rect 45292 19088 45332 19097
rect 45292 18929 45332 19048
rect 45771 19004 45813 19013
rect 45771 18964 45772 19004
rect 45812 18964 45813 19004
rect 45771 18955 45813 18964
rect 45291 18920 45333 18929
rect 45291 18880 45292 18920
rect 45332 18880 45333 18920
rect 45291 18871 45333 18880
rect 45195 18500 45237 18509
rect 45195 18460 45196 18500
rect 45236 18460 45237 18500
rect 45195 18451 45237 18460
rect 45387 18500 45429 18509
rect 45387 18460 45388 18500
rect 45428 18460 45429 18500
rect 45387 18451 45429 18460
rect 45099 18332 45141 18341
rect 45099 18292 45100 18332
rect 45140 18292 45141 18332
rect 45099 18283 45141 18292
rect 45100 17753 45140 18283
rect 45099 17744 45141 17753
rect 45099 17704 45100 17744
rect 45140 17704 45141 17744
rect 45099 17695 45141 17704
rect 45100 17610 45140 17695
rect 45004 17576 45044 17585
rect 45004 16997 45044 17536
rect 45003 16988 45045 16997
rect 45003 16948 45004 16988
rect 45044 16948 45045 16988
rect 45003 16939 45045 16948
rect 45004 16409 45044 16939
rect 45388 16745 45428 18451
rect 45483 17072 45525 17081
rect 45483 17032 45484 17072
rect 45524 17032 45525 17072
rect 45483 17023 45525 17032
rect 45387 16736 45429 16745
rect 45387 16696 45388 16736
rect 45428 16696 45429 16736
rect 45387 16687 45429 16696
rect 45484 16484 45524 17023
rect 45772 16988 45812 18955
rect 46060 17576 46100 19384
rect 46156 19375 46196 19384
rect 46444 19256 46484 19265
rect 46347 18920 46389 18929
rect 46347 18880 46348 18920
rect 46388 18880 46389 18920
rect 46444 18920 46484 19216
rect 46540 19256 46580 19459
rect 46540 19207 46580 19216
rect 46636 19181 46676 20056
rect 46828 19685 46868 20812
rect 47211 20768 47253 20777
rect 47211 20728 47212 20768
rect 47252 20728 47253 20768
rect 47211 20719 47253 20728
rect 47787 20768 47829 20777
rect 47787 20728 47788 20768
rect 47828 20728 47829 20768
rect 47787 20719 47829 20728
rect 47212 20634 47252 20719
rect 47116 20600 47156 20609
rect 46827 19676 46869 19685
rect 46827 19636 46828 19676
rect 46868 19636 46869 19676
rect 46827 19627 46869 19636
rect 47116 19433 47156 20560
rect 47788 20012 47828 20719
rect 47884 20189 47924 20896
rect 48556 20768 48596 21568
rect 48844 20768 48884 20777
rect 48556 20728 48844 20768
rect 48844 20719 48884 20728
rect 47883 20180 47925 20189
rect 47883 20140 47884 20180
rect 47924 20140 47925 20180
rect 47883 20131 47925 20140
rect 47499 19592 47541 19601
rect 47499 19552 47500 19592
rect 47540 19552 47541 19592
rect 47499 19543 47541 19552
rect 47211 19508 47253 19517
rect 47211 19468 47212 19508
rect 47252 19468 47253 19508
rect 47211 19459 47253 19468
rect 46731 19424 46773 19433
rect 46731 19384 46732 19424
rect 46772 19384 46773 19424
rect 46731 19375 46773 19384
rect 47115 19424 47157 19433
rect 47115 19384 47116 19424
rect 47156 19384 47157 19424
rect 47115 19375 47157 19384
rect 46732 19265 46772 19375
rect 46731 19256 46773 19265
rect 46731 19216 46732 19256
rect 46772 19216 46773 19256
rect 46731 19207 46773 19216
rect 46924 19256 46964 19265
rect 46635 19172 46677 19181
rect 46635 19132 46636 19172
rect 46676 19132 46677 19172
rect 46635 19123 46677 19132
rect 46636 19030 46676 19039
rect 46732 19004 46772 19207
rect 46676 18990 46772 19004
rect 46636 18964 46772 18990
rect 46828 19088 46868 19097
rect 46828 18920 46868 19048
rect 46924 18929 46964 19216
rect 47020 19256 47060 19267
rect 47020 19181 47060 19216
rect 47116 19256 47156 19265
rect 47212 19256 47252 19459
rect 47500 19340 47540 19543
rect 47500 19291 47540 19300
rect 47156 19216 47252 19256
rect 47788 19256 47828 19972
rect 47019 19172 47061 19181
rect 47019 19132 47020 19172
rect 47060 19132 47061 19172
rect 47019 19123 47061 19132
rect 46444 18880 46868 18920
rect 46923 18920 46965 18929
rect 46923 18880 46924 18920
rect 46964 18880 46965 18920
rect 46347 18871 46389 18880
rect 46923 18871 46965 18880
rect 46348 18752 46388 18871
rect 46539 18752 46581 18761
rect 46348 18712 46484 18752
rect 46348 18584 46388 18593
rect 46252 18544 46348 18584
rect 46155 18332 46197 18341
rect 46155 18292 46156 18332
rect 46196 18292 46197 18332
rect 46155 18283 46197 18292
rect 46156 18198 46196 18283
rect 46252 18080 46292 18544
rect 46348 18535 46388 18544
rect 46156 18040 46292 18080
rect 46156 17744 46196 18040
rect 46444 17753 46484 18712
rect 46539 18712 46540 18752
rect 46580 18712 46581 18752
rect 46539 18703 46581 18712
rect 46156 17695 46196 17704
rect 46252 17744 46292 17753
rect 46252 17576 46292 17704
rect 46060 17536 46292 17576
rect 46348 17744 46388 17753
rect 46348 17501 46388 17704
rect 46443 17744 46485 17753
rect 46443 17704 46444 17744
rect 46484 17704 46485 17744
rect 46443 17695 46485 17704
rect 46444 17610 46484 17695
rect 46347 17492 46389 17501
rect 46347 17452 46348 17492
rect 46388 17452 46389 17492
rect 46347 17443 46389 17452
rect 46540 17324 46580 18703
rect 46732 18584 46772 18593
rect 47019 18584 47061 18593
rect 46772 18544 47020 18584
rect 47060 18544 47061 18584
rect 46732 18535 46772 18544
rect 47019 18535 47061 18544
rect 46731 17744 46773 17753
rect 46731 17704 46732 17744
rect 46772 17704 46773 17744
rect 46731 17695 46773 17704
rect 46156 17284 46580 17324
rect 46156 17072 46196 17284
rect 46156 17023 46196 17032
rect 46251 17072 46293 17081
rect 46251 17032 46252 17072
rect 46292 17032 46293 17072
rect 46251 17023 46293 17032
rect 46348 17072 46388 17081
rect 45484 16435 45524 16444
rect 45580 16820 45620 16829
rect 45003 16400 45045 16409
rect 45003 16360 45004 16400
rect 45044 16360 45045 16400
rect 45003 16351 45045 16360
rect 45580 16073 45620 16780
rect 45579 16064 45621 16073
rect 45579 16024 45580 16064
rect 45620 16024 45621 16064
rect 45579 16015 45621 16024
rect 45772 15728 45812 16948
rect 46252 16938 46292 17023
rect 45964 16829 46004 16914
rect 45963 16820 46005 16829
rect 45963 16780 45964 16820
rect 46004 16780 46005 16820
rect 45963 16771 46005 16780
rect 45963 16568 46005 16577
rect 45963 16528 45964 16568
rect 46004 16528 46005 16568
rect 45963 16519 46005 16528
rect 45964 16232 46004 16519
rect 46348 16400 46388 17032
rect 46059 16316 46101 16325
rect 46059 16276 46060 16316
rect 46100 16276 46101 16316
rect 46059 16267 46101 16276
rect 45867 16064 45909 16073
rect 45867 16020 45868 16064
rect 45908 16020 45909 16064
rect 45867 16015 45909 16020
rect 45868 15905 45908 16015
rect 45867 15896 45909 15905
rect 45867 15856 45868 15896
rect 45908 15856 45909 15896
rect 45964 15896 46004 16192
rect 46060 16232 46100 16267
rect 46060 16181 46100 16192
rect 46251 16232 46293 16241
rect 46251 16192 46252 16232
rect 46292 16192 46293 16232
rect 46251 16183 46293 16192
rect 45964 15856 46100 15896
rect 45867 15847 45909 15856
rect 45772 15688 46004 15728
rect 45676 15560 45716 15569
rect 45716 15520 45812 15560
rect 45676 15511 45716 15520
rect 45003 15308 45045 15317
rect 45003 15268 45004 15308
rect 45044 15268 45045 15308
rect 45003 15259 45045 15268
rect 45004 15174 45044 15259
rect 45675 14804 45717 14813
rect 45675 14764 45676 14804
rect 45716 14764 45717 14804
rect 45675 14755 45717 14764
rect 45484 14720 45524 14729
rect 45387 14636 45429 14645
rect 45387 14596 45388 14636
rect 45428 14596 45429 14636
rect 45387 14587 45429 14596
rect 45388 14502 45428 14587
rect 45484 14477 45524 14680
rect 45579 14720 45621 14729
rect 45579 14680 45580 14720
rect 45620 14680 45621 14720
rect 45579 14671 45621 14680
rect 45676 14720 45716 14755
rect 45580 14586 45620 14671
rect 45676 14669 45716 14680
rect 45483 14468 45525 14477
rect 45483 14428 45484 14468
rect 45524 14428 45525 14468
rect 45483 14419 45525 14428
rect 45772 14393 45812 15520
rect 45867 14636 45909 14645
rect 45867 14596 45868 14636
rect 45908 14596 45909 14636
rect 45867 14587 45909 14596
rect 45868 14502 45908 14587
rect 45771 14384 45813 14393
rect 45771 14344 45772 14384
rect 45812 14344 45813 14384
rect 45771 14335 45813 14344
rect 45195 14216 45237 14225
rect 45195 14176 45196 14216
rect 45236 14176 45237 14216
rect 45195 14167 45237 14176
rect 45292 14220 45332 14229
rect 45332 14180 45524 14220
rect 45292 14171 45332 14180
rect 45099 14132 45141 14141
rect 45099 14092 45100 14132
rect 45140 14092 45141 14132
rect 45099 14083 45141 14092
rect 45100 14048 45140 14083
rect 45100 13997 45140 14008
rect 45196 14048 45236 14167
rect 45196 13999 45236 14008
rect 44908 13840 45140 13880
rect 44044 13124 44084 13133
rect 43756 13040 43796 13049
rect 43756 12545 43796 13000
rect 44044 12713 44084 13084
rect 44619 13124 44661 13133
rect 44619 13084 44620 13124
rect 44660 13084 44661 13124
rect 44619 13075 44661 13084
rect 44043 12704 44085 12713
rect 44043 12664 44044 12704
rect 44084 12664 44085 12704
rect 44043 12655 44085 12664
rect 44619 12704 44661 12713
rect 44619 12664 44620 12704
rect 44660 12664 44661 12704
rect 44619 12655 44661 12664
rect 43947 12620 43989 12629
rect 43947 12580 43948 12620
rect 43988 12580 43989 12620
rect 44427 12620 44469 12629
rect 43947 12578 43989 12580
rect 44044 12578 44084 12587
rect 44427 12580 44428 12620
rect 44468 12580 44469 12620
rect 43947 12571 44044 12578
rect 43755 12536 43797 12545
rect 43755 12496 43756 12536
rect 43796 12496 43797 12536
rect 43755 12487 43797 12496
rect 43852 12536 43892 12545
rect 43948 12538 44044 12571
rect 44084 12538 44180 12578
rect 44427 12571 44469 12580
rect 44044 12529 44084 12538
rect 43756 12402 43796 12487
rect 43852 12293 43892 12496
rect 44044 12377 44084 12462
rect 44043 12368 44085 12377
rect 44043 12328 44044 12368
rect 44084 12328 44085 12368
rect 44043 12319 44085 12328
rect 43851 12284 43893 12293
rect 43851 12244 43852 12284
rect 43892 12244 43893 12284
rect 43851 12235 43893 12244
rect 43660 12076 43988 12116
rect 43563 12067 43605 12076
rect 43659 11780 43701 11789
rect 43659 11740 43660 11780
rect 43700 11740 43796 11780
rect 43659 11731 43701 11740
rect 43660 11646 43700 11731
rect 43275 11360 43317 11369
rect 43275 11320 43276 11360
rect 43316 11320 43317 11360
rect 43275 11311 43317 11320
rect 43756 11276 43796 11740
rect 43851 11528 43893 11537
rect 43851 11488 43852 11528
rect 43892 11488 43893 11528
rect 43851 11479 43893 11488
rect 43852 11394 43892 11479
rect 43756 11236 43892 11276
rect 43468 11196 43508 11205
rect 42795 11108 42837 11117
rect 42795 11068 42796 11108
rect 42836 11068 42837 11108
rect 42795 11059 42837 11068
rect 43275 11108 43317 11117
rect 43275 11068 43276 11108
rect 43316 11068 43317 11108
rect 43275 11059 43317 11068
rect 42700 10975 42740 10984
rect 42796 11024 42836 11059
rect 42604 10890 42644 10975
rect 42796 10973 42836 10984
rect 42987 11024 43029 11033
rect 42987 10984 42988 11024
rect 43028 10984 43029 11024
rect 42987 10975 43029 10984
rect 43276 11024 43316 11059
rect 42988 10772 43028 10975
rect 43276 10973 43316 10984
rect 43372 11024 43412 11035
rect 43372 10949 43412 10984
rect 43371 10940 43413 10949
rect 43371 10900 43372 10940
rect 43412 10900 43413 10940
rect 43371 10891 43413 10900
rect 42988 10688 43028 10732
rect 43371 10772 43413 10781
rect 43371 10732 43372 10772
rect 43412 10732 43413 10772
rect 43371 10723 43413 10732
rect 42988 10648 43221 10688
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 42603 10352 42645 10361
rect 42603 10312 42604 10352
rect 42644 10312 42645 10352
rect 42603 10303 42645 10312
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 42604 9596 42644 10303
rect 43181 10278 43221 10648
rect 43275 10352 43317 10361
rect 43275 10312 43276 10352
rect 43316 10312 43317 10352
rect 43275 10303 43317 10312
rect 43181 10229 43221 10238
rect 43276 10218 43316 10303
rect 43372 10268 43412 10723
rect 43468 10688 43508 11156
rect 43659 11108 43701 11117
rect 43659 11068 43660 11108
rect 43700 11068 43701 11108
rect 43659 11059 43701 11068
rect 43660 10974 43700 11059
rect 43755 11024 43797 11033
rect 43755 10984 43756 11024
rect 43796 10984 43797 11024
rect 43755 10975 43797 10984
rect 43852 11024 43892 11236
rect 43852 10975 43892 10984
rect 43948 11024 43988 12076
rect 43948 10975 43988 10984
rect 44140 11024 44180 12538
rect 44428 12536 44468 12571
rect 44428 12485 44468 12496
rect 44524 12452 44564 12461
rect 44427 12368 44469 12377
rect 44524 12368 44564 12412
rect 44427 12328 44428 12368
rect 44468 12328 44564 12368
rect 44620 12368 44660 12655
rect 44716 12452 44756 13840
rect 44812 13831 44852 13840
rect 45003 13208 45045 13217
rect 45003 13168 45004 13208
rect 45044 13168 45045 13208
rect 45003 13159 45045 13168
rect 44907 13124 44949 13133
rect 44907 13084 44908 13124
rect 44948 13084 44949 13124
rect 44907 13075 44949 13084
rect 44811 13040 44853 13049
rect 44811 13000 44812 13040
rect 44852 13000 44853 13040
rect 44811 12991 44853 13000
rect 44812 12536 44852 12991
rect 44812 12487 44852 12496
rect 44716 12403 44756 12412
rect 44427 12319 44469 12328
rect 44620 12319 44660 12328
rect 44715 12284 44757 12293
rect 44715 12244 44716 12284
rect 44756 12244 44757 12284
rect 44715 12235 44757 12244
rect 44619 12116 44661 12125
rect 44619 12076 44620 12116
rect 44660 12076 44661 12116
rect 44619 12067 44661 12076
rect 44427 11528 44469 11537
rect 44427 11488 44428 11528
rect 44468 11488 44469 11528
rect 44427 11479 44469 11488
rect 44331 11276 44373 11285
rect 44331 11236 44332 11276
rect 44372 11236 44373 11276
rect 44331 11227 44373 11236
rect 44140 10975 44180 10984
rect 44332 11024 44372 11227
rect 44428 11117 44468 11479
rect 44427 11108 44469 11117
rect 44427 11068 44428 11108
rect 44468 11068 44469 11108
rect 44427 11059 44469 11068
rect 43756 10890 43796 10975
rect 44139 10772 44181 10781
rect 44139 10732 44140 10772
rect 44180 10732 44181 10772
rect 44139 10723 44181 10732
rect 43468 10648 43604 10688
rect 43372 10219 43412 10228
rect 43467 10268 43509 10277
rect 43467 10228 43468 10268
rect 43508 10228 43509 10268
rect 43467 10219 43509 10228
rect 43083 10184 43125 10193
rect 43083 10144 43084 10184
rect 43124 10144 43125 10184
rect 43083 10135 43125 10144
rect 43468 10184 43508 10219
rect 43564 10193 43604 10648
rect 44140 10638 44180 10723
rect 43084 10050 43124 10135
rect 43468 10133 43508 10144
rect 43563 10184 43605 10193
rect 43563 10144 43564 10184
rect 43604 10144 43605 10184
rect 43563 10135 43605 10144
rect 44043 10184 44085 10193
rect 44140 10184 44180 10193
rect 44043 10144 44044 10184
rect 44084 10144 44140 10184
rect 44043 10135 44085 10144
rect 44140 10135 44180 10144
rect 44235 10184 44277 10193
rect 44235 10144 44236 10184
rect 44276 10144 44277 10184
rect 44235 10135 44277 10144
rect 43851 10100 43893 10109
rect 43851 10060 43852 10100
rect 43892 10060 43893 10100
rect 43851 10051 43893 10060
rect 42987 10016 43029 10025
rect 42987 9976 42988 10016
rect 43028 9976 43029 10016
rect 42987 9967 43029 9976
rect 42604 9547 42644 9556
rect 42988 9512 43028 9967
rect 42988 9463 43028 9472
rect 43852 9512 43892 10051
rect 44236 10050 44276 10135
rect 43852 9463 43892 9472
rect 29451 9428 29493 9437
rect 29451 9388 29452 9428
rect 29492 9388 29493 9428
rect 29451 9379 29493 9388
rect 31755 9428 31797 9437
rect 31755 9388 31756 9428
rect 31796 9388 31797 9428
rect 31755 9379 31797 9388
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 44332 8840 44372 10984
rect 44428 11024 44468 11059
rect 44428 10974 44468 10984
rect 44524 10268 44564 10296
rect 44620 10268 44660 12067
rect 44564 10228 44660 10268
rect 44524 10219 44564 10228
rect 44620 9353 44660 10228
rect 44716 10436 44756 12235
rect 44619 9344 44661 9353
rect 44619 9304 44620 9344
rect 44660 9304 44661 9344
rect 44619 9295 44661 9304
rect 44716 9176 44756 10396
rect 44811 10184 44853 10193
rect 44811 10144 44812 10184
rect 44852 10144 44853 10184
rect 44811 10135 44853 10144
rect 44908 10184 44948 13075
rect 45004 11696 45044 13159
rect 45004 11647 45044 11656
rect 45100 10361 45140 13840
rect 45291 13208 45333 13217
rect 45291 13168 45292 13208
rect 45332 13168 45333 13208
rect 45291 13159 45333 13168
rect 45292 13074 45332 13159
rect 45484 13049 45524 14180
rect 45579 14048 45621 14057
rect 45579 14008 45580 14048
rect 45620 14008 45621 14048
rect 45579 13999 45621 14008
rect 45580 13914 45620 13999
rect 45772 13796 45812 14335
rect 45868 13796 45908 13805
rect 45772 13756 45868 13796
rect 45868 13217 45908 13756
rect 45867 13208 45909 13217
rect 45867 13168 45868 13208
rect 45908 13168 45909 13208
rect 45867 13159 45909 13168
rect 45483 13040 45525 13049
rect 45483 13000 45484 13040
rect 45524 13000 45525 13040
rect 45483 12991 45525 13000
rect 45867 13040 45909 13049
rect 45867 13000 45868 13040
rect 45908 13000 45909 13040
rect 45867 12991 45909 13000
rect 45387 12788 45429 12797
rect 45387 12748 45388 12788
rect 45428 12748 45429 12788
rect 45387 12739 45429 12748
rect 45099 10352 45141 10361
rect 45099 10312 45100 10352
rect 45140 10312 45141 10352
rect 45099 10303 45141 10312
rect 45388 10277 45428 12739
rect 45484 12704 45524 12991
rect 45580 12704 45620 12713
rect 45484 12664 45580 12704
rect 45580 12655 45620 12664
rect 45676 12536 45716 12545
rect 45868 12536 45908 12991
rect 45964 12797 46004 15688
rect 46060 14225 46100 15856
rect 46252 14720 46292 16183
rect 46348 15485 46388 16360
rect 46444 17072 46484 17081
rect 46444 16232 46484 17032
rect 46636 17072 46676 17081
rect 46636 16325 46676 17032
rect 46732 17072 46772 17695
rect 46923 17408 46965 17417
rect 46923 17368 46924 17408
rect 46964 17368 46965 17408
rect 46923 17359 46965 17368
rect 46635 16316 46677 16325
rect 46635 16276 46636 16316
rect 46676 16276 46677 16316
rect 46635 16267 46677 16276
rect 46540 16232 46580 16241
rect 46444 16192 46540 16232
rect 46540 16183 46580 16192
rect 46732 16148 46772 17032
rect 46828 17072 46868 17083
rect 46828 16997 46868 17032
rect 46924 17072 46964 17359
rect 46827 16988 46869 16997
rect 46827 16948 46828 16988
rect 46868 16948 46869 16988
rect 46827 16939 46869 16948
rect 46924 16577 46964 17032
rect 47020 16913 47060 18535
rect 47116 17417 47156 19216
rect 47788 19207 47828 19216
rect 47884 19256 47924 20131
rect 48364 20096 48404 20105
rect 48747 20096 48789 20105
rect 48404 20056 48500 20096
rect 48364 20047 48404 20056
rect 47979 20012 48021 20021
rect 47979 19972 47980 20012
rect 48020 19972 48021 20012
rect 47979 19963 48021 19972
rect 47884 19207 47924 19216
rect 47499 19172 47541 19181
rect 47499 19132 47500 19172
rect 47540 19132 47541 19172
rect 47499 19123 47541 19132
rect 47308 19088 47348 19097
rect 47308 18593 47348 19048
rect 47307 18584 47349 18593
rect 47307 18544 47308 18584
rect 47348 18544 47349 18584
rect 47307 18535 47349 18544
rect 47211 18332 47253 18341
rect 47211 18292 47212 18332
rect 47252 18292 47253 18332
rect 47211 18283 47253 18292
rect 47115 17408 47157 17417
rect 47115 17368 47116 17408
rect 47156 17368 47157 17408
rect 47115 17359 47157 17368
rect 47019 16904 47061 16913
rect 47019 16864 47020 16904
rect 47060 16864 47061 16904
rect 47019 16855 47061 16864
rect 46923 16568 46965 16577
rect 46923 16528 46924 16568
rect 46964 16528 46965 16568
rect 46923 16519 46965 16528
rect 46923 16232 46965 16241
rect 47020 16232 47060 16855
rect 47115 16820 47157 16829
rect 47115 16780 47116 16820
rect 47156 16780 47157 16820
rect 47115 16771 47157 16780
rect 46923 16192 46924 16232
rect 46964 16192 47060 16232
rect 46923 16183 46965 16192
rect 46636 16108 46772 16148
rect 46636 15653 46676 16108
rect 46924 16098 46964 16183
rect 46731 15896 46773 15905
rect 46731 15856 46732 15896
rect 46772 15856 46773 15896
rect 46731 15847 46773 15856
rect 46635 15644 46677 15653
rect 46635 15604 46636 15644
rect 46676 15604 46677 15644
rect 46635 15595 46677 15604
rect 46347 15476 46389 15485
rect 46347 15436 46348 15476
rect 46388 15436 46389 15476
rect 46347 15427 46389 15436
rect 46636 14813 46676 15595
rect 46732 15560 46772 15847
rect 46732 15511 46772 15520
rect 47116 15573 47156 16771
rect 47212 16661 47252 18283
rect 47500 17753 47540 19123
rect 47595 19088 47637 19097
rect 47595 19048 47596 19088
rect 47636 19048 47637 19088
rect 47595 19039 47637 19048
rect 47596 18584 47636 19039
rect 47636 18544 47828 18584
rect 47596 18535 47636 18544
rect 47499 17744 47541 17753
rect 47499 17704 47500 17744
rect 47540 17704 47541 17744
rect 47499 17695 47541 17704
rect 47500 17610 47540 17695
rect 47404 17576 47444 17587
rect 47404 17501 47444 17536
rect 47403 17492 47445 17501
rect 47403 17452 47404 17492
rect 47444 17452 47445 17492
rect 47403 17443 47445 17452
rect 47307 17072 47349 17081
rect 47307 17032 47308 17072
rect 47348 17032 47349 17072
rect 47307 17023 47349 17032
rect 47404 17072 47444 17081
rect 47308 16820 47348 17023
rect 47404 16997 47444 17032
rect 47403 16988 47445 16997
rect 47403 16948 47404 16988
rect 47444 16948 47445 16988
rect 47403 16939 47445 16948
rect 47211 16652 47253 16661
rect 47211 16612 47212 16652
rect 47252 16612 47253 16652
rect 47211 16603 47253 16612
rect 47308 16325 47348 16780
rect 47307 16316 47349 16325
rect 47307 16276 47308 16316
rect 47348 16276 47349 16316
rect 47307 16267 47349 16276
rect 47404 16073 47444 16939
rect 47692 16820 47732 16829
rect 47596 16780 47692 16820
rect 47596 16241 47636 16780
rect 47692 16771 47732 16780
rect 47595 16232 47637 16241
rect 47595 16192 47596 16232
rect 47636 16192 47637 16232
rect 47595 16183 47637 16192
rect 47788 16232 47828 18544
rect 47980 17669 48020 19963
rect 48076 19508 48116 19517
rect 48116 19468 48404 19508
rect 48076 19459 48116 19468
rect 48267 19340 48309 19349
rect 48267 19300 48268 19340
rect 48308 19300 48309 19340
rect 48267 19291 48309 19300
rect 48364 19340 48404 19468
rect 48460 19424 48500 20056
rect 48747 20056 48748 20096
rect 48788 20056 48789 20096
rect 48747 20047 48789 20056
rect 48748 19962 48788 20047
rect 48460 19375 48500 19384
rect 48364 19291 48404 19300
rect 48555 19340 48597 19349
rect 48555 19300 48556 19340
rect 48596 19300 48597 19340
rect 48555 19291 48597 19300
rect 48075 19256 48117 19265
rect 48075 19207 48076 19256
rect 48116 19207 48117 19256
rect 48268 19256 48308 19291
rect 48268 19205 48308 19216
rect 48556 19206 48596 19291
rect 48652 19256 48692 19265
rect 48076 19121 48116 19202
rect 48652 18845 48692 19216
rect 48843 19088 48885 19097
rect 48843 19048 48844 19088
rect 48884 19048 48885 19088
rect 48843 19039 48885 19048
rect 48651 18836 48693 18845
rect 48651 18796 48652 18836
rect 48692 18796 48693 18836
rect 48651 18787 48693 18796
rect 48555 18584 48597 18593
rect 48555 18544 48556 18584
rect 48596 18544 48597 18584
rect 48555 18535 48597 18544
rect 48556 18089 48596 18535
rect 48748 18332 48788 18341
rect 48652 18292 48748 18332
rect 48555 18080 48597 18089
rect 48555 18040 48556 18080
rect 48596 18040 48597 18080
rect 48555 18031 48597 18040
rect 48556 17828 48596 17837
rect 47979 17660 48021 17669
rect 47979 17620 47980 17660
rect 48020 17620 48021 17660
rect 47979 17611 48021 17620
rect 48556 17585 48596 17788
rect 48652 17753 48692 18292
rect 48748 18283 48788 18292
rect 48747 18080 48789 18089
rect 48747 18040 48748 18080
rect 48788 18040 48789 18080
rect 48747 18031 48789 18040
rect 48748 17996 48788 18031
rect 48748 17921 48788 17956
rect 48747 17912 48789 17921
rect 48747 17872 48748 17912
rect 48788 17872 48789 17912
rect 48747 17863 48789 17872
rect 48748 17832 48788 17863
rect 48651 17744 48693 17753
rect 48651 17704 48652 17744
rect 48692 17704 48693 17744
rect 48651 17695 48693 17704
rect 48555 17576 48597 17585
rect 48555 17536 48556 17576
rect 48596 17536 48597 17576
rect 48555 17527 48597 17536
rect 47788 16183 47828 16192
rect 47403 16064 47445 16073
rect 47403 16024 47404 16064
rect 47444 16024 47445 16064
rect 47403 16015 47445 16024
rect 47308 15573 47348 15600
rect 47116 15560 47348 15573
rect 47156 15533 47308 15560
rect 47116 15511 47156 15520
rect 47308 15485 47348 15520
rect 47499 15560 47541 15569
rect 47499 15520 47500 15560
rect 47540 15520 47541 15560
rect 47499 15511 47541 15520
rect 47596 15560 47636 16183
rect 47596 15511 47636 15520
rect 47787 15560 47829 15569
rect 47787 15520 47788 15560
rect 47828 15520 47829 15560
rect 47787 15511 47829 15520
rect 48267 15560 48309 15569
rect 48267 15520 48268 15560
rect 48308 15520 48309 15560
rect 48267 15511 48309 15520
rect 46827 15476 46869 15485
rect 46827 15436 46828 15476
rect 46868 15436 46869 15476
rect 46827 15427 46869 15436
rect 47020 15476 47060 15485
rect 46828 15342 46868 15427
rect 46923 15392 46965 15401
rect 46923 15352 46924 15392
rect 46964 15352 46965 15392
rect 46923 15343 46965 15352
rect 46924 15258 46964 15343
rect 47020 15308 47060 15436
rect 47307 15476 47349 15485
rect 47307 15436 47308 15476
rect 47348 15436 47349 15476
rect 47307 15427 47349 15436
rect 47500 15426 47540 15511
rect 47788 15426 47828 15511
rect 48075 15476 48117 15485
rect 48075 15436 48076 15476
rect 48116 15436 48117 15476
rect 48075 15427 48117 15436
rect 47883 15392 47925 15401
rect 47883 15352 47884 15392
rect 47924 15352 47925 15392
rect 47883 15343 47925 15352
rect 47308 15308 47348 15317
rect 47020 15268 47308 15308
rect 47308 15259 47348 15268
rect 47884 15258 47924 15343
rect 46635 14804 46677 14813
rect 46635 14764 46636 14804
rect 46676 14764 46677 14804
rect 46635 14755 46677 14764
rect 46827 14804 46869 14813
rect 46827 14764 46828 14804
rect 46868 14764 46869 14804
rect 46827 14755 46869 14764
rect 46252 14309 46292 14680
rect 46251 14300 46293 14309
rect 46251 14260 46252 14300
rect 46292 14260 46293 14300
rect 46251 14251 46293 14260
rect 46059 14216 46101 14225
rect 46059 14176 46060 14216
rect 46100 14176 46101 14216
rect 46059 14167 46101 14176
rect 46347 14216 46389 14225
rect 46347 14176 46348 14216
rect 46388 14176 46389 14216
rect 46347 14167 46389 14176
rect 46155 12872 46197 12881
rect 46155 12832 46156 12872
rect 46196 12832 46197 12872
rect 46155 12823 46197 12832
rect 45963 12788 46005 12797
rect 45963 12748 45964 12788
rect 46004 12748 46005 12788
rect 45963 12739 46005 12748
rect 45963 12620 46005 12629
rect 45963 12580 45964 12620
rect 46004 12580 46005 12620
rect 45963 12571 46005 12580
rect 45716 12496 45868 12536
rect 45676 12487 45716 12496
rect 45868 12487 45908 12496
rect 45964 12536 46004 12571
rect 45964 12485 46004 12496
rect 46059 12536 46101 12545
rect 46059 12496 46060 12536
rect 46100 12496 46101 12536
rect 46059 12487 46101 12496
rect 46156 12536 46196 12823
rect 46348 12536 46388 14167
rect 46731 14132 46773 14141
rect 46731 14092 46732 14132
rect 46772 14092 46773 14132
rect 46731 14083 46773 14092
rect 46539 14048 46581 14057
rect 46539 14008 46540 14048
rect 46580 14008 46581 14048
rect 46539 13999 46581 14008
rect 46540 13914 46580 13999
rect 46732 13998 46772 14083
rect 46828 14048 46868 14755
rect 47116 14720 47156 14729
rect 46923 14384 46965 14393
rect 46923 14344 46924 14384
rect 46964 14344 46965 14384
rect 46923 14335 46965 14344
rect 46828 13460 46868 14008
rect 46924 14048 46964 14335
rect 47019 14216 47061 14225
rect 47019 14176 47020 14216
rect 47060 14176 47061 14216
rect 47019 14167 47061 14176
rect 46924 13999 46964 14008
rect 47020 14048 47060 14167
rect 47116 14057 47156 14680
rect 47211 14300 47253 14309
rect 47211 14260 47212 14300
rect 47252 14260 47253 14300
rect 47211 14251 47253 14260
rect 47020 13999 47060 14008
rect 47115 14048 47157 14057
rect 47115 14008 47116 14048
rect 47156 14008 47157 14048
rect 47115 13999 47157 14008
rect 46828 13420 46964 13460
rect 46731 13376 46773 13385
rect 46731 13336 46732 13376
rect 46772 13336 46773 13376
rect 46731 13327 46773 13336
rect 46732 13208 46772 13327
rect 46732 13159 46772 13168
rect 46827 13208 46869 13217
rect 46827 13168 46828 13208
rect 46868 13168 46869 13208
rect 46827 13159 46869 13168
rect 46924 13208 46964 13420
rect 47019 13376 47061 13385
rect 47019 13336 47020 13376
rect 47060 13336 47061 13376
rect 47019 13327 47061 13336
rect 46444 13049 46484 13134
rect 46539 13124 46581 13133
rect 46539 13084 46540 13124
rect 46580 13084 46581 13124
rect 46539 13075 46581 13084
rect 46443 13040 46485 13049
rect 46443 13000 46444 13040
rect 46484 13000 46485 13040
rect 46443 12991 46485 13000
rect 46540 12788 46580 13075
rect 46828 13074 46868 13159
rect 46636 13040 46676 13049
rect 46636 12980 46676 13000
rect 46636 12940 46868 12980
rect 46196 12496 46292 12536
rect 46156 12487 46196 12496
rect 46060 12368 46100 12487
rect 45868 12328 46100 12368
rect 45771 11864 45813 11873
rect 45771 11824 45772 11864
rect 45812 11824 45813 11864
rect 45771 11815 45813 11824
rect 45675 11024 45717 11033
rect 45675 10984 45676 11024
rect 45716 10984 45717 11024
rect 45675 10975 45717 10984
rect 45676 10890 45716 10975
rect 45772 10940 45812 11815
rect 45868 11696 45908 12328
rect 46156 12284 46196 12293
rect 45868 11647 45908 11656
rect 45964 12244 46156 12284
rect 45867 11528 45909 11537
rect 45867 11488 45868 11528
rect 45908 11488 45909 11528
rect 45867 11479 45909 11488
rect 45772 10891 45812 10900
rect 45868 10856 45908 11479
rect 45964 10940 46004 12244
rect 46156 12235 46196 12244
rect 46252 12116 46292 12496
rect 46060 12076 46292 12116
rect 46060 11024 46100 12076
rect 46348 11696 46388 12496
rect 46444 12748 46580 12788
rect 46444 12536 46484 12748
rect 46444 12487 46484 12496
rect 46540 12664 46772 12704
rect 46540 12536 46580 12664
rect 46540 12487 46580 12496
rect 46636 12536 46676 12545
rect 46540 11696 46580 11705
rect 46348 11656 46540 11696
rect 46540 11647 46580 11656
rect 46636 11696 46676 12496
rect 46732 12452 46772 12664
rect 46828 12620 46868 12940
rect 46828 12571 46868 12580
rect 46924 12452 46964 13168
rect 46732 12412 46964 12452
rect 46923 11864 46965 11873
rect 47020 11864 47060 13327
rect 47212 12545 47252 14251
rect 47979 14048 48021 14057
rect 47979 14008 47980 14048
rect 48020 14008 48021 14048
rect 47979 13999 48021 14008
rect 48076 14048 48116 15427
rect 48268 14972 48308 15511
rect 48268 14923 48308 14932
rect 48268 14552 48308 14561
rect 48268 14393 48308 14512
rect 48267 14384 48309 14393
rect 48267 14344 48268 14384
rect 48308 14344 48309 14384
rect 48267 14335 48309 14344
rect 48652 14309 48692 17695
rect 48844 17072 48884 19039
rect 48940 17837 48980 23071
rect 49036 19256 49076 25843
rect 49131 25556 49173 25565
rect 49131 25516 49132 25556
rect 49172 25516 49173 25556
rect 49131 25507 49173 25516
rect 49132 25422 49172 25507
rect 49227 25304 49269 25313
rect 49227 25264 49228 25304
rect 49268 25264 49269 25304
rect 49227 25255 49269 25264
rect 49131 25220 49173 25229
rect 49131 25180 49132 25220
rect 49172 25180 49173 25220
rect 49131 25171 49173 25180
rect 49132 23129 49172 25171
rect 49228 25170 49268 25255
rect 49420 24809 49460 27103
rect 49803 26564 49845 26573
rect 49803 26524 49804 26564
rect 49844 26524 49845 26564
rect 49803 26515 49845 26524
rect 49804 25481 49844 26515
rect 49900 25565 49940 29044
rect 49996 28916 50036 28925
rect 49996 28337 50036 28876
rect 50380 28916 50420 28925
rect 50380 28673 50420 28876
rect 50379 28664 50421 28673
rect 50379 28624 50380 28664
rect 50420 28624 50421 28664
rect 50379 28615 50421 28624
rect 49995 28328 50037 28337
rect 49995 28288 49996 28328
rect 50036 28288 50037 28328
rect 49995 28279 50037 28288
rect 49996 27656 50036 28279
rect 49996 26153 50036 27616
rect 50283 27320 50325 27329
rect 50283 27280 50284 27320
rect 50324 27280 50325 27320
rect 50283 27271 50325 27280
rect 49995 26144 50037 26153
rect 49995 26104 49996 26144
rect 50036 26104 50037 26144
rect 49995 26095 50037 26104
rect 49899 25556 49941 25565
rect 49899 25516 49900 25556
rect 49940 25516 49941 25556
rect 49899 25507 49941 25516
rect 49803 25472 49845 25481
rect 49803 25432 49804 25472
rect 49844 25432 49845 25472
rect 49803 25423 49845 25432
rect 49227 24800 49269 24809
rect 49227 24760 49228 24800
rect 49268 24760 49269 24800
rect 49227 24751 49269 24760
rect 49419 24800 49461 24809
rect 49419 24760 49420 24800
rect 49460 24760 49461 24800
rect 49419 24751 49461 24760
rect 49228 24632 49268 24751
rect 49228 24583 49268 24592
rect 49227 24296 49269 24305
rect 49227 24256 49228 24296
rect 49268 24256 49269 24296
rect 49227 24247 49269 24256
rect 49131 23120 49173 23129
rect 49131 23080 49132 23120
rect 49172 23080 49173 23120
rect 49131 23071 49173 23080
rect 49228 23120 49268 24247
rect 49323 24128 49365 24137
rect 49323 24088 49324 24128
rect 49364 24088 49365 24128
rect 49323 24079 49365 24088
rect 49324 23969 49364 24079
rect 49323 23960 49365 23969
rect 49323 23920 49324 23960
rect 49364 23920 49365 23960
rect 49323 23911 49365 23920
rect 49228 23071 49268 23080
rect 49324 23036 49364 23911
rect 49420 23549 49460 24751
rect 49996 24632 50036 26095
rect 50188 25892 50228 25901
rect 50092 25852 50188 25892
rect 50092 25313 50132 25852
rect 50188 25843 50228 25852
rect 50091 25304 50133 25313
rect 50091 25264 50092 25304
rect 50132 25264 50133 25304
rect 50091 25255 50133 25264
rect 50188 25304 50228 25313
rect 50284 25304 50324 27271
rect 50572 25901 50612 29128
rect 50764 29093 50804 29632
rect 50860 29168 50900 31086
rect 51052 30680 51092 31564
rect 51339 31564 51340 31604
rect 51380 31564 51764 31604
rect 51339 31555 51381 31564
rect 51052 30631 51092 30640
rect 51244 31352 51284 31361
rect 51244 30428 51284 31312
rect 51340 31352 51380 31555
rect 51340 31303 51380 31312
rect 51435 31352 51477 31361
rect 51435 31312 51436 31352
rect 51476 31312 51477 31352
rect 51435 31303 51477 31312
rect 51436 31126 51476 31303
rect 51436 31025 51476 31086
rect 51435 31016 51477 31025
rect 51435 30976 51436 31016
rect 51476 30976 51477 31016
rect 51435 30967 51477 30976
rect 51244 30388 51572 30428
rect 50955 30260 50997 30269
rect 50955 30220 50956 30260
rect 50996 30220 50997 30260
rect 50955 30211 50997 30220
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 50956 29840 50996 30211
rect 51532 30092 51572 30388
rect 51436 30052 51572 30092
rect 51148 29924 51188 29933
rect 50956 29800 51092 29840
rect 50955 29672 50997 29681
rect 50955 29632 50956 29672
rect 50996 29632 50997 29672
rect 50955 29623 50997 29632
rect 50956 29538 50996 29623
rect 51052 29336 51092 29800
rect 51148 29513 51188 29884
rect 51436 29840 51476 30052
rect 51627 29924 51669 29933
rect 51627 29884 51628 29924
rect 51668 29884 51669 29924
rect 51627 29875 51669 29884
rect 51436 29791 51476 29800
rect 51531 29840 51573 29849
rect 51531 29800 51532 29840
rect 51572 29800 51573 29840
rect 51531 29791 51573 29800
rect 51628 29840 51668 29875
rect 51532 29706 51572 29791
rect 51628 29789 51668 29800
rect 51724 29840 51764 31564
rect 51860 31564 51916 31604
rect 51956 31564 51957 31604
rect 51820 31555 51860 31564
rect 51915 31555 51957 31564
rect 51820 31363 51860 31372
rect 51819 31312 51820 31361
rect 51860 31312 51861 31361
rect 51819 31303 51861 31312
rect 52012 31352 52052 32563
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 52780 32201 52820 32656
rect 52779 32192 52821 32201
rect 52779 32152 52780 32192
rect 52820 32152 52821 32192
rect 52779 32143 52821 32152
rect 52972 31940 53012 31949
rect 51820 31228 51860 31303
rect 52012 31193 52052 31312
rect 52108 31900 52972 31940
rect 52108 31352 52148 31900
rect 52972 31891 53012 31900
rect 53068 31781 53108 32824
rect 53164 32864 53204 32875
rect 53164 32789 53204 32824
rect 53355 32864 53397 32873
rect 53355 32824 53356 32864
rect 53396 32824 53397 32864
rect 53355 32815 53397 32824
rect 53452 32864 53492 32873
rect 53163 32780 53205 32789
rect 53163 32740 53164 32780
rect 53204 32740 53205 32780
rect 53163 32731 53205 32740
rect 53067 31772 53109 31781
rect 53067 31732 53068 31772
rect 53108 31732 53109 31772
rect 53067 31723 53109 31732
rect 52395 31604 52437 31613
rect 52395 31564 52396 31604
rect 52436 31564 52437 31604
rect 52395 31555 52437 31564
rect 52396 31436 52436 31555
rect 52491 31520 52533 31529
rect 52491 31480 52492 31520
rect 52532 31480 52533 31520
rect 52491 31471 52533 31480
rect 52396 31387 52436 31396
rect 52492 31386 52532 31471
rect 52587 31436 52629 31445
rect 52587 31396 52588 31436
rect 52628 31396 52629 31436
rect 52587 31387 52629 31396
rect 52011 31184 52053 31193
rect 52011 31144 52012 31184
rect 52052 31144 52053 31184
rect 52011 31135 52053 31144
rect 51819 31100 51861 31109
rect 51819 31060 51820 31100
rect 51860 31060 51861 31100
rect 51819 31051 51861 31060
rect 51724 29791 51764 29800
rect 51147 29504 51189 29513
rect 51147 29464 51148 29504
rect 51188 29464 51189 29504
rect 51147 29455 51189 29464
rect 51820 29336 51860 31051
rect 52011 31016 52053 31025
rect 52011 30976 52012 31016
rect 52052 30976 52053 31016
rect 52011 30967 52053 30976
rect 51052 29287 51092 29296
rect 51148 29296 51820 29336
rect 50955 29168 50997 29177
rect 50860 29128 50956 29168
rect 50996 29128 50997 29168
rect 50955 29119 50997 29128
rect 51148 29168 51188 29296
rect 51820 29287 51860 29296
rect 51916 30680 51956 30689
rect 51148 29119 51188 29128
rect 51244 29168 51284 29177
rect 50763 29084 50805 29093
rect 50763 29044 50764 29084
rect 50804 29044 50805 29084
rect 50763 29035 50805 29044
rect 50956 29034 50996 29119
rect 51244 29009 51284 29128
rect 51435 29168 51477 29177
rect 51435 29128 51436 29168
rect 51476 29128 51477 29168
rect 51435 29119 51477 29128
rect 51243 29000 51285 29009
rect 51243 28960 51244 29000
rect 51284 28960 51285 29000
rect 51243 28951 51285 28960
rect 51436 29000 51476 29119
rect 51531 29084 51573 29093
rect 51531 29044 51532 29084
rect 51572 29044 51573 29084
rect 51531 29035 51573 29044
rect 51628 29084 51668 29093
rect 51436 28951 51476 28960
rect 50763 28832 50805 28841
rect 50763 28792 50764 28832
rect 50804 28792 50805 28832
rect 50763 28783 50805 28792
rect 50764 26237 50804 28783
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 50859 28664 50901 28673
rect 50859 28624 50860 28664
rect 50900 28624 50901 28664
rect 50859 28615 50901 28624
rect 50860 28328 50900 28615
rect 50860 28279 50900 28288
rect 51148 27404 51188 27413
rect 50956 27364 51148 27404
rect 50859 27068 50901 27077
rect 50859 27028 50860 27068
rect 50900 27028 50901 27068
rect 50859 27019 50901 27028
rect 50860 26934 50900 27019
rect 50956 26741 50996 27364
rect 51148 27355 51188 27364
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 50955 26732 50997 26741
rect 50955 26692 50956 26732
rect 50996 26692 50997 26732
rect 50955 26683 50997 26692
rect 50763 26228 50805 26237
rect 50763 26188 50764 26228
rect 50804 26188 50805 26228
rect 50763 26179 50805 26188
rect 50571 25892 50613 25901
rect 50571 25852 50572 25892
rect 50612 25852 50613 25892
rect 50571 25843 50613 25852
rect 50379 25808 50421 25817
rect 50379 25768 50380 25808
rect 50420 25768 50421 25808
rect 50379 25759 50421 25768
rect 50228 25264 50324 25304
rect 50380 25304 50420 25759
rect 50764 25556 50804 26179
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 50764 25507 50804 25516
rect 50571 25388 50613 25397
rect 50571 25348 50572 25388
rect 50612 25348 50613 25388
rect 50571 25339 50613 25348
rect 51244 25388 51284 25397
rect 51532 25388 51572 29035
rect 51628 28841 51668 29044
rect 51627 28832 51669 28841
rect 51627 28792 51628 28832
rect 51668 28792 51669 28832
rect 51627 28783 51669 28792
rect 51916 28673 51956 30640
rect 52012 29672 52052 30967
rect 52108 29840 52148 31312
rect 52300 31352 52340 31363
rect 52300 31277 52340 31312
rect 52588 31302 52628 31387
rect 52683 31352 52725 31361
rect 52683 31312 52684 31352
rect 52724 31312 52725 31352
rect 52683 31303 52725 31312
rect 52972 31352 53012 31361
rect 52299 31268 52341 31277
rect 52299 31228 52300 31268
rect 52340 31228 52341 31268
rect 52299 31219 52341 31228
rect 52684 31218 52724 31303
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 52972 30596 53012 31312
rect 52876 30556 53012 30596
rect 52204 29840 52244 29849
rect 52108 29800 52204 29840
rect 52204 29791 52244 29800
rect 52108 29672 52148 29681
rect 52012 29632 52108 29672
rect 52108 29623 52148 29632
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 52204 29168 52244 29177
rect 52012 29084 52052 29093
rect 51915 28664 51957 28673
rect 51915 28624 51916 28664
rect 51956 28624 51957 28664
rect 51915 28615 51957 28624
rect 51724 28328 51764 28337
rect 51724 27161 51764 28288
rect 51819 28328 51861 28337
rect 51819 28288 51820 28328
rect 51860 28288 51861 28328
rect 51819 28279 51861 28288
rect 51723 27152 51765 27161
rect 51723 27112 51724 27152
rect 51764 27112 51765 27152
rect 51723 27103 51765 27112
rect 51723 26648 51765 26657
rect 51723 26608 51724 26648
rect 51764 26608 51765 26648
rect 51723 26599 51765 26608
rect 51284 25348 51572 25388
rect 50420 25264 50516 25304
rect 50092 25170 50132 25255
rect 50092 24632 50132 24641
rect 49996 24592 50092 24632
rect 50092 24583 50132 24592
rect 49803 24548 49845 24557
rect 49803 24508 49804 24548
rect 49844 24508 49845 24548
rect 49803 24499 49845 24508
rect 49804 23792 49844 24499
rect 50188 24464 50228 25264
rect 50380 25255 50420 25264
rect 50284 25136 50324 25145
rect 50324 25096 50420 25136
rect 50284 25087 50324 25096
rect 50283 24800 50325 24809
rect 50283 24760 50284 24800
rect 50324 24760 50325 24800
rect 50283 24751 50325 24760
rect 49996 24424 50228 24464
rect 49804 23743 49844 23752
rect 49900 23792 49940 23801
rect 49996 23792 50036 24424
rect 49940 23752 50036 23792
rect 50092 23792 50132 23801
rect 50284 23792 50324 24751
rect 50380 23876 50420 25096
rect 50476 24809 50516 25264
rect 50572 25254 50612 25339
rect 50667 25304 50709 25313
rect 50667 25264 50668 25304
rect 50708 25264 50709 25304
rect 50667 25255 50709 25264
rect 51052 25304 51092 25313
rect 50475 24800 50517 24809
rect 50475 24760 50476 24800
rect 50516 24760 50517 24800
rect 50475 24751 50517 24760
rect 50475 24464 50517 24473
rect 50475 24424 50476 24464
rect 50516 24424 50517 24464
rect 50475 24415 50517 24424
rect 50476 24002 50516 24415
rect 50668 24137 50708 25255
rect 50763 25136 50805 25145
rect 50956 25136 50996 25145
rect 50763 25096 50764 25136
rect 50804 25096 50805 25136
rect 50763 25087 50805 25096
rect 50860 25096 50956 25136
rect 50764 25002 50804 25087
rect 50667 24128 50709 24137
rect 50667 24088 50668 24128
rect 50708 24088 50709 24128
rect 50667 24079 50709 24088
rect 50571 24044 50613 24053
rect 50571 24004 50572 24044
rect 50612 24004 50613 24044
rect 50571 23995 50613 24004
rect 50476 23953 50516 23962
rect 50380 23827 50420 23836
rect 50572 23876 50612 23995
rect 50572 23827 50612 23836
rect 50132 23752 50284 23792
rect 49419 23540 49461 23549
rect 49419 23500 49420 23540
rect 49460 23500 49461 23540
rect 49419 23491 49461 23500
rect 49900 23381 49940 23752
rect 49996 23624 50036 23633
rect 49899 23372 49941 23381
rect 49899 23332 49900 23372
rect 49940 23332 49941 23372
rect 49899 23323 49941 23332
rect 49324 22987 49364 22996
rect 49708 23120 49748 23129
rect 49323 22448 49365 22457
rect 49323 22408 49324 22448
rect 49364 22408 49365 22448
rect 49708 22448 49748 23080
rect 49804 23036 49844 23045
rect 49804 22625 49844 22996
rect 49996 23036 50036 23584
rect 50092 23120 50132 23752
rect 50284 23288 50324 23752
rect 50475 23792 50517 23801
rect 50475 23752 50476 23792
rect 50516 23752 50517 23792
rect 50475 23743 50517 23752
rect 50668 23750 50708 23759
rect 50379 23540 50421 23549
rect 50379 23500 50380 23540
rect 50420 23500 50421 23540
rect 50379 23491 50421 23500
rect 50284 23239 50324 23248
rect 50092 23071 50132 23080
rect 49996 22987 50036 22996
rect 49900 22952 49940 22961
rect 49803 22616 49845 22625
rect 49803 22576 49804 22616
rect 49844 22576 49845 22616
rect 49803 22567 49845 22576
rect 49708 22408 49844 22448
rect 49323 22399 49365 22408
rect 49324 22314 49364 22399
rect 49611 22280 49653 22289
rect 49611 22240 49612 22280
rect 49652 22240 49653 22280
rect 49611 22231 49653 22240
rect 49708 22280 49748 22289
rect 49612 22146 49652 22231
rect 49708 22121 49748 22240
rect 49707 22112 49749 22121
rect 49707 22072 49708 22112
rect 49748 22072 49749 22112
rect 49707 22063 49749 22072
rect 49804 22054 49844 22408
rect 49804 21944 49844 22014
rect 49708 21904 49844 21944
rect 49420 21608 49460 21617
rect 49132 20768 49172 20777
rect 49132 20189 49172 20728
rect 49131 20180 49173 20189
rect 49131 20140 49132 20180
rect 49172 20140 49173 20180
rect 49131 20131 49173 20140
rect 49420 20105 49460 21568
rect 49515 21356 49557 21365
rect 49515 21316 49516 21356
rect 49556 21316 49557 21356
rect 49515 21307 49557 21316
rect 49516 20768 49556 21307
rect 49612 21020 49652 21029
rect 49708 21020 49748 21904
rect 49804 21692 49844 21701
rect 49900 21692 49940 22912
rect 50091 22448 50133 22457
rect 50091 22408 50092 22448
rect 50132 22408 50133 22448
rect 50091 22399 50133 22408
rect 49996 22196 50036 22205
rect 49996 21776 50036 22156
rect 49996 21727 50036 21736
rect 49844 21652 49940 21692
rect 49804 21643 49844 21652
rect 50092 21608 50132 22399
rect 50380 22280 50420 23491
rect 50476 23036 50516 23743
rect 50668 23708 50708 23710
rect 50860 23708 50900 25096
rect 50956 25087 50996 25096
rect 51052 24884 51092 25264
rect 51147 25136 51189 25145
rect 51147 25096 51148 25136
rect 51188 25096 51189 25136
rect 51147 25087 51189 25096
rect 50956 24844 51092 24884
rect 50956 24557 50996 24844
rect 51148 24800 51188 25087
rect 51052 24760 51188 24800
rect 50955 24548 50997 24557
rect 50955 24508 50956 24548
rect 50996 24508 50997 24548
rect 50955 24499 50997 24508
rect 50955 24128 50997 24137
rect 50955 24088 50956 24128
rect 50996 24088 50997 24128
rect 50955 24079 50997 24088
rect 50668 23668 50900 23708
rect 50860 23620 50900 23668
rect 50860 23571 50900 23580
rect 50956 23792 50996 24079
rect 50859 23372 50901 23381
rect 50859 23332 50860 23372
rect 50900 23332 50901 23372
rect 50859 23323 50901 23332
rect 50860 23288 50900 23323
rect 50860 23237 50900 23248
rect 50476 22987 50516 22996
rect 50667 23036 50709 23045
rect 50667 22996 50668 23036
rect 50708 22996 50709 23036
rect 50667 22987 50709 22996
rect 50668 22902 50708 22987
rect 50956 22877 50996 23752
rect 51052 23792 51092 24760
rect 51244 24716 51284 25348
rect 51724 25304 51764 26599
rect 51820 25472 51860 28279
rect 51916 27413 51956 28615
rect 52012 27833 52052 29044
rect 52204 29009 52244 29128
rect 52203 29000 52245 29009
rect 52203 28960 52204 29000
rect 52244 28960 52245 29000
rect 52203 28951 52245 28960
rect 52300 28916 52340 28925
rect 52108 28244 52148 28253
rect 52011 27824 52053 27833
rect 52011 27784 52012 27824
rect 52052 27784 52053 27824
rect 52011 27775 52053 27784
rect 52108 27740 52148 28204
rect 52300 28160 52340 28876
rect 52876 28748 52916 30556
rect 53068 30428 53108 30437
rect 53068 29933 53108 30388
rect 53067 29924 53109 29933
rect 53067 29884 53068 29924
rect 53108 29884 53109 29924
rect 53067 29875 53109 29884
rect 53164 29849 53204 32731
rect 53356 32730 53396 32815
rect 53452 32789 53492 32824
rect 53547 32864 53589 32873
rect 53547 32824 53548 32864
rect 53588 32824 53589 32864
rect 53547 32815 53589 32824
rect 53644 32864 53684 32899
rect 53451 32780 53493 32789
rect 53451 32740 53452 32780
rect 53492 32740 53493 32780
rect 53451 32731 53493 32740
rect 53452 32537 53492 32731
rect 53548 32730 53588 32815
rect 53644 32705 53684 32824
rect 53836 32864 53876 32873
rect 53643 32696 53685 32705
rect 53643 32656 53644 32696
rect 53684 32656 53685 32696
rect 53643 32647 53685 32656
rect 53451 32528 53493 32537
rect 53451 32488 53452 32528
rect 53492 32488 53493 32528
rect 53451 32479 53493 32488
rect 53355 32444 53397 32453
rect 53355 32404 53356 32444
rect 53396 32404 53397 32444
rect 53355 32395 53397 32404
rect 53356 32201 53396 32395
rect 53355 32192 53397 32201
rect 53355 32152 53356 32192
rect 53396 32152 53397 32192
rect 53355 32143 53397 32152
rect 53356 32058 53396 32143
rect 53643 31520 53685 31529
rect 53643 31480 53644 31520
rect 53684 31480 53685 31520
rect 53643 31471 53685 31480
rect 53644 30764 53684 31471
rect 53836 31277 53876 32824
rect 54028 32864 54068 32899
rect 54028 32621 54068 32824
rect 54124 32864 54164 33403
rect 54603 33368 54645 33377
rect 54603 33328 54604 33368
rect 54644 33328 54645 33368
rect 54603 33319 54645 33328
rect 54411 33116 54453 33125
rect 54411 33076 54412 33116
rect 54452 33076 54453 33116
rect 54411 33067 54453 33076
rect 54412 32873 54452 33067
rect 54124 32815 54164 32824
rect 54411 32864 54453 32873
rect 54411 32824 54412 32864
rect 54452 32824 54453 32864
rect 54411 32815 54453 32824
rect 54604 32864 54644 33319
rect 54700 33209 54740 33496
rect 54796 33461 54836 33664
rect 54795 33452 54837 33461
rect 54795 33412 54796 33452
rect 54836 33412 54837 33452
rect 54795 33403 54837 33412
rect 54988 33452 55028 33461
rect 54699 33200 54741 33209
rect 54699 33160 54700 33200
rect 54740 33160 54741 33200
rect 54699 33151 54741 33160
rect 54988 32873 55028 33412
rect 54604 32815 54644 32824
rect 54699 32864 54741 32873
rect 54699 32824 54700 32864
rect 54740 32824 54741 32864
rect 54699 32815 54741 32824
rect 54796 32864 54836 32873
rect 54027 32612 54069 32621
rect 54027 32572 54028 32612
rect 54068 32572 54069 32612
rect 54027 32563 54069 32572
rect 54412 31604 54452 32815
rect 54700 32730 54740 32815
rect 54603 32444 54645 32453
rect 54603 32404 54604 32444
rect 54644 32404 54645 32444
rect 54603 32395 54645 32404
rect 54508 31940 54548 31949
rect 54508 31781 54548 31900
rect 54507 31772 54549 31781
rect 54507 31732 54508 31772
rect 54548 31732 54549 31772
rect 54507 31723 54549 31732
rect 54604 31604 54644 32395
rect 54796 31865 54836 32824
rect 54892 32864 54932 32873
rect 54795 31856 54837 31865
rect 54795 31816 54796 31856
rect 54836 31816 54837 31856
rect 54795 31807 54837 31816
rect 54412 31564 54548 31604
rect 53931 31436 53973 31445
rect 53931 31396 53932 31436
rect 53972 31396 53973 31436
rect 53931 31387 53973 31396
rect 53835 31268 53877 31277
rect 53835 31228 53836 31268
rect 53876 31228 53877 31268
rect 53835 31219 53877 31228
rect 53644 30715 53684 30724
rect 53836 30605 53876 31219
rect 53835 30596 53877 30605
rect 53835 30556 53836 30596
rect 53876 30556 53877 30596
rect 53835 30547 53877 30556
rect 53932 30269 53972 31387
rect 54123 31352 54165 31361
rect 54123 31312 54124 31352
rect 54164 31312 54165 31352
rect 54123 31303 54165 31312
rect 54028 30680 54068 30689
rect 54028 30353 54068 30640
rect 54027 30344 54069 30353
rect 54027 30304 54028 30344
rect 54068 30304 54069 30344
rect 54027 30295 54069 30304
rect 53355 30260 53397 30269
rect 53355 30220 53356 30260
rect 53396 30220 53397 30260
rect 53355 30211 53397 30220
rect 53931 30260 53973 30269
rect 53931 30220 53932 30260
rect 53972 30220 53973 30260
rect 53931 30211 53973 30220
rect 53163 29840 53205 29849
rect 53163 29800 53164 29840
rect 53204 29800 53205 29840
rect 53163 29791 53205 29800
rect 53164 29168 53204 29791
rect 53356 29168 53396 30211
rect 53932 30092 53972 30211
rect 53932 30043 53972 30052
rect 53164 29119 53204 29128
rect 53260 29126 53300 29135
rect 53259 29086 53260 29093
rect 53356 29119 53396 29128
rect 53452 29168 53492 29177
rect 53644 29168 53684 29177
rect 53492 29128 53644 29168
rect 53452 29119 53492 29128
rect 53644 29119 53684 29128
rect 54028 29168 54068 30295
rect 54124 29672 54164 31303
rect 54219 30176 54261 30185
rect 54219 30136 54220 30176
rect 54260 30136 54261 30176
rect 54219 30127 54261 30136
rect 54220 29840 54260 30127
rect 54316 29849 54356 29934
rect 54220 29791 54260 29800
rect 54315 29840 54357 29849
rect 54315 29800 54316 29840
rect 54356 29800 54357 29840
rect 54315 29791 54357 29800
rect 54412 29672 54452 29677
rect 54124 29668 54452 29672
rect 54124 29632 54412 29668
rect 54412 29619 54452 29628
rect 54028 29119 54068 29128
rect 53300 29086 53301 29093
rect 53259 29084 53301 29086
rect 53259 29044 53260 29084
rect 53300 29044 53301 29084
rect 53259 29035 53301 29044
rect 53260 28991 53300 29035
rect 54315 28916 54357 28925
rect 54315 28876 54316 28916
rect 54356 28876 54357 28916
rect 54315 28867 54357 28876
rect 52876 28708 52964 28748
rect 52780 28505 52820 28590
rect 52779 28496 52821 28505
rect 52492 28421 52532 28465
rect 52779 28456 52780 28496
rect 52820 28456 52821 28496
rect 52779 28447 52821 28456
rect 52491 28412 52533 28421
rect 52491 28372 52492 28412
rect 52532 28372 52533 28412
rect 52491 28370 52533 28372
rect 52491 28363 52492 28370
rect 52395 28328 52437 28337
rect 52395 28288 52396 28328
rect 52436 28288 52437 28328
rect 52532 28363 52533 28370
rect 52492 28321 52532 28330
rect 52924 28328 52964 28708
rect 53067 28496 53109 28505
rect 53067 28456 53068 28496
rect 53108 28456 53109 28496
rect 53067 28447 53109 28456
rect 52395 28279 52437 28288
rect 52780 28288 52964 28328
rect 53068 28328 53108 28447
rect 52396 28194 52436 28279
rect 52204 28156 52340 28160
rect 52204 28120 52300 28156
rect 52204 27828 52244 28120
rect 52780 28160 52820 28288
rect 53068 28279 53108 28288
rect 53164 28328 53204 28337
rect 52972 28160 53012 28169
rect 53164 28160 53204 28288
rect 53260 28328 53300 28337
rect 53451 28328 53493 28337
rect 53300 28288 53396 28328
rect 53260 28279 53300 28288
rect 52780 28120 52868 28160
rect 52300 28107 52340 28116
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52828 27992 52868 28120
rect 53012 28120 53108 28160
rect 53164 28120 53300 28160
rect 52972 28111 53012 28120
rect 53068 28076 53108 28120
rect 53068 28036 53204 28076
rect 52828 27952 52964 27992
rect 52352 27943 52720 27952
rect 52204 27788 52436 27828
rect 52108 27700 52244 27740
rect 52011 27656 52053 27665
rect 52011 27616 52012 27656
rect 52052 27616 52053 27656
rect 52011 27607 52053 27616
rect 52012 27522 52052 27607
rect 52108 27572 52148 27583
rect 52108 27497 52148 27532
rect 52107 27488 52149 27497
rect 52107 27448 52108 27488
rect 52148 27448 52149 27488
rect 52107 27439 52149 27448
rect 52204 27488 52244 27700
rect 52396 27656 52436 27788
rect 52779 27824 52821 27833
rect 52779 27784 52780 27824
rect 52820 27784 52821 27824
rect 52924 27828 52964 27952
rect 52924 27824 53012 27828
rect 52924 27788 53060 27824
rect 52972 27784 53060 27788
rect 52779 27775 52821 27784
rect 52683 27656 52725 27665
rect 52396 27607 52436 27616
rect 52588 27645 52684 27656
rect 52628 27616 52684 27645
rect 52724 27616 52725 27656
rect 52683 27607 52725 27616
rect 52780 27656 52820 27775
rect 52588 27596 52628 27605
rect 52204 27439 52244 27448
rect 52300 27572 52340 27581
rect 51915 27404 51957 27413
rect 51915 27364 51916 27404
rect 51956 27364 51957 27404
rect 51915 27355 51957 27364
rect 51916 26816 51956 27355
rect 52300 27245 52340 27532
rect 52587 27488 52629 27497
rect 52587 27448 52588 27488
rect 52628 27448 52629 27488
rect 52587 27439 52629 27448
rect 52588 27354 52628 27439
rect 52299 27236 52341 27245
rect 52299 27196 52300 27236
rect 52340 27196 52341 27236
rect 52299 27187 52341 27196
rect 52107 27152 52149 27161
rect 52107 27112 52108 27152
rect 52148 27112 52149 27152
rect 52107 27103 52149 27112
rect 52012 26816 52052 26825
rect 51916 26776 52012 26816
rect 52012 26767 52052 26776
rect 52108 25556 52148 27103
rect 52684 26825 52724 27607
rect 52780 27329 52820 27616
rect 52876 27656 52916 27665
rect 52779 27320 52821 27329
rect 52779 27280 52780 27320
rect 52820 27280 52821 27320
rect 52779 27271 52821 27280
rect 52779 27152 52821 27161
rect 52779 27112 52780 27152
rect 52820 27112 52821 27152
rect 52779 27103 52821 27112
rect 52780 26993 52820 27103
rect 52876 27077 52916 27616
rect 53020 27572 53060 27784
rect 53164 27740 53204 28036
rect 53260 27917 53300 28120
rect 53259 27908 53301 27917
rect 53259 27868 53260 27908
rect 53300 27868 53301 27908
rect 53259 27859 53301 27868
rect 53164 27691 53204 27700
rect 53020 27532 53108 27572
rect 52875 27068 52917 27077
rect 52875 27028 52876 27068
rect 52916 27028 52917 27068
rect 52875 27019 52917 27028
rect 52779 26984 52821 26993
rect 52779 26944 52780 26984
rect 52820 26944 52821 26984
rect 52779 26935 52821 26944
rect 52683 26816 52725 26825
rect 52683 26776 52684 26816
rect 52724 26776 52725 26816
rect 52780 26816 52820 26935
rect 52876 26816 52916 26825
rect 52780 26776 52876 26816
rect 52683 26767 52725 26776
rect 52876 26767 52916 26776
rect 53068 26648 53108 27532
rect 52876 26608 53108 26648
rect 53260 26732 53300 26741
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 52299 25724 52341 25733
rect 52299 25684 52300 25724
rect 52340 25684 52341 25724
rect 52299 25675 52341 25684
rect 52300 25565 52340 25675
rect 52012 25516 52148 25556
rect 52299 25556 52341 25565
rect 52299 25516 52300 25556
rect 52340 25516 52341 25556
rect 51820 25432 51956 25472
rect 51916 25313 51956 25432
rect 51436 25264 51724 25304
rect 51436 25136 51476 25264
rect 51436 25087 51476 25096
rect 51531 25136 51573 25145
rect 51628 25136 51668 25145
rect 51531 25096 51532 25136
rect 51572 25096 51628 25136
rect 51531 25087 51573 25096
rect 51628 25087 51668 25096
rect 51148 24676 51284 24716
rect 51148 24473 51188 24676
rect 51436 24632 51476 24641
rect 51243 24548 51285 24557
rect 51243 24508 51244 24548
rect 51284 24508 51285 24548
rect 51243 24499 51285 24508
rect 51147 24464 51189 24473
rect 51147 24424 51148 24464
rect 51188 24424 51189 24464
rect 51147 24415 51189 24424
rect 51244 24414 51284 24499
rect 51147 24212 51189 24221
rect 51147 24172 51148 24212
rect 51188 24172 51189 24212
rect 51147 24163 51189 24172
rect 51052 23743 51092 23752
rect 50955 22868 50997 22877
rect 50955 22828 50956 22868
rect 50996 22828 50997 22868
rect 50955 22819 50997 22828
rect 50380 22231 50420 22240
rect 50475 22280 50517 22289
rect 50475 22240 50476 22280
rect 50516 22240 50517 22280
rect 50475 22231 50517 22240
rect 50092 21559 50132 21568
rect 50188 21608 50228 21619
rect 50188 21533 50228 21568
rect 50283 21608 50325 21617
rect 50283 21568 50284 21608
rect 50324 21568 50325 21608
rect 50283 21559 50325 21568
rect 50476 21608 50516 22231
rect 50956 22121 50996 22819
rect 50955 22112 50997 22121
rect 50955 22072 50956 22112
rect 50996 22072 50997 22112
rect 50955 22063 50997 22072
rect 50763 21944 50805 21953
rect 50763 21904 50764 21944
rect 50804 21904 50805 21944
rect 50763 21895 50805 21904
rect 50667 21692 50709 21701
rect 50667 21652 50668 21692
rect 50708 21652 50709 21692
rect 50667 21643 50709 21652
rect 50476 21559 50516 21568
rect 50571 21608 50613 21617
rect 50571 21568 50572 21608
rect 50612 21568 50613 21608
rect 50571 21559 50613 21568
rect 50668 21608 50708 21643
rect 50187 21524 50229 21533
rect 50187 21484 50188 21524
rect 50228 21484 50229 21524
rect 50187 21475 50229 21484
rect 50284 21474 50324 21559
rect 50572 21474 50612 21559
rect 50668 21557 50708 21568
rect 50764 21608 50804 21895
rect 51148 21776 51188 24163
rect 51243 24128 51285 24137
rect 51243 24088 51244 24128
rect 51284 24088 51285 24128
rect 51243 24079 51285 24088
rect 51244 23969 51284 24079
rect 51339 24044 51381 24053
rect 51339 24004 51340 24044
rect 51380 24004 51381 24044
rect 51339 23995 51381 24004
rect 51243 23960 51285 23969
rect 51243 23920 51244 23960
rect 51284 23920 51285 23960
rect 51243 23911 51285 23920
rect 51340 23910 51380 23995
rect 51436 23792 51476 24592
rect 51627 24044 51669 24053
rect 51627 24004 51628 24044
rect 51668 24004 51669 24044
rect 51627 23995 51669 24004
rect 51627 23962 51668 23995
rect 51627 23876 51667 23962
rect 51724 23886 51764 25264
rect 51820 25304 51860 25313
rect 51820 24809 51860 25264
rect 51915 25304 51957 25313
rect 51915 25264 51916 25304
rect 51956 25264 51957 25304
rect 51915 25255 51957 25264
rect 51916 25170 51956 25255
rect 51819 24800 51861 24809
rect 51819 24760 51820 24800
rect 51860 24760 51861 24800
rect 51819 24751 51861 24760
rect 51820 24632 51860 24641
rect 52012 24632 52052 25516
rect 52299 25507 52341 25516
rect 52300 25422 52340 25507
rect 52108 25388 52148 25397
rect 52108 25229 52148 25348
rect 52107 25220 52149 25229
rect 52107 25180 52108 25220
rect 52148 25180 52149 25220
rect 52107 25171 52149 25180
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 52299 24800 52341 24809
rect 52299 24760 52300 24800
rect 52340 24760 52341 24800
rect 52299 24751 52341 24760
rect 51860 24592 52052 24632
rect 51820 24583 51860 24592
rect 52300 24557 52340 24751
rect 52684 24632 52724 24641
rect 52588 24592 52684 24632
rect 52107 24548 52149 24557
rect 52107 24508 52108 24548
rect 52148 24508 52149 24548
rect 52107 24499 52149 24508
rect 52299 24548 52341 24557
rect 52299 24508 52300 24548
rect 52340 24508 52341 24548
rect 52299 24499 52341 24508
rect 52011 24212 52053 24221
rect 52011 24172 52012 24212
rect 52052 24172 52053 24212
rect 52011 24163 52053 24172
rect 51724 23876 51847 23886
rect 52012 23876 52052 24163
rect 51627 23836 51668 23876
rect 51724 23846 51860 23876
rect 51807 23836 51860 23846
rect 51628 23834 51668 23836
rect 51532 23792 51572 23801
rect 51436 23752 51532 23792
rect 51628 23785 51668 23794
rect 51724 23792 51764 23801
rect 51532 23743 51572 23752
rect 51724 23213 51764 23752
rect 51820 23800 51860 23836
rect 52108 23876 52148 24499
rect 52203 24464 52245 24473
rect 52203 24424 52204 24464
rect 52244 24424 52245 24464
rect 52203 24415 52245 24424
rect 52204 24044 52244 24415
rect 52204 23995 52244 24004
rect 52108 23836 52244 23876
rect 52012 23827 52052 23836
rect 51860 23792 51868 23800
rect 51860 23760 51956 23792
rect 51820 23752 51956 23760
rect 51820 23751 51860 23752
rect 51916 23549 51956 23752
rect 51915 23540 51957 23549
rect 51915 23500 51916 23540
rect 51956 23500 51957 23540
rect 51915 23491 51957 23500
rect 51723 23204 51765 23213
rect 51723 23164 51724 23204
rect 51764 23164 51765 23204
rect 51723 23155 51765 23164
rect 51532 23129 51572 23131
rect 51531 23120 51573 23129
rect 51531 23080 51532 23120
rect 51572 23080 51573 23120
rect 51531 23071 51573 23080
rect 51243 23036 51285 23045
rect 51243 22996 51244 23036
rect 51284 22996 51285 23036
rect 51243 22987 51285 22996
rect 51532 23036 51572 23071
rect 51532 22987 51572 22996
rect 51244 22280 51284 22987
rect 51339 22868 51381 22877
rect 51339 22828 51340 22868
rect 51380 22828 51381 22868
rect 51339 22819 51381 22828
rect 51531 22868 51573 22877
rect 51531 22828 51532 22868
rect 51572 22828 51573 22868
rect 51531 22819 51573 22828
rect 51340 22734 51380 22819
rect 51284 22240 51476 22280
rect 51244 22231 51284 22240
rect 51148 21736 51380 21776
rect 50764 21559 50804 21568
rect 51243 21608 51285 21617
rect 51243 21568 51244 21608
rect 51284 21568 51285 21608
rect 51243 21559 51285 21568
rect 51147 21524 51189 21533
rect 51147 21484 51148 21524
rect 51188 21484 51189 21524
rect 51147 21475 51189 21484
rect 51148 21390 51188 21475
rect 51244 21474 51284 21559
rect 49652 20980 49748 21020
rect 49612 20971 49652 20980
rect 49516 20719 49556 20728
rect 49996 20852 50036 20861
rect 49804 20600 49844 20609
rect 49611 20180 49653 20189
rect 49611 20140 49612 20180
rect 49652 20140 49653 20180
rect 49611 20131 49653 20140
rect 49419 20096 49461 20105
rect 49419 20056 49420 20096
rect 49460 20056 49461 20096
rect 49419 20047 49461 20056
rect 49612 20096 49652 20131
rect 49612 20045 49652 20056
rect 49611 19340 49653 19349
rect 49611 19300 49612 19340
rect 49652 19300 49653 19340
rect 49611 19291 49653 19300
rect 48939 17828 48981 17837
rect 48939 17788 48940 17828
rect 48980 17788 48981 17828
rect 48939 17779 48981 17788
rect 48939 17576 48981 17585
rect 48939 17536 48940 17576
rect 48980 17536 48981 17576
rect 48939 17527 48981 17536
rect 48844 17023 48884 17032
rect 48940 16316 48980 17527
rect 48844 16276 48980 16316
rect 48747 14720 48789 14729
rect 48747 14680 48748 14720
rect 48788 14680 48789 14720
rect 48747 14671 48789 14680
rect 48748 14586 48788 14671
rect 48651 14300 48693 14309
rect 48651 14260 48652 14300
rect 48692 14260 48693 14300
rect 48651 14251 48693 14260
rect 48363 14132 48405 14141
rect 48363 14092 48364 14132
rect 48404 14092 48405 14132
rect 48363 14083 48405 14092
rect 47787 13292 47829 13301
rect 47787 13252 47788 13292
rect 47828 13252 47829 13292
rect 47787 13243 47829 13252
rect 47691 13208 47733 13217
rect 47691 13168 47692 13208
rect 47732 13168 47733 13208
rect 47691 13159 47733 13168
rect 47692 13074 47732 13159
rect 47788 13158 47828 13243
rect 47980 12704 48020 13999
rect 48076 12881 48116 14008
rect 48172 13964 48212 13973
rect 48172 12980 48212 13924
rect 48364 13964 48404 14083
rect 48459 14048 48501 14057
rect 48459 14008 48460 14048
rect 48500 14008 48501 14048
rect 48459 13999 48501 14008
rect 48652 14048 48692 14057
rect 48364 13915 48404 13924
rect 48460 13914 48500 13999
rect 48268 13880 48308 13889
rect 48268 13796 48308 13840
rect 48652 13796 48692 14008
rect 48268 13756 48692 13796
rect 48172 12940 48308 12980
rect 48075 12872 48117 12881
rect 48075 12832 48076 12872
rect 48116 12832 48212 12872
rect 48075 12823 48117 12832
rect 48075 12704 48117 12713
rect 47980 12664 48076 12704
rect 48116 12664 48117 12704
rect 48075 12655 48117 12664
rect 47211 12536 47253 12545
rect 47211 12496 47212 12536
rect 47252 12496 47253 12536
rect 47211 12487 47253 12496
rect 48076 12536 48116 12655
rect 48172 12629 48212 12832
rect 48268 12797 48308 12940
rect 48267 12788 48309 12797
rect 48267 12748 48268 12788
rect 48308 12748 48309 12788
rect 48267 12739 48309 12748
rect 48171 12620 48213 12629
rect 48171 12580 48172 12620
rect 48212 12580 48213 12620
rect 48171 12571 48213 12580
rect 48076 12487 48116 12496
rect 48651 12536 48693 12545
rect 48651 12496 48652 12536
rect 48692 12496 48693 12536
rect 48651 12487 48693 12496
rect 47212 12402 47252 12487
rect 46923 11824 46924 11864
rect 46964 11824 47060 11864
rect 46923 11815 46965 11824
rect 46924 11730 46964 11815
rect 46636 11647 46676 11656
rect 48652 11696 48692 12487
rect 48652 11647 48692 11656
rect 46251 11612 46293 11621
rect 46251 11572 46252 11612
rect 46292 11572 46293 11612
rect 46251 11563 46293 11572
rect 48268 11612 48308 11621
rect 46252 11478 46292 11563
rect 46444 11470 46484 11479
rect 46348 11192 46388 11201
rect 46444 11192 46484 11430
rect 47115 11276 47157 11285
rect 47115 11236 47116 11276
rect 47156 11236 47157 11276
rect 47115 11227 47157 11236
rect 46388 11152 46484 11192
rect 46251 11108 46293 11117
rect 46251 11068 46252 11108
rect 46292 11068 46293 11108
rect 46251 11059 46293 11068
rect 46060 10975 46100 10984
rect 46252 11024 46292 11059
rect 46348 11033 46388 11152
rect 46252 10973 46292 10984
rect 46347 11024 46389 11033
rect 46347 10984 46348 11024
rect 46388 10984 46389 11024
rect 46347 10975 46389 10984
rect 45964 10891 46004 10900
rect 45868 10807 45908 10816
rect 45771 10352 45813 10361
rect 45771 10312 45772 10352
rect 45812 10312 45813 10352
rect 45771 10303 45813 10312
rect 45387 10268 45429 10277
rect 45387 10228 45388 10268
rect 45428 10228 45429 10268
rect 45387 10219 45429 10228
rect 44620 9136 44756 9176
rect 44812 9764 44852 10135
rect 44908 9941 44948 10144
rect 45003 10184 45045 10193
rect 45003 10144 45004 10184
rect 45044 10144 45045 10184
rect 45003 10135 45045 10144
rect 45100 10184 45140 10193
rect 45004 10050 45044 10135
rect 44907 9932 44949 9941
rect 44907 9892 44908 9932
rect 44948 9892 44949 9932
rect 44907 9883 44949 9892
rect 44812 9724 45044 9764
rect 44427 8840 44469 8849
rect 44332 8800 44428 8840
rect 44468 8800 44469 8840
rect 44427 8791 44469 8800
rect 44428 8706 44468 8791
rect 44620 8756 44660 9136
rect 44620 8707 44660 8716
rect 44812 8672 44852 9724
rect 45004 9680 45044 9724
rect 45100 9680 45140 10144
rect 45772 10184 45812 10303
rect 45963 10268 46005 10277
rect 45963 10228 45964 10268
rect 46004 10228 46005 10268
rect 45963 10219 46005 10228
rect 45196 10100 45236 10109
rect 45388 10100 45428 10109
rect 45236 10060 45388 10100
rect 45196 10051 45236 10060
rect 45388 10051 45428 10060
rect 45772 9857 45812 10144
rect 45771 9848 45813 9857
rect 45771 9808 45772 9848
rect 45812 9808 45813 9848
rect 45771 9799 45813 9808
rect 45100 9640 45908 9680
rect 45004 9631 45044 9640
rect 45483 9428 45525 9437
rect 45483 9388 45484 9428
rect 45524 9388 45525 9428
rect 45483 9379 45525 9388
rect 45291 9344 45333 9353
rect 45291 9304 45292 9344
rect 45332 9304 45333 9344
rect 45291 9295 45333 9304
rect 45292 9210 45332 9295
rect 45484 9294 45524 9379
rect 45100 8924 45140 8933
rect 45140 8884 45428 8924
rect 45100 8875 45140 8884
rect 44907 8840 44949 8849
rect 44907 8800 44908 8840
rect 44948 8800 44949 8840
rect 44907 8791 44949 8800
rect 44812 8623 44852 8632
rect 44908 8672 44948 8791
rect 45099 8756 45141 8765
rect 45099 8716 45100 8756
rect 45140 8716 45141 8756
rect 45099 8707 45141 8716
rect 45388 8756 45428 8884
rect 45388 8707 45428 8716
rect 45484 8840 45524 8849
rect 44908 8623 44948 8632
rect 45100 8672 45140 8707
rect 45100 8621 45140 8632
rect 45291 8672 45333 8681
rect 45291 8632 45292 8672
rect 45332 8632 45333 8672
rect 45291 8630 45333 8632
rect 45291 8623 45292 8630
rect 45332 8623 45333 8630
rect 45292 8537 45332 8590
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 45196 8084 45236 8093
rect 45484 8084 45524 8800
rect 45580 8756 45620 9640
rect 45771 9428 45813 9437
rect 45771 9388 45772 9428
rect 45812 9388 45813 9428
rect 45771 9379 45813 9388
rect 45580 8707 45620 8716
rect 45676 8672 45716 8681
rect 45676 8597 45716 8632
rect 45675 8588 45717 8597
rect 45675 8548 45676 8588
rect 45716 8548 45717 8588
rect 45675 8539 45717 8548
rect 45579 8504 45621 8513
rect 45579 8464 45580 8504
rect 45620 8464 45621 8504
rect 45579 8455 45621 8464
rect 45236 8044 45524 8084
rect 45196 8035 45236 8044
rect 45580 8000 45620 8455
rect 45580 7951 45620 7960
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 45676 7421 45716 8539
rect 45675 7412 45717 7421
rect 45675 7372 45676 7412
rect 45716 7372 45717 7412
rect 45675 7363 45717 7372
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 45772 4985 45812 9379
rect 45868 9344 45908 9640
rect 45868 9295 45908 9304
rect 45964 8765 46004 10219
rect 46636 10184 46676 10195
rect 47116 10193 47156 11227
rect 48268 10865 48308 11572
rect 48844 10949 48884 16276
rect 48940 16073 48980 16158
rect 48939 16064 48981 16073
rect 48939 16024 48940 16064
rect 48980 16024 48981 16064
rect 48939 16015 48981 16024
rect 49036 15896 49076 19216
rect 49419 19088 49461 19097
rect 49419 19048 49420 19088
rect 49460 19048 49461 19088
rect 49419 19039 49461 19048
rect 49420 18954 49460 19039
rect 49612 18761 49652 19291
rect 49611 18752 49653 18761
rect 49611 18712 49612 18752
rect 49652 18712 49653 18752
rect 49611 18703 49653 18712
rect 49131 18584 49173 18593
rect 49131 18544 49132 18584
rect 49172 18544 49173 18584
rect 49131 18535 49173 18544
rect 49324 18584 49364 18593
rect 49132 18450 49172 18535
rect 49324 18425 49364 18544
rect 49420 18584 49460 18595
rect 49420 18509 49460 18544
rect 49419 18500 49461 18509
rect 49419 18460 49420 18500
rect 49460 18460 49461 18500
rect 49419 18451 49461 18460
rect 49323 18416 49365 18425
rect 49323 18376 49324 18416
rect 49364 18376 49365 18416
rect 49323 18367 49365 18376
rect 49612 18416 49652 18703
rect 49612 18367 49652 18376
rect 49131 18332 49173 18341
rect 49131 18292 49132 18332
rect 49172 18292 49173 18332
rect 49131 18283 49173 18292
rect 49707 18332 49749 18341
rect 49707 18292 49708 18332
rect 49748 18292 49749 18332
rect 49707 18283 49749 18292
rect 49132 18198 49172 18283
rect 49323 18164 49365 18173
rect 49323 18124 49324 18164
rect 49364 18124 49365 18164
rect 49323 18115 49365 18124
rect 49131 17828 49173 17837
rect 49131 17788 49132 17828
rect 49172 17788 49173 17828
rect 49131 17779 49173 17788
rect 49324 17828 49364 18115
rect 49708 18080 49748 18283
rect 49804 18164 49844 20560
rect 49899 20180 49941 20189
rect 49899 20140 49900 20180
rect 49940 20140 49941 20180
rect 49899 20131 49941 20140
rect 49900 19256 49940 20131
rect 49996 19685 50036 20812
rect 50380 20852 50420 20861
rect 50188 20600 50228 20609
rect 49995 19676 50037 19685
rect 49995 19636 49996 19676
rect 50036 19636 50037 19676
rect 49995 19627 50037 19636
rect 49900 19207 49940 19216
rect 50091 18836 50133 18845
rect 50091 18787 50092 18836
rect 50132 18787 50133 18836
rect 50092 18701 50132 18770
rect 49899 18584 49941 18593
rect 49899 18544 49900 18584
rect 49940 18544 49941 18584
rect 49899 18535 49941 18544
rect 49996 18584 50036 18593
rect 50188 18584 50228 20560
rect 50380 19937 50420 20812
rect 50571 20852 50613 20861
rect 50571 20812 50572 20852
rect 50612 20812 50613 20852
rect 50571 20803 50613 20812
rect 50572 20718 50612 20803
rect 50764 20600 50804 20609
rect 50764 20012 50804 20560
rect 50956 20012 50996 20021
rect 50764 19972 50956 20012
rect 50379 19928 50421 19937
rect 50379 19888 50380 19928
rect 50420 19888 50421 19928
rect 50379 19879 50421 19888
rect 50284 19172 50324 19181
rect 50284 18752 50324 19132
rect 50380 18929 50420 19879
rect 50764 19844 50804 19853
rect 50804 19804 50900 19844
rect 50764 19795 50804 19804
rect 50763 19676 50805 19685
rect 50763 19636 50764 19676
rect 50804 19636 50805 19676
rect 50763 19627 50805 19636
rect 50667 19256 50709 19265
rect 50667 19216 50668 19256
rect 50708 19216 50709 19256
rect 50667 19207 50709 19216
rect 50668 19122 50708 19207
rect 50379 18920 50421 18929
rect 50379 18880 50380 18920
rect 50420 18880 50421 18920
rect 50379 18871 50421 18880
rect 50284 18703 50324 18712
rect 50379 18752 50421 18761
rect 50379 18712 50380 18752
rect 50420 18712 50421 18752
rect 50379 18703 50421 18712
rect 50036 18544 50228 18584
rect 49996 18535 50036 18544
rect 49900 18450 49940 18535
rect 50188 18173 50228 18544
rect 50380 18584 50420 18703
rect 50380 18535 50420 18544
rect 50476 18584 50516 18593
rect 50476 18341 50516 18544
rect 50572 18584 50612 18593
rect 50572 18425 50612 18544
rect 50571 18416 50613 18425
rect 50571 18376 50572 18416
rect 50612 18376 50613 18416
rect 50571 18367 50613 18376
rect 50475 18332 50517 18341
rect 50475 18292 50476 18332
rect 50516 18292 50517 18332
rect 50475 18283 50517 18292
rect 49899 18164 49941 18173
rect 49804 18124 49900 18164
rect 49940 18124 49941 18164
rect 49899 18115 49941 18124
rect 50187 18164 50229 18173
rect 50187 18124 50188 18164
rect 50228 18124 50229 18164
rect 50187 18115 50229 18124
rect 49708 18040 49844 18080
rect 49419 17912 49461 17921
rect 49419 17872 49420 17912
rect 49460 17872 49461 17912
rect 49419 17863 49461 17872
rect 49707 17912 49749 17921
rect 49707 17872 49708 17912
rect 49748 17872 49749 17912
rect 49707 17863 49749 17872
rect 49132 17694 49172 17779
rect 48940 15856 49076 15896
rect 48940 13973 48980 15856
rect 49324 15737 49364 17788
rect 49323 15728 49365 15737
rect 49323 15688 49324 15728
rect 49364 15688 49365 15728
rect 49323 15679 49365 15688
rect 49035 15644 49077 15653
rect 49035 15604 49036 15644
rect 49076 15604 49077 15644
rect 49035 15595 49077 15604
rect 49036 15560 49076 15595
rect 49036 15509 49076 15520
rect 49131 15560 49173 15569
rect 49131 15520 49132 15560
rect 49172 15520 49173 15560
rect 49131 15511 49173 15520
rect 49228 15560 49268 15569
rect 49132 15426 49172 15511
rect 49132 14720 49172 14729
rect 49036 14680 49132 14720
rect 49036 14048 49076 14680
rect 49132 14671 49172 14680
rect 49131 14216 49173 14225
rect 49131 14176 49132 14216
rect 49172 14176 49173 14216
rect 49131 14167 49173 14176
rect 48939 13964 48981 13973
rect 48939 13924 48940 13964
rect 48980 13924 48981 13964
rect 48939 13915 48981 13924
rect 49036 13805 49076 14008
rect 49035 13796 49077 13805
rect 49035 13756 49036 13796
rect 49076 13756 49077 13796
rect 49035 13747 49077 13756
rect 49132 13217 49172 14167
rect 49228 14132 49268 15520
rect 49324 15560 49364 15569
rect 49324 14729 49364 15520
rect 49420 14981 49460 17863
rect 49611 17744 49653 17753
rect 49611 17704 49612 17744
rect 49652 17704 49653 17744
rect 49611 17695 49653 17704
rect 49708 17744 49748 17863
rect 49804 17828 49844 18040
rect 49804 17779 49844 17788
rect 49900 17912 49940 17921
rect 49708 17695 49748 17704
rect 49515 17576 49557 17585
rect 49515 17536 49516 17576
rect 49556 17536 49557 17576
rect 49515 17527 49557 17536
rect 49516 17442 49556 17527
rect 49612 16400 49652 17695
rect 49803 17408 49845 17417
rect 49803 17368 49804 17408
rect 49844 17368 49845 17408
rect 49803 17359 49845 17368
rect 49708 17072 49748 17081
rect 49708 16913 49748 17032
rect 49707 16904 49749 16913
rect 49707 16864 49708 16904
rect 49748 16864 49749 16904
rect 49707 16855 49749 16864
rect 49516 16360 49652 16400
rect 49516 15896 49556 16360
rect 49708 16316 49748 16325
rect 49804 16316 49844 17359
rect 49900 17156 49940 17872
rect 49995 17828 50037 17837
rect 49995 17788 49996 17828
rect 50036 17788 50037 17828
rect 49995 17779 50037 17788
rect 49996 17694 50036 17779
rect 50188 17753 50228 18115
rect 50092 17744 50132 17753
rect 50092 17417 50132 17704
rect 50187 17744 50229 17753
rect 50187 17704 50188 17744
rect 50228 17704 50229 17744
rect 50187 17695 50229 17704
rect 50572 17744 50612 18367
rect 50764 17921 50804 19627
rect 50860 18509 50900 19804
rect 50956 18761 50996 19972
rect 51340 20012 51380 21736
rect 51436 20189 51476 22240
rect 51532 21608 51572 22819
rect 51916 21785 51956 23491
rect 52011 23372 52053 23381
rect 52011 23332 52012 23372
rect 52052 23332 52053 23372
rect 52011 23323 52053 23332
rect 52012 23120 52052 23323
rect 52108 23129 52148 23214
rect 52012 23071 52052 23080
rect 52107 23120 52149 23129
rect 52107 23080 52108 23120
rect 52148 23080 52149 23120
rect 52107 23071 52149 23080
rect 52204 22280 52244 23836
rect 52300 23540 52340 24499
rect 52491 23876 52533 23885
rect 52491 23836 52492 23876
rect 52532 23836 52533 23876
rect 52491 23827 52533 23836
rect 52299 23500 52340 23540
rect 52299 23456 52339 23500
rect 52299 23416 52340 23456
rect 52300 23372 52340 23416
rect 52492 23381 52532 23827
rect 52299 23332 52340 23372
rect 52491 23372 52533 23381
rect 52491 23332 52492 23372
rect 52532 23332 52533 23372
rect 52299 23288 52339 23332
rect 52491 23323 52533 23332
rect 52299 23248 52340 23288
rect 52300 23120 52340 23248
rect 52395 23204 52437 23213
rect 52395 23164 52396 23204
rect 52436 23164 52437 23204
rect 52395 23155 52437 23164
rect 52300 23071 52340 23080
rect 52396 23070 52436 23155
rect 52588 23045 52628 24592
rect 52684 24583 52724 24592
rect 52684 23120 52724 23129
rect 52587 23036 52629 23045
rect 52587 22996 52588 23036
rect 52628 22996 52629 23036
rect 52587 22987 52629 22996
rect 52587 22868 52629 22877
rect 52587 22828 52588 22868
rect 52628 22828 52629 22868
rect 52587 22819 52629 22828
rect 52588 22734 52628 22819
rect 52684 22793 52724 23080
rect 52683 22784 52725 22793
rect 52683 22744 52684 22784
rect 52724 22744 52725 22784
rect 52683 22735 52725 22744
rect 52395 22532 52437 22541
rect 52395 22492 52396 22532
rect 52436 22492 52437 22532
rect 52395 22483 52437 22492
rect 52684 22532 52724 22735
rect 52684 22483 52724 22492
rect 52396 22398 52436 22483
rect 52588 22280 52628 22289
rect 52204 22240 52588 22280
rect 52628 22240 52724 22280
rect 52588 22231 52628 22240
rect 52396 22112 52436 22121
rect 51915 21776 51957 21785
rect 51915 21736 51916 21776
rect 51956 21736 51957 21776
rect 51915 21727 51957 21736
rect 52396 21701 52436 22072
rect 52395 21692 52437 21701
rect 52395 21652 52396 21692
rect 52436 21652 52437 21692
rect 52395 21643 52437 21652
rect 51532 20945 51572 21568
rect 51820 21608 51860 21617
rect 52203 21608 52245 21617
rect 51627 21356 51669 21365
rect 51627 21316 51628 21356
rect 51668 21316 51669 21356
rect 51627 21307 51669 21316
rect 51628 21222 51668 21307
rect 51820 21281 51860 21568
rect 52108 21568 52204 21608
rect 52244 21568 52245 21608
rect 51915 21356 51957 21365
rect 51915 21316 51916 21356
rect 51956 21316 51957 21356
rect 51915 21307 51957 21316
rect 51819 21272 51861 21281
rect 51819 21232 51820 21272
rect 51860 21232 51861 21272
rect 51819 21223 51861 21232
rect 51916 21222 51956 21307
rect 51531 20936 51573 20945
rect 51531 20896 51532 20936
rect 51572 20896 51573 20936
rect 51531 20887 51573 20896
rect 52108 20525 52148 21568
rect 52203 21559 52245 21568
rect 52491 21608 52533 21617
rect 52491 21568 52492 21608
rect 52532 21568 52533 21608
rect 52491 21559 52533 21568
rect 52204 21474 52244 21559
rect 52300 21356 52340 21365
rect 52300 21029 52340 21316
rect 52492 21113 52532 21559
rect 52587 21440 52629 21449
rect 52587 21400 52588 21440
rect 52628 21400 52629 21440
rect 52587 21391 52629 21400
rect 52588 21306 52628 21391
rect 52491 21104 52533 21113
rect 52491 21064 52492 21104
rect 52532 21064 52533 21104
rect 52491 21055 52533 21064
rect 52299 21020 52341 21029
rect 52299 20980 52300 21020
rect 52340 20980 52341 21020
rect 52299 20971 52341 20980
rect 52491 20936 52533 20945
rect 52491 20896 52492 20936
rect 52532 20896 52533 20936
rect 52491 20887 52533 20896
rect 52492 20802 52532 20887
rect 52588 20777 52628 20862
rect 52203 20768 52245 20777
rect 52203 20728 52204 20768
rect 52244 20728 52245 20768
rect 52203 20719 52245 20728
rect 52587 20768 52629 20777
rect 52587 20728 52588 20768
rect 52628 20728 52629 20768
rect 52587 20719 52629 20728
rect 52107 20516 52149 20525
rect 52107 20476 52108 20516
rect 52148 20476 52149 20516
rect 52107 20467 52149 20476
rect 52204 20189 52244 20719
rect 52299 20600 52341 20609
rect 52684 20600 52724 22240
rect 52299 20560 52300 20600
rect 52340 20560 52341 20600
rect 52299 20551 52341 20560
rect 52588 20560 52724 20600
rect 52300 20466 52340 20551
rect 51435 20180 51477 20189
rect 51435 20140 51436 20180
rect 51476 20140 51477 20180
rect 51435 20131 51477 20140
rect 52203 20180 52245 20189
rect 52203 20140 52204 20180
rect 52244 20140 52245 20180
rect 52203 20131 52245 20140
rect 51340 19963 51380 19972
rect 51147 19928 51189 19937
rect 51147 19888 51148 19928
rect 51188 19888 51189 19928
rect 51147 19879 51189 19888
rect 51148 19794 51188 19879
rect 51436 19256 51476 20131
rect 51915 20012 51957 20021
rect 51915 19972 51916 20012
rect 51956 19972 51957 20012
rect 51915 19963 51957 19972
rect 51916 19878 51956 19963
rect 51532 19844 51572 19853
rect 51532 19685 51572 19804
rect 51724 19844 51764 19853
rect 51531 19676 51573 19685
rect 51531 19636 51532 19676
rect 51572 19636 51573 19676
rect 51531 19627 51573 19636
rect 51532 19256 51572 19265
rect 51436 19216 51532 19256
rect 51339 18836 51381 18845
rect 51339 18796 51340 18836
rect 51380 18796 51381 18836
rect 51339 18787 51381 18796
rect 50955 18752 50997 18761
rect 50955 18712 50956 18752
rect 50996 18712 50997 18752
rect 50955 18703 50997 18712
rect 51147 18668 51189 18677
rect 51147 18628 51148 18668
rect 51188 18628 51189 18668
rect 51147 18619 51189 18628
rect 50955 18584 50997 18593
rect 50955 18544 50956 18584
rect 50996 18544 50997 18584
rect 50955 18535 50997 18544
rect 51052 18584 51092 18593
rect 50859 18500 50901 18509
rect 50859 18460 50860 18500
rect 50900 18460 50901 18500
rect 50859 18451 50901 18460
rect 50763 17912 50805 17921
rect 50763 17872 50764 17912
rect 50804 17872 50805 17912
rect 50763 17863 50805 17872
rect 50572 17585 50612 17704
rect 50668 17744 50708 17753
rect 50476 17576 50516 17585
rect 50188 17536 50476 17576
rect 50091 17408 50133 17417
rect 50091 17368 50092 17408
rect 50132 17368 50133 17408
rect 50091 17359 50133 17368
rect 50092 17156 50132 17165
rect 49900 17116 50092 17156
rect 50092 17107 50132 17116
rect 50091 16988 50133 16997
rect 50091 16948 50092 16988
rect 50132 16948 50133 16988
rect 50091 16939 50133 16948
rect 50092 16400 50132 16939
rect 49748 16276 49844 16316
rect 49708 16267 49748 16276
rect 49611 16232 49653 16241
rect 49611 16192 49612 16232
rect 49652 16192 49653 16232
rect 49611 16183 49653 16192
rect 49612 16098 49652 16183
rect 49804 16064 49844 16276
rect 49996 16360 50132 16400
rect 49996 16241 50036 16360
rect 49995 16232 50037 16241
rect 49995 16192 49996 16232
rect 50036 16192 50037 16232
rect 49995 16183 50037 16192
rect 50092 16232 50132 16241
rect 50188 16232 50228 17536
rect 50476 17527 50516 17536
rect 50571 17576 50613 17585
rect 50571 17536 50572 17576
rect 50612 17536 50613 17576
rect 50571 17527 50613 17536
rect 50284 17072 50324 17081
rect 50324 17032 50420 17072
rect 50284 17023 50324 17032
rect 50283 16820 50325 16829
rect 50283 16780 50284 16820
rect 50324 16780 50325 16820
rect 50283 16771 50325 16780
rect 50284 16316 50324 16771
rect 50380 16745 50420 17032
rect 50572 16904 50612 17527
rect 50668 17240 50708 17704
rect 50763 17744 50805 17753
rect 50763 17704 50764 17744
rect 50804 17704 50805 17744
rect 50860 17744 50900 18451
rect 50956 18450 50996 18535
rect 51052 18425 51092 18544
rect 51148 18584 51188 18619
rect 51148 18533 51188 18544
rect 51244 18584 51284 18593
rect 51051 18416 51093 18425
rect 51051 18376 51052 18416
rect 51092 18376 51093 18416
rect 51051 18367 51093 18376
rect 51244 18173 51284 18544
rect 51243 18164 51285 18173
rect 51243 18124 51244 18164
rect 51284 18124 51285 18164
rect 51243 18115 51285 18124
rect 51052 17996 51092 18005
rect 51340 17996 51380 18787
rect 51435 18500 51477 18509
rect 51435 18460 51436 18500
rect 51476 18460 51477 18500
rect 51435 18451 51477 18460
rect 51092 17956 51380 17996
rect 51052 17947 51092 17956
rect 51051 17828 51093 17837
rect 51051 17788 51052 17828
rect 51092 17788 51093 17828
rect 51051 17779 51093 17788
rect 50956 17744 50996 17753
rect 50860 17704 50956 17744
rect 50763 17695 50805 17704
rect 50956 17695 50996 17704
rect 50764 17610 50804 17695
rect 51052 17576 51092 17779
rect 51340 17744 51380 17753
rect 50956 17536 51092 17576
rect 51244 17576 51284 17585
rect 50668 17200 50804 17240
rect 50476 16864 50612 16904
rect 50668 17072 50708 17081
rect 50379 16736 50421 16745
rect 50379 16696 50380 16736
rect 50420 16696 50421 16736
rect 50379 16687 50421 16696
rect 50379 16568 50421 16577
rect 50379 16528 50380 16568
rect 50420 16528 50421 16568
rect 50379 16519 50421 16528
rect 50380 16484 50420 16519
rect 50380 16433 50420 16444
rect 50284 16276 50420 16316
rect 50132 16192 50228 16232
rect 50092 16183 50132 16192
rect 49996 16098 50036 16183
rect 49900 16064 49940 16069
rect 49804 16060 49940 16064
rect 49804 16024 49900 16060
rect 49900 16011 49940 16020
rect 49516 15856 50036 15896
rect 49803 15644 49845 15653
rect 49803 15604 49804 15644
rect 49844 15604 49845 15644
rect 49803 15595 49845 15604
rect 49708 15560 49748 15569
rect 49612 15520 49708 15560
rect 49419 14972 49461 14981
rect 49419 14932 49420 14972
rect 49460 14932 49461 14972
rect 49419 14923 49461 14932
rect 49323 14720 49365 14729
rect 49323 14680 49324 14720
rect 49364 14680 49365 14720
rect 49323 14671 49365 14680
rect 49515 14300 49557 14309
rect 49515 14260 49516 14300
rect 49556 14260 49557 14300
rect 49515 14251 49557 14260
rect 49516 14141 49556 14251
rect 49323 14132 49365 14141
rect 49228 14092 49324 14132
rect 49364 14092 49365 14132
rect 49323 14083 49365 14092
rect 49515 14132 49557 14141
rect 49515 14092 49516 14132
rect 49556 14092 49557 14132
rect 49515 14083 49557 14092
rect 49324 13460 49364 14083
rect 49419 13544 49461 13553
rect 49419 13504 49420 13544
rect 49460 13504 49461 13544
rect 49419 13495 49461 13504
rect 49324 13411 49364 13420
rect 49131 13208 49173 13217
rect 49131 13168 49132 13208
rect 49172 13168 49173 13208
rect 49131 13159 49173 13168
rect 49132 12704 49172 13159
rect 49228 12704 49268 12713
rect 49132 12664 49228 12704
rect 49228 12655 49268 12664
rect 48939 12284 48981 12293
rect 48939 12244 48940 12284
rect 48980 12244 48981 12284
rect 48939 12235 48981 12244
rect 48843 10940 48885 10949
rect 48843 10900 48844 10940
rect 48884 10900 48885 10940
rect 48843 10891 48885 10900
rect 48267 10856 48309 10865
rect 48267 10816 48268 10856
rect 48308 10816 48309 10856
rect 48267 10807 48309 10816
rect 48940 10445 48980 12235
rect 49420 11192 49460 13495
rect 49612 13208 49652 15520
rect 49708 15511 49748 15520
rect 49804 15560 49844 15595
rect 49804 15509 49844 15520
rect 49900 15560 49940 15571
rect 49900 15485 49940 15520
rect 49996 15560 50036 15856
rect 50036 15520 50132 15560
rect 49996 15511 50036 15520
rect 49899 15476 49941 15485
rect 49899 15436 49900 15476
rect 49940 15436 49941 15476
rect 49899 15427 49941 15436
rect 49995 14720 50037 14729
rect 49995 14680 49996 14720
rect 50036 14680 50037 14720
rect 49995 14671 50037 14680
rect 49996 14586 50036 14671
rect 50092 14309 50132 15520
rect 49707 14300 49749 14309
rect 49707 14260 49708 14300
rect 49748 14260 49749 14300
rect 49707 14251 49749 14260
rect 50091 14300 50133 14309
rect 50091 14260 50092 14300
rect 50132 14260 50133 14300
rect 50091 14251 50133 14260
rect 49612 13159 49652 13168
rect 49708 13208 49748 14251
rect 49803 14048 49845 14057
rect 49803 14008 49804 14048
rect 49844 14008 49845 14048
rect 49803 13999 49845 14008
rect 49900 14048 49940 14057
rect 49804 13385 49844 13999
rect 49803 13376 49845 13385
rect 49803 13336 49804 13376
rect 49844 13336 49845 13376
rect 49803 13327 49845 13336
rect 49708 13159 49748 13168
rect 49804 13036 49844 13327
rect 49804 12987 49844 12996
rect 49803 12788 49845 12797
rect 49803 12748 49804 12788
rect 49844 12748 49845 12788
rect 49803 12739 49845 12748
rect 49515 12704 49557 12713
rect 49515 12664 49516 12704
rect 49556 12664 49557 12704
rect 49515 12655 49557 12664
rect 49804 12704 49844 12739
rect 49900 12713 49940 14008
rect 50187 13880 50229 13889
rect 50187 13840 50188 13880
rect 50228 13840 50229 13880
rect 50187 13831 50229 13840
rect 49516 11696 49556 12655
rect 49804 12653 49844 12664
rect 49899 12704 49941 12713
rect 49899 12664 49900 12704
rect 49940 12664 49941 12704
rect 49899 12655 49941 12664
rect 49707 12620 49749 12629
rect 49707 12580 49708 12620
rect 49748 12580 49749 12620
rect 49707 12571 49749 12580
rect 49708 12536 49748 12571
rect 49708 12485 49748 12496
rect 49900 12536 49940 12545
rect 49900 12461 49940 12496
rect 49995 12536 50037 12545
rect 49995 12496 49996 12536
rect 50036 12496 50037 12536
rect 49995 12487 50037 12496
rect 49899 12452 49941 12461
rect 49899 12412 49900 12452
rect 49940 12412 49941 12452
rect 49899 12403 49941 12412
rect 49516 11647 49556 11656
rect 49420 11143 49460 11152
rect 49323 11108 49365 11117
rect 49323 11068 49324 11108
rect 49364 11068 49365 11108
rect 49323 11059 49365 11068
rect 49324 11024 49364 11059
rect 47787 10436 47829 10445
rect 47787 10396 47788 10436
rect 47828 10396 47829 10436
rect 47787 10387 47829 10396
rect 48939 10436 48981 10445
rect 48939 10396 48940 10436
rect 48980 10396 48981 10436
rect 48939 10387 48981 10396
rect 47788 10302 47828 10387
rect 46636 10109 46676 10144
rect 47115 10184 47157 10193
rect 47115 10144 47116 10184
rect 47156 10144 47157 10184
rect 47115 10135 47157 10144
rect 48364 10184 48404 10193
rect 49228 10184 49268 10193
rect 48404 10144 48500 10184
rect 48364 10135 48404 10144
rect 46443 10100 46485 10109
rect 46443 10060 46444 10100
rect 46484 10060 46485 10100
rect 46443 10051 46485 10060
rect 46635 10100 46677 10109
rect 46635 10060 46636 10100
rect 46676 10060 46677 10100
rect 46635 10051 46677 10060
rect 47019 10100 47061 10109
rect 47019 10060 47020 10100
rect 47060 10060 47061 10100
rect 47019 10051 47061 10060
rect 46251 10016 46293 10025
rect 46251 9976 46252 10016
rect 46292 9976 46293 10016
rect 46251 9967 46293 9976
rect 46059 9848 46101 9857
rect 46059 9808 46060 9848
rect 46100 9808 46101 9848
rect 46059 9799 46101 9808
rect 45963 8756 46005 8765
rect 45963 8716 45964 8756
rect 46004 8716 46005 8756
rect 45963 8707 46005 8716
rect 46060 8681 46100 9799
rect 46252 9605 46292 9967
rect 46348 9684 46388 9693
rect 46251 9596 46293 9605
rect 46251 9556 46252 9596
rect 46292 9556 46293 9596
rect 46251 9547 46293 9556
rect 46155 9512 46197 9521
rect 46155 9472 46156 9512
rect 46196 9472 46197 9512
rect 46155 9463 46197 9472
rect 46252 9512 46292 9547
rect 46156 9378 46196 9463
rect 46252 9462 46292 9472
rect 46059 8672 46101 8681
rect 46059 8632 46060 8672
rect 46100 8632 46101 8672
rect 46059 8623 46101 8632
rect 46348 8597 46388 9644
rect 46444 8681 46484 10051
rect 46635 9932 46677 9941
rect 46635 9892 46636 9932
rect 46676 9892 46677 9932
rect 46635 9883 46677 9892
rect 46539 9512 46581 9521
rect 46539 9472 46540 9512
rect 46580 9472 46581 9512
rect 46539 9463 46581 9472
rect 46636 9512 46676 9883
rect 47020 9605 47060 10051
rect 47116 9680 47156 10135
rect 47980 10100 48020 10109
rect 47116 9631 47156 9640
rect 47788 10016 47828 10025
rect 46827 9596 46869 9605
rect 46827 9556 46828 9596
rect 46868 9556 46869 9596
rect 46827 9547 46869 9556
rect 47019 9596 47061 9605
rect 47019 9556 47020 9596
rect 47060 9556 47061 9596
rect 47019 9547 47061 9556
rect 46636 9463 46676 9472
rect 46731 9512 46773 9521
rect 46731 9472 46732 9512
rect 46772 9472 46773 9512
rect 46731 9463 46773 9472
rect 46828 9512 46868 9547
rect 47788 9521 47828 9976
rect 47980 9680 48020 10060
rect 48363 9932 48405 9941
rect 48363 9892 48364 9932
rect 48404 9892 48405 9932
rect 48363 9883 48405 9892
rect 48267 9764 48309 9773
rect 48267 9724 48268 9764
rect 48308 9724 48309 9764
rect 48267 9715 48309 9724
rect 48076 9680 48116 9689
rect 47980 9640 48076 9680
rect 48076 9631 48116 9640
rect 46540 9378 46580 9463
rect 46732 9378 46772 9463
rect 46828 9461 46868 9472
rect 47211 9512 47253 9521
rect 47211 9472 47212 9512
rect 47252 9472 47253 9512
rect 47211 9463 47253 9472
rect 47787 9512 47829 9521
rect 47787 9472 47788 9512
rect 47828 9472 47829 9512
rect 47787 9463 47829 9472
rect 48172 9512 48212 9521
rect 47212 9378 47252 9463
rect 47595 8840 47637 8849
rect 47595 8800 47596 8840
rect 47636 8800 47637 8840
rect 47595 8791 47637 8800
rect 46443 8672 46485 8681
rect 46443 8632 46444 8672
rect 46484 8632 46485 8672
rect 46443 8623 46485 8632
rect 47500 8672 47540 8681
rect 46347 8588 46389 8597
rect 46347 8548 46348 8588
rect 46388 8548 46389 8588
rect 46347 8539 46389 8548
rect 46444 8000 46484 8623
rect 47500 8168 47540 8632
rect 47596 8672 47636 8791
rect 47787 8756 47829 8765
rect 47787 8716 47788 8756
rect 47828 8716 47829 8756
rect 47787 8707 47829 8716
rect 48172 8756 48212 9472
rect 48268 9512 48308 9715
rect 48268 9463 48308 9472
rect 48364 9512 48404 9883
rect 48460 9857 48500 10144
rect 49036 10144 49228 10184
rect 48459 9848 48501 9857
rect 48459 9808 48460 9848
rect 48500 9808 48501 9848
rect 48459 9799 48501 9808
rect 48364 9017 48404 9472
rect 48363 9008 48405 9017
rect 48363 8968 48364 9008
rect 48404 8968 48405 9008
rect 48363 8959 48405 8968
rect 48364 8840 48404 8849
rect 48364 8756 48404 8800
rect 48172 8716 48404 8756
rect 47596 8623 47636 8632
rect 47788 8672 47828 8707
rect 47788 8621 47828 8632
rect 47692 8504 47732 8513
rect 47732 8464 47828 8504
rect 47692 8455 47732 8464
rect 47596 8168 47636 8177
rect 47500 8128 47596 8168
rect 47596 8119 47636 8128
rect 46444 7951 46484 7960
rect 46923 7748 46965 7757
rect 46923 7708 46924 7748
rect 46964 7708 46965 7748
rect 46923 7699 46965 7708
rect 47595 7748 47637 7757
rect 47595 7708 47596 7748
rect 47636 7708 47637 7748
rect 47595 7699 47637 7708
rect 46827 7412 46869 7421
rect 46827 7372 46828 7412
rect 46868 7372 46869 7412
rect 46827 7363 46869 7372
rect 46828 7278 46868 7363
rect 46924 7160 46964 7699
rect 47596 7614 47636 7699
rect 47788 7496 47828 8464
rect 47884 8000 47924 8009
rect 47884 7673 47924 7960
rect 47883 7664 47925 7673
rect 47883 7624 47884 7664
rect 47924 7624 47925 7664
rect 47883 7615 47925 7624
rect 48075 7580 48117 7589
rect 48075 7540 48076 7580
rect 48116 7540 48117 7580
rect 48075 7531 48117 7540
rect 47788 7456 48020 7496
rect 47980 7244 48020 7456
rect 48076 7328 48116 7531
rect 48076 7279 48116 7288
rect 47980 7195 48020 7204
rect 48172 7244 48212 8716
rect 48363 8588 48405 8597
rect 48363 8548 48364 8588
rect 48404 8548 48405 8588
rect 48363 8539 48405 8548
rect 48267 8000 48309 8009
rect 48267 7960 48268 8000
rect 48308 7960 48309 8000
rect 48267 7951 48309 7960
rect 48268 7866 48308 7951
rect 48172 7195 48212 7204
rect 46924 7111 46964 7120
rect 47883 7160 47925 7169
rect 47883 7120 47884 7160
rect 47924 7120 47925 7160
rect 47883 7111 47925 7120
rect 48268 7160 48308 7169
rect 48364 7160 48404 8539
rect 48460 8009 48500 9799
rect 48747 9596 48789 9605
rect 48747 9556 48748 9596
rect 48788 9556 48789 9596
rect 48747 9547 48789 9556
rect 48748 8765 48788 9547
rect 49036 9521 49076 10144
rect 49228 10135 49268 10144
rect 49324 10016 49364 10984
rect 49900 10856 49940 12403
rect 49996 12402 50036 12487
rect 50188 11285 50228 13831
rect 50380 13805 50420 16276
rect 50476 15653 50516 16864
rect 50668 16829 50708 17032
rect 50667 16820 50709 16829
rect 50667 16780 50668 16820
rect 50708 16780 50709 16820
rect 50667 16771 50709 16780
rect 50764 16745 50804 17200
rect 50571 16736 50613 16745
rect 50571 16696 50572 16736
rect 50612 16696 50613 16736
rect 50571 16687 50613 16696
rect 50763 16736 50805 16745
rect 50763 16696 50764 16736
rect 50804 16696 50805 16736
rect 50763 16687 50805 16696
rect 50572 16232 50612 16687
rect 50859 16652 50901 16661
rect 50859 16612 50860 16652
rect 50900 16612 50901 16652
rect 50859 16603 50901 16612
rect 50667 16568 50709 16577
rect 50667 16528 50668 16568
rect 50708 16528 50709 16568
rect 50667 16519 50709 16528
rect 50572 16183 50612 16192
rect 50668 16232 50708 16519
rect 50860 16484 50900 16603
rect 50668 16183 50708 16192
rect 50764 16444 50900 16484
rect 50764 16232 50804 16444
rect 50764 16183 50804 16192
rect 50860 16232 50900 16241
rect 50571 16064 50613 16073
rect 50571 16024 50572 16064
rect 50612 16024 50613 16064
rect 50571 16015 50613 16024
rect 50475 15644 50517 15653
rect 50475 15604 50476 15644
rect 50516 15604 50517 15644
rect 50475 15595 50517 15604
rect 50379 13796 50421 13805
rect 50379 13756 50380 13796
rect 50420 13756 50421 13796
rect 50379 13747 50421 13756
rect 50283 13376 50325 13385
rect 50283 13336 50284 13376
rect 50324 13336 50325 13376
rect 50283 13327 50325 13336
rect 50284 13242 50324 13327
rect 50379 13208 50421 13217
rect 50379 13168 50380 13208
rect 50420 13168 50421 13208
rect 50379 13159 50421 13168
rect 50380 13074 50420 13159
rect 50283 13040 50325 13049
rect 50283 13000 50284 13040
rect 50324 13000 50325 13040
rect 50283 12991 50325 13000
rect 50187 11276 50229 11285
rect 50187 11236 50188 11276
rect 50228 11236 50229 11276
rect 50187 11227 50229 11236
rect 50284 11108 50324 12991
rect 50572 12980 50612 16015
rect 50860 15653 50900 16192
rect 50956 16073 50996 17536
rect 51244 16661 51284 17536
rect 51340 16745 51380 17704
rect 51339 16736 51381 16745
rect 51339 16696 51340 16736
rect 51380 16696 51381 16736
rect 51339 16687 51381 16696
rect 51243 16652 51285 16661
rect 51243 16612 51244 16652
rect 51284 16612 51285 16652
rect 51243 16603 51285 16612
rect 51052 16232 51092 16243
rect 51052 16157 51092 16192
rect 51051 16148 51093 16157
rect 51051 16108 51052 16148
rect 51092 16108 51093 16148
rect 51051 16099 51093 16108
rect 50955 16064 50997 16073
rect 50955 16024 50956 16064
rect 50996 16024 50997 16064
rect 50955 16015 50997 16024
rect 50859 15644 50901 15653
rect 50859 15604 50860 15644
rect 50900 15604 50901 15644
rect 50859 15595 50901 15604
rect 50860 14477 50900 15595
rect 51052 15485 51092 16099
rect 51147 16064 51189 16073
rect 51147 16024 51148 16064
rect 51188 16024 51189 16064
rect 51147 16015 51189 16024
rect 51148 15930 51188 16015
rect 51436 15905 51476 18451
rect 51532 17072 51572 19216
rect 51627 19256 51669 19265
rect 51627 19216 51628 19256
rect 51668 19216 51669 19256
rect 51627 19207 51669 19216
rect 51628 18752 51668 19207
rect 51628 18703 51668 18712
rect 51724 18509 51764 19804
rect 52011 19004 52053 19013
rect 52011 18964 52012 19004
rect 52052 18964 52053 19004
rect 52011 18955 52053 18964
rect 51819 18668 51861 18677
rect 51819 18628 51820 18668
rect 51860 18628 51861 18668
rect 51819 18619 51861 18628
rect 51820 18584 51860 18619
rect 51820 18533 51860 18544
rect 51723 18500 51765 18509
rect 51723 18460 51724 18500
rect 51764 18460 51765 18500
rect 51723 18451 51765 18460
rect 51819 18416 51861 18425
rect 51819 18376 51820 18416
rect 51860 18376 51861 18416
rect 51819 18367 51861 18376
rect 51532 17023 51572 17032
rect 51628 18332 51668 18341
rect 51628 16829 51668 18292
rect 51627 16820 51669 16829
rect 51627 16780 51628 16820
rect 51668 16780 51669 16820
rect 51627 16771 51669 16780
rect 51627 16232 51669 16241
rect 51627 16192 51628 16232
rect 51668 16192 51669 16232
rect 51627 16183 51669 16192
rect 51435 15896 51477 15905
rect 51435 15856 51436 15896
rect 51476 15856 51477 15896
rect 51435 15847 51477 15856
rect 51051 15476 51093 15485
rect 51051 15436 51052 15476
rect 51092 15436 51093 15476
rect 51051 15427 51093 15436
rect 51052 15308 51092 15427
rect 50956 15268 51092 15308
rect 50956 14972 50996 15268
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 51148 14972 51188 14981
rect 50956 14932 51148 14972
rect 51148 14923 51188 14932
rect 51531 14888 51573 14897
rect 51531 14848 51532 14888
rect 51572 14848 51573 14888
rect 51531 14839 51573 14848
rect 51339 14720 51381 14729
rect 51339 14680 51340 14720
rect 51380 14680 51381 14720
rect 51339 14671 51381 14680
rect 51340 14586 51380 14671
rect 50859 14468 50901 14477
rect 50859 14428 50860 14468
rect 50900 14428 50901 14468
rect 50859 14419 50901 14428
rect 51532 14132 51572 14839
rect 51628 14813 51668 16183
rect 51820 15149 51860 18367
rect 51915 18332 51957 18341
rect 51915 18292 51916 18332
rect 51956 18292 51957 18332
rect 51915 18283 51957 18292
rect 51916 15821 51956 18283
rect 52012 16829 52052 18955
rect 52396 17744 52436 17753
rect 52588 17744 52628 20560
rect 52684 19088 52724 19097
rect 52684 18677 52724 19048
rect 52683 18668 52725 18677
rect 52683 18628 52684 18668
rect 52724 18628 52725 18668
rect 52683 18619 52725 18628
rect 52684 17744 52724 17753
rect 52588 17704 52684 17744
rect 52300 17576 52340 17585
rect 52396 17576 52436 17704
rect 52684 17695 52724 17704
rect 52588 17576 52628 17585
rect 52396 17536 52588 17576
rect 52300 16913 52340 17536
rect 52588 16997 52628 17536
rect 52876 17249 52916 26608
rect 53260 26405 53300 26692
rect 53356 26657 53396 28288
rect 53451 28288 53452 28328
rect 53492 28288 53493 28328
rect 53451 28279 53493 28288
rect 53452 26816 53492 28279
rect 53548 27656 53588 27665
rect 53548 27329 53588 27616
rect 53547 27320 53589 27329
rect 53547 27280 53548 27320
rect 53588 27280 53589 27320
rect 53547 27271 53589 27280
rect 53548 26993 53588 27271
rect 53547 26984 53589 26993
rect 53547 26944 53548 26984
rect 53588 26944 53589 26984
rect 53547 26935 53589 26944
rect 53740 26944 54260 26984
rect 53452 26767 53492 26776
rect 53548 26816 53588 26825
rect 53548 26657 53588 26776
rect 53644 26816 53684 26825
rect 53355 26648 53397 26657
rect 53355 26608 53356 26648
rect 53396 26608 53397 26648
rect 53355 26599 53397 26608
rect 53547 26648 53589 26657
rect 53547 26608 53548 26648
rect 53588 26608 53589 26648
rect 53547 26599 53589 26608
rect 53644 26489 53684 26776
rect 53740 26816 53780 26944
rect 53740 26767 53780 26776
rect 53931 26816 53973 26825
rect 53931 26776 53932 26816
rect 53972 26776 53973 26816
rect 53931 26767 53973 26776
rect 53355 26480 53397 26489
rect 53355 26440 53356 26480
rect 53396 26440 53397 26480
rect 53355 26431 53397 26440
rect 53643 26480 53685 26489
rect 53643 26440 53644 26480
rect 53684 26440 53685 26480
rect 53643 26431 53685 26440
rect 53259 26396 53301 26405
rect 53259 26356 53260 26396
rect 53300 26356 53301 26396
rect 53259 26347 53301 26356
rect 53163 26144 53205 26153
rect 53163 26104 53164 26144
rect 53204 26104 53205 26144
rect 53163 26095 53205 26104
rect 53356 26144 53396 26431
rect 53835 26396 53877 26405
rect 53835 26356 53836 26396
rect 53876 26356 53877 26396
rect 53932 26396 53972 26767
rect 54027 26648 54069 26657
rect 54027 26608 54028 26648
rect 54068 26608 54069 26648
rect 54027 26599 54069 26608
rect 54028 26514 54068 26599
rect 54123 26480 54165 26489
rect 54123 26440 54124 26480
rect 54164 26440 54165 26480
rect 54123 26431 54165 26440
rect 53932 26356 54068 26396
rect 53835 26347 53877 26356
rect 53356 26095 53396 26104
rect 53452 26144 53492 26153
rect 53644 26144 53684 26153
rect 53492 26104 53644 26144
rect 53452 26095 53492 26104
rect 53164 26010 53204 26095
rect 53067 25892 53109 25901
rect 53067 25852 53068 25892
rect 53108 25852 53109 25892
rect 53067 25843 53109 25852
rect 53068 25229 53108 25843
rect 53067 25220 53109 25229
rect 53067 25180 53068 25220
rect 53108 25180 53109 25220
rect 53067 25171 53109 25180
rect 53644 25132 53684 26104
rect 53740 26060 53780 26069
rect 53740 25556 53780 26020
rect 53836 25976 53876 26347
rect 54028 26144 54068 26356
rect 54124 26153 54164 26431
rect 53932 26060 53972 26071
rect 53932 25985 53972 26020
rect 53836 25927 53876 25936
rect 53931 25976 53973 25985
rect 53931 25936 53932 25976
rect 53972 25936 53973 25976
rect 53931 25927 53973 25936
rect 54028 25901 54068 26104
rect 54123 26144 54165 26153
rect 54123 26104 54124 26144
rect 54164 26104 54165 26144
rect 54123 26095 54165 26104
rect 54220 25976 54260 26944
rect 54316 26060 54356 28867
rect 54411 28328 54453 28337
rect 54411 28288 54412 28328
rect 54452 28288 54453 28328
rect 54411 28279 54453 28288
rect 54412 27656 54452 28279
rect 54412 27413 54452 27616
rect 54411 27404 54453 27413
rect 54411 27364 54412 27404
rect 54452 27364 54453 27404
rect 54411 27355 54453 27364
rect 54412 26060 54452 26069
rect 54316 26020 54412 26060
rect 54412 26011 54452 26020
rect 54220 25936 54356 25976
rect 54027 25892 54069 25901
rect 54027 25852 54028 25892
rect 54068 25852 54069 25892
rect 54027 25843 54069 25852
rect 54124 25556 54164 25565
rect 53740 25516 54124 25556
rect 54124 25507 54164 25516
rect 54219 25472 54261 25481
rect 54219 25432 54220 25472
rect 54260 25432 54261 25472
rect 54219 25423 54261 25432
rect 53739 25304 53781 25313
rect 53739 25264 53740 25304
rect 53780 25264 53781 25304
rect 53739 25255 53781 25264
rect 53836 25304 53876 25313
rect 54220 25304 54260 25423
rect 54316 25313 54356 25936
rect 54508 25649 54548 31564
rect 54604 31555 54644 31564
rect 54892 31520 54932 32824
rect 54987 32864 55029 32873
rect 54987 32824 54988 32864
rect 55028 32824 55029 32864
rect 54987 32815 55029 32824
rect 55084 32864 55124 33823
rect 55276 33704 55316 33916
rect 55468 33881 55508 33967
rect 55467 33876 55509 33881
rect 55467 33832 55468 33876
rect 55508 33832 55509 33876
rect 55467 33823 55509 33832
rect 55276 33655 55316 33664
rect 55372 33704 55412 33713
rect 55275 33452 55317 33461
rect 55275 33412 55276 33452
rect 55316 33412 55317 33452
rect 55275 33403 55317 33412
rect 55276 33032 55316 33403
rect 55372 33293 55412 33664
rect 55660 33704 55700 33713
rect 55467 33620 55509 33629
rect 55467 33580 55468 33620
rect 55508 33580 55509 33620
rect 55467 33571 55509 33580
rect 55371 33284 55413 33293
rect 55371 33244 55372 33284
rect 55412 33244 55413 33284
rect 55371 33235 55413 33244
rect 55276 32983 55316 32992
rect 55371 33032 55413 33041
rect 55371 32992 55372 33032
rect 55412 32992 55413 33032
rect 55371 32983 55413 32992
rect 55180 32948 55220 32959
rect 55180 32873 55220 32908
rect 55372 32948 55412 32983
rect 55372 32897 55412 32908
rect 55084 32815 55124 32824
rect 55179 32864 55221 32873
rect 55179 32824 55180 32864
rect 55220 32824 55221 32864
rect 55179 32815 55221 32824
rect 55468 32864 55508 33571
rect 55660 33377 55700 33664
rect 55755 33704 55797 33713
rect 55755 33664 55756 33704
rect 55796 33664 55797 33704
rect 55755 33655 55797 33664
rect 56044 33704 56084 34075
rect 56044 33655 56084 33664
rect 55659 33368 55701 33377
rect 55659 33328 55660 33368
rect 55700 33328 55701 33368
rect 55659 33319 55701 33328
rect 55756 33140 55796 33655
rect 55083 32696 55125 32705
rect 55083 32656 55084 32696
rect 55124 32656 55125 32696
rect 55083 32647 55125 32656
rect 54796 31480 54932 31520
rect 54603 30176 54645 30185
rect 54603 30136 54604 30176
rect 54644 30136 54645 30176
rect 54603 30127 54645 30136
rect 54604 29840 54644 30127
rect 54699 30092 54741 30101
rect 54796 30092 54836 31480
rect 54891 30680 54933 30689
rect 54891 30640 54892 30680
rect 54932 30640 54933 30680
rect 54891 30631 54933 30640
rect 54892 30546 54932 30631
rect 54699 30052 54700 30092
rect 54740 30052 54836 30092
rect 54699 30043 54741 30052
rect 54604 29791 54644 29800
rect 54700 29840 54740 30043
rect 55084 29924 55124 32647
rect 55275 31352 55317 31361
rect 55275 31312 55276 31352
rect 55316 31312 55317 31352
rect 55275 31303 55317 31312
rect 55372 31352 55412 31361
rect 55276 31218 55316 31303
rect 55372 30857 55412 31312
rect 55371 30848 55413 30857
rect 55371 30808 55372 30848
rect 55412 30808 55413 30848
rect 55371 30799 55413 30808
rect 55468 30260 55508 32824
rect 55660 33100 55796 33140
rect 55660 32192 55700 33100
rect 55851 33032 55893 33041
rect 55851 32992 55852 33032
rect 55892 32992 55893 33032
rect 55851 32983 55893 32992
rect 55852 32898 55892 32983
rect 56043 32864 56085 32873
rect 55852 32822 55892 32831
rect 55851 32782 55852 32789
rect 56043 32824 56044 32864
rect 56084 32824 56085 32864
rect 56043 32815 56085 32824
rect 56140 32864 56180 32873
rect 55892 32782 55893 32789
rect 55851 32780 55893 32782
rect 55851 32740 55852 32780
rect 55892 32740 55893 32780
rect 55851 32731 55893 32740
rect 55852 32687 55892 32731
rect 56044 32730 56084 32815
rect 55660 30689 55700 32152
rect 56140 31781 56180 32824
rect 56139 31772 56181 31781
rect 56139 31732 56140 31772
rect 56180 31732 56181 31772
rect 56139 31723 56181 31732
rect 56332 31604 56372 34588
rect 56428 33713 56468 35176
rect 56427 33704 56469 33713
rect 56427 33664 56428 33704
rect 56468 33664 56469 33704
rect 56427 33655 56469 33664
rect 56427 32780 56469 32789
rect 56427 32740 56428 32780
rect 56468 32740 56469 32780
rect 56427 32731 56469 32740
rect 56140 31564 56372 31604
rect 56043 30848 56085 30857
rect 56043 30808 56044 30848
rect 56084 30808 56085 30848
rect 56043 30799 56085 30808
rect 56044 30714 56084 30799
rect 55659 30680 55701 30689
rect 55659 30640 55660 30680
rect 55700 30640 55701 30680
rect 55659 30631 55701 30640
rect 55084 29875 55124 29884
rect 55372 30220 55508 30260
rect 56044 30428 56084 30437
rect 54700 29791 54740 29800
rect 54796 29840 54836 29849
rect 54796 28757 54836 29800
rect 54891 29840 54933 29849
rect 54891 29800 54892 29840
rect 54932 29800 54933 29840
rect 54891 29791 54933 29800
rect 54892 29513 54932 29791
rect 55276 29672 55316 29681
rect 55276 29513 55316 29632
rect 54891 29504 54933 29513
rect 54891 29464 54892 29504
rect 54932 29464 54933 29504
rect 54891 29455 54933 29464
rect 55275 29504 55317 29513
rect 55275 29464 55276 29504
rect 55316 29464 55317 29504
rect 55275 29455 55317 29464
rect 54892 29168 54932 29177
rect 54795 28748 54837 28757
rect 54795 28708 54796 28748
rect 54836 28708 54837 28748
rect 54795 28699 54837 28708
rect 54892 28337 54932 29128
rect 55179 29084 55221 29093
rect 55179 29044 55180 29084
rect 55220 29044 55221 29084
rect 55179 29035 55221 29044
rect 55083 28748 55125 28757
rect 55083 28708 55084 28748
rect 55124 28708 55125 28748
rect 55083 28699 55125 28708
rect 54891 28328 54933 28337
rect 54891 28288 54892 28328
rect 54932 28288 54933 28328
rect 54891 28279 54933 28288
rect 55084 28328 55124 28699
rect 55180 28580 55220 29035
rect 55180 28531 55220 28540
rect 55084 28279 55124 28288
rect 55275 28328 55317 28337
rect 55275 28288 55276 28328
rect 55316 28288 55317 28328
rect 55275 28279 55317 28288
rect 55180 28160 55220 28169
rect 55180 28001 55220 28120
rect 55179 27992 55221 28001
rect 55179 27952 55180 27992
rect 55220 27952 55221 27992
rect 55179 27943 55221 27952
rect 54987 27236 55029 27245
rect 54987 27196 54988 27236
rect 55028 27196 55029 27236
rect 54987 27187 55029 27196
rect 54603 26816 54645 26825
rect 54603 26776 54604 26816
rect 54644 26776 54645 26816
rect 54603 26767 54645 26776
rect 54604 26312 54644 26767
rect 54795 26396 54837 26405
rect 54795 26356 54796 26396
rect 54836 26356 54837 26396
rect 54795 26347 54837 26356
rect 54604 26263 54644 26272
rect 54796 26237 54836 26347
rect 54988 26237 55028 27187
rect 55180 26816 55220 26825
rect 55276 26816 55316 28279
rect 55220 26776 55316 26816
rect 55180 26767 55220 26776
rect 55083 26648 55125 26657
rect 55083 26608 55084 26648
rect 55124 26608 55125 26648
rect 55083 26599 55125 26608
rect 54795 26228 54837 26237
rect 54795 26188 54796 26228
rect 54836 26188 54837 26228
rect 54795 26179 54837 26188
rect 54987 26228 55029 26237
rect 54987 26188 54988 26228
rect 55028 26188 55029 26228
rect 54987 26179 55029 26188
rect 54796 26144 54836 26179
rect 54796 26093 54836 26104
rect 54988 26144 55028 26179
rect 55084 26153 55124 26599
rect 55372 26405 55412 30220
rect 55467 30092 55509 30101
rect 55467 30052 55468 30092
rect 55508 30052 55509 30092
rect 55467 30043 55509 30052
rect 55468 29958 55508 30043
rect 55660 29924 55700 29933
rect 55660 29345 55700 29884
rect 56044 29840 56084 30388
rect 56140 30101 56180 31564
rect 56428 30848 56468 32731
rect 56428 30799 56468 30808
rect 56524 32192 56564 32201
rect 56620 32192 56660 35587
rect 56812 34301 56852 35587
rect 57196 34553 57236 35848
rect 57292 35888 57332 35932
rect 57292 35839 57332 35848
rect 57388 35867 57428 35876
rect 57388 35645 57428 35827
rect 57387 35636 57429 35645
rect 57387 35596 57388 35636
rect 57428 35596 57429 35636
rect 57387 35587 57429 35596
rect 57484 35384 57524 35932
rect 57580 35888 57620 36931
rect 57675 35888 57717 35897
rect 57580 35848 57676 35888
rect 57716 35848 57717 35888
rect 57675 35839 57717 35848
rect 57868 35888 57908 35897
rect 57484 35335 57524 35344
rect 57484 34964 57524 34973
rect 57291 34628 57333 34637
rect 57291 34588 57292 34628
rect 57332 34588 57333 34628
rect 57291 34579 57333 34588
rect 57195 34544 57237 34553
rect 57100 34504 57196 34544
rect 57236 34504 57237 34544
rect 56811 34292 56853 34301
rect 56811 34252 56812 34292
rect 56852 34252 56853 34292
rect 56811 34243 56853 34252
rect 56564 32152 56660 32192
rect 56235 30596 56277 30605
rect 56235 30556 56236 30596
rect 56276 30556 56277 30596
rect 56235 30547 56277 30556
rect 56236 30462 56276 30547
rect 56428 30428 56468 30437
rect 56332 30388 56428 30428
rect 56139 30092 56181 30101
rect 56139 30052 56140 30092
rect 56180 30052 56181 30092
rect 56139 30043 56181 30052
rect 56044 29791 56084 29800
rect 56140 29840 56180 29849
rect 56140 29597 56180 29800
rect 56332 29840 56372 30388
rect 56428 30379 56468 30388
rect 56524 30353 56564 32152
rect 56812 31361 56852 34243
rect 56907 33704 56949 33713
rect 56907 33664 56908 33704
rect 56948 33664 56949 33704
rect 56907 33655 56949 33664
rect 56908 33570 56948 33655
rect 57100 32537 57140 34504
rect 57195 34495 57237 34504
rect 57292 34494 57332 34579
rect 57196 34376 57236 34385
rect 57196 34049 57236 34336
rect 57291 34208 57333 34217
rect 57291 34168 57292 34208
rect 57332 34168 57333 34208
rect 57291 34159 57333 34168
rect 57292 34074 57332 34159
rect 57484 34049 57524 34924
rect 57195 34040 57237 34049
rect 57195 34000 57196 34040
rect 57236 34000 57237 34040
rect 57195 33991 57237 34000
rect 57483 34040 57525 34049
rect 57483 34000 57484 34040
rect 57524 34000 57525 34040
rect 57483 33991 57525 34000
rect 57676 32789 57716 35839
rect 57771 35804 57813 35813
rect 57771 35764 57772 35804
rect 57812 35764 57813 35804
rect 57771 35755 57813 35764
rect 57772 35670 57812 35755
rect 57868 35729 57908 35848
rect 57964 35888 58004 37183
rect 58540 36560 58580 38200
rect 59692 38200 59884 38240
rect 58636 37400 58676 37409
rect 58636 36737 58676 37360
rect 59403 37400 59445 37409
rect 59403 37360 59404 37400
rect 59444 37360 59445 37400
rect 59403 37351 59445 37360
rect 59500 37400 59540 37411
rect 58827 37148 58869 37157
rect 58827 37108 58828 37148
rect 58868 37108 58869 37148
rect 58827 37099 58869 37108
rect 58635 36728 58677 36737
rect 58635 36688 58636 36728
rect 58676 36688 58677 36728
rect 58635 36679 58677 36688
rect 58828 36644 58868 37099
rect 59404 36896 59444 37351
rect 59500 37325 59540 37360
rect 59499 37316 59541 37325
rect 59499 37276 59500 37316
rect 59540 37276 59541 37316
rect 59499 37267 59541 37276
rect 59692 37241 59732 38200
rect 59884 38191 59924 38200
rect 61228 38240 61268 38249
rect 61420 38240 61460 38249
rect 61268 38200 61364 38240
rect 61228 38191 61268 38200
rect 59980 37988 60020 37997
rect 59884 37316 59924 37325
rect 59788 37276 59884 37316
rect 59691 37232 59733 37241
rect 59691 37192 59692 37232
rect 59732 37192 59733 37232
rect 59691 37183 59733 37192
rect 59404 36847 59444 36856
rect 59691 36896 59733 36905
rect 59691 36856 59692 36896
rect 59732 36856 59733 36896
rect 59691 36847 59733 36856
rect 59596 36728 59636 36737
rect 59212 36644 59252 36653
rect 58828 36595 58868 36604
rect 59116 36604 59212 36644
rect 58636 36560 58676 36569
rect 57964 35839 58004 35848
rect 58156 36520 58636 36560
rect 58156 35888 58196 36520
rect 58636 36511 58676 36520
rect 59020 36476 59060 36504
rect 59116 36476 59156 36604
rect 59212 36595 59252 36604
rect 59596 36485 59636 36688
rect 59692 36644 59732 36847
rect 59692 36595 59732 36604
rect 59788 36560 59828 37276
rect 59884 37267 59924 37276
rect 59980 36896 60020 37948
rect 61228 37988 61268 37997
rect 60268 37484 60308 37493
rect 60308 37444 60500 37484
rect 60268 37435 60308 37444
rect 60076 37232 60116 37243
rect 60076 37157 60116 37192
rect 60075 37148 60117 37157
rect 60075 37108 60076 37148
rect 60116 37108 60117 37148
rect 60075 37099 60117 37108
rect 60172 36900 60212 36909
rect 59980 36860 60172 36896
rect 59980 36856 60212 36860
rect 59980 36728 60020 36856
rect 60172 36851 60212 36856
rect 59980 36679 60020 36688
rect 60268 36728 60308 36737
rect 59883 36644 59925 36653
rect 59883 36604 59884 36644
rect 59924 36604 59925 36644
rect 59883 36595 59925 36604
rect 59788 36511 59828 36520
rect 59884 36510 59924 36595
rect 59060 36436 59156 36476
rect 59020 36427 59060 36436
rect 59019 36056 59061 36065
rect 59019 36016 59020 36056
rect 59060 36016 59061 36056
rect 59019 36007 59061 36016
rect 58444 35897 58484 35982
rect 58156 35839 58196 35848
rect 58252 35888 58292 35897
rect 58252 35729 58292 35848
rect 58443 35888 58485 35897
rect 58443 35848 58444 35888
rect 58484 35848 58485 35888
rect 58443 35839 58485 35848
rect 59020 35888 59060 36007
rect 59020 35839 59060 35848
rect 58636 35804 58676 35813
rect 58540 35764 58636 35804
rect 57867 35720 57909 35729
rect 57867 35680 57868 35720
rect 57908 35680 57909 35720
rect 57867 35671 57909 35680
rect 58251 35720 58293 35729
rect 58251 35680 58252 35720
rect 58292 35680 58293 35720
rect 58251 35671 58293 35680
rect 58348 35720 58388 35729
rect 58388 35680 58484 35720
rect 58348 35671 58388 35680
rect 57868 32873 57908 35671
rect 58348 35216 58388 35225
rect 58059 34376 58101 34385
rect 58059 34336 58060 34376
rect 58100 34336 58101 34376
rect 58059 34327 58101 34336
rect 58060 33872 58100 34327
rect 58060 33823 58100 33832
rect 58348 33629 58388 35176
rect 58444 35132 58484 35680
rect 58444 35083 58484 35092
rect 58540 35048 58580 35764
rect 58636 35755 58676 35764
rect 58731 35384 58773 35393
rect 58731 35344 58732 35384
rect 58772 35344 58773 35384
rect 58731 35335 58773 35344
rect 58732 35216 58772 35335
rect 58732 35167 58772 35176
rect 58540 34999 58580 35008
rect 58636 35132 58676 35141
rect 58636 35048 58676 35092
rect 58924 35048 58964 35057
rect 58636 35008 58924 35048
rect 58636 34796 58676 35008
rect 58924 34999 58964 35008
rect 58540 34756 58676 34796
rect 58540 34376 58580 34756
rect 58636 34385 58676 34470
rect 59116 34469 59156 36436
rect 59404 36476 59444 36485
rect 59404 36065 59444 36436
rect 59595 36476 59637 36485
rect 59595 36436 59596 36476
rect 59636 36436 59637 36476
rect 59595 36427 59637 36436
rect 59403 36056 59445 36065
rect 59403 36016 59404 36056
rect 59444 36016 59445 36056
rect 59403 36007 59445 36016
rect 59884 35888 59924 35897
rect 59404 35393 59444 35479
rect 59403 35388 59445 35393
rect 59403 35344 59404 35388
rect 59444 35344 59445 35388
rect 59403 35335 59445 35344
rect 59884 35225 59924 35848
rect 60268 35813 60308 36688
rect 60363 36728 60405 36737
rect 60363 36688 60364 36728
rect 60404 36688 60405 36728
rect 60363 36679 60405 36688
rect 60364 36594 60404 36679
rect 60267 35804 60309 35813
rect 60267 35764 60268 35804
rect 60308 35764 60309 35804
rect 60267 35755 60309 35764
rect 60171 35384 60213 35393
rect 60171 35344 60172 35384
rect 60212 35344 60213 35384
rect 60171 35335 60213 35344
rect 60172 35250 60212 35335
rect 60267 35300 60309 35309
rect 60267 35260 60268 35300
rect 60308 35260 60309 35300
rect 60267 35251 60309 35260
rect 59212 35216 59252 35225
rect 59115 34460 59157 34469
rect 58732 34420 59060 34460
rect 58540 34327 58580 34336
rect 58635 34376 58677 34385
rect 58635 34336 58636 34376
rect 58676 34336 58677 34376
rect 58635 34327 58677 34336
rect 58732 34376 58772 34420
rect 58732 34327 58772 34336
rect 58924 34292 58964 34301
rect 58444 34208 58484 34217
rect 58924 34208 58964 34252
rect 58484 34168 58964 34208
rect 58444 34159 58484 34168
rect 59020 33629 59060 34420
rect 59115 34420 59116 34460
rect 59156 34420 59157 34460
rect 59115 34411 59157 34420
rect 59212 33872 59252 35176
rect 59308 35216 59348 35225
rect 59883 35216 59925 35225
rect 59348 35176 59444 35216
rect 59308 35167 59348 35176
rect 59307 34460 59349 34469
rect 59307 34420 59308 34460
rect 59348 34420 59349 34460
rect 59307 34411 59349 34420
rect 59308 34376 59348 34411
rect 59308 34325 59348 34336
rect 59404 33965 59444 35176
rect 59883 35176 59884 35216
rect 59924 35176 59925 35216
rect 59883 35167 59925 35176
rect 60268 35216 60308 35251
rect 59884 34376 59924 35167
rect 60268 35165 60308 35176
rect 60460 35048 60500 37444
rect 60939 37400 60981 37409
rect 60939 37360 60940 37400
rect 60980 37360 60981 37400
rect 60939 37351 60981 37360
rect 60556 37316 60596 37325
rect 60596 37276 60884 37316
rect 60556 37267 60596 37276
rect 60844 36896 60884 37276
rect 60940 37266 60980 37351
rect 61228 36905 61268 37948
rect 60844 36847 60884 36856
rect 61227 36896 61269 36905
rect 61227 36856 61228 36896
rect 61268 36856 61269 36896
rect 61227 36847 61269 36856
rect 60940 36728 60980 36739
rect 60940 36653 60980 36688
rect 61036 36728 61076 36737
rect 60651 36644 60693 36653
rect 60651 36604 60652 36644
rect 60692 36604 60693 36644
rect 60651 36595 60693 36604
rect 60939 36644 60981 36653
rect 60939 36604 60940 36644
rect 60980 36604 60981 36644
rect 60939 36595 60981 36604
rect 60652 36560 60692 36595
rect 60652 36509 60692 36520
rect 60939 36476 60981 36485
rect 60939 36436 60940 36476
rect 60980 36436 60981 36476
rect 60939 36427 60981 36436
rect 60843 35888 60885 35897
rect 60843 35848 60844 35888
rect 60884 35848 60885 35888
rect 60843 35839 60885 35848
rect 60268 35008 60500 35048
rect 60172 34376 60212 34385
rect 59884 34336 60172 34376
rect 60172 34327 60212 34336
rect 59691 34208 59733 34217
rect 59691 34168 59692 34208
rect 59732 34168 59733 34208
rect 59691 34159 59733 34168
rect 59979 34208 60021 34217
rect 59979 34168 59980 34208
rect 60020 34168 60021 34208
rect 59979 34159 60021 34168
rect 59403 33956 59445 33965
rect 59403 33916 59404 33956
rect 59444 33916 59445 33956
rect 59403 33907 59445 33916
rect 59308 33872 59348 33881
rect 59212 33832 59308 33872
rect 59308 33823 59348 33832
rect 59595 33788 59637 33797
rect 59595 33748 59596 33788
rect 59636 33748 59637 33788
rect 59595 33739 59637 33748
rect 59404 33704 59444 33713
rect 58347 33620 58389 33629
rect 58347 33580 58348 33620
rect 58388 33580 58389 33620
rect 58347 33571 58389 33580
rect 59019 33620 59061 33629
rect 59019 33580 59020 33620
rect 59060 33580 59061 33620
rect 59019 33571 59061 33580
rect 59404 33545 59444 33664
rect 59499 33704 59541 33713
rect 59499 33664 59500 33704
rect 59540 33664 59541 33704
rect 59499 33655 59541 33664
rect 59596 33704 59636 33739
rect 59500 33570 59540 33655
rect 59596 33653 59636 33664
rect 59403 33536 59445 33545
rect 59403 33496 59404 33536
rect 59444 33496 59445 33536
rect 59403 33487 59445 33496
rect 58060 33452 58100 33461
rect 58060 33140 58100 33412
rect 57964 33100 58100 33140
rect 57867 32864 57909 32873
rect 57867 32824 57868 32864
rect 57908 32824 57909 32864
rect 57867 32815 57909 32824
rect 57675 32780 57717 32789
rect 57675 32740 57676 32780
rect 57716 32740 57717 32780
rect 57675 32731 57717 32740
rect 57099 32528 57141 32537
rect 57099 32488 57100 32528
rect 57140 32488 57141 32528
rect 57099 32479 57141 32488
rect 56908 32320 57428 32360
rect 56908 32276 56948 32320
rect 56908 32227 56948 32236
rect 57196 32192 57236 32201
rect 57099 31772 57141 31781
rect 57099 31732 57100 31772
rect 57140 31732 57141 31772
rect 57099 31723 57141 31732
rect 56811 31352 56853 31361
rect 56811 31312 56812 31352
rect 56852 31312 56853 31352
rect 56811 31303 56853 31312
rect 57100 31352 57140 31723
rect 57196 31604 57236 32152
rect 57292 32117 57332 32202
rect 57291 32108 57333 32117
rect 57291 32068 57292 32108
rect 57332 32068 57333 32108
rect 57291 32059 57333 32068
rect 57388 32024 57428 32320
rect 57676 32201 57716 32731
rect 57580 32192 57620 32201
rect 57675 32192 57717 32201
rect 57620 32152 57676 32192
rect 57716 32152 57717 32192
rect 57580 32143 57620 32152
rect 57675 32143 57717 32152
rect 57483 32108 57525 32117
rect 57483 32068 57484 32108
rect 57524 32068 57525 32108
rect 57483 32059 57525 32068
rect 57388 31975 57428 31984
rect 57484 31974 57524 32059
rect 57676 32058 57716 32143
rect 57867 32024 57909 32033
rect 57867 31984 57868 32024
rect 57908 31984 57909 32024
rect 57867 31975 57909 31984
rect 57771 31940 57813 31949
rect 57771 31900 57772 31940
rect 57812 31900 57813 31940
rect 57771 31891 57813 31900
rect 57772 31806 57812 31891
rect 57196 31555 57236 31564
rect 57868 31604 57908 31975
rect 57868 31555 57908 31564
rect 57484 31361 57524 31446
rect 57100 31303 57140 31312
rect 57483 31352 57525 31361
rect 57483 31312 57484 31352
rect 57524 31312 57525 31352
rect 57483 31303 57525 31312
rect 57580 31352 57620 31361
rect 57675 31352 57717 31361
rect 57620 31312 57676 31352
rect 57716 31312 57717 31352
rect 57580 31303 57620 31312
rect 57675 31303 57717 31312
rect 56523 30344 56565 30353
rect 56523 30304 56524 30344
rect 56564 30304 56565 30344
rect 56523 30295 56565 30304
rect 56236 29672 56276 29681
rect 56139 29588 56181 29597
rect 56139 29548 56140 29588
rect 56180 29548 56181 29588
rect 56139 29539 56181 29548
rect 55659 29336 55701 29345
rect 55659 29296 55660 29336
rect 55700 29296 55701 29336
rect 55659 29287 55701 29296
rect 56139 29336 56181 29345
rect 56139 29296 56140 29336
rect 56180 29296 56181 29336
rect 56139 29287 56181 29296
rect 56044 28916 56084 28925
rect 56044 28757 56084 28876
rect 56043 28748 56085 28757
rect 56043 28708 56044 28748
rect 56084 28708 56085 28748
rect 56043 28699 56085 28708
rect 56140 28328 56180 29287
rect 56236 29000 56276 29632
rect 56332 29168 56372 29800
rect 56620 29756 56660 29765
rect 56428 29168 56468 29177
rect 56332 29128 56428 29168
rect 56428 29119 56468 29128
rect 56524 29084 56564 29093
rect 56524 29000 56564 29044
rect 56236 28960 56564 29000
rect 56620 29000 56660 29716
rect 56812 29513 56852 31303
rect 57772 31226 57812 31235
rect 57196 31184 57236 31193
rect 57388 31184 57428 31189
rect 57236 31180 57428 31184
rect 57236 31144 57388 31180
rect 57196 31135 57236 31144
rect 57388 31131 57428 31140
rect 57483 31184 57525 31193
rect 57772 31184 57812 31186
rect 57483 31144 57484 31184
rect 57524 31144 57525 31184
rect 57483 31135 57525 31144
rect 57580 31144 57812 31184
rect 57964 31184 58004 33100
rect 58827 32864 58869 32873
rect 58827 32824 58828 32864
rect 58868 32824 58869 32864
rect 58827 32815 58869 32824
rect 58155 32528 58197 32537
rect 58155 32488 58156 32528
rect 58196 32488 58197 32528
rect 58155 32479 58197 32488
rect 58060 31361 58100 31446
rect 58059 31352 58101 31361
rect 58059 31312 58060 31352
rect 58100 31312 58101 31352
rect 58059 31303 58101 31312
rect 58156 31352 58196 32479
rect 58539 32192 58581 32201
rect 58539 32152 58540 32192
rect 58580 32152 58581 32192
rect 58539 32143 58581 32152
rect 58443 31688 58485 31697
rect 58443 31648 58444 31688
rect 58484 31648 58485 31688
rect 58443 31639 58485 31648
rect 58347 31436 58389 31445
rect 58347 31396 58348 31436
rect 58388 31396 58389 31436
rect 58347 31387 58389 31396
rect 58156 31303 58196 31312
rect 58251 31352 58293 31361
rect 58251 31312 58252 31352
rect 58292 31312 58293 31352
rect 58251 31303 58293 31312
rect 58348 31352 58388 31387
rect 58252 31218 58292 31303
rect 58348 31301 58388 31312
rect 57964 31144 58100 31184
rect 57388 30680 57428 30689
rect 57003 30344 57045 30353
rect 57003 30304 57004 30344
rect 57044 30304 57045 30344
rect 57003 30295 57045 30304
rect 57004 29840 57044 30295
rect 57388 30260 57428 30640
rect 57484 30680 57524 31135
rect 57484 30631 57524 30640
rect 57580 30680 57620 31144
rect 57676 30848 57716 30857
rect 57716 30808 57908 30848
rect 57676 30799 57716 30808
rect 57868 30764 57908 30808
rect 57868 30715 57908 30724
rect 57580 30631 57620 30640
rect 57771 30680 57813 30689
rect 57771 30640 57772 30680
rect 57812 30640 57813 30680
rect 57771 30631 57813 30640
rect 57388 30220 57620 30260
rect 57580 30101 57620 30220
rect 57579 30092 57621 30101
rect 57579 30052 57580 30092
rect 57620 30052 57621 30092
rect 57579 30043 57621 30052
rect 57004 29791 57044 29800
rect 56811 29504 56853 29513
rect 56811 29464 56812 29504
rect 56852 29464 56853 29504
rect 56811 29455 56853 29464
rect 57387 29504 57429 29513
rect 57387 29464 57388 29504
rect 57428 29464 57429 29504
rect 57387 29455 57429 29464
rect 56811 29336 56853 29345
rect 56811 29296 56812 29336
rect 56852 29296 56853 29336
rect 56811 29287 56853 29296
rect 56812 29168 56852 29287
rect 56812 29119 56852 29128
rect 57292 29168 57332 29177
rect 56620 28951 56660 28960
rect 56716 29084 56756 29093
rect 56716 29000 56756 29044
rect 57004 29000 57044 29009
rect 56716 28960 57004 29000
rect 56716 28748 56756 28960
rect 57004 28951 57044 28960
rect 56332 28708 56756 28748
rect 56140 28279 56180 28288
rect 56236 28328 56276 28337
rect 55755 28076 55797 28085
rect 55755 28036 55756 28076
rect 55796 28036 55797 28076
rect 55755 28027 55797 28036
rect 55564 27404 55604 27413
rect 55564 27245 55604 27364
rect 55563 27236 55605 27245
rect 55563 27196 55564 27236
rect 55604 27196 55605 27236
rect 55563 27187 55605 27196
rect 55564 26489 55604 27187
rect 55563 26480 55605 26489
rect 55563 26440 55564 26480
rect 55604 26440 55605 26480
rect 55563 26431 55605 26440
rect 55371 26396 55413 26405
rect 55371 26356 55372 26396
rect 55412 26356 55413 26396
rect 55371 26347 55413 26356
rect 54988 26093 55028 26104
rect 55083 26144 55125 26153
rect 55083 26104 55084 26144
rect 55124 26104 55125 26144
rect 55083 26095 55125 26104
rect 55084 26010 55124 26095
rect 54795 25976 54837 25985
rect 54795 25936 54796 25976
rect 54836 25936 54837 25976
rect 54795 25927 54837 25936
rect 54604 25892 54644 25901
rect 54644 25852 54740 25892
rect 54604 25843 54644 25852
rect 54507 25640 54549 25649
rect 54507 25600 54508 25640
rect 54548 25600 54549 25640
rect 54507 25591 54549 25600
rect 54603 25472 54645 25481
rect 54603 25432 54604 25472
rect 54644 25432 54645 25472
rect 54603 25423 54645 25432
rect 54508 25313 54548 25398
rect 53876 25264 54260 25304
rect 54315 25304 54357 25313
rect 54315 25264 54316 25304
rect 54356 25264 54357 25304
rect 53836 25255 53876 25264
rect 54315 25255 54357 25264
rect 54412 25304 54452 25313
rect 53740 25170 53780 25255
rect 54124 25178 54164 25187
rect 53644 25083 53684 25092
rect 54316 25170 54356 25255
rect 54028 24632 54068 24641
rect 53835 24548 53877 24557
rect 53835 24508 53836 24548
rect 53876 24508 53877 24548
rect 53835 24499 53877 24508
rect 53836 24414 53876 24499
rect 54028 24212 54068 24592
rect 53836 24172 54068 24212
rect 53067 24044 53109 24053
rect 53067 24004 53068 24044
rect 53108 24004 53109 24044
rect 53067 23995 53109 24004
rect 53068 23910 53108 23995
rect 53163 23792 53205 23801
rect 53163 23752 53164 23792
rect 53204 23752 53205 23792
rect 53163 23743 53205 23752
rect 53836 23792 53876 24172
rect 54124 24044 54164 25138
rect 54412 25052 54452 25264
rect 54507 25304 54549 25313
rect 54507 25264 54508 25304
rect 54548 25264 54549 25304
rect 54507 25255 54549 25264
rect 54604 25304 54644 25423
rect 54604 25255 54644 25264
rect 54316 25012 54452 25052
rect 54316 24137 54356 25012
rect 54412 24632 54452 24641
rect 54700 24632 54740 25852
rect 54796 25842 54836 25927
rect 54795 25304 54837 25313
rect 54795 25264 54796 25304
rect 54836 25264 54837 25304
rect 54795 25255 54837 25264
rect 54452 24592 54740 24632
rect 54412 24583 54452 24592
rect 54796 24473 54836 25255
rect 55083 24800 55125 24809
rect 55083 24760 55084 24800
rect 55124 24760 55125 24800
rect 55083 24751 55125 24760
rect 55084 24641 55124 24751
rect 55083 24632 55125 24641
rect 55083 24592 55084 24632
rect 55124 24592 55125 24632
rect 55083 24583 55125 24592
rect 55275 24632 55317 24641
rect 55275 24592 55276 24632
rect 55316 24592 55317 24632
rect 55275 24583 55317 24592
rect 55276 24498 55316 24583
rect 54795 24464 54837 24473
rect 54795 24424 54796 24464
rect 54836 24424 54837 24464
rect 54795 24415 54837 24424
rect 54315 24128 54357 24137
rect 54315 24088 54316 24128
rect 54356 24088 54357 24128
rect 54315 24079 54357 24088
rect 53836 23743 53876 23752
rect 53932 24004 54164 24044
rect 54219 24044 54261 24053
rect 54219 24004 54220 24044
rect 54260 24004 54261 24044
rect 53932 23792 53972 24004
rect 54219 23995 54261 24004
rect 54220 23801 54260 23995
rect 54796 23801 54836 24415
rect 55083 24128 55125 24137
rect 55083 24088 55084 24128
rect 55124 24088 55125 24128
rect 55083 24079 55125 24088
rect 54987 24044 55029 24053
rect 54987 24004 54988 24044
rect 55028 24004 55029 24044
rect 54987 23995 55029 24004
rect 54988 23910 55028 23995
rect 53932 23743 53972 23752
rect 54027 23792 54069 23801
rect 54027 23752 54028 23792
rect 54068 23752 54069 23792
rect 54027 23743 54069 23752
rect 54124 23792 54164 23801
rect 53164 23658 53204 23743
rect 54028 23658 54068 23743
rect 54124 23549 54164 23752
rect 54219 23792 54261 23801
rect 54219 23752 54220 23792
rect 54260 23752 54261 23792
rect 54219 23743 54261 23752
rect 54795 23792 54837 23801
rect 54795 23752 54796 23792
rect 54836 23752 54837 23792
rect 54795 23743 54837 23752
rect 55084 23792 55124 24079
rect 55756 24044 55796 28027
rect 55947 27572 55989 27581
rect 55947 27532 55948 27572
rect 55988 27532 55989 27572
rect 55947 27523 55989 27532
rect 55851 26144 55893 26153
rect 55851 26104 55852 26144
rect 55892 26104 55893 26144
rect 55948 26144 55988 27523
rect 56236 27413 56276 28288
rect 56332 28328 56372 28708
rect 57292 28412 57332 29128
rect 57388 29168 57428 29455
rect 57484 29345 57524 29431
rect 57483 29340 57525 29345
rect 57483 29296 57484 29340
rect 57524 29296 57525 29340
rect 57483 29287 57525 29296
rect 57388 29119 57428 29128
rect 57292 28372 57524 28412
rect 56332 28279 56372 28288
rect 57004 28328 57044 28337
rect 56428 28244 56468 28253
rect 56620 28244 56660 28253
rect 56468 28204 56620 28244
rect 56428 28195 56468 28204
rect 56620 28195 56660 28204
rect 56235 27404 56277 27413
rect 56235 27364 56236 27404
rect 56276 27364 56277 27404
rect 56235 27355 56277 27364
rect 57004 26825 57044 28288
rect 57484 27824 57524 28372
rect 57484 27775 57524 27784
rect 57580 27656 57620 30043
rect 57772 29840 57812 30631
rect 57868 29840 57908 29849
rect 57772 29800 57868 29840
rect 57868 29791 57908 29800
rect 57963 29588 58005 29597
rect 57963 29548 57964 29588
rect 58004 29548 58005 29588
rect 57963 29539 58005 29548
rect 57867 28328 57909 28337
rect 57867 28288 57868 28328
rect 57908 28288 57909 28328
rect 57867 28279 57909 28288
rect 57868 28194 57908 28279
rect 57675 27740 57717 27749
rect 57675 27700 57676 27740
rect 57716 27700 57717 27740
rect 57675 27691 57717 27700
rect 57580 27607 57620 27616
rect 57676 27656 57716 27691
rect 57676 27605 57716 27616
rect 57772 27656 57812 27665
rect 56043 26816 56085 26825
rect 56043 26776 56044 26816
rect 56084 26776 56085 26816
rect 56043 26767 56085 26776
rect 57003 26816 57045 26825
rect 57003 26776 57004 26816
rect 57044 26776 57140 26816
rect 57003 26767 57045 26776
rect 56044 26682 56084 26767
rect 56428 26732 56468 26741
rect 56428 26228 56468 26692
rect 56523 26396 56565 26405
rect 56523 26356 56524 26396
rect 56564 26356 56565 26396
rect 56523 26347 56565 26356
rect 56332 26188 56468 26228
rect 56140 26144 56180 26153
rect 55948 26104 56084 26144
rect 55851 26095 55893 26104
rect 55852 26010 55892 26095
rect 55947 25976 55989 25985
rect 55947 25936 55948 25976
rect 55988 25936 55989 25976
rect 55947 25927 55989 25936
rect 55948 25842 55988 25927
rect 55948 24044 55988 24053
rect 55756 24004 55948 24044
rect 55948 23995 55988 24004
rect 55659 23960 55701 23969
rect 55659 23920 55660 23960
rect 55700 23920 55701 23960
rect 55659 23911 55701 23920
rect 55084 23743 55124 23752
rect 55660 23792 55700 23911
rect 55563 23708 55605 23717
rect 55563 23668 55564 23708
rect 55604 23668 55605 23708
rect 55563 23659 55605 23668
rect 55564 23574 55604 23659
rect 54123 23540 54165 23549
rect 54123 23500 54124 23540
rect 54164 23500 54165 23540
rect 54123 23491 54165 23500
rect 54027 23372 54069 23381
rect 54027 23332 54028 23372
rect 54068 23332 54069 23372
rect 54027 23323 54069 23332
rect 54028 23060 54068 23323
rect 55660 23129 55700 23752
rect 56044 23792 56084 26104
rect 56140 25985 56180 26104
rect 56235 26060 56277 26069
rect 56235 26020 56236 26060
rect 56276 26020 56277 26060
rect 56235 26011 56277 26020
rect 56139 25976 56181 25985
rect 56139 25936 56140 25976
rect 56180 25936 56181 25976
rect 56139 25927 56181 25936
rect 56236 25926 56276 26011
rect 56332 25976 56372 26188
rect 56524 26144 56564 26347
rect 56524 26095 56564 26104
rect 56332 25927 56372 25936
rect 56428 26060 56468 26069
rect 56428 25565 56468 26020
rect 57003 26060 57045 26069
rect 57003 26020 57004 26060
rect 57044 26020 57045 26060
rect 57003 26011 57045 26020
rect 56523 25976 56565 25985
rect 56523 25936 56524 25976
rect 56564 25936 56565 25976
rect 56523 25927 56565 25936
rect 56427 25556 56469 25565
rect 56427 25516 56428 25556
rect 56468 25516 56469 25556
rect 56427 25507 56469 25516
rect 56524 25132 56564 25927
rect 56716 25892 56756 25901
rect 56619 25640 56661 25649
rect 56619 25600 56620 25640
rect 56660 25600 56661 25640
rect 56619 25591 56661 25600
rect 56620 25304 56660 25591
rect 56716 25481 56756 25852
rect 57004 25556 57044 26011
rect 56908 25516 57004 25556
rect 56715 25472 56757 25481
rect 56715 25432 56716 25472
rect 56756 25432 56757 25472
rect 56715 25423 56757 25432
rect 56620 25255 56660 25264
rect 56716 25304 56756 25313
rect 56756 25264 56852 25304
rect 56716 25255 56756 25264
rect 56524 25083 56564 25092
rect 56715 24968 56757 24977
rect 56715 24928 56716 24968
rect 56756 24928 56757 24968
rect 56715 24919 56757 24928
rect 56620 24632 56660 24641
rect 56428 24548 56468 24557
rect 56468 24508 56564 24548
rect 56428 24499 56468 24508
rect 56427 24212 56469 24221
rect 56427 24172 56428 24212
rect 56468 24172 56469 24212
rect 56427 24163 56469 24172
rect 56428 24044 56468 24163
rect 56524 24137 56564 24508
rect 56523 24128 56565 24137
rect 56523 24088 56524 24128
rect 56564 24088 56565 24128
rect 56523 24079 56565 24088
rect 56428 23995 56468 24004
rect 55948 23624 55988 23633
rect 55659 23120 55701 23129
rect 55659 23080 55660 23120
rect 55700 23080 55701 23120
rect 55659 23071 55701 23080
rect 53067 23036 53109 23045
rect 53067 22996 53068 23036
rect 53108 22996 53109 23036
rect 53067 22987 53109 22996
rect 53548 23020 53695 23060
rect 53068 21617 53108 22987
rect 53259 22952 53301 22961
rect 53548 22952 53588 23020
rect 53259 22912 53260 22952
rect 53300 22912 53588 22952
rect 53259 22903 53301 22912
rect 53544 22784 53586 22793
rect 53544 22744 53545 22784
rect 53585 22744 53586 22784
rect 53544 22735 53586 22744
rect 53545 22596 53585 22735
rect 53655 22596 53695 23020
rect 53944 23036 53986 23045
rect 53944 22996 53945 23036
rect 53985 22996 53986 23036
rect 54028 23020 54095 23060
rect 55948 23045 55988 23584
rect 53944 22987 53986 22996
rect 53945 22596 53985 22987
rect 54055 22596 54095 23020
rect 55254 23036 55296 23045
rect 55254 22996 55255 23036
rect 55295 22996 55296 23036
rect 55254 22987 55296 22996
rect 55947 23036 55989 23045
rect 55947 22996 55948 23036
rect 55988 22996 55989 23036
rect 55947 22987 55989 22996
rect 54454 22952 54496 22961
rect 54454 22912 54455 22952
rect 54495 22912 54496 22952
rect 54454 22903 54496 22912
rect 54744 22952 54786 22961
rect 54744 22912 54745 22952
rect 54785 22912 54786 22952
rect 54744 22903 54786 22912
rect 55144 22952 55186 22961
rect 55144 22912 55145 22952
rect 55185 22912 55186 22952
rect 55144 22903 55186 22912
rect 54344 22868 54386 22877
rect 54344 22828 54345 22868
rect 54385 22828 54386 22868
rect 54344 22819 54386 22828
rect 54345 22596 54385 22819
rect 54455 22596 54495 22903
rect 54745 22596 54785 22903
rect 54854 22784 54896 22793
rect 54854 22744 54855 22784
rect 54895 22744 54896 22784
rect 54854 22735 54896 22744
rect 54855 22596 54895 22735
rect 55145 22596 55185 22903
rect 55255 22596 55295 22987
rect 55755 22952 55797 22961
rect 56044 22952 56084 23752
rect 56332 23792 56372 23801
rect 56139 23708 56181 23717
rect 56139 23668 56140 23708
rect 56180 23668 56181 23708
rect 56139 23659 56181 23668
rect 56140 23060 56180 23659
rect 56332 23381 56372 23752
rect 56524 23717 56564 24079
rect 56620 23792 56660 24592
rect 56620 23743 56660 23752
rect 56716 23792 56756 24919
rect 56812 24464 56852 25264
rect 56908 24977 56948 25516
rect 57004 25507 57044 25516
rect 57100 25388 57140 26776
rect 57675 26228 57717 26237
rect 57675 26188 57676 26228
rect 57716 26188 57717 26228
rect 57675 26179 57717 26188
rect 57676 25985 57716 26179
rect 57675 25976 57717 25985
rect 57675 25936 57676 25976
rect 57716 25936 57717 25976
rect 57675 25927 57717 25936
rect 57387 25892 57429 25901
rect 57387 25852 57388 25892
rect 57428 25852 57429 25892
rect 57387 25843 57429 25852
rect 57291 25640 57333 25649
rect 57291 25600 57292 25640
rect 57332 25600 57333 25640
rect 57291 25591 57333 25600
rect 57004 25348 57140 25388
rect 56907 24968 56949 24977
rect 56907 24928 56908 24968
rect 56948 24928 56949 24968
rect 56907 24919 56949 24928
rect 57004 24632 57044 25348
rect 57292 25052 57332 25591
rect 57388 25304 57428 25843
rect 57483 25556 57525 25565
rect 57483 25516 57484 25556
rect 57524 25516 57525 25556
rect 57483 25507 57525 25516
rect 57484 25422 57524 25507
rect 57484 25304 57524 25313
rect 57388 25264 57484 25304
rect 57484 25255 57524 25264
rect 57676 25304 57716 25927
rect 57772 25649 57812 27616
rect 57868 26144 57908 26153
rect 57868 25901 57908 26104
rect 57964 25985 58004 29539
rect 58060 27908 58100 31144
rect 58252 30680 58292 30689
rect 58444 30680 58484 31639
rect 58540 31352 58580 32143
rect 58635 32108 58677 32117
rect 58635 32068 58636 32108
rect 58676 32068 58677 32108
rect 58635 32059 58677 32068
rect 58636 31604 58676 32059
rect 58636 31555 58676 31564
rect 58636 31352 58676 31361
rect 58540 31312 58636 31352
rect 58636 31303 58676 31312
rect 58828 31352 58868 32815
rect 58924 32192 58964 32201
rect 58964 32152 59060 32192
rect 58924 32143 58964 32152
rect 58923 31940 58965 31949
rect 58923 31900 58924 31940
rect 58964 31900 58965 31940
rect 58923 31891 58965 31900
rect 58828 31303 58868 31312
rect 58924 31352 58964 31891
rect 58924 31303 58964 31312
rect 58292 30640 58484 30680
rect 59020 30680 59060 32152
rect 59307 32108 59349 32117
rect 59307 32068 59308 32108
rect 59348 32068 59349 32108
rect 59307 32059 59349 32068
rect 59211 31352 59253 31361
rect 59211 31312 59212 31352
rect 59252 31312 59253 31352
rect 59211 31303 59253 31312
rect 59115 31184 59157 31193
rect 59115 31144 59116 31184
rect 59156 31144 59157 31184
rect 59115 31135 59157 31144
rect 59116 31050 59156 31135
rect 59115 30680 59157 30689
rect 59020 30640 59116 30680
rect 59156 30640 59157 30680
rect 58252 30353 58292 30640
rect 59115 30631 59157 30640
rect 59116 30546 59156 30631
rect 59212 30353 59252 31303
rect 58251 30344 58293 30353
rect 58251 30304 58252 30344
rect 58292 30304 58293 30344
rect 58251 30295 58293 30304
rect 59211 30344 59253 30353
rect 59211 30304 59212 30344
rect 59252 30304 59253 30344
rect 59211 30295 59253 30304
rect 59212 30092 59252 30101
rect 59308 30092 59348 32059
rect 59252 30052 59348 30092
rect 59403 30092 59445 30101
rect 59403 30052 59404 30092
rect 59444 30052 59445 30092
rect 59212 30043 59252 30052
rect 59403 30043 59445 30052
rect 59595 30092 59637 30101
rect 59595 30052 59596 30092
rect 59636 30052 59637 30092
rect 59595 30043 59637 30052
rect 59404 29924 59444 30043
rect 59596 29958 59636 30043
rect 59404 29875 59444 29884
rect 59020 29672 59060 29681
rect 59212 29672 59252 29681
rect 58828 29632 59020 29672
rect 58155 29336 58197 29345
rect 58155 29296 58156 29336
rect 58196 29296 58197 29336
rect 58155 29287 58197 29296
rect 58156 29202 58196 29287
rect 58828 29177 58868 29632
rect 59020 29623 59060 29632
rect 59116 29632 59212 29672
rect 58923 29504 58965 29513
rect 58923 29464 58924 29504
rect 58964 29464 58965 29504
rect 58923 29455 58965 29464
rect 58251 29168 58293 29177
rect 58251 29128 58252 29168
rect 58292 29128 58293 29168
rect 58251 29119 58293 29128
rect 58827 29168 58869 29177
rect 58827 29128 58828 29168
rect 58868 29128 58869 29168
rect 58827 29119 58869 29128
rect 58924 29168 58964 29455
rect 59116 29168 59156 29632
rect 59212 29623 59252 29632
rect 59692 29513 59732 34159
rect 59883 34124 59925 34133
rect 59883 34084 59884 34124
rect 59924 34084 59925 34124
rect 59883 34075 59925 34084
rect 59884 33713 59924 34075
rect 59980 33872 60020 34159
rect 59980 33823 60020 33832
rect 59883 33704 59925 33713
rect 59883 33664 59884 33704
rect 59924 33664 59925 33704
rect 59883 33655 59925 33664
rect 59884 33570 59924 33655
rect 59980 33452 60020 33461
rect 59788 32192 59828 32201
rect 59788 31781 59828 32152
rect 59980 31781 60020 33412
rect 60171 32696 60213 32705
rect 60171 32656 60172 32696
rect 60212 32656 60213 32696
rect 60171 32647 60213 32656
rect 60172 32562 60212 32647
rect 60171 32192 60213 32201
rect 60171 32152 60172 32192
rect 60212 32152 60213 32192
rect 60171 32143 60213 32152
rect 60172 32058 60212 32143
rect 59787 31772 59829 31781
rect 59787 31732 59788 31772
rect 59828 31732 59829 31772
rect 59787 31723 59829 31732
rect 59979 31772 60021 31781
rect 59979 31732 59980 31772
rect 60020 31732 60021 31772
rect 59979 31723 60021 31732
rect 60268 30596 60308 35008
rect 60459 34040 60501 34049
rect 60459 34000 60460 34040
rect 60500 34000 60501 34040
rect 60459 33991 60501 34000
rect 60460 32369 60500 33991
rect 60651 33956 60693 33965
rect 60651 33916 60652 33956
rect 60692 33916 60693 33956
rect 60651 33907 60693 33916
rect 60459 32360 60501 32369
rect 60459 32320 60460 32360
rect 60500 32320 60501 32360
rect 60459 32311 60501 32320
rect 60364 32192 60404 32201
rect 60364 31949 60404 32152
rect 60363 31940 60405 31949
rect 60363 31900 60364 31940
rect 60404 31900 60405 31940
rect 60363 31891 60405 31900
rect 60460 31940 60500 31951
rect 60460 31865 60500 31900
rect 60459 31856 60501 31865
rect 60459 31816 60460 31856
rect 60500 31816 60501 31856
rect 60459 31807 60501 31816
rect 60555 31688 60597 31697
rect 60555 31648 60556 31688
rect 60596 31648 60597 31688
rect 60555 31639 60597 31648
rect 60556 30689 60596 31639
rect 60555 30680 60597 30689
rect 60555 30640 60556 30680
rect 60596 30640 60597 30680
rect 60555 30631 60597 30640
rect 60172 30556 60308 30596
rect 60172 30017 60212 30556
rect 60268 30428 60308 30439
rect 60268 30353 60308 30388
rect 60267 30344 60309 30353
rect 60267 30304 60268 30344
rect 60308 30304 60309 30344
rect 60267 30295 60309 30304
rect 60171 30008 60213 30017
rect 60171 29968 60172 30008
rect 60212 29968 60213 30008
rect 60171 29959 60213 29968
rect 59788 29924 59828 29933
rect 59691 29504 59733 29513
rect 59691 29464 59692 29504
rect 59732 29464 59733 29504
rect 59691 29455 59733 29464
rect 59788 29429 59828 29884
rect 59787 29420 59829 29429
rect 59787 29380 59788 29420
rect 59828 29380 59829 29420
rect 59787 29371 59829 29380
rect 60075 29420 60117 29429
rect 60075 29380 60076 29420
rect 60116 29380 60117 29420
rect 60075 29371 60117 29380
rect 59692 29177 59732 29262
rect 58924 29119 58964 29128
rect 59020 29128 59116 29168
rect 58252 29034 58292 29119
rect 58828 29034 58868 29119
rect 58923 28496 58965 28505
rect 58923 28456 58924 28496
rect 58964 28456 58965 28496
rect 58923 28447 58965 28456
rect 58827 27908 58869 27917
rect 58060 27868 58292 27908
rect 58059 27740 58101 27749
rect 58059 27700 58060 27740
rect 58100 27700 58101 27740
rect 58059 27691 58101 27700
rect 58060 27656 58100 27691
rect 58060 27605 58100 27616
rect 58155 27404 58197 27413
rect 58155 27364 58156 27404
rect 58196 27364 58197 27404
rect 58155 27355 58197 27364
rect 58156 27270 58196 27355
rect 57963 25976 58005 25985
rect 57963 25936 57964 25976
rect 58004 25936 58005 25976
rect 57963 25927 58005 25936
rect 57867 25892 57909 25901
rect 57867 25852 57868 25892
rect 57908 25852 57909 25892
rect 57867 25843 57909 25852
rect 57771 25640 57813 25649
rect 57771 25600 57772 25640
rect 57812 25600 57813 25640
rect 57771 25591 57813 25600
rect 57771 25472 57813 25481
rect 57771 25432 57772 25472
rect 57812 25432 57813 25472
rect 57771 25423 57813 25432
rect 57676 25255 57716 25264
rect 57772 25304 57812 25423
rect 57772 25255 57812 25264
rect 57292 25012 57428 25052
rect 57004 24583 57044 24592
rect 56812 24424 57140 24464
rect 56811 23960 56853 23969
rect 56811 23920 56812 23960
rect 56852 23920 56853 23960
rect 56811 23911 56853 23920
rect 56716 23743 56756 23752
rect 56812 23792 56852 23911
rect 56812 23743 56852 23752
rect 56907 23792 56949 23801
rect 56907 23752 56908 23792
rect 56948 23752 56949 23792
rect 56907 23743 56949 23752
rect 57100 23792 57140 24424
rect 57100 23743 57140 23752
rect 57196 23792 57236 23801
rect 56523 23708 56565 23717
rect 56523 23668 56524 23708
rect 56564 23668 56565 23708
rect 56523 23659 56565 23668
rect 56908 23658 56948 23743
rect 57196 23549 57236 23752
rect 57291 23792 57333 23801
rect 57291 23752 57292 23792
rect 57332 23752 57333 23792
rect 57291 23743 57333 23752
rect 57388 23792 57428 25012
rect 57483 24716 57525 24725
rect 57483 24676 57484 24716
rect 57524 24676 57525 24716
rect 57483 24667 57525 24676
rect 57388 23743 57428 23752
rect 57292 23658 57332 23743
rect 57195 23540 57237 23549
rect 57195 23500 57196 23540
rect 57236 23500 57237 23540
rect 57195 23491 57237 23500
rect 56331 23372 56373 23381
rect 56331 23332 56332 23372
rect 56372 23332 56373 23372
rect 56331 23323 56373 23332
rect 57099 23288 57141 23297
rect 57099 23248 57100 23288
rect 57140 23248 57141 23288
rect 57099 23239 57141 23248
rect 57100 23060 57140 23239
rect 57484 23060 57524 24667
rect 57868 24641 57908 25843
rect 58059 24884 58101 24893
rect 58059 24844 58060 24884
rect 58100 24844 58101 24884
rect 58059 24835 58101 24844
rect 57867 24632 57909 24641
rect 57867 24592 57868 24632
rect 57908 24592 57909 24632
rect 57867 24583 57909 24592
rect 57868 24498 57908 24583
rect 57867 24212 57909 24221
rect 57867 24172 57868 24212
rect 57908 24172 57909 24212
rect 57867 24163 57909 24172
rect 57771 23960 57813 23969
rect 57771 23920 57772 23960
rect 57812 23920 57813 23960
rect 57771 23911 57813 23920
rect 57772 23826 57812 23911
rect 57868 23801 57908 24163
rect 57867 23792 57909 23801
rect 57867 23752 57868 23792
rect 57908 23752 57909 23792
rect 57867 23743 57909 23752
rect 57868 23658 57908 23743
rect 58060 23060 58100 24835
rect 58252 24473 58292 27868
rect 58827 27868 58828 27908
rect 58868 27868 58869 27908
rect 58827 27859 58869 27868
rect 58539 27656 58581 27665
rect 58539 27616 58540 27656
rect 58580 27616 58581 27656
rect 58539 27607 58581 27616
rect 58443 26900 58485 26909
rect 58443 26860 58444 26900
rect 58484 26860 58485 26900
rect 58443 26851 58485 26860
rect 58444 26766 58484 26851
rect 58540 26312 58580 27607
rect 58828 27572 58868 27859
rect 58828 27523 58868 27532
rect 58731 27320 58773 27329
rect 58731 27280 58732 27320
rect 58772 27280 58773 27320
rect 58731 27271 58773 27280
rect 58636 26648 58676 26657
rect 58636 26489 58676 26608
rect 58635 26480 58677 26489
rect 58635 26440 58636 26480
rect 58676 26440 58677 26480
rect 58635 26431 58677 26440
rect 58540 26272 58676 26312
rect 58347 26144 58389 26153
rect 58347 26104 58348 26144
rect 58388 26104 58389 26144
rect 58347 26095 58389 26104
rect 58251 24464 58293 24473
rect 58251 24424 58252 24464
rect 58292 24424 58293 24464
rect 58251 24415 58293 24424
rect 58251 23876 58293 23885
rect 58251 23836 58252 23876
rect 58292 23836 58293 23876
rect 58251 23827 58293 23836
rect 58252 23297 58292 23827
rect 58251 23288 58293 23297
rect 58251 23248 58252 23288
rect 58292 23248 58293 23288
rect 58251 23239 58293 23248
rect 56140 23020 56385 23060
rect 55755 22912 55756 22952
rect 55796 22912 55892 22952
rect 56044 22912 56180 22952
rect 55755 22903 55797 22912
rect 55654 22868 55696 22877
rect 55654 22828 55655 22868
rect 55695 22828 55696 22868
rect 55852 22868 55892 22912
rect 55852 22828 56095 22868
rect 55654 22819 55696 22828
rect 55544 22784 55586 22793
rect 55544 22744 55545 22784
rect 55585 22744 55586 22784
rect 55544 22735 55586 22744
rect 55545 22596 55585 22735
rect 55655 22596 55695 22819
rect 55755 22784 55797 22793
rect 55755 22744 55756 22784
rect 55796 22744 55985 22784
rect 55755 22735 55797 22744
rect 55945 22596 55985 22744
rect 56055 22596 56095 22828
rect 56140 22793 56180 22912
rect 56139 22784 56181 22793
rect 56139 22744 56140 22784
rect 56180 22744 56181 22784
rect 56139 22735 56181 22744
rect 56345 22596 56385 23020
rect 56454 23036 56496 23045
rect 56454 22996 56455 23036
rect 56495 22996 56496 23036
rect 57100 23020 57185 23060
rect 56454 22987 56496 22996
rect 56455 22596 56495 22987
rect 56744 22952 56786 22961
rect 56744 22912 56745 22952
rect 56785 22912 56786 22952
rect 56744 22903 56786 22912
rect 56745 22596 56785 22903
rect 56854 22784 56896 22793
rect 56854 22744 56855 22784
rect 56895 22744 56896 22784
rect 56854 22735 56896 22744
rect 56855 22596 56895 22735
rect 57145 22596 57185 23020
rect 57255 23020 57524 23060
rect 58055 23020 58100 23060
rect 58348 23060 58388 26095
rect 58443 25472 58485 25481
rect 58443 25432 58444 25472
rect 58484 25432 58485 25472
rect 58443 25423 58485 25432
rect 58444 25304 58484 25423
rect 58444 25255 58484 25264
rect 58539 25136 58581 25145
rect 58539 25096 58540 25136
rect 58580 25096 58581 25136
rect 58539 25087 58581 25096
rect 58540 25002 58580 25087
rect 58636 23060 58676 26272
rect 58732 26144 58772 27271
rect 58828 26648 58868 26657
rect 58828 26153 58868 26608
rect 58732 26095 58772 26104
rect 58827 26144 58869 26153
rect 58827 26104 58828 26144
rect 58868 26104 58869 26144
rect 58827 26095 58869 26104
rect 58924 25976 58964 28447
rect 59020 28337 59060 29128
rect 59116 29119 59156 29128
rect 59308 29168 59348 29177
rect 59308 29000 59348 29128
rect 59691 29168 59733 29177
rect 59691 29128 59692 29168
rect 59732 29128 59733 29168
rect 59691 29119 59733 29128
rect 59308 28960 60020 29000
rect 59116 28916 59156 28925
rect 59156 28876 59924 28916
rect 59116 28867 59156 28876
rect 59115 28748 59157 28757
rect 59115 28708 59116 28748
rect 59156 28708 59157 28748
rect 59115 28699 59157 28708
rect 59403 28748 59445 28757
rect 59403 28708 59404 28748
rect 59444 28708 59445 28748
rect 59403 28699 59445 28708
rect 59019 28328 59061 28337
rect 59019 28288 59020 28328
rect 59060 28288 59061 28328
rect 59019 28279 59061 28288
rect 59020 28160 59060 28169
rect 59020 27749 59060 28120
rect 59019 27740 59061 27749
rect 59019 27700 59020 27740
rect 59060 27700 59061 27740
rect 59019 27691 59061 27700
rect 59020 27404 59060 27413
rect 59020 26909 59060 27364
rect 59116 27077 59156 28699
rect 59307 27992 59349 28001
rect 59307 27952 59308 27992
rect 59348 27952 59349 27992
rect 59307 27943 59349 27952
rect 59212 27572 59252 27581
rect 59115 27068 59157 27077
rect 59115 27028 59116 27068
rect 59156 27028 59157 27068
rect 59115 27019 59157 27028
rect 59019 26900 59061 26909
rect 59019 26860 59020 26900
rect 59060 26860 59061 26900
rect 59019 26851 59061 26860
rect 59212 26573 59252 27532
rect 59211 26564 59253 26573
rect 59211 26524 59212 26564
rect 59252 26524 59253 26564
rect 59211 26515 59253 26524
rect 59308 26396 59348 27943
rect 59404 27824 59444 28699
rect 59884 28412 59924 28876
rect 59980 28496 60020 28960
rect 60076 28841 60116 29371
rect 60556 29168 60596 30631
rect 60652 29882 60692 33907
rect 60844 33545 60884 35839
rect 60940 35141 60980 36427
rect 61036 35981 61076 36688
rect 61132 36728 61172 36737
rect 61035 35972 61077 35981
rect 61035 35932 61036 35972
rect 61076 35932 61077 35972
rect 61035 35923 61077 35932
rect 61132 35897 61172 36688
rect 61227 36728 61269 36737
rect 61227 36688 61228 36728
rect 61268 36688 61269 36728
rect 61227 36679 61269 36688
rect 61131 35888 61173 35897
rect 61131 35848 61132 35888
rect 61172 35848 61173 35888
rect 61131 35839 61173 35848
rect 61228 35888 61268 36679
rect 61324 36485 61364 38200
rect 61323 36476 61365 36485
rect 61323 36436 61324 36476
rect 61364 36436 61365 36476
rect 61323 36427 61365 36436
rect 61420 36065 61460 38200
rect 61516 38240 61556 38249
rect 61516 36476 61556 38200
rect 64684 38240 64724 38251
rect 65260 38240 65300 38249
rect 64684 38165 64724 38200
rect 65164 38200 65260 38240
rect 63819 38156 63861 38165
rect 63819 38116 63820 38156
rect 63860 38116 63861 38156
rect 63819 38107 63861 38116
rect 64683 38156 64725 38165
rect 64683 38116 64684 38156
rect 64724 38116 64725 38156
rect 64683 38107 64725 38116
rect 64876 38156 64916 38165
rect 62283 38072 62325 38081
rect 62283 38032 62284 38072
rect 62324 38032 62325 38072
rect 62283 38023 62325 38032
rect 61804 37400 61844 37409
rect 62187 37400 62229 37409
rect 61844 37360 61940 37400
rect 61804 37351 61844 37360
rect 61708 36476 61748 36485
rect 61516 36436 61708 36476
rect 61708 36317 61748 36436
rect 61707 36308 61749 36317
rect 61707 36268 61708 36308
rect 61748 36268 61749 36308
rect 61707 36259 61749 36268
rect 61419 36056 61461 36065
rect 61419 36016 61420 36056
rect 61460 36016 61461 36056
rect 61419 36007 61461 36016
rect 61803 35972 61845 35981
rect 61803 35932 61804 35972
rect 61844 35932 61845 35972
rect 61803 35923 61845 35932
rect 61228 35839 61268 35848
rect 61323 35888 61365 35897
rect 61323 35848 61324 35888
rect 61364 35848 61365 35888
rect 61323 35839 61365 35848
rect 61420 35888 61460 35897
rect 61036 35729 61076 35814
rect 61324 35754 61364 35839
rect 61035 35720 61077 35729
rect 61035 35680 61036 35720
rect 61076 35680 61077 35720
rect 61035 35671 61077 35680
rect 61227 35552 61269 35561
rect 61227 35512 61228 35552
rect 61268 35512 61269 35552
rect 61227 35503 61269 35512
rect 61132 35216 61172 35225
rect 60939 35132 60981 35141
rect 60939 35092 60940 35132
rect 60980 35092 60981 35132
rect 60939 35083 60981 35092
rect 61035 35048 61077 35057
rect 61132 35048 61172 35176
rect 61035 35008 61036 35048
rect 61076 35008 61172 35048
rect 61228 35216 61268 35503
rect 61420 35477 61460 35848
rect 61516 35888 61556 35897
rect 61516 35813 61556 35848
rect 61708 35877 61748 35886
rect 61515 35804 61557 35813
rect 61708 35804 61748 35837
rect 61515 35764 61516 35804
rect 61556 35764 61557 35804
rect 61515 35755 61557 35764
rect 61612 35764 61748 35804
rect 61419 35468 61461 35477
rect 61419 35428 61420 35468
rect 61460 35428 61461 35468
rect 61419 35419 61461 35428
rect 61035 34999 61077 35008
rect 61228 34964 61268 35176
rect 61420 35216 61460 35227
rect 61420 35141 61460 35176
rect 61419 35132 61461 35141
rect 61419 35092 61420 35132
rect 61460 35092 61461 35132
rect 61419 35083 61461 35092
rect 61132 34924 61268 34964
rect 61419 34964 61461 34973
rect 61419 34924 61420 34964
rect 61460 34924 61461 34964
rect 61132 33881 61172 34924
rect 61419 34915 61461 34924
rect 61420 34830 61460 34915
rect 61419 34712 61461 34721
rect 61419 34672 61420 34712
rect 61460 34672 61461 34712
rect 61419 34663 61461 34672
rect 61323 34208 61365 34217
rect 61323 34168 61324 34208
rect 61364 34168 61365 34208
rect 61323 34159 61365 34168
rect 61324 34074 61364 34159
rect 61131 33872 61173 33881
rect 61131 33832 61132 33872
rect 61172 33832 61173 33872
rect 61131 33823 61173 33832
rect 61323 33788 61365 33797
rect 61323 33748 61324 33788
rect 61364 33748 61365 33788
rect 61323 33739 61365 33748
rect 60843 33536 60885 33545
rect 60843 33496 60844 33536
rect 60884 33496 60885 33536
rect 60843 33487 60885 33496
rect 61324 33209 61364 33739
rect 61420 33452 61460 34663
rect 61516 33797 61556 35755
rect 61612 35477 61652 35764
rect 61804 35720 61844 35923
rect 61611 35468 61653 35477
rect 61611 35428 61612 35468
rect 61652 35428 61653 35468
rect 61611 35419 61653 35428
rect 61612 35216 61652 35227
rect 61612 35141 61652 35176
rect 61611 35132 61653 35141
rect 61611 35092 61612 35132
rect 61652 35092 61653 35132
rect 61611 35083 61653 35092
rect 61804 34721 61844 35680
rect 61900 35225 61940 37360
rect 62187 37360 62188 37400
rect 62228 37360 62229 37400
rect 62187 37351 62229 37360
rect 62188 36233 62228 37351
rect 62187 36224 62229 36233
rect 62187 36184 62188 36224
rect 62228 36184 62229 36224
rect 62187 36175 62229 36184
rect 61899 35216 61941 35225
rect 61899 35176 61900 35216
rect 61940 35176 61941 35216
rect 61899 35167 61941 35176
rect 61996 35216 62036 35225
rect 62188 35216 62228 36175
rect 62036 35176 62228 35216
rect 61996 35167 62036 35176
rect 61803 34712 61845 34721
rect 61803 34672 61804 34712
rect 61844 34672 61845 34712
rect 61803 34663 61845 34672
rect 61803 34544 61845 34553
rect 61803 34504 61804 34544
rect 61844 34504 61845 34544
rect 61803 34495 61845 34504
rect 61515 33788 61557 33797
rect 61515 33748 61516 33788
rect 61556 33748 61557 33788
rect 61515 33739 61557 33748
rect 61804 33620 61844 34495
rect 62091 34208 62133 34217
rect 62091 34168 62092 34208
rect 62132 34168 62133 34208
rect 62091 34159 62133 34168
rect 61995 33872 62037 33881
rect 61995 33832 61996 33872
rect 62036 33832 62037 33872
rect 61995 33823 62037 33832
rect 61996 33738 62036 33823
rect 61611 33536 61653 33545
rect 61611 33496 61612 33536
rect 61652 33496 61653 33536
rect 61611 33487 61653 33496
rect 61420 33412 61556 33452
rect 61516 33284 61556 33412
rect 61516 33244 61560 33284
rect 61323 33200 61365 33209
rect 61520 33200 61560 33244
rect 61323 33160 61324 33200
rect 61364 33160 61365 33200
rect 61323 33151 61365 33160
rect 61516 33160 61560 33200
rect 61324 33032 61364 33151
rect 61228 32992 61364 33032
rect 60748 32192 60788 32201
rect 60748 31865 60788 32152
rect 60939 32192 60981 32201
rect 60939 32152 60940 32192
rect 60980 32152 60981 32192
rect 60939 32143 60981 32152
rect 61132 32192 61172 32203
rect 60844 32108 60884 32117
rect 60747 31856 60789 31865
rect 60747 31816 60748 31856
rect 60788 31816 60789 31856
rect 60747 31807 60789 31816
rect 60844 31520 60884 32068
rect 60940 32024 60980 32143
rect 61036 32108 61076 32119
rect 61132 32117 61172 32152
rect 61036 32033 61076 32068
rect 61131 32108 61173 32117
rect 61131 32068 61132 32108
rect 61172 32068 61173 32108
rect 61131 32059 61173 32068
rect 60940 31975 60980 31984
rect 61035 32024 61077 32033
rect 61035 31984 61036 32024
rect 61076 31984 61077 32024
rect 61035 31975 61077 31984
rect 61035 31856 61077 31865
rect 61035 31816 61036 31856
rect 61076 31816 61077 31856
rect 61035 31807 61077 31816
rect 60748 31480 60844 31520
rect 60748 30680 60788 31480
rect 60844 31471 60884 31480
rect 61036 31184 61076 31807
rect 61131 31520 61173 31529
rect 61131 31480 61132 31520
rect 61172 31480 61173 31520
rect 61131 31471 61173 31480
rect 61132 31352 61172 31471
rect 61228 31445 61268 32992
rect 61324 32864 61364 32873
rect 61324 31697 61364 32824
rect 61516 32201 61556 33160
rect 61515 32192 61557 32201
rect 61515 32152 61516 32192
rect 61556 32152 61557 32192
rect 61515 32143 61557 32152
rect 61515 32024 61557 32033
rect 61515 31984 61516 32024
rect 61556 31984 61557 32024
rect 61515 31975 61557 31984
rect 61516 31890 61556 31975
rect 61323 31688 61365 31697
rect 61323 31648 61324 31688
rect 61364 31648 61365 31688
rect 61323 31639 61365 31648
rect 61515 31520 61557 31529
rect 61515 31480 61516 31520
rect 61556 31480 61557 31520
rect 61515 31471 61557 31480
rect 61227 31436 61269 31445
rect 61227 31396 61228 31436
rect 61268 31396 61269 31436
rect 61227 31387 61269 31396
rect 61419 31436 61461 31445
rect 61419 31396 61420 31436
rect 61460 31396 61461 31436
rect 61419 31387 61461 31396
rect 61132 31303 61172 31312
rect 61228 31352 61268 31387
rect 61228 31302 61268 31312
rect 61324 31184 61364 31189
rect 61036 31180 61364 31184
rect 61036 31144 61324 31180
rect 61324 31131 61364 31140
rect 60844 30848 60884 30857
rect 60884 30808 61364 30848
rect 60844 30799 60884 30808
rect 61324 30764 61364 30808
rect 61324 30715 61364 30724
rect 60940 30680 60980 30689
rect 60748 30640 60940 30680
rect 60940 30631 60980 30640
rect 61036 30680 61076 30689
rect 60939 30428 60981 30437
rect 60939 30388 60940 30428
rect 60980 30388 60981 30428
rect 60939 30379 60981 30388
rect 60940 30092 60980 30379
rect 60940 30043 60980 30052
rect 60747 29924 60789 29933
rect 60747 29884 60748 29924
rect 60788 29884 60789 29924
rect 60747 29882 60789 29884
rect 60652 29875 60789 29882
rect 60652 29842 60788 29875
rect 60748 29790 60788 29842
rect 60747 29672 60789 29681
rect 60747 29632 60748 29672
rect 60788 29632 60789 29672
rect 60747 29623 60789 29632
rect 60940 29672 60980 29681
rect 60556 29119 60596 29128
rect 60459 28916 60501 28925
rect 60459 28876 60460 28916
rect 60500 28876 60501 28916
rect 60459 28867 60501 28876
rect 60075 28832 60117 28841
rect 60075 28792 60076 28832
rect 60116 28792 60117 28832
rect 60075 28783 60117 28792
rect 59980 28447 60020 28456
rect 59884 28363 59924 28372
rect 60075 28412 60117 28421
rect 60075 28372 60076 28412
rect 60116 28372 60117 28412
rect 60075 28363 60117 28372
rect 59787 28328 59829 28337
rect 59787 28288 59788 28328
rect 59828 28288 59829 28328
rect 59787 28279 59829 28288
rect 59788 28194 59828 28279
rect 60076 28278 60116 28363
rect 60171 28328 60213 28337
rect 60171 28288 60172 28328
rect 60212 28288 60213 28328
rect 60171 28279 60213 28288
rect 60172 28194 60212 28279
rect 59979 28160 60021 28169
rect 59979 28120 59980 28160
rect 60020 28120 60021 28160
rect 59979 28111 60021 28120
rect 59444 27784 59636 27824
rect 59404 27775 59444 27784
rect 59596 27572 59636 27784
rect 59596 27523 59636 27532
rect 59980 27572 60020 28111
rect 59980 27523 60020 27532
rect 59788 27404 59828 27413
rect 59212 26356 59348 26396
rect 59692 27364 59788 27404
rect 59019 26312 59061 26321
rect 59019 26272 59020 26312
rect 59060 26272 59061 26312
rect 59019 26263 59061 26272
rect 58828 25936 58964 25976
rect 58731 25388 58773 25397
rect 58731 25348 58732 25388
rect 58772 25348 58773 25388
rect 58731 25339 58773 25348
rect 58732 25254 58772 25339
rect 58828 23060 58868 25936
rect 58924 25472 58964 25483
rect 58924 25397 58964 25432
rect 58923 25388 58965 25397
rect 58923 25348 58924 25388
rect 58964 25348 58965 25388
rect 58923 25339 58965 25348
rect 59020 24548 59060 26263
rect 59115 26228 59157 26237
rect 59115 26188 59116 26228
rect 59156 26188 59157 26228
rect 59115 26179 59157 26188
rect 59116 26094 59156 26179
rect 59212 25733 59252 26356
rect 59692 26237 59732 27364
rect 59788 27355 59828 27364
rect 60172 27404 60212 27413
rect 59980 26816 60020 26825
rect 59884 26776 59980 26816
rect 59499 26228 59541 26237
rect 59499 26188 59500 26228
rect 59540 26188 59541 26228
rect 59499 26179 59541 26188
rect 59691 26228 59733 26237
rect 59691 26188 59692 26228
rect 59732 26188 59733 26228
rect 59691 26179 59733 26188
rect 59308 26144 59348 26153
rect 59308 25817 59348 26104
rect 59404 26060 59444 26069
rect 59307 25808 59349 25817
rect 59307 25768 59308 25808
rect 59348 25768 59349 25808
rect 59307 25759 59349 25768
rect 59211 25724 59253 25733
rect 59211 25684 59212 25724
rect 59252 25684 59253 25724
rect 59211 25675 59253 25684
rect 58924 24508 59060 24548
rect 59116 25472 59156 25481
rect 59404 25472 59444 26020
rect 59500 25976 59540 26179
rect 59692 26144 59732 26179
rect 59692 26094 59732 26104
rect 59596 26060 59636 26071
rect 59596 25985 59636 26020
rect 59500 25927 59540 25936
rect 59595 25976 59637 25985
rect 59595 25936 59596 25976
rect 59636 25936 59637 25976
rect 59595 25927 59637 25936
rect 59884 25901 59924 26776
rect 59980 26767 60020 26776
rect 60075 26732 60117 26741
rect 60075 26692 60076 26732
rect 60116 26692 60117 26732
rect 60075 26683 60117 26692
rect 59979 26228 60021 26237
rect 59979 26188 59980 26228
rect 60020 26188 60021 26228
rect 59979 26179 60021 26188
rect 59980 26144 60020 26179
rect 60076 26144 60116 26683
rect 60172 26573 60212 27364
rect 60267 26816 60309 26825
rect 60267 26776 60268 26816
rect 60308 26776 60309 26816
rect 60267 26767 60309 26776
rect 60171 26564 60213 26573
rect 60171 26524 60172 26564
rect 60212 26524 60213 26564
rect 60171 26515 60213 26524
rect 60268 26153 60308 26767
rect 60460 26732 60500 28867
rect 60555 28328 60597 28337
rect 60555 28288 60556 28328
rect 60596 28288 60597 28328
rect 60555 28279 60597 28288
rect 60652 28328 60692 28339
rect 60556 28194 60596 28279
rect 60652 28253 60692 28288
rect 60651 28244 60693 28253
rect 60651 28204 60652 28244
rect 60692 28204 60693 28244
rect 60651 28195 60693 28204
rect 60748 27908 60788 29623
rect 60940 28505 60980 29632
rect 60939 28496 60981 28505
rect 60939 28456 60940 28496
rect 60980 28456 60981 28496
rect 61036 28496 61076 30640
rect 61132 30680 61172 30691
rect 61132 30605 61172 30640
rect 61131 30596 61173 30605
rect 61131 30556 61132 30596
rect 61172 30556 61173 30596
rect 61131 30547 61173 30556
rect 61420 30437 61460 31387
rect 61516 31352 61556 31471
rect 61612 31361 61652 33487
rect 61707 33452 61749 33461
rect 61707 33412 61708 33452
rect 61748 33412 61749 33452
rect 61707 33403 61749 33412
rect 61708 32192 61748 33403
rect 61804 33377 61844 33580
rect 61995 33452 62037 33461
rect 61995 33412 61996 33452
rect 62036 33412 62037 33452
rect 61995 33403 62037 33412
rect 61803 33368 61845 33377
rect 61803 33328 61804 33368
rect 61844 33328 61845 33368
rect 61803 33319 61845 33328
rect 61996 33318 62036 33403
rect 61803 32696 61845 32705
rect 61803 32656 61804 32696
rect 61844 32656 61845 32696
rect 61803 32647 61845 32656
rect 61708 32143 61748 32152
rect 61804 32192 61844 32647
rect 61804 32143 61844 32152
rect 62092 31613 62132 34159
rect 62188 32864 62228 35176
rect 62284 34553 62324 38023
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 62763 37400 62805 37409
rect 62763 37360 62764 37400
rect 62804 37360 62805 37400
rect 62763 37351 62805 37360
rect 62475 35132 62517 35141
rect 62475 35092 62476 35132
rect 62516 35092 62517 35132
rect 62475 35083 62517 35092
rect 62379 34964 62421 34973
rect 62379 34924 62380 34964
rect 62420 34924 62421 34964
rect 62379 34915 62421 34924
rect 62283 34544 62325 34553
rect 62283 34504 62284 34544
rect 62324 34504 62325 34544
rect 62283 34495 62325 34504
rect 62380 34460 62420 34915
rect 62476 34544 62516 35083
rect 62476 34495 62516 34504
rect 62380 34411 62420 34420
rect 62571 34460 62613 34469
rect 62571 34420 62572 34460
rect 62612 34420 62613 34460
rect 62571 34411 62613 34420
rect 62284 34376 62324 34385
rect 62284 34124 62324 34336
rect 62572 34326 62612 34411
rect 62667 34376 62709 34385
rect 62667 34336 62668 34376
rect 62708 34336 62709 34376
rect 62667 34327 62709 34336
rect 62764 34376 62804 37351
rect 62956 37232 62996 37241
rect 62860 36728 62900 36737
rect 62860 35981 62900 36688
rect 62859 35972 62901 35981
rect 62859 35932 62860 35972
rect 62900 35932 62901 35972
rect 62859 35923 62901 35932
rect 62860 35225 62900 35923
rect 62956 35477 62996 37192
rect 63724 36728 63764 36737
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 63724 36233 63764 36688
rect 63723 36224 63765 36233
rect 63723 36184 63724 36224
rect 63764 36184 63765 36224
rect 63723 36175 63765 36184
rect 63820 36056 63860 38107
rect 64204 37484 64244 37493
rect 64108 37442 64148 37451
rect 64108 37400 64148 37402
rect 63916 37360 64148 37400
rect 63916 36140 63956 37360
rect 64204 37316 64244 37444
rect 64395 37484 64437 37493
rect 64395 37444 64396 37484
rect 64436 37444 64437 37484
rect 64395 37435 64437 37444
rect 64396 37350 64436 37435
rect 64491 37400 64533 37409
rect 64491 37360 64492 37400
rect 64532 37360 64533 37400
rect 64491 37351 64533 37360
rect 63916 36091 63956 36100
rect 64012 37276 64244 37316
rect 63724 36016 63860 36056
rect 63724 35636 63764 36016
rect 64012 35897 64052 37276
rect 64300 37274 64340 37283
rect 64492 37266 64532 37351
rect 64300 37174 64340 37234
rect 64779 37232 64821 37241
rect 64779 37192 64780 37232
rect 64820 37192 64821 37232
rect 64779 37183 64821 37192
rect 64204 37134 64340 37174
rect 64108 36812 64148 36821
rect 64204 36812 64244 37134
rect 64780 37098 64820 37183
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 64148 36772 64244 36812
rect 64108 36763 64148 36772
rect 64299 36728 64341 36737
rect 64299 36688 64300 36728
rect 64340 36688 64341 36728
rect 64299 36679 64341 36688
rect 64684 36728 64724 36737
rect 64300 36594 64340 36679
rect 64684 36149 64724 36688
rect 64779 36728 64821 36737
rect 64779 36688 64780 36728
rect 64820 36688 64821 36728
rect 64779 36679 64821 36688
rect 64683 36140 64725 36149
rect 64683 36100 64684 36140
rect 64724 36100 64725 36140
rect 64683 36091 64725 36100
rect 64299 36056 64341 36065
rect 64299 36016 64300 36056
rect 64340 36016 64341 36056
rect 64299 36007 64341 36016
rect 64588 36056 64628 36065
rect 63819 35888 63861 35897
rect 63819 35848 63820 35888
rect 63860 35848 63861 35888
rect 63819 35839 63861 35848
rect 64011 35888 64053 35897
rect 64011 35848 64012 35888
rect 64052 35848 64053 35888
rect 64011 35839 64053 35848
rect 64204 35888 64244 35897
rect 63820 35754 63860 35839
rect 63916 35720 63956 35729
rect 64108 35720 64148 35725
rect 63956 35716 64148 35720
rect 63956 35680 64108 35716
rect 63916 35671 63956 35680
rect 64108 35667 64148 35676
rect 63724 35596 63860 35636
rect 62955 35468 62997 35477
rect 62955 35428 62956 35468
rect 62996 35428 62997 35468
rect 62955 35419 62997 35428
rect 62859 35216 62901 35225
rect 62859 35176 62860 35216
rect 62900 35176 62901 35216
rect 62859 35167 62901 35176
rect 62860 35082 62900 35167
rect 63531 34964 63573 34973
rect 63531 34924 63532 34964
rect 63572 34924 63573 34964
rect 63531 34915 63573 34924
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 63532 34628 63572 34915
rect 63350 34588 63572 34628
rect 63350 34395 63390 34588
rect 63627 34460 63669 34469
rect 63627 34420 63628 34460
rect 63668 34420 63669 34460
rect 63627 34411 63669 34420
rect 63052 34376 63092 34385
rect 62764 34336 63052 34376
rect 62668 34242 62708 34327
rect 62764 34124 62804 34336
rect 63052 34327 63092 34336
rect 63244 34376 63284 34385
rect 63148 34208 63188 34217
rect 62284 34084 62804 34124
rect 62956 34168 63148 34208
rect 62091 31604 62133 31613
rect 62091 31564 62092 31604
rect 62132 31564 62133 31604
rect 62091 31555 62133 31564
rect 61707 31520 61749 31529
rect 61707 31480 61708 31520
rect 61748 31480 61749 31520
rect 61707 31471 61749 31480
rect 61516 31303 61556 31312
rect 61611 31352 61653 31361
rect 61611 31312 61612 31352
rect 61652 31312 61653 31352
rect 61611 31303 61653 31312
rect 61708 31352 61748 31471
rect 61803 31436 61845 31445
rect 61803 31396 61804 31436
rect 61844 31396 61845 31436
rect 61803 31387 61845 31396
rect 61708 31303 61748 31312
rect 61804 31352 61844 31387
rect 61612 31218 61652 31303
rect 61804 31301 61844 31312
rect 61708 30680 61748 30689
rect 62188 30680 62228 32824
rect 61748 30640 62228 30680
rect 61708 30631 61748 30640
rect 61611 30596 61653 30605
rect 61611 30556 61612 30596
rect 61652 30556 61653 30596
rect 61611 30547 61653 30556
rect 61419 30428 61461 30437
rect 61419 30388 61420 30428
rect 61460 30388 61461 30428
rect 61419 30379 61461 30388
rect 61227 30260 61269 30269
rect 61227 30220 61228 30260
rect 61268 30220 61269 30260
rect 61227 30211 61269 30220
rect 61132 29924 61172 29933
rect 61132 29597 61172 29884
rect 61131 29588 61173 29597
rect 61131 29548 61132 29588
rect 61172 29548 61173 29588
rect 61131 29539 61173 29548
rect 61036 28456 61172 28496
rect 60939 28447 60981 28456
rect 60843 28328 60885 28337
rect 60843 28288 60844 28328
rect 60884 28288 60885 28328
rect 60843 28279 60885 28288
rect 60940 28328 60980 28447
rect 60940 28279 60980 28288
rect 61035 28328 61077 28337
rect 61035 28288 61036 28328
rect 61076 28288 61077 28328
rect 61035 28279 61077 28288
rect 60844 28156 60884 28279
rect 61036 28194 61076 28279
rect 60844 28107 60884 28116
rect 60556 27868 60788 27908
rect 60556 26993 60596 27868
rect 60843 27824 60885 27833
rect 60652 27784 60844 27824
rect 60884 27784 60885 27824
rect 60652 27656 60692 27784
rect 60843 27775 60885 27784
rect 60555 26984 60597 26993
rect 60555 26944 60556 26984
rect 60596 26944 60597 26984
rect 60555 26935 60597 26944
rect 60460 26692 60596 26732
rect 60459 26564 60501 26573
rect 60459 26524 60460 26564
rect 60500 26524 60501 26564
rect 60459 26515 60501 26524
rect 60172 26144 60212 26153
rect 60076 26104 60172 26144
rect 59980 26093 60020 26104
rect 60172 26095 60212 26104
rect 60267 26144 60309 26153
rect 60267 26104 60268 26144
rect 60308 26104 60309 26144
rect 60267 26095 60309 26104
rect 60268 26010 60308 26095
rect 60460 26060 60500 26515
rect 60556 26060 60596 26692
rect 60652 26321 60692 27616
rect 61035 27656 61077 27665
rect 61035 27616 61036 27656
rect 61076 27616 61077 27656
rect 61035 27607 61077 27616
rect 60748 27572 60788 27581
rect 60748 27161 60788 27532
rect 60844 27497 60884 27582
rect 60940 27572 60980 27581
rect 60843 27488 60885 27497
rect 60843 27448 60844 27488
rect 60884 27448 60885 27488
rect 60843 27439 60885 27448
rect 60747 27152 60789 27161
rect 60747 27112 60748 27152
rect 60788 27112 60789 27152
rect 60747 27103 60789 27112
rect 60747 26984 60789 26993
rect 60747 26944 60748 26984
rect 60788 26944 60789 26984
rect 60747 26935 60789 26944
rect 60651 26312 60693 26321
rect 60651 26272 60652 26312
rect 60692 26272 60693 26312
rect 60651 26263 60693 26272
rect 60556 26020 60692 26060
rect 60460 26011 60500 26020
rect 59979 25976 60021 25985
rect 59979 25936 59980 25976
rect 60020 25936 60021 25976
rect 59979 25927 60021 25936
rect 60652 25976 60692 26020
rect 59883 25892 59925 25901
rect 59883 25852 59884 25892
rect 59924 25852 59925 25892
rect 59883 25843 59925 25852
rect 59595 25808 59637 25817
rect 59595 25768 59596 25808
rect 59636 25768 59637 25808
rect 59595 25759 59637 25768
rect 59156 25432 59444 25472
rect 58924 24044 58964 24508
rect 59020 24380 59060 24389
rect 59020 24221 59060 24340
rect 59019 24212 59061 24221
rect 59019 24172 59020 24212
rect 59060 24172 59061 24212
rect 59019 24163 59061 24172
rect 58924 24004 59060 24044
rect 59020 23129 59060 24004
rect 59116 23801 59156 25432
rect 59211 25304 59253 25313
rect 59211 25264 59212 25304
rect 59252 25264 59253 25304
rect 59211 25255 59253 25264
rect 59404 25304 59444 25313
rect 59115 23792 59157 23801
rect 59115 23752 59116 23792
rect 59156 23752 59157 23792
rect 59115 23743 59157 23752
rect 59019 23120 59061 23129
rect 59019 23080 59020 23120
rect 59060 23080 59061 23120
rect 59019 23071 59061 23080
rect 59212 23060 59252 25255
rect 59404 24893 59444 25264
rect 59499 25304 59541 25313
rect 59499 25264 59500 25304
rect 59540 25264 59541 25304
rect 59499 25255 59541 25264
rect 59500 25170 59540 25255
rect 59596 25145 59636 25759
rect 59595 25136 59637 25145
rect 59788 25136 59828 25145
rect 59595 25092 59596 25136
rect 59636 25092 59637 25136
rect 59595 25087 59637 25092
rect 59692 25096 59788 25136
rect 59596 25001 59636 25087
rect 59403 24884 59445 24893
rect 59692 24884 59732 25096
rect 59788 25087 59828 25096
rect 59403 24844 59404 24884
rect 59444 24844 59445 24884
rect 59403 24835 59445 24844
rect 59596 24844 59732 24884
rect 59787 24884 59829 24893
rect 59787 24844 59788 24884
rect 59828 24844 59829 24884
rect 59500 24632 59540 24641
rect 59308 24592 59500 24632
rect 59308 23792 59348 24592
rect 59500 24583 59540 24592
rect 59596 23885 59636 24844
rect 59787 24835 59829 24844
rect 59691 24380 59733 24389
rect 59691 24340 59692 24380
rect 59732 24340 59733 24380
rect 59691 24331 59733 24340
rect 59595 23876 59637 23885
rect 59595 23836 59596 23876
rect 59636 23836 59637 23876
rect 59595 23827 59637 23836
rect 59308 23743 59348 23752
rect 59403 23792 59445 23801
rect 59403 23752 59404 23792
rect 59444 23752 59445 23792
rect 59403 23743 59445 23752
rect 59500 23792 59540 23801
rect 59404 23658 59444 23743
rect 59500 23624 59540 23752
rect 59596 23792 59636 23827
rect 59596 23743 59636 23752
rect 59595 23624 59637 23633
rect 59500 23584 59596 23624
rect 59636 23584 59637 23624
rect 59595 23575 59637 23584
rect 59499 23456 59541 23465
rect 59499 23416 59500 23456
rect 59540 23416 59541 23456
rect 59499 23407 59541 23416
rect 59500 23060 59540 23407
rect 59692 23060 59732 24331
rect 59788 23792 59828 24835
rect 59884 24809 59924 25843
rect 59980 25842 60020 25927
rect 60555 25892 60597 25901
rect 60555 25852 60556 25892
rect 60596 25852 60597 25892
rect 60555 25843 60597 25852
rect 60267 25724 60309 25733
rect 60267 25684 60268 25724
rect 60308 25684 60309 25724
rect 60267 25675 60309 25684
rect 59979 25556 60021 25565
rect 59979 25516 59980 25556
rect 60020 25516 60021 25556
rect 59979 25507 60021 25516
rect 59980 25388 60020 25507
rect 59980 25339 60020 25348
rect 60171 25388 60213 25397
rect 60171 25348 60172 25388
rect 60212 25348 60213 25388
rect 60171 25339 60213 25348
rect 60075 25304 60117 25313
rect 60075 25264 60076 25304
rect 60116 25264 60117 25304
rect 60075 25255 60117 25264
rect 59883 24800 59925 24809
rect 59883 24760 59884 24800
rect 59924 24760 59925 24800
rect 59883 24751 59925 24760
rect 59883 24632 59925 24641
rect 59883 24592 59884 24632
rect 59924 24592 59925 24632
rect 59883 24583 59925 24592
rect 59884 24498 59924 24583
rect 59883 23876 59925 23885
rect 59883 23836 59884 23876
rect 59924 23836 59925 23876
rect 59883 23827 59925 23836
rect 59788 23743 59828 23752
rect 59884 23792 59924 23827
rect 59980 23801 60020 23886
rect 59884 23741 59924 23752
rect 59979 23792 60021 23801
rect 59979 23752 59980 23792
rect 60020 23752 60021 23792
rect 59979 23743 60021 23752
rect 60076 23792 60116 25255
rect 60172 25254 60212 25339
rect 60171 24968 60213 24977
rect 60171 24928 60172 24968
rect 60212 24928 60213 24968
rect 60171 24919 60213 24928
rect 60076 23743 60116 23752
rect 59978 23120 60020 23129
rect 59978 23080 59979 23120
rect 60019 23080 60020 23120
rect 59978 23071 60020 23080
rect 58348 23020 58495 23060
rect 58636 23020 58785 23060
rect 58828 23020 58895 23060
rect 59212 23020 59295 23060
rect 59500 23020 59585 23060
rect 57255 22596 57295 23020
rect 57544 22868 57586 22877
rect 57544 22828 57545 22868
rect 57585 22828 57586 22868
rect 57544 22819 57586 22828
rect 57944 22868 57986 22877
rect 57944 22828 57945 22868
rect 57985 22828 57986 22868
rect 57944 22819 57986 22828
rect 57545 22596 57585 22819
rect 57654 22784 57696 22793
rect 57654 22744 57655 22784
rect 57695 22744 57696 22784
rect 57654 22735 57696 22744
rect 57655 22596 57695 22735
rect 57945 22596 57985 22819
rect 58055 22596 58095 23020
rect 58344 22952 58386 22961
rect 58344 22912 58345 22952
rect 58385 22912 58386 22952
rect 58344 22903 58386 22912
rect 58345 22596 58385 22903
rect 58455 22596 58495 23020
rect 58745 22596 58785 23020
rect 58855 22596 58895 23020
rect 59144 22784 59186 22793
rect 59144 22744 59145 22784
rect 59185 22744 59186 22784
rect 59144 22735 59186 22744
rect 59145 22596 59185 22735
rect 59255 22596 59295 23020
rect 59545 22596 59585 23020
rect 59655 23020 59732 23060
rect 59980 23060 60020 23071
rect 59980 23020 60095 23060
rect 59655 22596 59695 23020
rect 59944 22952 59986 22961
rect 59944 22912 59945 22952
rect 59985 22912 59986 22952
rect 59944 22903 59986 22912
rect 59945 22596 59985 22903
rect 60055 22596 60095 23020
rect 60172 22784 60212 24919
rect 60268 24893 60308 25675
rect 60363 25556 60405 25565
rect 60363 25516 60364 25556
rect 60404 25516 60405 25556
rect 60363 25507 60405 25516
rect 60556 25556 60596 25843
rect 60364 25422 60404 25507
rect 60556 25313 60596 25516
rect 60652 25388 60692 25936
rect 60748 25817 60788 26935
rect 60844 26909 60884 26940
rect 60843 26900 60885 26909
rect 60843 26860 60844 26900
rect 60884 26860 60885 26900
rect 60843 26851 60885 26860
rect 60844 26816 60884 26851
rect 60747 25808 60789 25817
rect 60747 25768 60748 25808
rect 60788 25768 60789 25808
rect 60747 25759 60789 25768
rect 60748 25565 60788 25759
rect 60747 25556 60789 25565
rect 60747 25516 60748 25556
rect 60788 25516 60789 25556
rect 60747 25507 60789 25516
rect 60748 25388 60788 25397
rect 60652 25348 60748 25388
rect 60748 25339 60788 25348
rect 60844 25313 60884 26776
rect 60940 25976 60980 27532
rect 61036 27522 61076 27607
rect 60980 25936 61076 25976
rect 60940 25927 60980 25936
rect 60555 25304 60597 25313
rect 60555 25264 60556 25304
rect 60596 25264 60597 25304
rect 60555 25255 60597 25264
rect 60843 25304 60885 25313
rect 60843 25264 60844 25304
rect 60884 25264 60885 25304
rect 60843 25255 60885 25264
rect 60940 25220 60980 25229
rect 60267 24884 60309 24893
rect 60267 24844 60268 24884
rect 60308 24844 60309 24884
rect 60267 24835 60309 24844
rect 60747 24800 60789 24809
rect 60747 24760 60748 24800
rect 60788 24760 60789 24800
rect 60747 24751 60789 24760
rect 60555 24716 60597 24725
rect 60555 24676 60556 24716
rect 60596 24676 60597 24716
rect 60555 24667 60597 24676
rect 60363 23792 60405 23801
rect 60363 23752 60364 23792
rect 60404 23752 60405 23792
rect 60363 23743 60405 23752
rect 60267 23624 60309 23633
rect 60267 23584 60268 23624
rect 60308 23584 60309 23624
rect 60267 23575 60309 23584
rect 60268 22961 60308 23575
rect 60364 23465 60404 23743
rect 60363 23456 60405 23465
rect 60363 23416 60364 23456
rect 60404 23416 60405 23456
rect 60363 23407 60405 23416
rect 60267 22952 60309 22961
rect 60267 22912 60268 22952
rect 60308 22912 60309 22952
rect 60267 22903 60309 22912
rect 60556 22868 60596 24667
rect 60748 24632 60788 24751
rect 60748 24583 60788 24592
rect 60940 23792 60980 25180
rect 60940 23743 60980 23752
rect 61036 23792 61076 25936
rect 61132 24389 61172 28456
rect 61228 27992 61268 30211
rect 61324 30092 61364 30101
rect 61612 30092 61652 30547
rect 61364 30052 61652 30092
rect 61324 30043 61364 30052
rect 61708 29924 61748 29933
rect 61324 29672 61364 29681
rect 61324 28673 61364 29632
rect 61516 29672 61556 29683
rect 61708 29681 61748 29884
rect 61516 29597 61556 29632
rect 61707 29672 61749 29681
rect 61707 29632 61708 29672
rect 61748 29632 61749 29672
rect 61707 29623 61749 29632
rect 61515 29588 61557 29597
rect 61515 29548 61516 29588
rect 61556 29548 61557 29588
rect 61515 29539 61557 29548
rect 61804 29345 61844 30640
rect 62476 30101 62516 34084
rect 62764 32864 62804 32875
rect 62764 32789 62804 32824
rect 62572 32780 62612 32789
rect 62572 31940 62612 32740
rect 62763 32780 62805 32789
rect 62763 32740 62764 32780
rect 62804 32740 62805 32780
rect 62763 32731 62805 32740
rect 62860 32705 62900 32790
rect 62859 32696 62901 32705
rect 62859 32656 62860 32696
rect 62900 32656 62901 32696
rect 62859 32647 62901 32656
rect 62956 32528 62996 34168
rect 63148 34159 63188 34168
rect 63244 33881 63284 34336
rect 63350 33956 63390 34355
rect 63531 34376 63573 34385
rect 63531 34336 63532 34376
rect 63572 34336 63573 34376
rect 63531 34327 63573 34336
rect 63628 34376 63668 34411
rect 63532 34150 63572 34327
rect 63350 33916 63476 33956
rect 63243 33872 63285 33881
rect 63243 33832 63244 33872
rect 63284 33832 63285 33872
rect 63243 33823 63285 33832
rect 63244 33461 63284 33823
rect 63436 33704 63476 33916
rect 63532 33872 63572 34110
rect 63628 33965 63668 34336
rect 63724 34376 63764 34385
rect 63627 33956 63669 33965
rect 63627 33916 63628 33956
rect 63668 33916 63669 33956
rect 63627 33907 63669 33916
rect 63724 33881 63764 34336
rect 63532 33823 63572 33832
rect 63723 33872 63765 33881
rect 63723 33832 63724 33872
rect 63764 33832 63765 33872
rect 63723 33823 63765 33832
rect 63628 33704 63668 33713
rect 63436 33664 63628 33704
rect 63628 33655 63668 33664
rect 63243 33452 63285 33461
rect 63243 33412 63244 33452
rect 63284 33412 63285 33452
rect 63243 33403 63285 33412
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 63820 33140 63860 35596
rect 64011 34964 64053 34973
rect 64011 34924 64012 34964
rect 64052 34924 64053 34964
rect 64011 34915 64053 34924
rect 64012 34830 64052 34915
rect 64011 34544 64053 34553
rect 63916 34504 64012 34544
rect 64052 34504 64053 34544
rect 63916 33704 63956 34504
rect 64011 34495 64053 34504
rect 64012 34410 64052 34495
rect 64204 34469 64244 35848
rect 64300 35888 64340 36007
rect 64588 35897 64628 36016
rect 64300 35839 64340 35848
rect 64587 35888 64629 35897
rect 64587 35848 64588 35888
rect 64628 35848 64629 35888
rect 64587 35839 64629 35848
rect 64780 35888 64820 36679
rect 64876 36233 64916 38116
rect 65068 37988 65108 37997
rect 64875 36224 64917 36233
rect 64875 36184 64876 36224
rect 64916 36184 64917 36224
rect 64875 36175 64917 36184
rect 65068 36149 65108 37948
rect 65164 37409 65204 38200
rect 65260 38191 65300 38200
rect 65452 38240 65492 38249
rect 65452 38081 65492 38200
rect 65548 38240 65588 38249
rect 65740 38240 65780 38249
rect 65588 38200 65740 38240
rect 65451 38072 65493 38081
rect 65451 38032 65452 38072
rect 65492 38032 65493 38072
rect 65451 38023 65493 38032
rect 65260 37988 65300 37997
rect 65260 37493 65300 37948
rect 65548 37904 65588 38200
rect 65740 38191 65780 38200
rect 66892 38240 66932 38249
rect 66892 38081 66932 38200
rect 68331 38240 68373 38249
rect 68331 38200 68332 38240
rect 68372 38200 68373 38240
rect 68331 38191 68373 38200
rect 68716 38240 68756 38249
rect 67755 38156 67797 38165
rect 67755 38116 67756 38156
rect 67796 38116 67797 38156
rect 67755 38107 67797 38116
rect 66507 38072 66549 38081
rect 66507 38032 66508 38072
rect 66548 38032 66549 38072
rect 66507 38023 66549 38032
rect 66891 38072 66933 38081
rect 66891 38032 66892 38072
rect 66932 38032 66933 38072
rect 66891 38023 66933 38032
rect 67756 38072 67796 38107
rect 68332 38106 68372 38191
rect 65835 37988 65877 37997
rect 65835 37948 65836 37988
rect 65876 37948 65877 37988
rect 65835 37939 65877 37948
rect 65452 37864 65588 37904
rect 65259 37484 65301 37493
rect 65259 37444 65260 37484
rect 65300 37444 65301 37484
rect 65259 37435 65301 37444
rect 65163 37400 65205 37409
rect 65163 37360 65164 37400
rect 65204 37360 65205 37400
rect 65163 37351 65205 37360
rect 65452 37241 65492 37864
rect 65836 37854 65876 37939
rect 65547 37400 65589 37409
rect 65547 37360 65548 37400
rect 65588 37360 65589 37400
rect 65547 37351 65589 37360
rect 65931 37400 65973 37409
rect 65931 37360 65932 37400
rect 65972 37360 65973 37400
rect 65931 37351 65973 37360
rect 65451 37232 65493 37241
rect 65451 37192 65452 37232
rect 65492 37192 65493 37232
rect 65451 37183 65493 37192
rect 65548 36728 65588 37351
rect 65932 37266 65972 37351
rect 65588 36688 65684 36728
rect 65548 36679 65588 36688
rect 65163 36224 65205 36233
rect 65163 36184 65164 36224
rect 65204 36184 65205 36224
rect 65163 36175 65205 36184
rect 65067 36140 65109 36149
rect 65067 36100 65068 36140
rect 65108 36100 65109 36140
rect 65067 36091 65109 36100
rect 64780 35839 64820 35848
rect 64875 35888 64917 35897
rect 64875 35848 64876 35888
rect 64916 35848 64917 35888
rect 64875 35839 64917 35848
rect 64972 35888 65012 35897
rect 64876 35754 64916 35839
rect 64972 35729 65012 35848
rect 65068 35888 65108 35897
rect 64971 35720 65013 35729
rect 64971 35680 64972 35720
rect 65012 35680 65013 35720
rect 64971 35671 65013 35680
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 64203 34460 64245 34469
rect 64203 34420 64204 34460
rect 64244 34420 64245 34460
rect 64203 34411 64245 34420
rect 64779 34460 64821 34469
rect 64779 34420 64780 34460
rect 64820 34420 64821 34460
rect 64779 34411 64821 34420
rect 64683 34376 64725 34385
rect 64683 34336 64684 34376
rect 64724 34336 64725 34376
rect 64683 34327 64725 34336
rect 64300 34292 64340 34301
rect 64012 34252 64300 34292
rect 64012 33872 64052 34252
rect 64300 34243 64340 34252
rect 64684 34242 64724 34327
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 64012 33823 64052 33832
rect 64491 33872 64533 33881
rect 64491 33832 64492 33872
rect 64532 33832 64533 33872
rect 64491 33823 64533 33832
rect 64299 33788 64341 33797
rect 64299 33748 64300 33788
rect 64340 33748 64341 33788
rect 64299 33739 64341 33748
rect 64108 33704 64148 33713
rect 63916 33664 64108 33704
rect 64108 33655 64148 33664
rect 64204 33704 64244 33713
rect 63915 33536 63957 33545
rect 63915 33496 63916 33536
rect 63956 33496 63957 33536
rect 63915 33487 63957 33496
rect 63147 33116 63189 33125
rect 63147 33076 63148 33116
rect 63188 33076 63189 33116
rect 63147 33067 63189 33076
rect 63628 33100 63860 33140
rect 63148 32864 63188 33067
rect 63532 33032 63572 33041
rect 63148 32815 63188 32824
rect 63244 32864 63284 32873
rect 63284 32824 63476 32864
rect 63244 32815 63284 32824
rect 63051 32696 63093 32705
rect 63051 32652 63052 32696
rect 63092 32652 63093 32696
rect 63051 32647 63093 32652
rect 62860 32488 62996 32528
rect 63052 32528 63092 32647
rect 63052 32488 63188 32528
rect 62763 32192 62805 32201
rect 62763 32152 62764 32192
rect 62804 32152 62805 32192
rect 62763 32143 62805 32152
rect 62764 32058 62804 32143
rect 62860 32108 62900 32488
rect 63148 32192 63188 32488
rect 63148 32143 63188 32152
rect 63339 32192 63381 32201
rect 63339 32152 63340 32192
rect 63380 32152 63381 32192
rect 63339 32143 63381 32152
rect 62860 32059 62900 32068
rect 63051 32108 63093 32117
rect 63051 32068 63052 32108
rect 63092 32068 63093 32108
rect 63051 32059 63093 32068
rect 62956 32024 62996 32033
rect 62956 31940 62996 31984
rect 63052 31974 63092 32059
rect 63340 32058 63380 32143
rect 63436 31949 63476 32824
rect 63532 32117 63572 32992
rect 63531 32108 63573 32117
rect 63531 32068 63532 32108
rect 63572 32068 63573 32108
rect 63531 32059 63573 32068
rect 62572 31900 62996 31940
rect 63435 31940 63477 31949
rect 63435 31900 63436 31940
rect 63476 31900 63477 31940
rect 63435 31891 63477 31900
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 63532 31604 63572 32059
rect 63340 31564 63572 31604
rect 63243 31436 63285 31445
rect 63243 31396 63244 31436
rect 63284 31396 63285 31436
rect 63243 31387 63285 31396
rect 63340 31394 63380 31564
rect 63244 31352 63284 31387
rect 63340 31345 63380 31354
rect 63436 31352 63476 31361
rect 63244 31301 63284 31312
rect 62571 30680 62613 30689
rect 62571 30640 62572 30680
rect 62612 30640 62613 30680
rect 62571 30631 62613 30640
rect 62572 30546 62612 30631
rect 63436 30521 63476 31312
rect 63531 31352 63573 31361
rect 63531 31312 63532 31352
rect 63572 31312 63573 31352
rect 63531 31303 63573 31312
rect 63532 31218 63572 31303
rect 63435 30512 63477 30521
rect 63435 30472 63436 30512
rect 63476 30472 63477 30512
rect 63435 30463 63477 30472
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 62475 30092 62517 30101
rect 62475 30052 62476 30092
rect 62516 30052 62517 30092
rect 62475 30043 62517 30052
rect 63531 30092 63573 30101
rect 63531 30052 63532 30092
rect 63572 30052 63573 30092
rect 63531 30043 63573 30052
rect 61899 30008 61941 30017
rect 61899 29968 61900 30008
rect 61940 29968 61941 30008
rect 61899 29959 61941 29968
rect 61900 29874 61940 29959
rect 62092 29924 62132 29933
rect 61803 29336 61845 29345
rect 61803 29296 61804 29336
rect 61844 29296 61845 29336
rect 61803 29287 61845 29296
rect 61900 29168 61940 29177
rect 61516 29128 61900 29168
rect 61323 28664 61365 28673
rect 61323 28624 61324 28664
rect 61364 28624 61365 28664
rect 61323 28615 61365 28624
rect 61324 28496 61364 28507
rect 61324 28421 61364 28456
rect 61323 28412 61365 28421
rect 61323 28372 61324 28412
rect 61364 28372 61365 28412
rect 61323 28363 61365 28372
rect 61516 28328 61556 29128
rect 61900 29119 61940 29128
rect 62092 28925 62132 29884
rect 62283 29168 62325 29177
rect 62283 29128 62284 29168
rect 62324 29128 62325 29168
rect 62283 29119 62325 29128
rect 62284 29034 62324 29119
rect 62476 29093 62516 30043
rect 63148 29168 63188 29177
rect 62956 29128 63148 29168
rect 62475 29084 62517 29093
rect 62475 29044 62476 29084
rect 62516 29044 62517 29084
rect 62475 29035 62517 29044
rect 61708 28916 61748 28925
rect 62091 28916 62133 28925
rect 61748 28876 61940 28916
rect 61708 28867 61748 28876
rect 61803 28664 61845 28673
rect 61803 28624 61804 28664
rect 61844 28624 61845 28664
rect 61803 28615 61845 28624
rect 61611 28412 61653 28421
rect 61611 28372 61612 28412
rect 61652 28372 61653 28412
rect 61611 28363 61653 28372
rect 61516 28279 61556 28288
rect 61612 28328 61652 28363
rect 61612 28277 61652 28288
rect 61708 28328 61748 28337
rect 61708 28169 61748 28288
rect 61804 28328 61844 28615
rect 61804 28279 61844 28288
rect 61900 28253 61940 28876
rect 62091 28876 62092 28916
rect 62132 28876 62133 28916
rect 62091 28867 62133 28876
rect 62091 28664 62133 28673
rect 62091 28624 62092 28664
rect 62132 28624 62133 28664
rect 62091 28615 62133 28624
rect 61995 28328 62037 28337
rect 61995 28288 61996 28328
rect 62036 28288 62037 28328
rect 61995 28279 62037 28288
rect 62092 28328 62132 28615
rect 62283 28496 62325 28505
rect 62283 28456 62284 28496
rect 62324 28456 62325 28496
rect 62283 28447 62325 28456
rect 62187 28412 62229 28421
rect 62187 28372 62188 28412
rect 62228 28372 62229 28412
rect 62187 28363 62229 28372
rect 62092 28279 62132 28288
rect 62188 28328 62228 28363
rect 61899 28244 61941 28253
rect 61899 28204 61900 28244
rect 61940 28204 61941 28244
rect 61899 28195 61941 28204
rect 61707 28160 61749 28169
rect 61707 28120 61708 28160
rect 61748 28120 61749 28160
rect 61707 28111 61749 28120
rect 61228 27952 61460 27992
rect 61227 27824 61269 27833
rect 61227 27784 61228 27824
rect 61268 27784 61269 27824
rect 61227 27775 61269 27784
rect 61228 27656 61268 27775
rect 61228 27607 61268 27616
rect 61420 27656 61460 27952
rect 61900 27833 61940 28195
rect 61996 28194 62036 28279
rect 62188 28277 62228 28288
rect 62284 28328 62324 28447
rect 62859 28412 62901 28421
rect 62859 28372 62860 28412
rect 62900 28372 62901 28412
rect 62859 28363 62901 28372
rect 62284 28279 62324 28288
rect 62860 28328 62900 28363
rect 62956 28337 62996 29128
rect 63148 29119 63188 29128
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 63051 28580 63093 28589
rect 63051 28540 63052 28580
rect 63092 28540 63093 28580
rect 63051 28531 63093 28540
rect 62860 28277 62900 28288
rect 62955 28328 62997 28337
rect 62955 28288 62956 28328
rect 62996 28288 62997 28328
rect 62955 28279 62997 28288
rect 63052 28328 63092 28531
rect 63052 28279 63092 28288
rect 63436 28328 63476 28337
rect 63532 28328 63572 30043
rect 63476 28288 63572 28328
rect 63436 28279 63476 28288
rect 62763 28160 62805 28169
rect 62763 28120 62764 28160
rect 62804 28120 62900 28160
rect 62763 28111 62805 28120
rect 62764 28026 62804 28111
rect 61515 27824 61557 27833
rect 61515 27784 61516 27824
rect 61556 27784 61557 27824
rect 61515 27775 61557 27784
rect 61899 27824 61941 27833
rect 61899 27784 61900 27824
rect 61940 27784 61941 27824
rect 61899 27775 61941 27784
rect 61323 27488 61365 27497
rect 61323 27448 61324 27488
rect 61364 27448 61365 27488
rect 61323 27439 61365 27448
rect 61228 27404 61268 27413
rect 61228 27161 61268 27364
rect 61227 27152 61269 27161
rect 61227 27112 61228 27152
rect 61268 27112 61269 27152
rect 61227 27103 61269 27112
rect 61228 26816 61268 26825
rect 61324 26816 61364 27439
rect 61268 26776 61364 26816
rect 61420 27068 61460 27616
rect 61516 27656 61556 27775
rect 61516 27607 61556 27616
rect 61899 27656 61941 27665
rect 61899 27616 61900 27656
rect 61940 27616 61941 27656
rect 61899 27607 61941 27616
rect 62380 27656 62420 27665
rect 61228 26767 61268 26776
rect 61420 26741 61460 27028
rect 61900 27068 61940 27607
rect 61900 27019 61940 27028
rect 62380 26993 62420 27616
rect 62764 27656 62804 27665
rect 62571 27236 62613 27245
rect 62571 27196 62572 27236
rect 62612 27196 62613 27236
rect 62571 27187 62613 27196
rect 62379 26984 62421 26993
rect 62379 26944 62380 26984
rect 62420 26944 62421 26984
rect 62379 26935 62421 26944
rect 61611 26900 61653 26909
rect 61611 26860 61612 26900
rect 61652 26860 61653 26900
rect 61611 26851 61653 26860
rect 62091 26900 62133 26909
rect 62091 26860 62092 26900
rect 62132 26860 62133 26900
rect 62091 26851 62133 26860
rect 61612 26766 61652 26851
rect 61803 26816 61845 26825
rect 61803 26776 61804 26816
rect 61844 26776 61845 26816
rect 61803 26767 61845 26776
rect 61419 26732 61461 26741
rect 61419 26692 61420 26732
rect 61460 26692 61461 26732
rect 61419 26683 61461 26692
rect 61804 26682 61844 26767
rect 61900 26648 61940 26657
rect 61900 26405 61940 26608
rect 61419 26396 61461 26405
rect 61419 26347 61420 26396
rect 61460 26347 61461 26396
rect 61899 26396 61941 26405
rect 61899 26356 61900 26396
rect 61940 26356 61941 26396
rect 61899 26347 61941 26356
rect 61420 26261 61460 26330
rect 61324 26153 61364 26238
rect 61228 26144 61268 26153
rect 61228 25976 61268 26104
rect 61323 26144 61365 26153
rect 61323 26104 61324 26144
rect 61364 26104 61365 26144
rect 61323 26095 61365 26104
rect 61708 26144 61748 26153
rect 61708 25976 61748 26104
rect 61228 25936 61748 25976
rect 61804 26144 61844 26153
rect 61323 25304 61365 25313
rect 61323 25264 61324 25304
rect 61364 25264 61365 25304
rect 61323 25255 61365 25264
rect 61324 24725 61364 25255
rect 61323 24716 61365 24725
rect 61323 24676 61324 24716
rect 61364 24676 61365 24716
rect 61323 24667 61365 24676
rect 61323 24548 61365 24557
rect 61323 24508 61324 24548
rect 61364 24508 61365 24548
rect 61323 24499 61365 24508
rect 61227 24464 61269 24473
rect 61227 24424 61228 24464
rect 61268 24424 61269 24464
rect 61227 24415 61269 24424
rect 61131 24380 61173 24389
rect 61131 24340 61132 24380
rect 61172 24340 61173 24380
rect 61131 24331 61173 24340
rect 61228 23885 61268 24415
rect 61227 23876 61269 23885
rect 61227 23836 61228 23876
rect 61268 23836 61269 23876
rect 61227 23827 61269 23836
rect 61036 23743 61076 23752
rect 61131 23792 61173 23801
rect 61131 23752 61132 23792
rect 61172 23752 61173 23792
rect 61131 23743 61173 23752
rect 61228 23792 61268 23827
rect 61132 23658 61172 23743
rect 61228 23742 61268 23752
rect 61131 23204 61173 23213
rect 61131 23164 61132 23204
rect 61172 23164 61173 23204
rect 61131 23155 61173 23164
rect 61132 23060 61172 23155
rect 61324 23060 61364 24499
rect 61804 24473 61844 26104
rect 61900 26144 61940 26153
rect 61900 24716 61940 26104
rect 61996 26144 62036 26153
rect 61996 25901 62036 26104
rect 61995 25892 62037 25901
rect 61995 25852 61996 25892
rect 62036 25852 62037 25892
rect 61995 25843 62037 25852
rect 61996 25145 62036 25843
rect 62092 25649 62132 26851
rect 62283 26648 62325 26657
rect 62283 26608 62284 26648
rect 62324 26608 62325 26648
rect 62283 26599 62325 26608
rect 62091 25640 62133 25649
rect 62091 25600 62092 25640
rect 62132 25600 62133 25640
rect 62091 25591 62133 25600
rect 62188 25304 62228 25313
rect 61995 25136 62037 25145
rect 61995 25096 61996 25136
rect 62036 25096 62037 25136
rect 61995 25087 62037 25096
rect 62188 24809 62228 25264
rect 62187 24800 62229 24809
rect 62187 24760 62188 24800
rect 62228 24760 62229 24800
rect 62187 24751 62229 24760
rect 61900 24676 62036 24716
rect 61900 24548 61940 24557
rect 61803 24464 61845 24473
rect 61803 24424 61804 24464
rect 61844 24424 61845 24464
rect 61803 24415 61845 24424
rect 61803 24128 61845 24137
rect 61803 24088 61804 24128
rect 61844 24088 61845 24128
rect 61803 24079 61845 24088
rect 61804 23633 61844 24079
rect 61803 23624 61845 23633
rect 61803 23584 61804 23624
rect 61844 23584 61845 23624
rect 61803 23575 61845 23584
rect 61900 23465 61940 24508
rect 61996 23885 62036 24676
rect 62187 24380 62229 24389
rect 62187 24340 62188 24380
rect 62228 24340 62229 24380
rect 62187 24331 62229 24340
rect 62091 24128 62133 24137
rect 62091 24088 62092 24128
rect 62132 24088 62133 24128
rect 62091 24079 62133 24088
rect 61995 23876 62037 23885
rect 61995 23836 61996 23876
rect 62036 23836 62037 23876
rect 61995 23827 62037 23836
rect 62092 23792 62132 24079
rect 62188 24044 62228 24331
rect 62188 23995 62228 24004
rect 62284 23876 62324 26599
rect 62475 24296 62517 24305
rect 62475 24256 62476 24296
rect 62516 24256 62517 24296
rect 62572 24296 62612 27187
rect 62764 26069 62804 27616
rect 62763 26060 62805 26069
rect 62763 26020 62764 26060
rect 62804 26020 62805 26060
rect 62763 26011 62805 26020
rect 62763 25808 62805 25817
rect 62763 25768 62764 25808
rect 62804 25768 62805 25808
rect 62763 25759 62805 25768
rect 62667 25220 62709 25229
rect 62667 25180 62668 25220
rect 62708 25180 62709 25220
rect 62667 25171 62709 25180
rect 62668 24548 62708 25171
rect 62764 24632 62804 25759
rect 62860 24809 62900 28120
rect 63628 27824 63668 33100
rect 63820 32948 63860 32957
rect 63916 32948 63956 33487
rect 64011 33368 64053 33377
rect 64011 33328 64012 33368
rect 64052 33328 64053 33368
rect 64011 33319 64053 33328
rect 63860 32908 63956 32948
rect 63820 32899 63860 32908
rect 64012 32864 64052 33319
rect 63916 32824 64052 32864
rect 63916 32780 63956 32824
rect 63820 32740 63956 32780
rect 63723 32192 63765 32201
rect 63723 32152 63724 32192
rect 63764 32152 63765 32192
rect 63723 32143 63765 32152
rect 63724 32058 63764 32143
rect 63723 31940 63765 31949
rect 63723 31900 63724 31940
rect 63764 31900 63765 31940
rect 63723 31891 63765 31900
rect 63724 31352 63764 31891
rect 63724 31303 63764 31312
rect 63820 31352 63860 32740
rect 64012 32696 64052 32705
rect 64012 31865 64052 32656
rect 64204 32360 64244 33664
rect 64300 33704 64340 33739
rect 64492 33738 64532 33823
rect 64300 33629 64340 33664
rect 64588 33704 64628 33715
rect 64588 33629 64628 33664
rect 64683 33704 64725 33713
rect 64683 33664 64684 33704
rect 64724 33664 64725 33704
rect 64683 33655 64725 33664
rect 64780 33704 64820 34411
rect 65068 33797 65108 35848
rect 65164 34385 65204 36175
rect 65259 36056 65301 36065
rect 65259 36016 65260 36056
rect 65300 36016 65301 36056
rect 65259 36007 65301 36016
rect 65260 35888 65300 36007
rect 65644 35981 65684 36688
rect 66219 36056 66261 36065
rect 66219 36016 66220 36056
rect 66260 36016 66261 36056
rect 66219 36007 66261 36016
rect 65643 35972 65685 35981
rect 65643 35932 65644 35972
rect 65684 35932 65685 35972
rect 65643 35923 65685 35932
rect 65260 35839 65300 35848
rect 65356 35888 65396 35897
rect 65163 34376 65205 34385
rect 65163 34336 65164 34376
rect 65204 34336 65205 34376
rect 65163 34327 65205 34336
rect 65356 34301 65396 35848
rect 65451 35888 65493 35897
rect 65451 35848 65452 35888
rect 65492 35848 65493 35888
rect 65451 35839 65493 35848
rect 65548 35888 65588 35897
rect 65452 35754 65492 35839
rect 65548 35645 65588 35848
rect 65547 35636 65589 35645
rect 65547 35596 65548 35636
rect 65588 35596 65589 35636
rect 65547 35587 65589 35596
rect 65548 34376 65588 34385
rect 65644 34376 65684 35923
rect 65835 35888 65877 35897
rect 65835 35848 65836 35888
rect 65876 35848 65877 35888
rect 65835 35839 65877 35848
rect 65836 35754 65876 35839
rect 65739 35720 65781 35729
rect 65739 35680 65740 35720
rect 65780 35680 65781 35720
rect 65739 35671 65781 35680
rect 65740 35057 65780 35671
rect 65739 35048 65781 35057
rect 65739 35008 65740 35048
rect 65780 35008 65781 35048
rect 65739 34999 65781 35008
rect 65588 34336 65684 34376
rect 65548 34327 65588 34336
rect 65355 34292 65397 34301
rect 65355 34252 65356 34292
rect 65396 34252 65397 34292
rect 65355 34243 65397 34252
rect 65067 33788 65109 33797
rect 65067 33748 65068 33788
rect 65108 33748 65109 33788
rect 65067 33739 65109 33748
rect 64299 33620 64341 33629
rect 64299 33580 64300 33620
rect 64340 33580 64341 33620
rect 64299 33571 64341 33580
rect 64587 33620 64629 33629
rect 64587 33580 64588 33620
rect 64628 33580 64629 33620
rect 64587 33571 64629 33580
rect 64300 33540 64340 33571
rect 64588 33377 64628 33571
rect 64684 33570 64724 33655
rect 64780 33545 64820 33664
rect 64779 33536 64821 33545
rect 64779 33496 64780 33536
rect 64820 33496 64821 33536
rect 64779 33487 64821 33496
rect 64587 33368 64629 33377
rect 64587 33328 64588 33368
rect 64628 33328 64629 33368
rect 64587 33319 64629 33328
rect 64875 33200 64917 33209
rect 64875 33160 64876 33200
rect 64916 33160 64917 33200
rect 64875 33151 64917 33160
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 64108 32320 64244 32360
rect 64011 31856 64053 31865
rect 64011 31816 64012 31856
rect 64052 31816 64053 31856
rect 64011 31807 64053 31816
rect 63820 31303 63860 31312
rect 63915 31352 63957 31361
rect 63915 31312 63916 31352
rect 63956 31312 63957 31352
rect 63915 31303 63957 31312
rect 64012 31352 64052 31807
rect 64012 31303 64052 31312
rect 63916 31218 63956 31303
rect 64012 30680 64052 30689
rect 63723 30428 63765 30437
rect 63723 30388 63724 30428
rect 63764 30388 63765 30428
rect 63723 30379 63765 30388
rect 63724 30294 63764 30379
rect 64012 30269 64052 30640
rect 64011 30260 64053 30269
rect 64011 30220 64012 30260
rect 64052 30220 64053 30260
rect 64011 30211 64053 30220
rect 63532 27784 63668 27824
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 63243 25976 63285 25985
rect 63243 25936 63244 25976
rect 63284 25936 63285 25976
rect 63243 25927 63285 25936
rect 63244 25842 63284 25927
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 63051 25472 63093 25481
rect 63051 25432 63052 25472
rect 63092 25432 63093 25472
rect 63051 25423 63093 25432
rect 62859 24800 62901 24809
rect 62859 24760 62860 24800
rect 62900 24760 62901 24800
rect 62859 24751 62901 24760
rect 62860 24632 62900 24641
rect 62764 24592 62860 24632
rect 62860 24583 62900 24592
rect 62956 24632 62996 24641
rect 62668 24508 62804 24548
rect 62667 24296 62709 24305
rect 62572 24256 62668 24296
rect 62708 24256 62709 24296
rect 62475 24247 62517 24256
rect 62667 24247 62709 24256
rect 62092 23743 62132 23752
rect 62188 23836 62324 23876
rect 61899 23456 61941 23465
rect 61899 23416 61900 23456
rect 61940 23416 61941 23456
rect 61899 23407 61941 23416
rect 61611 23372 61653 23381
rect 61611 23332 61612 23372
rect 61652 23332 61653 23372
rect 61611 23323 61653 23332
rect 60854 23036 60896 23045
rect 60854 22996 60855 23036
rect 60895 22996 60896 23036
rect 61132 23020 61185 23060
rect 60854 22987 60896 22996
rect 60747 22868 60789 22877
rect 60455 22828 60596 22868
rect 60745 22828 60748 22868
rect 60788 22828 60789 22868
rect 60172 22744 60385 22784
rect 60345 22596 60385 22744
rect 60455 22596 60495 22828
rect 60745 22819 60789 22828
rect 60745 22596 60785 22819
rect 60855 22596 60895 22987
rect 61145 22596 61185 23020
rect 61255 23020 61364 23060
rect 61612 23060 61652 23323
rect 62188 23060 62228 23836
rect 62379 23624 62421 23633
rect 62379 23584 62380 23624
rect 62420 23584 62421 23624
rect 62379 23575 62421 23584
rect 62380 23060 62420 23575
rect 61612 23020 61695 23060
rect 61255 22596 61295 23020
rect 61544 22784 61586 22793
rect 61544 22744 61545 22784
rect 61585 22744 61586 22784
rect 61544 22735 61586 22744
rect 61545 22596 61585 22735
rect 61655 22596 61695 23020
rect 62055 23020 62228 23060
rect 62345 23020 62420 23060
rect 62476 23060 62516 24247
rect 62667 23876 62709 23885
rect 62667 23836 62668 23876
rect 62708 23836 62709 23876
rect 62667 23827 62709 23836
rect 62571 23792 62613 23801
rect 62571 23752 62572 23792
rect 62612 23752 62613 23792
rect 62571 23743 62613 23752
rect 62668 23792 62708 23827
rect 62572 23658 62612 23743
rect 62668 23297 62708 23752
rect 62667 23288 62709 23297
rect 62667 23248 62668 23288
rect 62708 23248 62709 23288
rect 62667 23239 62709 23248
rect 62764 23060 62804 24508
rect 62859 24380 62901 24389
rect 62859 24340 62860 24380
rect 62900 24340 62901 24380
rect 62859 24331 62901 24340
rect 62860 24137 62900 24331
rect 62859 24128 62901 24137
rect 62859 24088 62860 24128
rect 62900 24088 62901 24128
rect 62859 24079 62901 24088
rect 62859 23876 62901 23885
rect 62859 23836 62860 23876
rect 62900 23836 62901 23876
rect 62859 23827 62901 23836
rect 62860 23633 62900 23827
rect 62859 23624 62901 23633
rect 62859 23584 62860 23624
rect 62900 23584 62901 23624
rect 62859 23575 62901 23584
rect 62956 23381 62996 24592
rect 63052 24632 63092 25423
rect 63340 25136 63380 25145
rect 63380 25096 63476 25136
rect 63340 25087 63380 25096
rect 63052 24583 63092 24592
rect 63148 24632 63188 24641
rect 63340 24632 63380 24641
rect 63188 24592 63340 24632
rect 63148 24583 63188 24592
rect 63340 24583 63380 24592
rect 63051 24296 63093 24305
rect 63051 24256 63052 24296
rect 63092 24256 63093 24296
rect 63051 24247 63093 24256
rect 62955 23372 62997 23381
rect 62955 23332 62956 23372
rect 62996 23332 62997 23372
rect 62955 23323 62997 23332
rect 62476 23020 62612 23060
rect 61944 22784 61986 22793
rect 61944 22744 61945 22784
rect 61985 22744 61986 22784
rect 61944 22735 61986 22744
rect 61945 22596 61985 22735
rect 62055 22596 62095 23020
rect 62345 22596 62385 23020
rect 62572 22784 62612 23020
rect 62455 22744 62612 22784
rect 62745 23020 62804 23060
rect 62455 22596 62495 22744
rect 62745 22596 62785 23020
rect 63052 22784 63092 24247
rect 63147 24044 63189 24053
rect 63147 24004 63148 24044
rect 63188 24004 63189 24044
rect 63147 23995 63189 24004
rect 63148 23060 63188 23995
rect 63244 23876 63284 23885
rect 63284 23836 63380 23876
rect 63244 23827 63284 23836
rect 63243 23708 63285 23717
rect 63243 23668 63244 23708
rect 63284 23668 63285 23708
rect 63243 23659 63285 23668
rect 62855 22744 63092 22784
rect 63145 23020 63188 23060
rect 63244 23060 63284 23659
rect 63340 23549 63380 23836
rect 63339 23540 63381 23549
rect 63339 23500 63340 23540
rect 63380 23500 63381 23540
rect 63339 23491 63381 23500
rect 63436 23297 63476 25096
rect 63532 24641 63572 27784
rect 63627 27656 63669 27665
rect 63627 27616 63628 27656
rect 63668 27616 63669 27656
rect 63627 27607 63669 27616
rect 63628 27522 63668 27607
rect 64108 26993 64148 32320
rect 64203 32192 64245 32201
rect 64203 32152 64204 32192
rect 64244 32152 64245 32192
rect 64203 32143 64245 32152
rect 64587 32192 64629 32201
rect 64587 32152 64588 32192
rect 64628 32152 64629 32192
rect 64587 32143 64629 32152
rect 64204 30680 64244 32143
rect 64588 32058 64628 32143
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 64396 30680 64436 30689
rect 64204 30640 64396 30680
rect 64396 30101 64436 30640
rect 64876 30185 64916 33151
rect 65068 33140 65108 33739
rect 65356 33629 65396 34243
rect 65355 33620 65397 33629
rect 65355 33580 65356 33620
rect 65396 33580 65397 33620
rect 65355 33571 65397 33580
rect 64972 33100 65108 33140
rect 64875 30176 64917 30185
rect 64875 30136 64876 30176
rect 64916 30136 64917 30176
rect 64875 30127 64917 30136
rect 64395 30092 64437 30101
rect 64395 30052 64396 30092
rect 64436 30052 64437 30092
rect 64395 30043 64437 30052
rect 64780 29840 64820 29849
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 64491 29336 64533 29345
rect 64491 29296 64492 29336
rect 64532 29296 64533 29336
rect 64491 29287 64533 29296
rect 64492 29168 64532 29287
rect 64780 29261 64820 29800
rect 64876 29840 64916 30127
rect 64876 29791 64916 29800
rect 64972 29597 65012 33100
rect 65644 32873 65684 34336
rect 65836 32957 65876 32988
rect 66220 32957 66260 36007
rect 66411 35804 66453 35813
rect 66411 35764 66412 35804
rect 66452 35764 66453 35804
rect 66411 35755 66453 35764
rect 66412 35670 66452 35755
rect 65835 32948 65877 32957
rect 65835 32908 65836 32948
rect 65876 32908 65877 32948
rect 65835 32899 65877 32908
rect 66219 32948 66261 32957
rect 66219 32908 66220 32948
rect 66260 32908 66261 32948
rect 66219 32899 66261 32908
rect 65643 32864 65685 32873
rect 65643 32824 65644 32864
rect 65684 32824 65685 32864
rect 65643 32815 65685 32824
rect 65836 32864 65876 32899
rect 65452 32780 65492 32789
rect 65452 32033 65492 32740
rect 65644 32201 65684 32815
rect 65836 32285 65876 32824
rect 66508 32453 66548 38023
rect 67756 38021 67796 38032
rect 66700 37988 66740 37997
rect 66700 37409 66740 37948
rect 67467 37988 67509 37997
rect 67467 37948 67468 37988
rect 67508 37948 67509 37988
rect 67467 37939 67509 37948
rect 67371 37484 67413 37493
rect 67371 37444 67372 37484
rect 67412 37444 67413 37484
rect 67371 37435 67413 37444
rect 67468 37484 67508 37939
rect 68427 37484 68469 37493
rect 67468 37444 67700 37484
rect 66699 37400 66741 37409
rect 66699 37360 66700 37400
rect 66740 37360 66741 37400
rect 66699 37351 66741 37360
rect 66796 37400 66836 37409
rect 66700 36476 66740 36485
rect 66604 36436 66700 36476
rect 66604 35897 66644 36436
rect 66700 36427 66740 36436
rect 66796 36065 66836 37360
rect 67372 37350 67412 37435
rect 67180 37316 67220 37325
rect 67220 37276 67316 37316
rect 67180 37267 67220 37276
rect 67083 36812 67125 36821
rect 67083 36772 67084 36812
rect 67124 36772 67125 36812
rect 67083 36763 67125 36772
rect 67084 36728 67124 36763
rect 66795 36056 66837 36065
rect 66795 36016 66796 36056
rect 66836 36016 66837 36056
rect 66795 36007 66837 36016
rect 66603 35888 66645 35897
rect 66603 35848 66604 35888
rect 66644 35848 66645 35888
rect 66603 35839 66645 35848
rect 66796 35888 66836 36007
rect 66796 35839 66836 35848
rect 66507 32444 66549 32453
rect 66507 32404 66508 32444
rect 66548 32404 66549 32444
rect 66507 32395 66549 32404
rect 66604 32285 66644 35839
rect 66987 34460 67029 34469
rect 66987 34420 66988 34460
rect 67028 34420 67029 34460
rect 66987 34411 67029 34420
rect 66795 34292 66837 34301
rect 66795 34252 66796 34292
rect 66836 34252 66837 34292
rect 66795 34243 66837 34252
rect 66700 34208 66740 34217
rect 66700 33713 66740 34168
rect 66699 33704 66741 33713
rect 66699 33664 66700 33704
rect 66740 33664 66741 33704
rect 66699 33655 66741 33664
rect 66796 33704 66836 34243
rect 66700 33368 66740 33655
rect 66796 33545 66836 33664
rect 66892 33704 66932 33715
rect 66892 33629 66932 33664
rect 66988 33704 67028 34411
rect 67084 34376 67124 36688
rect 67180 36644 67220 36655
rect 67180 36569 67220 36604
rect 67179 36560 67221 36569
rect 67179 36520 67180 36560
rect 67220 36520 67221 36560
rect 67179 36511 67221 36520
rect 67276 36560 67316 37276
rect 67371 36896 67413 36905
rect 67371 36856 67372 36896
rect 67412 36856 67413 36896
rect 67371 36847 67413 36856
rect 67372 36644 67412 36847
rect 67468 36728 67508 37444
rect 67564 37325 67604 37356
rect 67563 37316 67605 37325
rect 67563 37276 67564 37316
rect 67604 37276 67605 37316
rect 67563 37267 67605 37276
rect 67468 36679 67508 36688
rect 67564 37232 67604 37267
rect 67372 36595 67412 36604
rect 67276 36511 67316 36520
rect 67275 35804 67317 35813
rect 67275 35764 67276 35804
rect 67316 35764 67317 35804
rect 67275 35755 67317 35764
rect 67180 34553 67220 34597
rect 67179 34544 67221 34553
rect 67179 34504 67180 34544
rect 67220 34504 67221 34544
rect 67179 34502 67221 34504
rect 67179 34495 67180 34502
rect 67220 34495 67221 34502
rect 67276 34544 67316 35755
rect 67564 35720 67604 37192
rect 67660 36954 67700 37444
rect 68427 37444 68428 37484
rect 68468 37444 68469 37484
rect 68427 37435 68469 37444
rect 67755 37232 67797 37241
rect 67755 37192 67756 37232
rect 67796 37192 67797 37232
rect 67755 37183 67797 37192
rect 67756 37098 67796 37183
rect 67660 36905 67700 36914
rect 68139 36896 68181 36905
rect 68139 36856 68140 36896
rect 68180 36856 68181 36896
rect 68139 36847 68181 36856
rect 67756 36728 67796 36737
rect 67659 36056 67701 36065
rect 67659 36016 67660 36056
rect 67700 36016 67701 36056
rect 67659 36007 67701 36016
rect 67756 36056 67796 36688
rect 67851 36728 67893 36737
rect 67851 36688 67852 36728
rect 67892 36688 67893 36728
rect 67851 36679 67893 36688
rect 67852 36594 67892 36679
rect 68140 36560 68180 36847
rect 68235 36812 68277 36821
rect 68235 36772 68236 36812
rect 68276 36772 68372 36812
rect 68235 36763 68277 36772
rect 68332 36728 68372 36772
rect 68332 36679 68372 36688
rect 68140 36511 68180 36520
rect 68331 36560 68373 36569
rect 68331 36520 68332 36560
rect 68372 36520 68373 36560
rect 68331 36511 68373 36520
rect 68332 36426 68372 36511
rect 67756 36016 68084 36056
rect 67660 35888 67700 36007
rect 67660 35839 67700 35848
rect 67564 35680 67700 35720
rect 67660 34964 67700 35680
rect 67756 35645 67796 36016
rect 67851 35888 67893 35897
rect 67851 35848 67852 35888
rect 67892 35848 67893 35888
rect 67851 35839 67893 35848
rect 67755 35636 67797 35645
rect 67755 35596 67756 35636
rect 67796 35596 67797 35636
rect 67755 35587 67797 35596
rect 67660 34924 67796 34964
rect 67276 34495 67316 34504
rect 67372 34502 67412 34554
rect 67660 34544 67700 34553
rect 67660 34502 67700 34504
rect 67372 34469 67700 34502
rect 67180 34453 67220 34462
rect 67371 34462 67700 34469
rect 67371 34460 67413 34462
rect 67371 34420 67372 34460
rect 67412 34420 67413 34460
rect 67371 34411 67413 34420
rect 67468 34376 67508 34387
rect 67124 34336 67316 34376
rect 67084 34327 67124 34336
rect 66988 33655 67028 33664
rect 67083 33704 67125 33713
rect 67083 33664 67084 33704
rect 67124 33664 67125 33704
rect 67083 33655 67125 33664
rect 67276 33704 67316 34336
rect 67468 34301 67508 34336
rect 67563 34376 67605 34385
rect 67563 34336 67564 34376
rect 67604 34336 67605 34376
rect 67563 34327 67605 34336
rect 67467 34292 67509 34301
rect 67467 34252 67468 34292
rect 67508 34252 67509 34292
rect 67467 34243 67509 34252
rect 67564 33956 67604 34327
rect 67756 34049 67796 34924
rect 67755 34040 67797 34049
rect 67755 34000 67756 34040
rect 67796 34000 67797 34040
rect 67755 33991 67797 34000
rect 67391 33916 67604 33956
rect 67391 33881 67431 33916
rect 67372 33872 67431 33881
rect 67412 33832 67431 33872
rect 67372 33823 67412 33832
rect 67852 33797 67892 35839
rect 67947 34376 67989 34385
rect 67947 34336 67948 34376
rect 67988 34336 67989 34376
rect 67947 34327 67989 34336
rect 68044 34376 68084 36016
rect 68235 35720 68277 35729
rect 68235 35680 68236 35720
rect 68276 35680 68277 35720
rect 68235 35671 68277 35680
rect 68236 35216 68276 35671
rect 68236 35167 68276 35176
rect 68235 35048 68277 35057
rect 68235 35008 68236 35048
rect 68276 35008 68277 35048
rect 68235 34999 68277 35008
rect 67948 34242 67988 34327
rect 67467 33788 67509 33797
rect 67467 33748 67468 33788
rect 67508 33748 67509 33788
rect 67467 33739 67509 33748
rect 67851 33788 67893 33797
rect 67851 33748 67852 33788
rect 67892 33748 67893 33788
rect 67851 33739 67893 33748
rect 66891 33620 66933 33629
rect 66891 33580 66892 33620
rect 66932 33580 66933 33620
rect 66891 33571 66933 33580
rect 67084 33570 67124 33655
rect 66795 33536 66837 33545
rect 66795 33496 66796 33536
rect 66836 33496 66837 33536
rect 66795 33487 66837 33496
rect 66700 33328 67028 33368
rect 66699 32864 66741 32873
rect 66699 32824 66700 32864
rect 66740 32824 66741 32864
rect 66699 32815 66741 32824
rect 66700 32730 66740 32815
rect 66795 32696 66837 32705
rect 66795 32656 66796 32696
rect 66836 32656 66837 32696
rect 66795 32647 66837 32656
rect 65835 32276 65877 32285
rect 65835 32236 65836 32276
rect 65876 32236 65877 32276
rect 65835 32227 65877 32236
rect 66603 32276 66645 32285
rect 66603 32236 66604 32276
rect 66644 32236 66645 32276
rect 66603 32227 66645 32236
rect 65643 32192 65685 32201
rect 65643 32152 65644 32192
rect 65684 32152 65685 32192
rect 65643 32143 65685 32152
rect 66123 32192 66165 32201
rect 66123 32152 66124 32192
rect 66164 32152 66165 32192
rect 66123 32143 66165 32152
rect 66411 32192 66453 32201
rect 66411 32152 66412 32192
rect 66452 32152 66453 32192
rect 66411 32143 66453 32152
rect 66796 32192 66836 32647
rect 66796 32143 66836 32152
rect 65451 32024 65493 32033
rect 65451 31984 65452 32024
rect 65492 31984 65493 32024
rect 65451 31975 65493 31984
rect 65740 31940 65780 31949
rect 65355 31772 65397 31781
rect 65355 31732 65356 31772
rect 65396 31732 65397 31772
rect 65355 31723 65397 31732
rect 65260 30680 65300 30689
rect 65164 30640 65260 30680
rect 65068 30017 65108 30102
rect 65067 30008 65109 30017
rect 65067 29968 65068 30008
rect 65108 29968 65109 30008
rect 65067 29959 65109 29968
rect 65067 29840 65109 29849
rect 65067 29800 65068 29840
rect 65108 29800 65109 29840
rect 65067 29791 65109 29800
rect 65068 29706 65108 29791
rect 64971 29588 65013 29597
rect 64971 29548 64972 29588
rect 65012 29548 65013 29588
rect 64971 29539 65013 29548
rect 64779 29252 64821 29261
rect 64779 29212 64780 29252
rect 64820 29212 64821 29252
rect 64779 29203 64821 29212
rect 64492 29119 64532 29128
rect 64875 29168 64917 29177
rect 64875 29128 64876 29168
rect 64916 29128 64917 29168
rect 64875 29119 64917 29128
rect 64588 29084 64628 29093
rect 64300 28916 64340 28925
rect 64340 28876 64436 28916
rect 64300 28867 64340 28876
rect 64299 28748 64341 28757
rect 64299 28708 64300 28748
rect 64340 28708 64341 28748
rect 64299 28699 64341 28708
rect 64203 28328 64245 28337
rect 64300 28328 64340 28699
rect 64396 28337 64436 28876
rect 64203 28288 64204 28328
rect 64244 28288 64300 28328
rect 64203 28279 64245 28288
rect 64300 28279 64340 28288
rect 64395 28328 64437 28337
rect 64395 28288 64396 28328
rect 64436 28288 64437 28328
rect 64395 28279 64437 28288
rect 64204 27665 64244 28279
rect 64588 28160 64628 29044
rect 64780 29084 64820 29093
rect 64684 29000 64724 29009
rect 64684 28841 64724 28960
rect 64683 28832 64725 28841
rect 64683 28792 64684 28832
rect 64724 28792 64725 28832
rect 64683 28783 64725 28792
rect 64780 28244 64820 29044
rect 64876 29034 64916 29119
rect 65164 28757 65204 30640
rect 65260 30631 65300 30640
rect 65356 30512 65396 31723
rect 65740 31361 65780 31900
rect 66124 31781 66164 32143
rect 66412 32058 66452 32143
rect 66508 32108 66548 32117
rect 66123 31772 66165 31781
rect 66123 31732 66124 31772
rect 66164 31732 66165 31772
rect 66123 31723 66165 31732
rect 65739 31352 65781 31361
rect 65739 31312 65740 31352
rect 65780 31312 65781 31352
rect 66124 31352 66164 31723
rect 66508 31688 66548 32068
rect 66700 32108 66740 32117
rect 66603 32024 66645 32033
rect 66603 31984 66604 32024
rect 66644 31984 66645 32024
rect 66700 32024 66740 32068
rect 66795 32024 66837 32033
rect 66700 31984 66796 32024
rect 66836 31984 66837 32024
rect 66603 31975 66645 31984
rect 66795 31975 66837 31984
rect 66604 31890 66644 31975
rect 66891 31856 66933 31865
rect 66891 31816 66892 31856
rect 66932 31816 66933 31856
rect 66891 31807 66933 31816
rect 66220 31648 66548 31688
rect 66220 31604 66260 31648
rect 66220 31555 66260 31564
rect 66220 31352 66260 31361
rect 66412 31352 66452 31361
rect 66124 31312 66220 31352
rect 65739 31303 65781 31312
rect 66220 31303 66260 31312
rect 66316 31312 66412 31352
rect 65835 31184 65877 31193
rect 65835 31144 65836 31184
rect 65876 31144 65877 31184
rect 65835 31135 65877 31144
rect 65260 30472 65396 30512
rect 65260 29933 65300 30472
rect 65739 30344 65781 30353
rect 65739 30304 65740 30344
rect 65780 30304 65781 30344
rect 65739 30295 65781 30304
rect 65451 30260 65493 30269
rect 65451 30220 65452 30260
rect 65492 30220 65493 30260
rect 65451 30211 65493 30220
rect 65355 30008 65397 30017
rect 65355 29968 65356 30008
rect 65396 29968 65397 30008
rect 65355 29959 65397 29968
rect 65452 30008 65492 30211
rect 65452 29959 65492 29968
rect 65259 29924 65301 29933
rect 65259 29884 65260 29924
rect 65300 29884 65301 29924
rect 65259 29882 65301 29884
rect 65259 29875 65260 29882
rect 65300 29875 65301 29882
rect 65356 29924 65396 29959
rect 65356 29873 65396 29884
rect 65547 29924 65589 29933
rect 65547 29884 65548 29924
rect 65588 29884 65589 29924
rect 65547 29875 65589 29884
rect 65260 29833 65300 29842
rect 65451 29840 65493 29849
rect 65451 29800 65452 29840
rect 65492 29800 65493 29840
rect 65451 29791 65493 29800
rect 65452 29336 65492 29791
rect 65548 29790 65588 29875
rect 65644 29840 65684 29849
rect 65644 29681 65684 29800
rect 65643 29672 65685 29681
rect 65643 29632 65644 29672
rect 65684 29632 65685 29672
rect 65643 29623 65685 29632
rect 65547 29588 65589 29597
rect 65547 29548 65548 29588
rect 65588 29548 65589 29588
rect 65547 29539 65589 29548
rect 65452 29287 65492 29296
rect 65355 29252 65397 29261
rect 65355 29212 65356 29252
rect 65396 29212 65397 29252
rect 65355 29203 65397 29212
rect 65259 29084 65301 29093
rect 65259 29044 65260 29084
rect 65300 29044 65301 29084
rect 65259 29035 65301 29044
rect 65260 28950 65300 29035
rect 65259 28832 65301 28841
rect 65259 28792 65260 28832
rect 65300 28792 65301 28832
rect 65259 28783 65301 28792
rect 65163 28748 65205 28757
rect 65163 28708 65164 28748
rect 65204 28708 65205 28748
rect 65163 28699 65205 28708
rect 65260 28412 65300 28783
rect 65356 28580 65396 29203
rect 65451 29168 65493 29177
rect 65451 29128 65452 29168
rect 65492 29128 65493 29168
rect 65451 29119 65493 29128
rect 65452 28748 65492 29119
rect 65548 29093 65588 29539
rect 65740 29504 65780 30295
rect 65644 29464 65780 29504
rect 65547 29084 65589 29093
rect 65547 29044 65548 29084
rect 65588 29044 65589 29084
rect 65547 29035 65589 29044
rect 65644 28748 65684 29464
rect 65836 29345 65876 31135
rect 66316 30185 66356 31312
rect 66412 31303 66452 31312
rect 66508 31352 66548 31361
rect 66508 31016 66548 31312
rect 66412 30976 66548 31016
rect 66412 30848 66452 30976
rect 66412 30773 66452 30808
rect 66411 30764 66453 30773
rect 66411 30724 66412 30764
rect 66452 30724 66453 30764
rect 66411 30715 66453 30724
rect 66412 30684 66452 30715
rect 66604 30680 66644 30689
rect 66315 30176 66357 30185
rect 66315 30136 66316 30176
rect 66356 30136 66357 30176
rect 66315 30127 66357 30136
rect 65932 30008 65972 30017
rect 65932 29933 65972 29968
rect 65931 29924 65973 29933
rect 65931 29884 65932 29924
rect 65972 29884 65973 29924
rect 65931 29875 65973 29884
rect 66315 29924 66357 29933
rect 66315 29884 66316 29924
rect 66356 29884 66357 29924
rect 66315 29875 66357 29884
rect 65932 29588 65972 29875
rect 66219 29840 66261 29849
rect 66219 29800 66220 29840
rect 66260 29800 66261 29840
rect 66219 29791 66261 29800
rect 66316 29840 66356 29875
rect 66604 29849 66644 30640
rect 66699 30680 66741 30689
rect 66699 30640 66700 30680
rect 66740 30640 66741 30680
rect 66699 30631 66741 30640
rect 66796 30680 66836 30689
rect 66700 30546 66740 30631
rect 66220 29706 66260 29791
rect 66316 29789 66356 29800
rect 66603 29840 66645 29849
rect 66603 29800 66604 29840
rect 66644 29800 66645 29840
rect 66603 29791 66645 29800
rect 66700 29756 66740 29765
rect 66411 29672 66453 29681
rect 66411 29628 66412 29672
rect 66452 29628 66453 29672
rect 66411 29623 66453 29628
rect 65932 29548 66260 29588
rect 65835 29336 65877 29345
rect 65835 29296 65836 29336
rect 65876 29296 65877 29336
rect 65835 29287 65877 29296
rect 65836 29168 65876 29177
rect 65836 28925 65876 29128
rect 65932 29168 65972 29177
rect 65932 29009 65972 29128
rect 66028 29168 66068 29177
rect 65931 29000 65973 29009
rect 65931 28960 65932 29000
rect 65972 28960 65973 29000
rect 65931 28951 65973 28960
rect 65835 28916 65877 28925
rect 65835 28876 65836 28916
rect 65876 28876 65877 28916
rect 65835 28867 65877 28876
rect 65452 28708 65588 28748
rect 65644 28708 65876 28748
rect 65452 28580 65492 28589
rect 65356 28540 65452 28580
rect 65548 28580 65588 28708
rect 65740 28580 65780 28589
rect 65548 28540 65740 28580
rect 65452 28496 65492 28540
rect 65740 28531 65780 28540
rect 65452 28456 65684 28496
rect 65260 28372 65492 28412
rect 65259 28244 65301 28253
rect 64780 28204 65108 28244
rect 64588 28120 64820 28160
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 64780 27824 64820 28120
rect 64396 27784 64820 27824
rect 64203 27656 64245 27665
rect 64203 27616 64204 27656
rect 64244 27616 64245 27656
rect 64203 27607 64245 27616
rect 63915 26984 63957 26993
rect 63915 26944 63916 26984
rect 63956 26944 63957 26984
rect 63915 26935 63957 26944
rect 64107 26984 64149 26993
rect 64107 26944 64108 26984
rect 64148 26944 64149 26984
rect 64107 26935 64149 26944
rect 63820 26900 63860 26909
rect 63723 26816 63765 26825
rect 63723 26776 63724 26816
rect 63764 26776 63765 26816
rect 63723 26767 63765 26776
rect 63724 26682 63764 26767
rect 63627 26060 63669 26069
rect 63627 26020 63628 26060
rect 63668 26020 63669 26060
rect 63627 26011 63669 26020
rect 63628 25313 63668 26011
rect 63723 25472 63765 25481
rect 63820 25472 63860 26860
rect 63916 26850 63956 26935
rect 64012 26900 64052 26909
rect 63915 26732 63957 26741
rect 63915 26692 63916 26732
rect 63956 26692 63957 26732
rect 63915 26683 63957 26692
rect 63916 25892 63956 26683
rect 64012 25976 64052 26860
rect 64108 26816 64148 26825
rect 64108 26321 64148 26776
rect 64107 26312 64149 26321
rect 64107 26272 64108 26312
rect 64148 26272 64149 26312
rect 64107 26263 64149 26272
rect 64204 26144 64244 27607
rect 64396 27068 64436 27784
rect 65068 27665 65108 28204
rect 65259 28204 65260 28244
rect 65300 28204 65301 28244
rect 65259 28195 65301 28204
rect 65067 27656 65109 27665
rect 65067 27616 65068 27656
rect 65108 27616 65109 27656
rect 65067 27607 65109 27616
rect 65068 27488 65108 27607
rect 65068 27439 65108 27448
rect 64396 27019 64436 27028
rect 64780 27404 64820 27413
rect 64395 26900 64437 26909
rect 64395 26860 64396 26900
rect 64436 26860 64437 26900
rect 64395 26851 64437 26860
rect 64396 26816 64436 26851
rect 64396 26765 64436 26776
rect 64588 26816 64628 26825
rect 64588 26657 64628 26776
rect 64684 26816 64724 26825
rect 64780 26816 64820 27364
rect 64875 27404 64917 27413
rect 64875 27364 64876 27404
rect 64916 27364 65012 27404
rect 64875 27355 64917 27364
rect 64972 27320 65012 27364
rect 64972 27280 65108 27320
rect 64876 26816 64916 26844
rect 64724 26776 64876 26816
rect 64684 26767 64724 26776
rect 64876 26767 64916 26776
rect 64971 26816 65013 26825
rect 64971 26776 64972 26816
rect 65012 26776 65013 26816
rect 64971 26767 65013 26776
rect 64972 26682 65012 26767
rect 64587 26648 64629 26657
rect 64587 26608 64588 26648
rect 64628 26608 64820 26648
rect 64587 26599 64629 26608
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 64683 26312 64725 26321
rect 64683 26272 64684 26312
rect 64724 26272 64725 26312
rect 64683 26263 64725 26272
rect 64396 26144 64436 26153
rect 64204 26104 64396 26144
rect 64396 26095 64436 26104
rect 64012 25936 64628 25976
rect 63916 25852 64244 25892
rect 63723 25432 63724 25472
rect 63764 25432 63860 25472
rect 63723 25423 63765 25432
rect 63724 25338 63764 25423
rect 64108 25397 64148 25428
rect 64107 25388 64149 25397
rect 64107 25348 64108 25388
rect 64148 25348 64149 25388
rect 64107 25339 64149 25348
rect 63627 25304 63669 25313
rect 63627 25264 63628 25304
rect 63668 25264 63669 25304
rect 63627 25255 63669 25264
rect 64012 25304 64052 25313
rect 63531 24632 63573 24641
rect 63531 24592 63532 24632
rect 63572 24592 63573 24632
rect 63628 24632 63668 25255
rect 63724 24632 63764 24641
rect 63628 24592 63724 24632
rect 63531 24583 63573 24592
rect 63724 24583 63764 24592
rect 64012 24464 64052 25264
rect 64108 25304 64148 25339
rect 64108 25145 64148 25264
rect 64107 25136 64149 25145
rect 64107 25096 64108 25136
rect 64148 25096 64149 25136
rect 64107 25087 64149 25096
rect 64204 25132 64244 25852
rect 64588 25556 64628 25936
rect 64588 25507 64628 25516
rect 64588 25262 64628 25271
rect 64587 25222 64588 25229
rect 64628 25222 64629 25229
rect 64587 25220 64629 25222
rect 64684 25220 64724 26263
rect 64587 25180 64588 25220
rect 64628 25180 64724 25220
rect 64780 25304 64820 26608
rect 64971 26564 65013 26573
rect 64971 26524 64972 26564
rect 65012 26524 65013 26564
rect 64971 26515 65013 26524
rect 64875 25976 64917 25985
rect 64875 25936 64876 25976
rect 64916 25936 64917 25976
rect 64875 25927 64917 25936
rect 64587 25171 64629 25180
rect 64588 25127 64628 25171
rect 64780 25145 64820 25264
rect 64876 25304 64916 25927
rect 64876 25255 64916 25264
rect 64779 25136 64821 25145
rect 64108 24725 64148 25087
rect 64204 25083 64244 25092
rect 64779 25096 64780 25136
rect 64820 25096 64821 25136
rect 64779 25087 64821 25096
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 64683 24800 64725 24809
rect 64683 24760 64684 24800
rect 64724 24760 64725 24800
rect 64683 24751 64725 24760
rect 64107 24716 64149 24725
rect 64107 24676 64108 24716
rect 64148 24676 64149 24716
rect 64107 24667 64149 24676
rect 64491 24716 64533 24725
rect 64491 24676 64492 24716
rect 64532 24676 64533 24716
rect 64491 24667 64533 24676
rect 64299 24464 64341 24473
rect 64012 24424 64244 24464
rect 63627 24212 63669 24221
rect 63627 24172 63628 24212
rect 63668 24172 63669 24212
rect 63627 24163 63669 24172
rect 63531 23960 63573 23969
rect 63531 23920 63532 23960
rect 63572 23920 63573 23960
rect 63531 23911 63573 23920
rect 63435 23288 63477 23297
rect 63435 23248 63436 23288
rect 63476 23248 63477 23288
rect 63435 23239 63477 23248
rect 63532 23060 63572 23911
rect 63628 23060 63668 24163
rect 64011 24044 64053 24053
rect 64011 24004 64012 24044
rect 64052 24004 64053 24044
rect 64011 23995 64053 24004
rect 64012 23910 64052 23995
rect 63916 23792 63956 23803
rect 63916 23717 63956 23752
rect 64204 23792 64244 24424
rect 64299 24424 64300 24464
rect 64340 24424 64341 24464
rect 64299 24415 64341 24424
rect 64300 23885 64340 24415
rect 64299 23876 64341 23885
rect 64299 23836 64300 23876
rect 64340 23836 64341 23876
rect 64299 23827 64341 23836
rect 64204 23743 64244 23752
rect 64300 23792 64340 23827
rect 64300 23741 64340 23752
rect 64395 23792 64437 23801
rect 64395 23752 64396 23792
rect 64436 23752 64437 23792
rect 64395 23743 64437 23752
rect 64492 23792 64532 24667
rect 64587 24632 64629 24641
rect 64587 24592 64588 24632
rect 64628 24592 64629 24632
rect 64587 24583 64629 24592
rect 64588 24498 64628 24583
rect 64492 23743 64532 23752
rect 63915 23708 63957 23717
rect 63915 23668 63916 23708
rect 63956 23668 63957 23708
rect 63915 23659 63957 23668
rect 64396 23658 64436 23743
rect 64299 23624 64341 23633
rect 64299 23584 64300 23624
rect 64340 23584 64341 23624
rect 64299 23575 64341 23584
rect 64011 23456 64053 23465
rect 64011 23416 64012 23456
rect 64052 23416 64053 23456
rect 64011 23407 64053 23416
rect 64012 23060 64052 23407
rect 64300 23060 64340 23575
rect 64491 23288 64533 23297
rect 64491 23248 64492 23288
rect 64532 23248 64533 23288
rect 64491 23239 64533 23248
rect 64492 23060 64532 23239
rect 63244 23020 63295 23060
rect 63532 23020 63585 23060
rect 63628 23020 63695 23060
rect 64012 23020 64095 23060
rect 64300 23020 64385 23060
rect 62855 22596 62895 22744
rect 63145 22596 63185 23020
rect 63255 22596 63295 23020
rect 63545 22596 63585 23020
rect 63655 22596 63695 23020
rect 63944 22952 63986 22961
rect 63944 22912 63945 22952
rect 63985 22912 63986 22952
rect 63944 22903 63986 22912
rect 63945 22596 63985 22903
rect 64055 22596 64095 23020
rect 64345 22596 64385 23020
rect 64455 23020 64532 23060
rect 64684 23060 64724 24751
rect 64779 23792 64821 23801
rect 64779 23752 64780 23792
rect 64820 23752 64821 23792
rect 64779 23743 64821 23752
rect 64780 23658 64820 23743
rect 64876 23624 64916 23633
rect 64876 23381 64916 23584
rect 64875 23372 64917 23381
rect 64875 23332 64876 23372
rect 64916 23332 64917 23372
rect 64875 23323 64917 23332
rect 64972 23060 65012 26515
rect 64684 23020 64785 23060
rect 64455 22596 64495 23020
rect 64745 22596 64785 23020
rect 64855 23020 65012 23060
rect 65068 23060 65108 27280
rect 65163 26984 65205 26993
rect 65163 26944 65164 26984
rect 65204 26944 65205 26984
rect 65163 26935 65205 26944
rect 65164 24716 65204 26935
rect 65260 26573 65300 28195
rect 65355 28160 65397 28169
rect 65355 28120 65356 28160
rect 65396 28120 65397 28160
rect 65355 28111 65397 28120
rect 65356 27656 65396 28111
rect 65356 27607 65396 27616
rect 65452 27656 65492 28372
rect 65644 28328 65684 28456
rect 65836 28421 65876 28708
rect 65835 28412 65877 28421
rect 65835 28372 65836 28412
rect 65876 28372 65877 28412
rect 65835 28363 65877 28372
rect 65644 28279 65684 28288
rect 65932 28244 65972 28253
rect 65740 28160 65780 28169
rect 65548 28120 65740 28160
rect 65548 27882 65588 28120
rect 65740 28111 65780 28120
rect 65548 27833 65588 27842
rect 65932 27824 65972 28204
rect 66028 27992 66068 29128
rect 66124 29168 66164 29177
rect 66220 29168 66260 29548
rect 66412 29537 66452 29623
rect 66700 29420 66740 29716
rect 66796 29513 66836 30640
rect 66892 30680 66932 31807
rect 66988 30932 67028 33328
rect 67276 32201 67316 33664
rect 67468 33704 67508 33739
rect 67371 33536 67413 33545
rect 67371 33496 67372 33536
rect 67412 33496 67413 33536
rect 67371 33487 67413 33496
rect 67275 32192 67317 32201
rect 67275 32152 67276 32192
rect 67316 32152 67317 32192
rect 67275 32143 67317 32152
rect 67180 32033 67220 32064
rect 67179 32024 67221 32033
rect 67179 31984 67180 32024
rect 67220 31984 67221 32024
rect 67179 31975 67221 31984
rect 67180 31940 67220 31975
rect 67180 31352 67220 31900
rect 67276 31361 67316 31446
rect 67180 31303 67220 31312
rect 67275 31352 67317 31361
rect 67275 31312 67276 31352
rect 67316 31312 67317 31352
rect 67275 31303 67317 31312
rect 67372 31352 67412 33487
rect 67468 33209 67508 33664
rect 67564 33704 67604 33713
rect 67467 33200 67509 33209
rect 67467 33160 67468 33200
rect 67508 33160 67509 33200
rect 67467 33151 67509 33160
rect 67564 33140 67604 33664
rect 67755 33704 67797 33713
rect 67755 33664 67756 33704
rect 67796 33664 67797 33704
rect 67755 33655 67797 33664
rect 67756 33570 67796 33655
rect 68044 33536 68084 34336
rect 68140 34964 68180 34973
rect 68140 34301 68180 34924
rect 68139 34292 68181 34301
rect 68139 34252 68140 34292
rect 68180 34252 68181 34292
rect 68139 34243 68181 34252
rect 68140 34204 68180 34243
rect 68140 34155 68180 34164
rect 68139 34040 68181 34049
rect 68139 34000 68140 34040
rect 68180 34000 68181 34040
rect 68139 33991 68181 34000
rect 68140 33704 68180 33991
rect 68140 33655 68180 33664
rect 68044 33496 68180 33536
rect 67564 33116 67892 33140
rect 67564 33100 67852 33116
rect 67892 33076 68084 33116
rect 67852 33067 67892 33076
rect 67563 32864 67605 32873
rect 67563 32824 67564 32864
rect 67604 32824 67605 32864
rect 67563 32815 67605 32824
rect 68044 32864 68084 33076
rect 68140 32873 68180 33496
rect 68044 32815 68084 32824
rect 68139 32864 68181 32873
rect 68139 32824 68140 32864
rect 68180 32824 68181 32864
rect 68139 32815 68181 32824
rect 67468 32192 67508 32201
rect 67468 31781 67508 32152
rect 67564 32192 67604 32815
rect 67659 32696 67701 32705
rect 67659 32656 67660 32696
rect 67700 32656 67701 32696
rect 67659 32647 67701 32656
rect 68139 32696 68181 32705
rect 68139 32656 68140 32696
rect 68180 32656 68181 32696
rect 68139 32647 68181 32656
rect 67660 32418 67700 32647
rect 68140 32562 68180 32647
rect 67660 32369 67700 32378
rect 67659 32276 67701 32285
rect 67659 32236 67660 32276
rect 67700 32236 67701 32276
rect 67659 32227 67701 32236
rect 67564 31865 67604 32152
rect 67563 31856 67605 31865
rect 67563 31816 67564 31856
rect 67604 31816 67605 31856
rect 67563 31807 67605 31816
rect 67467 31772 67509 31781
rect 67467 31732 67468 31772
rect 67508 31732 67509 31772
rect 67467 31723 67509 31732
rect 67083 31184 67125 31193
rect 67083 31144 67084 31184
rect 67124 31144 67125 31184
rect 67083 31135 67125 31144
rect 67084 31050 67124 31135
rect 66988 30892 67316 30932
rect 67083 30764 67125 30773
rect 67083 30724 67084 30764
rect 67124 30724 67125 30764
rect 67083 30715 67125 30724
rect 66892 29933 66932 30640
rect 66987 30680 67029 30689
rect 66987 30640 66988 30680
rect 67028 30640 67029 30680
rect 66987 30631 67029 30640
rect 67084 30680 67124 30715
rect 66891 29924 66933 29933
rect 66891 29884 66892 29924
rect 66932 29884 66933 29924
rect 66891 29875 66933 29884
rect 66795 29504 66837 29513
rect 66795 29464 66796 29504
rect 66836 29464 66837 29504
rect 66795 29455 66837 29464
rect 66316 29380 66740 29420
rect 66316 29336 66356 29380
rect 66988 29336 67028 30631
rect 67084 30629 67124 30640
rect 67276 30512 67316 30892
rect 67372 30689 67412 31312
rect 67564 31268 67604 31277
rect 67467 31184 67509 31193
rect 67564 31184 67604 31228
rect 67467 31144 67468 31184
rect 67508 31144 67604 31184
rect 67467 31135 67509 31144
rect 67371 30680 67413 30689
rect 67371 30640 67372 30680
rect 67412 30640 67413 30680
rect 67371 30631 67413 30640
rect 67276 30472 67604 30512
rect 67180 30428 67220 30437
rect 67083 30092 67125 30101
rect 67083 30052 67084 30092
rect 67124 30052 67125 30092
rect 67083 30043 67125 30052
rect 67084 29840 67124 30043
rect 67084 29791 67124 29800
rect 67180 29681 67220 30388
rect 67179 29672 67221 29681
rect 67179 29632 67180 29672
rect 67220 29632 67221 29672
rect 67179 29623 67221 29632
rect 67371 29504 67413 29513
rect 67371 29464 67372 29504
rect 67412 29464 67413 29504
rect 67371 29455 67413 29464
rect 66316 29287 66356 29296
rect 66604 29296 66988 29336
rect 66412 29168 66452 29177
rect 66220 29128 66412 29168
rect 66124 28169 66164 29128
rect 66412 29119 66452 29128
rect 66508 29168 66548 29177
rect 66411 29000 66453 29009
rect 66411 28960 66412 29000
rect 66452 28960 66453 29000
rect 66411 28951 66453 28960
rect 66315 28664 66357 28673
rect 66315 28624 66316 28664
rect 66356 28624 66357 28664
rect 66315 28615 66357 28624
rect 66316 28328 66356 28615
rect 66123 28160 66165 28169
rect 66123 28120 66124 28160
rect 66164 28120 66165 28160
rect 66123 28111 66165 28120
rect 66028 27952 66260 27992
rect 66028 27824 66068 27833
rect 65932 27784 66028 27824
rect 66028 27775 66068 27784
rect 65740 27656 65780 27665
rect 65452 27607 65492 27616
rect 65548 27616 65740 27656
rect 65259 26564 65301 26573
rect 65259 26524 65260 26564
rect 65300 26524 65301 26564
rect 65259 26515 65301 26524
rect 65260 26144 65300 26155
rect 65260 26069 65300 26104
rect 65259 26060 65301 26069
rect 65259 26020 65260 26060
rect 65300 26020 65301 26060
rect 65259 26011 65301 26020
rect 65451 25976 65493 25985
rect 65451 25936 65452 25976
rect 65492 25936 65493 25976
rect 65451 25927 65493 25936
rect 65452 25304 65492 25927
rect 65548 25817 65588 27616
rect 65740 27607 65780 27616
rect 65836 27656 65876 27665
rect 65836 27413 65876 27616
rect 65931 27656 65973 27665
rect 65931 27616 65932 27656
rect 65972 27616 65973 27656
rect 65931 27607 65973 27616
rect 65932 27522 65972 27607
rect 65835 27404 65877 27413
rect 65835 27364 65836 27404
rect 65876 27364 65877 27404
rect 65835 27355 65877 27364
rect 65739 27068 65781 27077
rect 65739 27028 65740 27068
rect 65780 27028 65781 27068
rect 65739 27019 65781 27028
rect 65643 26144 65685 26153
rect 65643 26104 65644 26144
rect 65684 26104 65685 26144
rect 65643 26095 65685 26104
rect 65644 26010 65684 26095
rect 65547 25808 65589 25817
rect 65547 25768 65548 25808
rect 65588 25768 65589 25808
rect 65547 25759 65589 25768
rect 65740 25724 65780 27019
rect 65931 26144 65973 26153
rect 65931 26104 65932 26144
rect 65972 26104 65973 26144
rect 65931 26095 65973 26104
rect 66123 26144 66165 26153
rect 66123 26104 66124 26144
rect 66164 26104 66165 26144
rect 66123 26095 66165 26104
rect 65644 25684 65780 25724
rect 65452 25255 65492 25264
rect 65547 25304 65589 25313
rect 65547 25264 65548 25304
rect 65588 25264 65589 25304
rect 65547 25255 65589 25264
rect 65548 25170 65588 25255
rect 65547 24884 65589 24893
rect 65547 24844 65548 24884
rect 65588 24844 65589 24884
rect 65547 24835 65589 24844
rect 65164 24676 65300 24716
rect 65163 24296 65205 24305
rect 65163 24256 65164 24296
rect 65204 24256 65205 24296
rect 65163 24247 65205 24256
rect 65164 23792 65204 24247
rect 65260 24044 65300 24676
rect 65260 23995 65300 24004
rect 65451 23960 65493 23969
rect 65451 23920 65452 23960
rect 65492 23920 65493 23960
rect 65451 23911 65493 23920
rect 65452 23826 65492 23911
rect 65164 23743 65204 23752
rect 65260 23624 65300 23633
rect 65300 23584 65396 23624
rect 65260 23575 65300 23584
rect 65068 23020 65185 23060
rect 65356 23045 65396 23584
rect 65548 23060 65588 24835
rect 64855 22596 64895 23020
rect 65145 22596 65185 23020
rect 65254 23036 65296 23045
rect 65254 22996 65255 23036
rect 65295 22996 65296 23036
rect 65254 22987 65296 22996
rect 65355 23036 65397 23045
rect 65355 22996 65356 23036
rect 65396 22996 65397 23036
rect 65355 22987 65397 22996
rect 65545 23020 65588 23060
rect 65644 23060 65684 25684
rect 65835 25472 65877 25481
rect 65835 25432 65836 25472
rect 65876 25432 65877 25472
rect 65835 25423 65877 25432
rect 65932 25472 65972 26095
rect 66124 26010 66164 26095
rect 66220 25640 66260 27952
rect 66316 27917 66356 28288
rect 66412 27992 66452 28951
rect 66508 28841 66548 29128
rect 66604 29168 66644 29296
rect 66988 29287 67028 29296
rect 66604 29119 66644 29128
rect 67372 29168 67412 29455
rect 67372 29119 67412 29128
rect 66795 29084 66837 29093
rect 66795 29044 66796 29084
rect 66836 29044 66837 29084
rect 66795 29035 66837 29044
rect 66796 28950 66836 29035
rect 67468 28916 67508 28927
rect 67468 28841 67508 28876
rect 66507 28832 66549 28841
rect 66507 28792 66508 28832
rect 66548 28792 66549 28832
rect 66507 28783 66549 28792
rect 67467 28832 67509 28841
rect 67467 28792 67468 28832
rect 67508 28792 67509 28832
rect 67467 28783 67509 28792
rect 67179 28748 67221 28757
rect 67179 28708 67180 28748
rect 67220 28708 67221 28748
rect 67179 28699 67221 28708
rect 66891 28580 66933 28589
rect 66891 28540 66892 28580
rect 66932 28540 66933 28580
rect 66891 28531 66933 28540
rect 66507 27992 66549 28001
rect 66412 27952 66508 27992
rect 66548 27952 66549 27992
rect 66507 27943 66549 27952
rect 66315 27908 66357 27917
rect 66315 27868 66316 27908
rect 66356 27868 66357 27908
rect 66315 27859 66357 27868
rect 66508 27656 66548 27943
rect 66508 27607 66548 27616
rect 66603 27404 66645 27413
rect 66603 27364 66604 27404
rect 66644 27364 66645 27404
rect 66603 27355 66645 27364
rect 66508 26144 66548 26153
rect 66508 26069 66548 26104
rect 66507 26060 66549 26069
rect 66507 26020 66508 26060
rect 66548 26020 66549 26060
rect 66507 26011 66549 26020
rect 66220 25600 66452 25640
rect 65932 25423 65972 25432
rect 66316 25472 66356 25481
rect 65836 25388 65876 25423
rect 65836 25337 65876 25348
rect 66028 25388 66068 25397
rect 65740 25304 65780 25315
rect 65740 25229 65780 25264
rect 65739 25220 65781 25229
rect 65739 25180 65740 25220
rect 65780 25180 65781 25220
rect 65739 25171 65781 25180
rect 66028 25136 66068 25348
rect 66124 25313 66164 25398
rect 66123 25304 66165 25313
rect 66123 25264 66124 25304
rect 66164 25264 66165 25304
rect 66123 25255 66165 25264
rect 66316 25136 66356 25432
rect 66028 25096 66356 25136
rect 65740 24548 65780 24557
rect 65740 23801 65780 24508
rect 65931 24548 65973 24557
rect 65931 24508 65932 24548
rect 65972 24508 65973 24548
rect 65931 24499 65973 24508
rect 65932 23885 65972 24499
rect 66027 23960 66069 23969
rect 66027 23920 66028 23960
rect 66068 23920 66069 23960
rect 66027 23911 66069 23920
rect 65931 23876 65973 23885
rect 65931 23836 65932 23876
rect 65972 23836 65973 23876
rect 65931 23827 65973 23836
rect 65739 23792 65781 23801
rect 65739 23752 65740 23792
rect 65780 23752 65781 23792
rect 65739 23743 65781 23752
rect 65932 23792 65972 23827
rect 65740 23465 65780 23743
rect 65932 23742 65972 23752
rect 66028 23792 66068 23911
rect 66028 23743 66068 23752
rect 66124 23792 66164 25096
rect 66412 24557 66452 25600
rect 66411 24548 66453 24557
rect 66411 24508 66412 24548
rect 66452 24508 66453 24548
rect 66411 24499 66453 24508
rect 66508 23792 66548 26011
rect 66604 25565 66644 27355
rect 66603 25556 66645 25565
rect 66603 25516 66604 25556
rect 66644 25516 66645 25556
rect 66603 25507 66645 25516
rect 66699 25388 66741 25397
rect 66699 25348 66700 25388
rect 66740 25348 66741 25388
rect 66699 25339 66741 25348
rect 66604 25304 66644 25313
rect 66604 24473 66644 25264
rect 66700 25304 66740 25339
rect 66700 25253 66740 25264
rect 66795 25304 66837 25313
rect 66795 25264 66796 25304
rect 66836 25264 66837 25304
rect 66795 25255 66837 25264
rect 66796 25132 66836 25255
rect 66796 25083 66836 25092
rect 66892 24968 66932 28531
rect 66987 28412 67029 28421
rect 66987 28372 66988 28412
rect 67028 28372 67029 28412
rect 66987 28363 67029 28372
rect 66988 24977 67028 28363
rect 67180 28328 67220 28699
rect 67220 28288 67412 28328
rect 67180 28279 67220 28288
rect 67372 26144 67412 28288
rect 67372 26095 67412 26104
rect 67180 25481 67220 25566
rect 67179 25472 67221 25481
rect 67179 25432 67180 25472
rect 67220 25432 67221 25472
rect 67179 25423 67221 25432
rect 67275 25388 67317 25397
rect 67275 25348 67276 25388
rect 67316 25348 67317 25388
rect 67275 25339 67317 25348
rect 67179 25304 67221 25313
rect 67179 25264 67180 25304
rect 67220 25264 67221 25304
rect 67179 25255 67221 25264
rect 67180 25170 67220 25255
rect 66700 24928 66932 24968
rect 66987 24968 67029 24977
rect 66987 24928 66988 24968
rect 67028 24928 67029 24968
rect 66603 24464 66645 24473
rect 66603 24424 66604 24464
rect 66644 24424 66645 24464
rect 66603 24415 66645 24424
rect 66700 24212 66740 24928
rect 66987 24919 67029 24928
rect 66988 24632 67028 24641
rect 66988 24473 67028 24592
rect 67084 24632 67124 24643
rect 67084 24557 67124 24592
rect 67180 24632 67220 24641
rect 67083 24548 67125 24557
rect 67083 24508 67084 24548
rect 67124 24508 67125 24548
rect 67083 24499 67125 24508
rect 66987 24464 67029 24473
rect 66987 24424 66988 24464
rect 67028 24424 67029 24464
rect 66987 24415 67029 24424
rect 66700 24172 66932 24212
rect 66796 23792 66836 23801
rect 66508 23752 66796 23792
rect 66124 23743 66164 23752
rect 66796 23743 66836 23752
rect 66220 23708 66260 23717
rect 66412 23708 66452 23717
rect 66260 23668 66412 23708
rect 66220 23659 66260 23668
rect 66412 23659 66452 23668
rect 65739 23456 65781 23465
rect 65739 23416 65740 23456
rect 65780 23416 65781 23456
rect 65739 23407 65781 23416
rect 66027 23204 66069 23213
rect 66027 23164 66028 23204
rect 66068 23164 66069 23204
rect 66027 23155 66069 23164
rect 66028 23060 66068 23155
rect 66892 23060 66932 24172
rect 67180 24053 67220 24592
rect 67276 24632 67316 25339
rect 67372 25304 67412 25313
rect 67372 25145 67412 25264
rect 67467 25304 67509 25313
rect 67467 25264 67468 25304
rect 67508 25264 67509 25304
rect 67467 25255 67509 25264
rect 67468 25170 67508 25255
rect 67564 25229 67604 30472
rect 67563 25220 67605 25229
rect 67563 25180 67564 25220
rect 67604 25180 67605 25220
rect 67563 25171 67605 25180
rect 67371 25136 67413 25145
rect 67371 25096 67372 25136
rect 67412 25096 67413 25136
rect 67371 25087 67413 25096
rect 67660 25052 67700 32227
rect 68236 32108 68276 34999
rect 68331 34712 68373 34721
rect 68331 34672 68332 34712
rect 68372 34672 68373 34712
rect 68331 34663 68373 34672
rect 67852 32068 68276 32108
rect 67755 31940 67797 31949
rect 67755 31900 67756 31940
rect 67796 31900 67797 31940
rect 67755 31891 67797 31900
rect 67756 27329 67796 31891
rect 67755 27320 67797 27329
rect 67755 27280 67756 27320
rect 67796 27280 67797 27320
rect 67755 27271 67797 27280
rect 67468 25012 67700 25052
rect 67371 24968 67413 24977
rect 67371 24928 67372 24968
rect 67412 24928 67413 24968
rect 67371 24919 67413 24928
rect 67276 24583 67316 24592
rect 67275 24464 67317 24473
rect 67275 24424 67276 24464
rect 67316 24424 67317 24464
rect 67275 24415 67317 24424
rect 67276 24305 67316 24415
rect 67275 24296 67317 24305
rect 67275 24256 67276 24296
rect 67316 24256 67317 24296
rect 67275 24247 67317 24256
rect 67179 24044 67221 24053
rect 67179 24004 67180 24044
rect 67220 24004 67221 24044
rect 67179 23995 67221 24004
rect 67372 23060 67412 24919
rect 67468 23297 67508 25012
rect 67659 24632 67701 24641
rect 67659 24592 67660 24632
rect 67700 24592 67701 24632
rect 67659 24583 67701 24592
rect 67563 24128 67605 24137
rect 67563 24088 67564 24128
rect 67604 24088 67605 24128
rect 67563 24079 67605 24088
rect 67467 23288 67509 23297
rect 67467 23248 67468 23288
rect 67508 23248 67509 23288
rect 67467 23239 67509 23248
rect 65644 23020 65695 23060
rect 66028 23020 66095 23060
rect 66892 23020 67185 23060
rect 65255 22596 65295 22987
rect 65545 22596 65585 23020
rect 65655 22596 65695 23020
rect 65944 22952 65986 22961
rect 65944 22912 65945 22952
rect 65985 22912 65986 22952
rect 65944 22903 65986 22912
rect 65945 22596 65985 22903
rect 66055 22596 66095 23020
rect 66744 22952 66786 22961
rect 66744 22912 66745 22952
rect 66785 22912 66786 22952
rect 66744 22903 66786 22912
rect 66454 22868 66496 22877
rect 66454 22828 66455 22868
rect 66495 22828 66496 22868
rect 66454 22819 66496 22828
rect 66344 22784 66386 22793
rect 66344 22744 66345 22784
rect 66385 22744 66386 22784
rect 66344 22735 66386 22744
rect 66345 22596 66385 22735
rect 66455 22596 66495 22819
rect 66745 22596 66785 22903
rect 66854 22868 66896 22877
rect 66854 22828 66855 22868
rect 66895 22828 66896 22868
rect 66854 22819 66896 22828
rect 66855 22596 66895 22819
rect 67145 22596 67185 23020
rect 67276 23020 67412 23060
rect 67276 22784 67316 23020
rect 67564 22784 67604 24079
rect 67660 23792 67700 24583
rect 67660 23743 67700 23752
rect 67852 23549 67892 32068
rect 68332 32024 68372 34663
rect 68428 34637 68468 37435
rect 68524 36728 68564 36737
rect 68524 35897 68564 36688
rect 68620 36728 68660 36737
rect 68523 35888 68565 35897
rect 68523 35848 68524 35888
rect 68564 35848 68565 35888
rect 68523 35839 68565 35848
rect 68620 35813 68660 36688
rect 68619 35804 68661 35813
rect 68619 35764 68620 35804
rect 68660 35764 68661 35804
rect 68619 35755 68661 35764
rect 68716 35300 68756 38200
rect 69580 38240 69620 38359
rect 69580 38081 69620 38200
rect 69579 38072 69621 38081
rect 69579 38032 69580 38072
rect 69620 38032 69621 38072
rect 69579 38023 69621 38032
rect 69387 37568 69429 37577
rect 69387 37528 69388 37568
rect 69428 37528 69429 37568
rect 69387 37519 69429 37528
rect 68907 37400 68949 37409
rect 68907 37360 68908 37400
rect 68948 37360 68949 37400
rect 68907 37351 68949 37360
rect 68908 37266 68948 37351
rect 69003 37232 69045 37241
rect 69003 37192 69004 37232
rect 69044 37192 69045 37232
rect 69003 37183 69045 37192
rect 69004 36737 69044 37183
rect 69388 36896 69428 37519
rect 69772 37400 69812 37411
rect 69772 37325 69812 37360
rect 69771 37316 69813 37325
rect 69771 37276 69772 37316
rect 69812 37276 69813 37316
rect 69771 37267 69813 37276
rect 69868 36905 69908 38368
rect 69964 38240 70004 38249
rect 69388 36847 69428 36856
rect 69867 36896 69909 36905
rect 69867 36856 69868 36896
rect 69908 36856 69909 36896
rect 69867 36847 69909 36856
rect 68811 36728 68853 36737
rect 68811 36688 68812 36728
rect 68852 36688 68853 36728
rect 68811 36679 68853 36688
rect 68908 36728 68948 36737
rect 68812 36594 68852 36679
rect 68811 35720 68853 35729
rect 68811 35680 68812 35720
rect 68852 35680 68853 35720
rect 68811 35671 68853 35680
rect 68812 35586 68852 35671
rect 68524 35260 68756 35300
rect 68427 34628 68469 34637
rect 68427 34588 68428 34628
rect 68468 34588 68469 34628
rect 68427 34579 68469 34588
rect 68427 33284 68469 33293
rect 68427 33244 68428 33284
rect 68468 33244 68469 33284
rect 68427 33235 68469 33244
rect 68428 32360 68468 33235
rect 68428 32311 68468 32320
rect 68044 31984 68372 32024
rect 67947 31352 67989 31361
rect 67947 31312 67948 31352
rect 67988 31312 67989 31352
rect 67947 31303 67989 31312
rect 67948 31218 67988 31303
rect 68044 30512 68084 31984
rect 68428 31940 68468 31949
rect 68332 31900 68428 31940
rect 68139 31856 68181 31865
rect 68139 31816 68140 31856
rect 68180 31816 68181 31856
rect 68139 31807 68181 31816
rect 68140 30680 68180 31807
rect 68235 31604 68277 31613
rect 68235 31564 68236 31604
rect 68276 31564 68277 31604
rect 68235 31555 68277 31564
rect 68236 31193 68276 31555
rect 68235 31184 68277 31193
rect 68235 31144 68236 31184
rect 68276 31144 68277 31184
rect 68235 31135 68277 31144
rect 68140 30631 68180 30640
rect 68235 30680 68277 30689
rect 68235 30640 68236 30680
rect 68276 30640 68277 30680
rect 68235 30631 68277 30640
rect 68332 30680 68372 31900
rect 68428 31891 68468 31900
rect 68427 31772 68469 31781
rect 68427 31732 68428 31772
rect 68468 31732 68469 31772
rect 68427 31723 68469 31732
rect 68428 30848 68468 31723
rect 68524 31352 68564 35260
rect 68908 35132 68948 36688
rect 69003 36728 69045 36737
rect 69003 36688 69004 36728
rect 69044 36688 69045 36728
rect 69003 36679 69045 36688
rect 69100 36728 69140 36737
rect 69004 36594 69044 36679
rect 69003 36056 69045 36065
rect 69003 36016 69004 36056
rect 69044 36016 69045 36056
rect 69003 36007 69045 36016
rect 68716 35092 68948 35132
rect 68619 34376 68661 34385
rect 68619 34336 68620 34376
rect 68660 34336 68661 34376
rect 68619 34327 68661 34336
rect 68716 34376 68756 35092
rect 68907 34544 68949 34553
rect 68907 34504 68908 34544
rect 68948 34504 68949 34544
rect 68907 34495 68949 34504
rect 68620 34242 68660 34327
rect 68716 33293 68756 34336
rect 68811 34376 68853 34385
rect 68811 34336 68812 34376
rect 68852 34336 68853 34376
rect 68811 34327 68853 34336
rect 68908 34376 68948 34495
rect 68908 34327 68948 34336
rect 68812 34242 68852 34327
rect 68811 34124 68853 34133
rect 68811 34084 68812 34124
rect 68852 34084 68853 34124
rect 68811 34075 68853 34084
rect 68715 33284 68757 33293
rect 68715 33244 68716 33284
rect 68756 33244 68757 33284
rect 68715 33235 68757 33244
rect 68812 32360 68852 34075
rect 69004 33704 69044 36007
rect 69100 35813 69140 36688
rect 69291 36728 69333 36737
rect 69291 36688 69292 36728
rect 69332 36688 69333 36728
rect 69291 36679 69333 36688
rect 69099 35804 69141 35813
rect 69099 35764 69100 35804
rect 69140 35764 69141 35804
rect 69099 35755 69141 35764
rect 69099 34964 69141 34973
rect 69099 34924 69100 34964
rect 69140 34924 69141 34964
rect 69099 34915 69141 34924
rect 69100 34830 69140 34915
rect 69099 34628 69141 34637
rect 69099 34588 69100 34628
rect 69140 34588 69141 34628
rect 69099 34579 69141 34588
rect 69004 33655 69044 33664
rect 69100 33140 69140 34579
rect 68620 32320 68812 32360
rect 68620 32108 68660 32320
rect 68812 32311 68852 32320
rect 68908 33100 69140 33140
rect 69292 33140 69332 36679
rect 69580 36476 69620 36485
rect 69580 35897 69620 36436
rect 69579 35888 69621 35897
rect 69579 35848 69580 35888
rect 69620 35848 69621 35888
rect 69579 35839 69621 35848
rect 69964 35636 70004 38200
rect 70060 38240 70100 38249
rect 70060 37577 70100 38200
rect 70156 38240 70196 38368
rect 74188 38368 74420 38408
rect 70156 38191 70196 38200
rect 70252 38240 70292 38249
rect 70059 37568 70101 37577
rect 70059 37528 70060 37568
rect 70100 37528 70101 37568
rect 70059 37519 70101 37528
rect 69868 35596 70004 35636
rect 69771 35468 69813 35477
rect 69771 35428 69772 35468
rect 69812 35428 69813 35468
rect 69771 35419 69813 35428
rect 69675 34376 69717 34385
rect 69675 34336 69676 34376
rect 69716 34336 69717 34376
rect 69675 34327 69717 34336
rect 69580 34208 69620 34217
rect 69580 33629 69620 34168
rect 69579 33620 69621 33629
rect 69579 33580 69580 33620
rect 69620 33580 69621 33620
rect 69579 33571 69621 33580
rect 69580 33140 69620 33571
rect 69292 33100 69428 33140
rect 68620 32059 68660 32068
rect 68812 31352 68852 31361
rect 68524 31312 68812 31352
rect 68523 31184 68565 31193
rect 68523 31144 68524 31184
rect 68564 31144 68565 31184
rect 68523 31135 68565 31144
rect 68428 30799 68468 30808
rect 68332 30631 68372 30640
rect 68236 30546 68276 30631
rect 68044 30472 68180 30512
rect 67948 29840 67988 29849
rect 67948 28757 67988 29800
rect 67947 28748 67989 28757
rect 67947 28708 67948 28748
rect 67988 28708 67989 28748
rect 67947 28699 67989 28708
rect 68043 26648 68085 26657
rect 68043 26608 68044 26648
rect 68084 26608 68085 26648
rect 68043 26599 68085 26608
rect 68044 26514 68084 26599
rect 68140 24305 68180 30472
rect 68427 28916 68469 28925
rect 68427 28876 68428 28916
rect 68468 28876 68469 28916
rect 68427 28867 68469 28876
rect 68428 28782 68468 28867
rect 68332 28160 68372 28169
rect 68332 28001 68372 28120
rect 68331 27992 68373 28001
rect 68331 27952 68332 27992
rect 68372 27952 68373 27992
rect 68331 27943 68373 27952
rect 68427 27572 68469 27581
rect 68427 27532 68428 27572
rect 68468 27532 68469 27572
rect 68427 27523 68469 27532
rect 68428 27438 68468 27523
rect 68524 27245 68564 31135
rect 68619 31100 68661 31109
rect 68619 31060 68620 31100
rect 68660 31060 68661 31100
rect 68619 31051 68661 31060
rect 68523 27236 68565 27245
rect 68523 27196 68524 27236
rect 68564 27196 68565 27236
rect 68523 27187 68565 27196
rect 68620 27068 68660 31051
rect 68812 28757 68852 31312
rect 68811 28748 68853 28757
rect 68811 28708 68812 28748
rect 68852 28708 68853 28748
rect 68811 28699 68853 28708
rect 68908 28412 68948 33100
rect 69004 32108 69044 32117
rect 69004 31109 69044 32068
rect 69099 31268 69141 31277
rect 69099 31228 69100 31268
rect 69140 31228 69141 31268
rect 69099 31219 69141 31228
rect 69003 31100 69045 31109
rect 69003 31060 69004 31100
rect 69044 31060 69045 31100
rect 69003 31051 69045 31060
rect 69100 30848 69140 31219
rect 69100 30799 69140 30808
rect 69003 30680 69045 30689
rect 69003 30640 69004 30680
rect 69044 30640 69045 30680
rect 69003 30631 69045 30640
rect 69004 30546 69044 30631
rect 69100 30428 69140 30437
rect 69100 29840 69140 30388
rect 69291 30428 69333 30437
rect 69291 30388 69292 30428
rect 69332 30388 69333 30428
rect 69291 30379 69333 30388
rect 69292 30294 69332 30379
rect 69100 29800 69332 29840
rect 69100 29672 69140 29681
rect 69100 29513 69140 29632
rect 69099 29504 69141 29513
rect 69099 29464 69100 29504
rect 69140 29464 69141 29504
rect 69099 29455 69141 29464
rect 69100 29177 69140 29455
rect 69195 29420 69237 29429
rect 69195 29380 69196 29420
rect 69236 29380 69237 29420
rect 69195 29371 69237 29380
rect 69099 29168 69141 29177
rect 69099 29128 69100 29168
rect 69140 29128 69141 29168
rect 69099 29119 69141 29128
rect 69100 28412 69140 28421
rect 68908 28372 69100 28412
rect 68907 28160 68949 28169
rect 68907 28120 68908 28160
rect 68948 28120 68949 28160
rect 68907 28111 68949 28120
rect 68908 28026 68948 28111
rect 69100 28085 69140 28372
rect 69099 28076 69141 28085
rect 69099 28036 69100 28076
rect 69140 28036 69141 28076
rect 69099 28027 69141 28036
rect 69196 27908 69236 29371
rect 69100 27868 69236 27908
rect 69100 27329 69140 27868
rect 69195 27656 69237 27665
rect 69195 27616 69196 27656
rect 69236 27616 69237 27656
rect 69195 27607 69237 27616
rect 69099 27320 69141 27329
rect 69099 27280 69100 27320
rect 69140 27280 69141 27320
rect 69099 27271 69141 27280
rect 68428 27028 68660 27068
rect 68428 25061 68468 27028
rect 69196 26816 69236 27607
rect 69196 26767 69236 26776
rect 69292 26321 69332 29800
rect 69291 26312 69333 26321
rect 69291 26272 69292 26312
rect 69332 26272 69333 26312
rect 69291 26263 69333 26272
rect 69195 26228 69237 26237
rect 69195 26188 69196 26228
rect 69236 26188 69237 26228
rect 69195 26179 69237 26188
rect 68812 26144 68852 26153
rect 68524 25892 68564 25901
rect 68524 25313 68564 25852
rect 68812 25565 68852 26104
rect 69003 26144 69045 26153
rect 69003 26104 69004 26144
rect 69044 26104 69045 26144
rect 69003 26095 69045 26104
rect 69196 26144 69236 26179
rect 69388 26153 69428 33100
rect 69484 33100 69620 33140
rect 69484 27404 69524 33100
rect 69580 29168 69620 29177
rect 69580 28757 69620 29128
rect 69579 28748 69621 28757
rect 69579 28708 69580 28748
rect 69620 28708 69621 28748
rect 69579 28699 69621 28708
rect 69580 27665 69620 28699
rect 69579 27656 69621 27665
rect 69579 27616 69580 27656
rect 69620 27616 69621 27656
rect 69579 27607 69621 27616
rect 69580 27522 69620 27607
rect 69484 27364 69620 27404
rect 69483 26228 69525 26237
rect 69483 26188 69484 26228
rect 69524 26188 69525 26228
rect 69483 26179 69525 26188
rect 68908 26060 68948 26069
rect 68716 25556 68756 25565
rect 68811 25556 68853 25565
rect 68756 25516 68812 25556
rect 68852 25516 68853 25556
rect 68716 25507 68756 25516
rect 68811 25507 68853 25516
rect 68812 25422 68852 25507
rect 68908 25472 68948 26020
rect 69004 25976 69044 26095
rect 69196 26093 69236 26104
rect 69387 26144 69429 26153
rect 69387 26104 69388 26144
rect 69428 26104 69429 26144
rect 69387 26095 69429 26104
rect 69484 26144 69524 26179
rect 69484 26093 69524 26104
rect 69580 26069 69620 27364
rect 69676 26573 69716 34327
rect 69772 34040 69812 35419
rect 69868 34217 69908 35596
rect 69867 34208 69909 34217
rect 69867 34168 69868 34208
rect 69908 34168 69909 34208
rect 69867 34159 69909 34168
rect 69772 34000 69908 34040
rect 69771 32780 69813 32789
rect 69771 32740 69772 32780
rect 69812 32740 69813 32780
rect 69771 32731 69813 32740
rect 69772 32646 69812 32731
rect 69771 31856 69813 31865
rect 69771 31816 69772 31856
rect 69812 31816 69813 31856
rect 69771 31807 69813 31816
rect 69772 27329 69812 31807
rect 69771 27320 69813 27329
rect 69771 27280 69772 27320
rect 69812 27280 69813 27320
rect 69771 27271 69813 27280
rect 69771 26648 69813 26657
rect 69771 26608 69772 26648
rect 69812 26608 69813 26648
rect 69771 26599 69813 26608
rect 69675 26564 69717 26573
rect 69675 26524 69676 26564
rect 69716 26524 69717 26564
rect 69675 26515 69717 26524
rect 69675 26312 69717 26321
rect 69675 26272 69676 26312
rect 69716 26272 69717 26312
rect 69675 26263 69717 26272
rect 69676 26144 69716 26263
rect 69772 26153 69812 26599
rect 69100 26060 69140 26069
rect 69100 25976 69140 26020
rect 69579 26060 69621 26069
rect 69579 26020 69580 26060
rect 69620 26020 69621 26060
rect 69579 26011 69621 26020
rect 69484 25976 69524 25985
rect 69100 25936 69484 25976
rect 69004 25927 69044 25936
rect 69484 25927 69524 25936
rect 69676 25733 69716 26104
rect 69771 26144 69813 26153
rect 69771 26104 69772 26144
rect 69812 26104 69813 26144
rect 69771 26095 69813 26104
rect 69772 26010 69812 26095
rect 69868 25985 69908 34000
rect 70060 33032 70100 37519
rect 70156 37400 70196 37409
rect 70252 37400 70292 38200
rect 73996 38240 74036 38249
rect 74188 38240 74228 38368
rect 74036 38200 74132 38240
rect 73996 38191 74036 38200
rect 70196 37360 70292 37400
rect 70444 38156 70484 38165
rect 70156 37351 70196 37360
rect 70347 37232 70389 37241
rect 70347 37192 70348 37232
rect 70388 37192 70389 37232
rect 70347 37183 70389 37192
rect 70348 37098 70388 37183
rect 70444 37157 70484 38116
rect 71020 38156 71060 38165
rect 70636 37988 70676 37997
rect 70636 37493 70676 37948
rect 70828 37988 70868 37997
rect 70635 37484 70677 37493
rect 70635 37444 70636 37484
rect 70676 37444 70677 37484
rect 70635 37435 70677 37444
rect 70731 37400 70773 37409
rect 70731 37360 70732 37400
rect 70772 37360 70773 37400
rect 70731 37351 70773 37360
rect 70443 37148 70485 37157
rect 70443 37108 70444 37148
rect 70484 37108 70485 37148
rect 70443 37099 70485 37108
rect 70732 36737 70772 37351
rect 70251 36728 70293 36737
rect 70251 36688 70252 36728
rect 70292 36688 70293 36728
rect 70251 36679 70293 36688
rect 70731 36728 70773 36737
rect 70731 36688 70732 36728
rect 70772 36688 70773 36728
rect 70731 36679 70773 36688
rect 70252 36065 70292 36679
rect 70732 36594 70772 36679
rect 70828 36653 70868 37948
rect 71020 37325 71060 38116
rect 73996 37988 74036 37997
rect 73708 37948 73996 37988
rect 73132 37568 73172 37577
rect 71500 37400 71540 37409
rect 71019 37316 71061 37325
rect 71019 37276 71020 37316
rect 71060 37276 71061 37316
rect 71019 37267 71061 37276
rect 71020 36821 71060 37267
rect 71019 36812 71061 36821
rect 71019 36772 71020 36812
rect 71060 36772 71061 36812
rect 71019 36763 71061 36772
rect 71500 36737 71540 37360
rect 71595 37400 71637 37409
rect 71595 37360 71596 37400
rect 71636 37360 71637 37400
rect 71595 37351 71637 37360
rect 72363 37400 72405 37409
rect 72363 37360 72364 37400
rect 72404 37360 72405 37400
rect 72363 37351 72405 37360
rect 71499 36728 71541 36737
rect 71499 36688 71500 36728
rect 71540 36688 71541 36728
rect 71499 36679 71541 36688
rect 71596 36728 71636 37351
rect 72364 37266 72404 37351
rect 72748 37316 72788 37325
rect 72748 36989 72788 37276
rect 73035 37232 73077 37241
rect 73035 37192 73036 37232
rect 73076 37192 73077 37232
rect 73035 37183 73077 37192
rect 72747 36980 72789 36989
rect 72747 36940 72748 36980
rect 72788 36940 72789 36980
rect 72747 36931 72789 36940
rect 72268 36856 72692 36896
rect 71596 36653 71636 36688
rect 71980 36728 72020 36737
rect 70827 36644 70869 36653
rect 70827 36604 70828 36644
rect 70868 36604 70869 36644
rect 70827 36595 70869 36604
rect 71115 36644 71157 36653
rect 71115 36604 71116 36644
rect 71156 36604 71157 36644
rect 71115 36595 71157 36604
rect 71595 36644 71637 36653
rect 71595 36604 71596 36644
rect 71636 36604 71637 36644
rect 71595 36595 71637 36604
rect 70251 36056 70293 36065
rect 70251 36016 70252 36056
rect 70292 36016 70293 36056
rect 70251 36007 70293 36016
rect 70252 35216 70292 36007
rect 71116 35384 71156 36595
rect 71403 36560 71445 36569
rect 71403 36520 71404 36560
rect 71444 36520 71445 36560
rect 71403 36511 71445 36520
rect 71307 35888 71349 35897
rect 71307 35848 71308 35888
rect 71348 35848 71349 35888
rect 71307 35839 71349 35848
rect 71404 35888 71444 36511
rect 71980 36476 72020 36688
rect 72171 36728 72213 36737
rect 72171 36688 72172 36728
rect 72212 36688 72213 36728
rect 72171 36679 72213 36688
rect 72172 36594 72212 36679
rect 72268 36644 72308 36856
rect 72556 36728 72596 36737
rect 72268 36595 72308 36604
rect 72460 36644 72500 36653
rect 72364 36560 72404 36569
rect 72364 36476 72404 36520
rect 71980 36436 72404 36476
rect 72460 36401 72500 36604
rect 72459 36392 72501 36401
rect 72459 36352 72460 36392
rect 72500 36352 72501 36392
rect 72459 36343 72501 36352
rect 72556 36224 72596 36688
rect 72652 36560 72692 36856
rect 72748 36737 72788 36822
rect 73036 36737 73076 37183
rect 72747 36728 72789 36737
rect 72940 36728 72980 36737
rect 72747 36688 72748 36728
rect 72788 36688 72884 36728
rect 72747 36679 72789 36688
rect 72748 36560 72788 36569
rect 72652 36520 72748 36560
rect 72748 36511 72788 36520
rect 72172 36184 72596 36224
rect 72172 36140 72212 36184
rect 72172 36091 72212 36100
rect 71595 35972 71637 35981
rect 71595 35932 71596 35972
rect 71636 35932 71637 35972
rect 71595 35923 71637 35932
rect 72267 35972 72309 35981
rect 72267 35932 72268 35972
rect 72308 35932 72309 35972
rect 72267 35923 72309 35932
rect 71308 35754 71348 35839
rect 70252 35167 70292 35176
rect 70828 35344 71156 35384
rect 70155 34376 70197 34385
rect 70155 34336 70156 34376
rect 70196 34336 70197 34376
rect 70155 34327 70197 34336
rect 70156 33872 70196 34327
rect 70156 33823 70196 33832
rect 70060 32992 70484 33032
rect 70155 32864 70197 32873
rect 70155 32824 70156 32864
rect 70196 32824 70197 32864
rect 70155 32815 70197 32824
rect 70156 31361 70196 32815
rect 70444 31520 70484 32992
rect 70828 32873 70868 35344
rect 71019 35216 71061 35225
rect 71019 35176 71020 35216
rect 71060 35176 71061 35216
rect 71019 35167 71061 35176
rect 71116 35216 71156 35344
rect 71116 35167 71156 35176
rect 70923 34964 70965 34973
rect 70923 34924 70924 34964
rect 70964 34924 70965 34964
rect 70923 34915 70965 34924
rect 70924 34376 70964 34915
rect 71020 34628 71060 35167
rect 71404 34628 71444 35848
rect 71596 35888 71636 35923
rect 71596 35837 71636 35848
rect 72075 35888 72117 35897
rect 72075 35848 72076 35888
rect 72116 35848 72117 35888
rect 72075 35839 72117 35848
rect 72076 35754 72116 35839
rect 71500 35720 71540 35729
rect 71540 35680 71828 35720
rect 71500 35671 71540 35680
rect 71691 35384 71733 35393
rect 71691 35344 71692 35384
rect 71732 35344 71733 35384
rect 71691 35335 71733 35344
rect 71500 35216 71540 35225
rect 71692 35216 71732 35335
rect 71500 35057 71540 35176
rect 71596 35176 71692 35216
rect 71499 35048 71541 35057
rect 71499 35008 71500 35048
rect 71540 35008 71541 35048
rect 71499 34999 71541 35008
rect 71060 34588 71252 34628
rect 71404 34588 71540 34628
rect 71020 34579 71060 34588
rect 70964 34336 71156 34376
rect 70924 34327 70964 34336
rect 71116 33704 71156 34336
rect 71212 34204 71252 34588
rect 71307 34544 71349 34553
rect 71307 34504 71308 34544
rect 71348 34504 71349 34544
rect 71307 34495 71349 34504
rect 71212 34155 71252 34164
rect 71308 34376 71348 34495
rect 71404 34385 71444 34470
rect 71308 33881 71348 34336
rect 71403 34376 71445 34385
rect 71403 34336 71404 34376
rect 71444 34336 71445 34376
rect 71403 34327 71445 34336
rect 71500 34208 71540 34588
rect 71404 34168 71540 34208
rect 71307 33872 71349 33881
rect 71307 33832 71308 33872
rect 71348 33832 71349 33872
rect 71307 33823 71349 33832
rect 71308 33704 71348 33713
rect 71116 33664 71308 33704
rect 71308 33655 71348 33664
rect 71404 33704 71444 34168
rect 71596 33704 71636 35176
rect 71692 35167 71732 35176
rect 71788 35132 71828 35680
rect 72075 35216 72117 35225
rect 72075 35176 72076 35216
rect 72116 35176 72117 35216
rect 72075 35167 72117 35176
rect 71788 35083 71828 35092
rect 71980 35132 72020 35141
rect 71883 35048 71925 35057
rect 71883 35008 71884 35048
rect 71924 35008 71925 35048
rect 71883 34999 71925 35008
rect 71884 34914 71924 34999
rect 71692 34544 71732 34553
rect 71980 34544 72020 35092
rect 72076 35082 72116 35167
rect 72171 35132 72213 35141
rect 72171 35092 72172 35132
rect 72212 35092 72213 35132
rect 72171 35083 72213 35092
rect 71732 34504 72020 34544
rect 71692 34495 71732 34504
rect 71787 34376 71829 34385
rect 71787 34336 71788 34376
rect 71828 34336 71829 34376
rect 71787 34327 71829 34336
rect 71980 34376 72020 34504
rect 71980 34327 72020 34336
rect 72075 34376 72117 34385
rect 72075 34336 72076 34376
rect 72116 34336 72117 34376
rect 72075 34327 72117 34336
rect 72172 34376 72212 35083
rect 71788 33872 71828 34327
rect 71883 34292 71925 34301
rect 71883 34252 71884 34292
rect 71924 34252 71925 34292
rect 71883 34243 71925 34252
rect 71884 34158 71924 34243
rect 72076 34242 72116 34327
rect 72172 34133 72212 34336
rect 72171 34124 72213 34133
rect 72171 34084 72172 34124
rect 72212 34084 72213 34124
rect 72171 34075 72213 34084
rect 71788 33823 71828 33832
rect 72075 33872 72117 33881
rect 72075 33832 72076 33872
rect 72116 33832 72117 33872
rect 72075 33823 72117 33832
rect 71404 33536 71444 33664
rect 71308 33496 71444 33536
rect 71500 33664 71596 33704
rect 70827 32864 70869 32873
rect 70827 32824 70828 32864
rect 70868 32824 70869 32864
rect 70827 32815 70869 32824
rect 71019 32864 71061 32873
rect 71019 32824 71020 32864
rect 71060 32824 71061 32864
rect 71019 32815 71061 32824
rect 71020 32730 71060 32815
rect 71308 31613 71348 33496
rect 71500 33140 71540 33664
rect 71596 33655 71636 33664
rect 71884 33704 71924 33713
rect 71404 33100 71540 33140
rect 71596 33452 71636 33461
rect 71404 31688 71444 33100
rect 71499 32192 71541 32201
rect 71499 32152 71500 32192
rect 71540 32152 71541 32192
rect 71499 32143 71541 32152
rect 71500 32058 71540 32143
rect 71596 32108 71636 33412
rect 71884 33293 71924 33664
rect 71979 33704 72021 33713
rect 71979 33664 71980 33704
rect 72020 33664 72021 33704
rect 71979 33655 72021 33664
rect 72076 33704 72116 33823
rect 72076 33655 72116 33664
rect 71980 33570 72020 33655
rect 71883 33284 71925 33293
rect 71883 33244 71884 33284
rect 71924 33244 71925 33284
rect 71883 33235 71925 33244
rect 72268 33140 72308 35923
rect 72460 35716 72500 36184
rect 72651 36056 72693 36065
rect 72651 36016 72652 36056
rect 72692 36016 72693 36056
rect 72651 36007 72693 36016
rect 72460 35667 72500 35676
rect 72556 35888 72596 35897
rect 72459 34880 72501 34889
rect 72459 34840 72460 34880
rect 72500 34840 72501 34880
rect 72459 34831 72501 34840
rect 72363 34292 72405 34301
rect 72363 34252 72364 34292
rect 72404 34252 72405 34292
rect 72363 34243 72405 34252
rect 72364 34158 72404 34243
rect 72460 34040 72500 34831
rect 72076 33100 72308 33140
rect 72364 34000 72500 34040
rect 71691 32780 71733 32789
rect 71691 32740 71692 32780
rect 71732 32740 71733 32780
rect 71691 32731 71733 32740
rect 71596 32059 71636 32068
rect 71692 32024 71732 32731
rect 71883 32612 71925 32621
rect 71883 32572 71884 32612
rect 71924 32572 71925 32612
rect 71883 32563 71925 32572
rect 71884 32192 71924 32563
rect 72076 32201 72116 33100
rect 72364 32789 72404 34000
rect 72459 33872 72501 33881
rect 72556 33872 72596 35848
rect 72652 35888 72692 36007
rect 72844 35981 72884 36688
rect 72940 36569 72980 36688
rect 73035 36728 73077 36737
rect 73035 36688 73036 36728
rect 73076 36688 73077 36728
rect 73035 36679 73077 36688
rect 73036 36594 73076 36679
rect 73132 36653 73172 37528
rect 73419 37400 73461 37409
rect 73419 37360 73420 37400
rect 73460 37360 73461 37400
rect 73419 37351 73461 37360
rect 73516 37400 73556 37409
rect 73420 37266 73460 37351
rect 73516 37157 73556 37360
rect 73612 37174 73652 37183
rect 73515 37148 73557 37157
rect 73515 37108 73516 37148
rect 73556 37108 73557 37148
rect 73515 37099 73557 37108
rect 73612 36896 73652 37134
rect 73708 37148 73748 37948
rect 73996 37939 74036 37948
rect 74092 37820 74132 38200
rect 74188 38191 74228 38200
rect 74284 38240 74324 38249
rect 73900 37780 74132 37820
rect 73804 37325 73844 37410
rect 73803 37316 73845 37325
rect 73803 37276 73804 37316
rect 73844 37276 73845 37316
rect 73803 37267 73845 37276
rect 73708 37108 73844 37148
rect 73516 36856 73652 36896
rect 73707 36896 73749 36905
rect 73707 36856 73708 36896
rect 73748 36856 73749 36896
rect 73324 36812 73364 36821
rect 73516 36812 73556 36856
rect 73707 36847 73749 36856
rect 73364 36772 73556 36812
rect 73324 36763 73364 36772
rect 73227 36728 73269 36737
rect 73227 36688 73228 36728
rect 73268 36688 73269 36728
rect 73227 36679 73269 36688
rect 73516 36728 73556 36772
rect 73516 36679 73556 36688
rect 73131 36644 73173 36653
rect 73131 36604 73132 36644
rect 73172 36604 73173 36644
rect 73131 36595 73173 36604
rect 73228 36594 73268 36679
rect 73611 36644 73653 36653
rect 73611 36604 73612 36644
rect 73652 36604 73653 36644
rect 73611 36595 73653 36604
rect 72939 36560 72981 36569
rect 72939 36520 72940 36560
rect 72980 36520 72981 36560
rect 72939 36511 72981 36520
rect 73515 36560 73557 36569
rect 73515 36520 73516 36560
rect 73556 36520 73557 36560
rect 73515 36511 73557 36520
rect 72939 36392 72981 36401
rect 72939 36352 72940 36392
rect 72980 36352 72981 36392
rect 72939 36343 72981 36352
rect 72940 36140 72980 36343
rect 72843 35972 72885 35981
rect 72843 35932 72844 35972
rect 72884 35932 72885 35972
rect 72843 35923 72885 35932
rect 72652 35839 72692 35848
rect 72843 35300 72885 35309
rect 72843 35260 72844 35300
rect 72884 35260 72885 35300
rect 72843 35251 72885 35260
rect 72844 35166 72884 35251
rect 72940 35216 72980 36100
rect 73516 35972 73556 36511
rect 73612 36510 73652 36595
rect 73708 36560 73748 36847
rect 73804 36644 73844 37108
rect 73804 36595 73844 36604
rect 73900 36728 73940 37780
rect 74188 37400 74228 37409
rect 74091 37316 74133 37325
rect 74091 37276 74092 37316
rect 74132 37276 74133 37316
rect 74091 37267 74133 37276
rect 73995 37148 74037 37157
rect 73995 37108 73996 37148
rect 74036 37108 74037 37148
rect 73995 37099 74037 37108
rect 73996 36728 74036 37099
rect 74092 36896 74132 37267
rect 74188 36905 74228 37360
rect 74284 37325 74324 38200
rect 74283 37316 74325 37325
rect 74283 37276 74284 37316
rect 74324 37276 74325 37316
rect 74283 37267 74325 37276
rect 74092 36847 74132 36856
rect 74187 36896 74229 36905
rect 74187 36856 74188 36896
rect 74228 36856 74229 36896
rect 74380 36896 74420 38368
rect 75915 38368 75916 38408
rect 75956 38368 75957 38408
rect 75915 38359 75957 38368
rect 74476 38240 74516 38249
rect 74476 37409 74516 38200
rect 74572 38240 74612 38249
rect 74475 37400 74517 37409
rect 74475 37360 74476 37400
rect 74516 37360 74517 37400
rect 74475 37351 74517 37360
rect 74572 37064 74612 38200
rect 74668 38240 74708 38249
rect 74668 37493 74708 38200
rect 74764 38240 74804 38249
rect 74667 37484 74709 37493
rect 74667 37444 74668 37484
rect 74708 37444 74709 37484
rect 74667 37435 74709 37444
rect 74764 37241 74804 38200
rect 75628 38240 75668 38249
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 75628 37661 75668 38200
rect 75916 38240 75956 38359
rect 75916 38191 75956 38200
rect 77260 38156 77300 38165
rect 77068 38116 77260 38156
rect 76204 37988 76244 37997
rect 76204 37661 76244 37948
rect 75051 37652 75093 37661
rect 75051 37612 75052 37652
rect 75092 37612 75093 37652
rect 75051 37603 75093 37612
rect 75627 37652 75669 37661
rect 75627 37612 75628 37652
rect 75668 37612 75669 37652
rect 75627 37603 75669 37612
rect 76203 37652 76245 37661
rect 76203 37612 76204 37652
rect 76244 37612 76245 37652
rect 76203 37603 76245 37612
rect 75052 37400 75092 37603
rect 75339 37484 75381 37493
rect 75339 37444 75340 37484
rect 75380 37444 75381 37484
rect 75339 37435 75381 37444
rect 74956 37360 75052 37400
rect 74763 37232 74805 37241
rect 74763 37192 74764 37232
rect 74804 37192 74805 37232
rect 74763 37183 74805 37192
rect 74572 37024 74900 37064
rect 74571 36896 74613 36905
rect 74380 36856 74516 36896
rect 74187 36847 74229 36856
rect 74188 36728 74228 36739
rect 73996 36688 74132 36728
rect 73708 36511 73748 36520
rect 73900 36392 73940 36688
rect 73708 36352 73940 36392
rect 73516 35932 73652 35972
rect 73515 35804 73557 35813
rect 73515 35764 73516 35804
rect 73556 35764 73557 35804
rect 73515 35755 73557 35764
rect 73323 35300 73365 35309
rect 73323 35260 73324 35300
rect 73364 35260 73365 35300
rect 73323 35251 73365 35260
rect 72940 35167 72980 35176
rect 73036 35216 73076 35225
rect 72747 34544 72789 34553
rect 72747 34504 72748 34544
rect 72788 34504 72789 34544
rect 72747 34495 72789 34504
rect 72651 34376 72693 34385
rect 72651 34336 72652 34376
rect 72692 34336 72693 34376
rect 72651 34327 72693 34336
rect 72748 34376 72788 34495
rect 72748 34327 72788 34336
rect 72459 33832 72460 33872
rect 72500 33832 72596 33872
rect 72652 33872 72692 34327
rect 72459 33823 72501 33832
rect 72652 33823 72692 33832
rect 72460 33032 72500 33823
rect 72555 33704 72597 33713
rect 72555 33664 72556 33704
rect 72596 33664 72597 33704
rect 72555 33655 72597 33664
rect 72556 33570 72596 33655
rect 73036 33461 73076 35176
rect 73131 35216 73173 35225
rect 73131 35176 73132 35216
rect 73172 35176 73173 35216
rect 73131 35167 73173 35176
rect 73132 35082 73172 35167
rect 73324 35166 73364 35251
rect 72651 33452 72693 33461
rect 72651 33412 72652 33452
rect 72692 33412 72693 33452
rect 72651 33403 72693 33412
rect 73035 33452 73077 33461
rect 73035 33412 73036 33452
rect 73076 33412 73077 33452
rect 73035 33403 73077 33412
rect 72652 33318 72692 33403
rect 73035 33284 73077 33293
rect 73516 33284 73556 35755
rect 73612 35216 73652 35932
rect 73708 35393 73748 36352
rect 73803 36056 73845 36065
rect 73803 36016 73804 36056
rect 73844 36016 73845 36056
rect 73803 36007 73845 36016
rect 73804 35888 73844 36007
rect 73899 35972 73941 35981
rect 73899 35932 73900 35972
rect 73940 35932 73941 35972
rect 73899 35923 73941 35932
rect 73804 35839 73844 35848
rect 73900 35888 73940 35923
rect 73900 35837 73940 35848
rect 73996 35888 74036 35897
rect 73996 35393 74036 35848
rect 74092 35888 74132 36688
rect 74188 36653 74228 36688
rect 74284 36728 74324 36737
rect 74187 36644 74229 36653
rect 74187 36604 74188 36644
rect 74228 36604 74229 36644
rect 74187 36595 74229 36604
rect 74284 36485 74324 36688
rect 74380 36728 74420 36737
rect 74283 36476 74325 36485
rect 74283 36436 74284 36476
rect 74324 36436 74325 36476
rect 74283 36427 74325 36436
rect 74380 36065 74420 36688
rect 74379 36056 74421 36065
rect 74379 36016 74380 36056
rect 74420 36016 74421 36056
rect 74379 36007 74421 36016
rect 74092 35729 74132 35848
rect 74284 35972 74324 35981
rect 74284 35813 74324 35932
rect 74476 35888 74516 36856
rect 74571 36856 74572 36896
rect 74612 36856 74613 36896
rect 74571 36847 74613 36856
rect 74572 36644 74612 36847
rect 74572 36595 74612 36604
rect 74763 36560 74805 36569
rect 74763 36520 74764 36560
rect 74804 36520 74805 36560
rect 74763 36511 74805 36520
rect 74764 36426 74804 36511
rect 74668 35972 74708 35983
rect 74860 35981 74900 37024
rect 74668 35897 74708 35932
rect 74859 35972 74901 35981
rect 74859 35932 74860 35972
rect 74900 35932 74901 35972
rect 74859 35923 74901 35932
rect 74380 35848 74516 35888
rect 74667 35888 74709 35897
rect 74667 35848 74668 35888
rect 74708 35848 74709 35888
rect 74283 35804 74325 35813
rect 74283 35764 74284 35804
rect 74324 35764 74325 35804
rect 74283 35755 74325 35764
rect 74091 35720 74133 35729
rect 74091 35680 74092 35720
rect 74132 35680 74133 35720
rect 74091 35671 74133 35680
rect 73707 35384 73749 35393
rect 73707 35344 73708 35384
rect 73748 35344 73749 35384
rect 73707 35335 73749 35344
rect 73995 35384 74037 35393
rect 73995 35344 73996 35384
rect 74036 35344 74037 35384
rect 73995 35335 74037 35344
rect 73708 35216 73748 35225
rect 73612 35176 73708 35216
rect 73612 34553 73652 35176
rect 73708 35167 73748 35176
rect 73611 34544 73653 34553
rect 73611 34504 73612 34544
rect 73652 34504 73653 34544
rect 73611 34495 73653 34504
rect 73611 34376 73653 34385
rect 73611 34336 73612 34376
rect 73652 34336 73653 34376
rect 73611 34327 73653 34336
rect 74091 34376 74133 34385
rect 74091 34336 74092 34376
rect 74132 34336 74133 34376
rect 74091 34327 74133 34336
rect 73612 34242 73652 34327
rect 73995 33368 74037 33377
rect 73995 33328 73996 33368
rect 74036 33328 74037 33368
rect 73995 33319 74037 33328
rect 73035 33244 73036 33284
rect 73076 33244 73077 33284
rect 73035 33235 73077 33244
rect 73420 33244 73556 33284
rect 72843 33032 72885 33041
rect 72460 32992 72788 33032
rect 72460 32864 72500 32992
rect 72460 32815 72500 32824
rect 72556 32864 72596 32873
rect 72363 32780 72405 32789
rect 72363 32740 72364 32780
rect 72404 32740 72405 32780
rect 72363 32731 72405 32740
rect 72172 32696 72212 32705
rect 72212 32656 72308 32696
rect 72172 32647 72212 32656
rect 72268 32360 72308 32656
rect 72364 32638 72404 32647
rect 72363 32572 72364 32621
rect 72404 32572 72405 32621
rect 72363 32563 72405 32572
rect 72364 32503 72404 32563
rect 72556 32537 72596 32824
rect 72651 32612 72693 32621
rect 72651 32572 72652 32612
rect 72692 32572 72693 32612
rect 72651 32563 72693 32572
rect 72555 32528 72597 32537
rect 72555 32488 72556 32528
rect 72596 32488 72597 32528
rect 72555 32479 72597 32488
rect 72652 32360 72692 32563
rect 72268 32320 72404 32360
rect 71884 32143 71924 32152
rect 72075 32192 72117 32201
rect 72268 32192 72308 32201
rect 72075 32152 72076 32192
rect 72116 32152 72212 32192
rect 72075 32143 72117 32152
rect 71787 32108 71829 32117
rect 71787 32068 71788 32108
rect 71828 32068 71829 32108
rect 71787 32059 71829 32068
rect 71692 31975 71732 31984
rect 71788 31974 71828 32059
rect 72076 32058 72116 32143
rect 72076 31940 72116 31949
rect 71404 31648 71540 31688
rect 71307 31604 71349 31613
rect 71307 31564 71308 31604
rect 71348 31564 71349 31604
rect 71307 31555 71349 31564
rect 70252 31480 70444 31520
rect 70155 31352 70197 31361
rect 70155 31312 70156 31352
rect 70196 31312 70197 31352
rect 70155 31303 70197 31312
rect 69964 31184 70004 31193
rect 69964 30689 70004 31144
rect 70156 30689 70196 31303
rect 69963 30680 70005 30689
rect 69963 30640 69964 30680
rect 70004 30640 70005 30680
rect 69963 30631 70005 30640
rect 70155 30680 70197 30689
rect 70155 30640 70156 30680
rect 70196 30640 70197 30680
rect 70155 30631 70197 30640
rect 69964 30353 70004 30631
rect 69963 30344 70005 30353
rect 69963 30304 69964 30344
rect 70004 30304 70005 30344
rect 69963 30295 70005 30304
rect 70155 28496 70197 28505
rect 70155 28456 70156 28496
rect 70196 28456 70197 28496
rect 70155 28447 70197 28456
rect 70059 28160 70101 28169
rect 70059 28120 70060 28160
rect 70100 28120 70101 28160
rect 70059 28111 70101 28120
rect 69963 27236 70005 27245
rect 69963 27196 69964 27236
rect 70004 27196 70005 27236
rect 69963 27187 70005 27196
rect 69964 26489 70004 27187
rect 70060 26825 70100 28111
rect 70059 26816 70101 26825
rect 70059 26776 70060 26816
rect 70100 26776 70101 26816
rect 70059 26767 70101 26776
rect 69963 26480 70005 26489
rect 69963 26440 69964 26480
rect 70004 26440 70005 26480
rect 69963 26431 70005 26440
rect 69964 26312 70004 26323
rect 69964 26237 70004 26272
rect 69963 26228 70005 26237
rect 69963 26188 69964 26228
rect 70004 26188 70005 26228
rect 69963 26179 70005 26188
rect 69867 25976 69909 25985
rect 69867 25936 69868 25976
rect 69908 25936 69909 25976
rect 69867 25927 69909 25936
rect 69675 25724 69717 25733
rect 69675 25684 69676 25724
rect 69716 25684 69717 25724
rect 69675 25675 69717 25684
rect 70060 25640 70100 26767
rect 70156 26405 70196 28447
rect 70155 26396 70197 26405
rect 70155 26356 70156 26396
rect 70196 26356 70197 26396
rect 70155 26347 70197 26356
rect 70156 26060 70196 26347
rect 70156 26011 70196 26020
rect 70252 25892 70292 31480
rect 70444 31471 70484 31480
rect 71403 31520 71445 31529
rect 71403 31480 71404 31520
rect 71444 31480 71445 31520
rect 71403 31471 71445 31480
rect 71404 31436 71444 31471
rect 71404 31385 71444 31396
rect 71308 30689 71348 30774
rect 70444 30680 70484 30689
rect 70348 30640 70444 30680
rect 70348 27665 70388 30640
rect 70444 30631 70484 30640
rect 70539 30680 70581 30689
rect 70539 30640 70540 30680
rect 70580 30640 70581 30680
rect 70539 30631 70581 30640
rect 71307 30680 71349 30689
rect 71307 30640 71308 30680
rect 71348 30640 71349 30680
rect 71307 30631 71349 30640
rect 70443 29252 70485 29261
rect 70540 29252 70580 30631
rect 71307 30512 71349 30521
rect 71307 30472 71308 30512
rect 71348 30472 71349 30512
rect 71307 30463 71349 30472
rect 71115 30260 71157 30269
rect 71115 30220 71116 30260
rect 71156 30220 71157 30260
rect 71115 30211 71157 30220
rect 70923 30092 70965 30101
rect 70923 30052 70924 30092
rect 70964 30052 70965 30092
rect 70923 30043 70965 30052
rect 70924 29958 70964 30043
rect 70732 29924 70772 29933
rect 70443 29212 70444 29252
rect 70484 29212 70580 29252
rect 70636 29884 70732 29924
rect 70443 29203 70485 29212
rect 70444 29168 70484 29203
rect 70444 29117 70484 29128
rect 70443 28916 70485 28925
rect 70443 28876 70444 28916
rect 70484 28876 70485 28916
rect 70443 28867 70485 28876
rect 70444 28328 70484 28867
rect 70539 28580 70581 28589
rect 70539 28540 70540 28580
rect 70580 28540 70581 28580
rect 70539 28531 70581 28540
rect 70540 28342 70580 28531
rect 70636 28505 70676 29884
rect 70732 29875 70772 29884
rect 71116 29840 71156 30211
rect 71116 29791 71156 29800
rect 71308 29840 71348 30463
rect 71403 30428 71445 30437
rect 71403 30388 71404 30428
rect 71444 30388 71445 30428
rect 71403 30379 71445 30388
rect 71308 29791 71348 29800
rect 71404 29840 71444 30379
rect 71500 30101 71540 31648
rect 71595 31604 71637 31613
rect 71595 31564 71596 31604
rect 71636 31564 71637 31604
rect 71595 31555 71637 31564
rect 71596 31470 71636 31555
rect 71788 31352 71828 31361
rect 71596 31184 71636 31193
rect 71596 30521 71636 31144
rect 71691 30680 71733 30689
rect 71691 30640 71692 30680
rect 71732 30640 71733 30680
rect 71691 30631 71733 30640
rect 71692 30546 71732 30631
rect 71595 30512 71637 30521
rect 71595 30472 71596 30512
rect 71636 30472 71637 30512
rect 71595 30463 71637 30472
rect 71788 30437 71828 31312
rect 71884 31184 71924 31193
rect 71884 30680 71924 31144
rect 72076 30848 72116 31900
rect 72172 30932 72212 32152
rect 72268 31613 72308 32152
rect 72364 32192 72404 32320
rect 72652 32311 72692 32320
rect 72556 32192 72596 32201
rect 72748 32192 72788 32992
rect 72843 32992 72844 33032
rect 72884 32992 72885 33032
rect 72843 32983 72885 32992
rect 72844 32898 72884 32983
rect 72404 32152 72556 32192
rect 72364 32143 72404 32152
rect 72556 32143 72596 32152
rect 72652 32152 72788 32192
rect 72844 32192 72884 32201
rect 72267 31604 72309 31613
rect 72267 31564 72268 31604
rect 72308 31564 72309 31604
rect 72267 31555 72309 31564
rect 72460 31361 72500 31446
rect 72555 31436 72597 31445
rect 72555 31396 72556 31436
rect 72596 31396 72597 31436
rect 72555 31387 72597 31396
rect 72364 31352 72404 31361
rect 72267 31184 72309 31193
rect 72267 31144 72268 31184
rect 72308 31144 72309 31184
rect 72267 31135 72309 31144
rect 72268 31050 72308 31135
rect 72172 30892 72308 30932
rect 72076 30808 72212 30848
rect 71787 30428 71829 30437
rect 71787 30388 71788 30428
rect 71828 30388 71829 30428
rect 71884 30428 71924 30640
rect 71980 30605 72020 30690
rect 72075 30680 72117 30689
rect 72075 30640 72076 30680
rect 72116 30640 72117 30680
rect 72075 30631 72117 30640
rect 71979 30596 72021 30605
rect 71979 30556 71980 30596
rect 72020 30556 72021 30596
rect 71979 30547 72021 30556
rect 72076 30512 72116 30631
rect 72172 30596 72212 30808
rect 72172 30547 72212 30556
rect 72268 30680 72308 30892
rect 72076 30463 72116 30472
rect 71884 30388 72020 30428
rect 71787 30379 71829 30388
rect 71691 30344 71733 30353
rect 71691 30304 71692 30344
rect 71732 30304 71733 30344
rect 71691 30295 71733 30304
rect 71499 30092 71541 30101
rect 71499 30052 71500 30092
rect 71540 30052 71541 30092
rect 71499 30043 71541 30052
rect 71500 29924 71540 30043
rect 71596 29924 71636 29933
rect 71500 29884 71596 29924
rect 71404 29791 71444 29800
rect 71212 29672 71252 29681
rect 71115 29336 71157 29345
rect 71115 29296 71116 29336
rect 71156 29296 71157 29336
rect 71115 29287 71157 29296
rect 71116 29202 71156 29287
rect 70828 29168 70868 29177
rect 70828 28925 70868 29128
rect 71020 29168 71060 29179
rect 71020 29093 71060 29128
rect 71019 29084 71061 29093
rect 71019 29044 71020 29084
rect 71060 29044 71061 29084
rect 71019 29035 71061 29044
rect 70827 28916 70869 28925
rect 71116 28916 71156 28925
rect 70827 28876 70828 28916
rect 70868 28876 70869 28916
rect 70827 28867 70869 28876
rect 71020 28876 71116 28916
rect 71020 28664 71060 28876
rect 71116 28867 71156 28876
rect 71115 28748 71157 28757
rect 71115 28708 71116 28748
rect 71156 28708 71157 28748
rect 71115 28699 71157 28708
rect 70924 28624 71060 28664
rect 70743 28505 70783 28580
rect 70635 28496 70677 28505
rect 70635 28456 70636 28496
rect 70676 28456 70677 28496
rect 70635 28447 70677 28456
rect 70732 28496 70784 28505
rect 70783 28456 70784 28496
rect 70732 28447 70784 28456
rect 70540 28293 70580 28302
rect 70732 28342 70772 28348
rect 70732 28339 70785 28342
rect 70772 28299 70785 28339
rect 70732 28290 70785 28299
rect 70444 28279 70484 28288
rect 70443 28160 70485 28169
rect 70745 28160 70785 28290
rect 70924 28328 70964 28624
rect 71116 28496 71156 28699
rect 71116 28447 71156 28456
rect 71019 28412 71061 28421
rect 71019 28372 71020 28412
rect 71060 28372 71061 28412
rect 71019 28363 71061 28372
rect 71212 28412 71252 29632
rect 71596 29597 71636 29884
rect 71595 29588 71637 29597
rect 71595 29548 71596 29588
rect 71636 29548 71637 29588
rect 71595 29539 71637 29548
rect 71308 29345 71348 29431
rect 71307 29340 71349 29345
rect 71307 29296 71308 29340
rect 71348 29296 71349 29340
rect 71307 29287 71349 29296
rect 71403 29168 71445 29177
rect 71403 29128 71404 29168
rect 71444 29128 71445 29168
rect 71403 29119 71445 29128
rect 71500 29168 71540 29177
rect 71307 29084 71349 29093
rect 71307 29044 71308 29084
rect 71348 29044 71349 29084
rect 71307 29035 71349 29044
rect 71212 28363 71252 28372
rect 70924 28279 70964 28288
rect 71020 28278 71060 28363
rect 71308 28328 71348 29035
rect 71404 29034 71444 29119
rect 71403 28916 71445 28925
rect 71403 28876 71404 28916
rect 71444 28876 71445 28916
rect 71403 28867 71445 28876
rect 71308 28279 71348 28288
rect 71404 28160 71444 28867
rect 71500 28505 71540 29128
rect 71499 28496 71541 28505
rect 71499 28456 71500 28496
rect 71540 28456 71541 28496
rect 71499 28447 71541 28456
rect 70443 28120 70444 28160
rect 70484 28120 70485 28160
rect 70443 28111 70485 28120
rect 70732 28120 70785 28160
rect 71308 28120 71444 28160
rect 70347 27656 70389 27665
rect 70347 27616 70348 27656
rect 70388 27616 70389 27656
rect 70347 27607 70389 27616
rect 70444 27656 70484 28111
rect 70444 27607 70484 27616
rect 69964 25600 70100 25640
rect 70156 25852 70292 25892
rect 69483 25556 69525 25565
rect 69483 25516 69484 25556
rect 69524 25516 69525 25556
rect 69483 25507 69525 25516
rect 69004 25472 69044 25481
rect 68908 25432 69004 25472
rect 69044 25432 69236 25472
rect 69004 25423 69044 25432
rect 68523 25304 68565 25313
rect 68620 25304 68660 25313
rect 68523 25264 68524 25304
rect 68564 25264 68620 25304
rect 68523 25255 68565 25264
rect 68620 25255 68660 25264
rect 68524 25170 68564 25255
rect 68427 25052 68469 25061
rect 68427 25012 68428 25052
rect 68468 25012 68469 25052
rect 68427 25003 68469 25012
rect 68715 24884 68757 24893
rect 68715 24844 68716 24884
rect 68756 24844 68757 24884
rect 68715 24835 68757 24844
rect 68716 24548 68756 24835
rect 68716 24499 68756 24508
rect 69100 24632 69140 24641
rect 68427 24464 68469 24473
rect 68427 24424 68428 24464
rect 68468 24424 68469 24464
rect 68427 24415 68469 24424
rect 68139 24296 68181 24305
rect 68139 24256 68140 24296
rect 68180 24256 68181 24296
rect 68139 24247 68181 24256
rect 67947 24212 67989 24221
rect 67947 24172 67948 24212
rect 67988 24172 67989 24212
rect 67947 24163 67989 24172
rect 67851 23540 67893 23549
rect 67851 23500 67852 23540
rect 67892 23500 67893 23540
rect 67851 23491 67893 23500
rect 67659 23204 67701 23213
rect 67659 23164 67660 23204
rect 67700 23164 67701 23204
rect 67659 23155 67701 23164
rect 67660 23060 67700 23155
rect 67948 23060 67988 24163
rect 68043 23624 68085 23633
rect 68043 23584 68044 23624
rect 68084 23584 68085 23624
rect 68043 23575 68085 23584
rect 67660 23020 67725 23060
rect 67685 22952 67725 23020
rect 67660 22912 67725 22952
rect 67945 23020 67988 23060
rect 68044 23060 68084 23575
rect 68428 23060 68468 24415
rect 68908 24380 68948 24389
rect 68715 24212 68757 24221
rect 68715 24172 68716 24212
rect 68756 24172 68757 24212
rect 68715 24163 68757 24172
rect 68044 23020 68095 23060
rect 67660 22868 67700 22912
rect 67255 22744 67316 22784
rect 67545 22744 67604 22784
rect 67655 22828 67700 22868
rect 67255 22596 67295 22744
rect 67545 22596 67585 22744
rect 67655 22596 67695 22828
rect 67945 22596 67985 23020
rect 68055 22596 68095 23020
rect 68344 23036 68386 23045
rect 68344 22996 68345 23036
rect 68385 22996 68386 23036
rect 68428 23020 68495 23060
rect 68344 22987 68386 22996
rect 68345 22596 68385 22987
rect 68455 22596 68495 23020
rect 68716 22784 68756 24163
rect 68811 24044 68853 24053
rect 68811 24004 68812 24044
rect 68852 24004 68853 24044
rect 68811 23995 68853 24004
rect 68812 23910 68852 23995
rect 68908 23885 68948 24340
rect 68907 23876 68949 23885
rect 68907 23836 68908 23876
rect 68948 23836 68949 23876
rect 68907 23827 68949 23836
rect 68811 23792 68853 23801
rect 68811 23752 68812 23792
rect 68852 23752 68853 23792
rect 68811 23743 68853 23752
rect 69100 23792 69140 24592
rect 69100 23743 69140 23752
rect 69196 23792 69236 25432
rect 69292 25304 69332 25313
rect 69292 24464 69332 25264
rect 69388 25304 69428 25315
rect 69388 25229 69428 25264
rect 69387 25220 69429 25229
rect 69387 25180 69388 25220
rect 69428 25180 69429 25220
rect 69387 25171 69429 25180
rect 69484 25132 69524 25507
rect 69867 25388 69909 25397
rect 69867 25348 69868 25388
rect 69908 25348 69909 25388
rect 69867 25339 69909 25348
rect 69868 25254 69908 25339
rect 69675 25220 69717 25229
rect 69675 25180 69676 25220
rect 69716 25180 69717 25220
rect 69675 25171 69717 25180
rect 69484 25083 69524 25092
rect 69676 25136 69716 25171
rect 69676 25085 69716 25096
rect 69484 24632 69524 24641
rect 69964 24632 70004 25600
rect 70060 25397 70100 25482
rect 70059 25388 70101 25397
rect 70059 25348 70060 25388
rect 70100 25348 70101 25388
rect 70059 25339 70101 25348
rect 70059 25220 70101 25229
rect 70059 25180 70060 25220
rect 70100 25180 70101 25220
rect 70059 25171 70101 25180
rect 69524 24592 70004 24632
rect 69484 24583 69524 24592
rect 69292 24424 70004 24464
rect 69483 24296 69525 24305
rect 69483 24256 69484 24296
rect 69524 24256 69525 24296
rect 69483 24247 69525 24256
rect 69675 24296 69717 24305
rect 69675 24256 69676 24296
rect 69716 24256 69717 24296
rect 69675 24247 69717 24256
rect 69387 23876 69429 23885
rect 69387 23836 69388 23876
rect 69428 23836 69429 23876
rect 69387 23827 69429 23836
rect 69196 23743 69236 23752
rect 69292 23792 69332 23801
rect 68812 23060 68852 23743
rect 69292 23633 69332 23752
rect 69388 23792 69428 23827
rect 69388 23741 69428 23752
rect 69099 23624 69141 23633
rect 69099 23584 69100 23624
rect 69140 23584 69141 23624
rect 69099 23575 69141 23584
rect 69291 23624 69333 23633
rect 69291 23584 69292 23624
rect 69332 23584 69333 23624
rect 69291 23575 69333 23584
rect 69100 23060 69140 23575
rect 69291 23204 69333 23213
rect 69291 23164 69292 23204
rect 69332 23164 69333 23204
rect 69291 23155 69333 23164
rect 69292 23060 69332 23155
rect 68812 23020 68895 23060
rect 69100 23020 69185 23060
rect 68716 22744 68785 22784
rect 68745 22596 68785 22744
rect 68855 22596 68895 23020
rect 69145 22596 69185 23020
rect 69255 23020 69332 23060
rect 69484 23060 69524 24247
rect 69676 23060 69716 24247
rect 69964 23792 70004 24424
rect 70060 24380 70100 25171
rect 70156 24464 70196 25852
rect 70251 25724 70293 25733
rect 70251 25684 70252 25724
rect 70292 25684 70293 25724
rect 70251 25675 70293 25684
rect 70252 25556 70292 25675
rect 70252 25507 70292 25516
rect 70348 24632 70388 27607
rect 70732 27488 70772 28120
rect 71115 27824 71157 27833
rect 71115 27784 71116 27824
rect 71156 27784 71157 27824
rect 71115 27775 71157 27784
rect 71116 27690 71156 27775
rect 70828 27656 70868 27665
rect 71212 27656 71252 27667
rect 70868 27616 71060 27656
rect 70828 27607 70868 27616
rect 70732 27448 70868 27488
rect 70828 26816 70868 27448
rect 71020 26984 71060 27616
rect 71212 27581 71252 27616
rect 71211 27572 71253 27581
rect 71211 27532 71212 27572
rect 71252 27532 71253 27572
rect 71211 27523 71253 27532
rect 71116 27404 71156 27413
rect 71156 27364 71252 27404
rect 71116 27355 71156 27364
rect 71020 26935 71060 26944
rect 70923 26900 70965 26909
rect 70923 26860 70924 26900
rect 70964 26860 70965 26900
rect 70923 26851 70965 26860
rect 71115 26900 71157 26909
rect 71115 26860 71116 26900
rect 71156 26860 71157 26900
rect 71115 26851 71157 26860
rect 70444 26732 70484 26741
rect 70484 26692 70772 26732
rect 70444 26683 70484 26692
rect 70443 26564 70485 26573
rect 70443 26524 70444 26564
rect 70484 26524 70485 26564
rect 70443 26515 70485 26524
rect 70444 25976 70484 26515
rect 70539 26228 70581 26237
rect 70539 26188 70540 26228
rect 70580 26188 70581 26228
rect 70539 26186 70581 26188
rect 70539 26179 70540 26186
rect 70580 26179 70581 26186
rect 70540 26093 70580 26146
rect 70635 26060 70677 26069
rect 70635 26020 70636 26060
rect 70676 26020 70677 26060
rect 70635 26011 70677 26020
rect 70444 25936 70580 25976
rect 70443 25808 70485 25817
rect 70443 25768 70444 25808
rect 70484 25768 70485 25808
rect 70443 25759 70485 25768
rect 70348 24583 70388 24592
rect 70156 24424 70388 24464
rect 70060 24340 70292 24380
rect 70059 23876 70101 23885
rect 70059 23836 70060 23876
rect 70100 23836 70101 23876
rect 70059 23827 70101 23836
rect 69964 23743 70004 23752
rect 70060 23792 70100 23827
rect 70060 23741 70100 23752
rect 70156 23792 70196 23803
rect 70156 23717 70196 23752
rect 70252 23792 70292 24340
rect 70252 23743 70292 23752
rect 70155 23708 70197 23717
rect 70155 23668 70156 23708
rect 70196 23668 70197 23708
rect 70155 23659 70197 23668
rect 69963 23540 70005 23549
rect 69963 23500 69964 23540
rect 70004 23500 70005 23540
rect 69963 23491 70005 23500
rect 69964 23060 70004 23491
rect 70059 23288 70101 23297
rect 70059 23248 70060 23288
rect 70100 23248 70101 23288
rect 70059 23239 70101 23248
rect 70060 23060 70100 23239
rect 70348 23060 70388 24424
rect 69484 23020 69585 23060
rect 69255 22596 69295 23020
rect 69545 22596 69585 23020
rect 69655 23020 69716 23060
rect 69945 23020 70004 23060
rect 70055 23020 70100 23060
rect 70345 23020 70388 23060
rect 70444 23060 70484 25759
rect 70444 23020 70495 23060
rect 69655 22596 69695 23020
rect 69945 22596 69985 23020
rect 70055 22596 70095 23020
rect 70345 22596 70385 23020
rect 70455 22596 70495 23020
rect 70540 22793 70580 25936
rect 70636 25926 70676 26011
rect 70732 25976 70772 26692
rect 70828 26657 70868 26776
rect 70924 26766 70964 26851
rect 71116 26766 71156 26851
rect 71212 26816 71252 27364
rect 71212 26767 71252 26776
rect 70827 26648 70869 26657
rect 70827 26608 70828 26648
rect 70868 26608 70869 26648
rect 70827 26599 70869 26608
rect 70828 26237 70868 26599
rect 71212 26312 71252 26321
rect 70924 26272 71212 26312
rect 70827 26228 70869 26237
rect 70827 26188 70828 26228
rect 70868 26188 70869 26228
rect 70827 26179 70869 26188
rect 70924 26144 70964 26272
rect 70924 26095 70964 26104
rect 70732 25927 70772 25936
rect 70828 26060 70868 26069
rect 70731 25808 70773 25817
rect 70731 25768 70732 25808
rect 70772 25768 70773 25808
rect 70731 25759 70773 25768
rect 70732 23060 70772 25759
rect 70828 24968 70868 26020
rect 71020 25132 71060 26272
rect 71212 26263 71252 26272
rect 71115 26144 71157 26153
rect 71115 26104 71116 26144
rect 71156 26104 71157 26144
rect 71115 26095 71157 26104
rect 71116 26010 71156 26095
rect 71308 25640 71348 28120
rect 71692 28076 71732 30295
rect 71787 30260 71829 30269
rect 71787 30220 71788 30260
rect 71828 30220 71829 30260
rect 71787 30211 71829 30220
rect 71788 30092 71828 30211
rect 71788 30043 71828 30052
rect 71788 29672 71828 29681
rect 71788 29093 71828 29632
rect 71980 29668 72020 30388
rect 72268 30269 72308 30640
rect 72364 30596 72404 31312
rect 72459 31352 72501 31361
rect 72459 31312 72460 31352
rect 72500 31312 72501 31352
rect 72459 31303 72501 31312
rect 72556 31352 72596 31387
rect 72459 31184 72501 31193
rect 72459 31144 72460 31184
rect 72500 31144 72501 31184
rect 72459 31135 72501 31144
rect 72460 30764 72500 31135
rect 72460 30715 72500 30724
rect 72459 30596 72501 30605
rect 72364 30556 72460 30596
rect 72500 30556 72501 30596
rect 72459 30547 72501 30556
rect 72363 30428 72405 30437
rect 72363 30388 72364 30428
rect 72404 30388 72405 30428
rect 72363 30379 72405 30388
rect 72267 30260 72309 30269
rect 72267 30220 72268 30260
rect 72308 30220 72309 30260
rect 72267 30211 72309 30220
rect 72075 30008 72117 30017
rect 72075 29968 72076 30008
rect 72116 29968 72117 30008
rect 72075 29959 72117 29968
rect 72267 30008 72309 30017
rect 72267 29968 72268 30008
rect 72308 29968 72309 30008
rect 72267 29959 72309 29968
rect 72076 29840 72116 29959
rect 72076 29791 72116 29800
rect 72171 29840 72213 29849
rect 72171 29800 72172 29840
rect 72212 29800 72213 29840
rect 72171 29791 72213 29800
rect 72172 29706 72212 29791
rect 71980 29619 72020 29628
rect 72268 29177 72308 29959
rect 72172 29168 72212 29177
rect 71787 29084 71829 29093
rect 71787 29044 71788 29084
rect 71828 29044 71829 29084
rect 71787 29035 71829 29044
rect 71788 28916 71828 28925
rect 71828 28876 71924 28916
rect 71788 28867 71828 28876
rect 71884 28421 71924 28876
rect 71883 28412 71925 28421
rect 71883 28372 71884 28412
rect 71924 28372 71925 28412
rect 71883 28363 71925 28372
rect 72075 28412 72117 28421
rect 72075 28372 72076 28412
rect 72116 28372 72117 28412
rect 72075 28363 72117 28372
rect 71787 28328 71829 28337
rect 71787 28288 71788 28328
rect 71828 28288 71829 28328
rect 71787 28279 71829 28288
rect 71884 28328 71924 28363
rect 71788 28194 71828 28279
rect 71884 28278 71924 28288
rect 71980 28328 72020 28337
rect 71980 28169 72020 28288
rect 72076 28328 72116 28363
rect 72172 28337 72212 29128
rect 72267 29168 72309 29177
rect 72267 29128 72268 29168
rect 72308 29128 72309 29168
rect 72267 29119 72309 29128
rect 72268 28841 72308 29119
rect 72267 28832 72309 28841
rect 72267 28792 72268 28832
rect 72308 28792 72309 28832
rect 72267 28783 72309 28792
rect 72268 28580 72308 28783
rect 72268 28531 72308 28540
rect 72076 28277 72116 28288
rect 72171 28328 72213 28337
rect 72171 28288 72172 28328
rect 72212 28288 72213 28328
rect 72171 28279 72213 28288
rect 71979 28160 72021 28169
rect 71979 28120 71980 28160
rect 72020 28120 72021 28160
rect 71979 28111 72021 28120
rect 71692 28036 71828 28076
rect 71500 27833 71540 27837
rect 71499 27828 71541 27833
rect 71499 27784 71500 27828
rect 71540 27784 71541 27828
rect 71499 27775 71541 27784
rect 71500 27693 71540 27775
rect 71596 27656 71636 27665
rect 71403 27572 71445 27581
rect 71403 27532 71404 27572
rect 71444 27532 71445 27572
rect 71403 27523 71445 27532
rect 71404 26816 71444 27523
rect 71499 27488 71541 27497
rect 71499 27448 71500 27488
rect 71540 27448 71541 27488
rect 71499 27439 71541 27448
rect 71404 26767 71444 26776
rect 71500 26816 71540 27439
rect 71596 27161 71636 27616
rect 71692 27656 71732 27665
rect 71692 27413 71732 27616
rect 71691 27404 71733 27413
rect 71691 27364 71692 27404
rect 71732 27364 71733 27404
rect 71691 27355 71733 27364
rect 71788 27329 71828 28036
rect 72267 27992 72309 28001
rect 72267 27952 72268 27992
rect 72308 27952 72309 27992
rect 72267 27943 72309 27952
rect 71980 27404 72020 27413
rect 72020 27364 72116 27404
rect 71980 27355 72020 27364
rect 71787 27320 71829 27329
rect 71787 27280 71788 27320
rect 71828 27280 71829 27320
rect 71787 27271 71829 27280
rect 71595 27152 71637 27161
rect 71595 27112 71596 27152
rect 71636 27112 71637 27152
rect 71595 27103 71637 27112
rect 71691 26984 71733 26993
rect 71691 26944 71692 26984
rect 71732 26944 71733 26984
rect 71691 26935 71733 26944
rect 71500 26321 71540 26776
rect 71692 26816 71732 26935
rect 72076 26909 72116 27364
rect 72075 26900 72117 26909
rect 72075 26860 72076 26900
rect 72116 26860 72117 26900
rect 72075 26851 72117 26860
rect 71692 26767 71732 26776
rect 71980 26732 72020 26741
rect 71788 26692 71980 26732
rect 71596 26648 71636 26657
rect 71499 26312 71541 26321
rect 71499 26272 71500 26312
rect 71540 26272 71541 26312
rect 71499 26263 71541 26272
rect 71596 26069 71636 26608
rect 71788 26312 71828 26692
rect 71980 26683 72020 26692
rect 72076 26564 72116 26851
rect 71788 26263 71828 26272
rect 71884 26524 72116 26564
rect 72268 26564 72308 27943
rect 72364 26984 72404 30379
rect 72460 30092 72500 30547
rect 72460 30043 72500 30052
rect 72556 29840 72596 31312
rect 72652 30596 72692 32152
rect 72844 32108 72884 32152
rect 72748 32068 72884 32108
rect 72748 31352 72788 32068
rect 72843 31688 72885 31697
rect 72843 31648 72844 31688
rect 72884 31648 72885 31688
rect 72843 31639 72885 31648
rect 72748 31303 72788 31312
rect 72844 31352 72884 31639
rect 73036 31445 73076 33235
rect 73420 33140 73460 33244
rect 73324 33100 73460 33140
rect 73228 32192 73268 32201
rect 73132 32152 73228 32192
rect 73035 31436 73077 31445
rect 73035 31396 73036 31436
rect 73076 31396 73077 31436
rect 73035 31387 73077 31396
rect 72844 31303 72884 31312
rect 72940 31352 72980 31361
rect 72940 31193 72980 31312
rect 73036 31352 73076 31387
rect 73036 31302 73076 31312
rect 72939 31184 72981 31193
rect 72939 31144 72940 31184
rect 72980 31144 72981 31184
rect 72939 31135 72981 31144
rect 73132 31016 73172 32152
rect 73228 32143 73268 32152
rect 72844 30976 73172 31016
rect 73228 31436 73268 31445
rect 73324 31436 73364 33100
rect 73996 31697 74036 33319
rect 74092 32873 74132 34327
rect 74091 32864 74133 32873
rect 74091 32824 74092 32864
rect 74132 32824 74133 32864
rect 74091 32815 74133 32824
rect 74092 32192 74132 32815
rect 73995 31688 74037 31697
rect 73995 31648 73996 31688
rect 74036 31648 74037 31688
rect 73995 31639 74037 31648
rect 73708 31445 73748 31476
rect 73268 31396 73364 31436
rect 73707 31436 73749 31445
rect 73707 31396 73708 31436
rect 73748 31396 73749 31436
rect 72844 30689 72884 30976
rect 72843 30680 72885 30689
rect 72843 30640 72844 30680
rect 72884 30640 72885 30680
rect 72843 30631 72885 30640
rect 72652 30556 72788 30596
rect 72651 30260 72693 30269
rect 72651 30220 72652 30260
rect 72692 30220 72693 30260
rect 72651 30211 72693 30220
rect 72652 30092 72692 30211
rect 72652 30043 72692 30052
rect 72748 30017 72788 30556
rect 72844 30546 72884 30631
rect 73228 30269 73268 31396
rect 73707 31387 73749 31396
rect 73611 31352 73653 31361
rect 73611 31312 73612 31352
rect 73652 31312 73653 31352
rect 73611 31303 73653 31312
rect 73708 31352 73748 31387
rect 73900 31352 73940 31361
rect 73515 31268 73557 31277
rect 73515 31228 73516 31268
rect 73556 31228 73557 31268
rect 73515 31219 73557 31228
rect 73420 31184 73460 31193
rect 73420 31025 73460 31144
rect 73419 31016 73461 31025
rect 73419 30976 73420 31016
rect 73460 30976 73461 31016
rect 73419 30967 73461 30976
rect 73227 30260 73269 30269
rect 73227 30220 73228 30260
rect 73268 30220 73269 30260
rect 73227 30211 73269 30220
rect 73227 30092 73269 30101
rect 73227 30052 73228 30092
rect 73268 30052 73269 30092
rect 73227 30043 73269 30052
rect 72747 30008 72789 30017
rect 72747 29968 72748 30008
rect 72788 29968 72789 30008
rect 72747 29959 72789 29968
rect 72844 29924 72884 29933
rect 72884 29884 72980 29924
rect 72844 29875 72884 29884
rect 72556 29800 72788 29840
rect 72748 29756 72788 29800
rect 72748 29716 72884 29756
rect 72652 29672 72692 29681
rect 72460 29632 72652 29672
rect 72460 28412 72500 29632
rect 72652 29623 72692 29632
rect 72555 29168 72597 29177
rect 72555 29128 72556 29168
rect 72596 29128 72597 29168
rect 72555 29119 72597 29128
rect 72556 29034 72596 29119
rect 72747 28496 72789 28505
rect 72747 28456 72748 28496
rect 72788 28456 72789 28496
rect 72747 28447 72789 28456
rect 72460 28363 72500 28372
rect 72748 28328 72788 28447
rect 72844 28421 72884 29716
rect 72940 29588 72980 29884
rect 73131 29840 73173 29849
rect 73131 29800 73132 29840
rect 73172 29800 73173 29840
rect 73131 29791 73173 29800
rect 73228 29840 73268 30043
rect 73420 29933 73460 30967
rect 73516 30521 73556 31219
rect 73612 31218 73652 31303
rect 73708 31100 73748 31312
rect 73804 31331 73844 31340
rect 73804 31277 73844 31291
rect 73803 31268 73845 31277
rect 73803 31228 73804 31268
rect 73844 31228 73845 31268
rect 73803 31219 73845 31228
rect 73804 31196 73844 31219
rect 73612 31060 73748 31100
rect 73515 30512 73557 30521
rect 73515 30472 73516 30512
rect 73556 30472 73557 30512
rect 73515 30463 73557 30472
rect 73612 30101 73652 31060
rect 73900 31025 73940 31312
rect 73899 31016 73941 31025
rect 73899 30976 73900 31016
rect 73940 30976 73941 31016
rect 73899 30967 73941 30976
rect 74092 30932 74132 32152
rect 74187 31688 74229 31697
rect 74187 31648 74188 31688
rect 74228 31648 74229 31688
rect 74187 31639 74229 31648
rect 73996 30892 74132 30932
rect 73708 30680 73748 30689
rect 73708 30605 73748 30640
rect 73996 30605 74036 30892
rect 73707 30596 73749 30605
rect 73707 30556 73708 30596
rect 73748 30556 73749 30596
rect 73707 30547 73749 30556
rect 73995 30596 74037 30605
rect 73995 30556 73996 30596
rect 74036 30556 74037 30596
rect 73995 30547 74037 30556
rect 73611 30092 73653 30101
rect 73611 30052 73612 30092
rect 73652 30052 73653 30092
rect 73611 30043 73653 30052
rect 73612 29958 73652 30043
rect 73419 29924 73461 29933
rect 73419 29875 73420 29924
rect 73228 29791 73268 29800
rect 73323 29840 73365 29849
rect 73323 29800 73324 29840
rect 73364 29800 73365 29840
rect 73323 29791 73365 29800
rect 73460 29875 73461 29924
rect 73132 29706 73172 29791
rect 73324 29706 73364 29791
rect 73420 29790 73460 29845
rect 72940 29548 73172 29588
rect 73035 28832 73077 28841
rect 73035 28792 73036 28832
rect 73076 28792 73077 28832
rect 73035 28783 73077 28792
rect 72843 28412 72885 28421
rect 72843 28372 72844 28412
rect 72884 28372 72885 28412
rect 72843 28363 72885 28372
rect 72748 28279 72788 28288
rect 72844 28328 72884 28363
rect 72844 28278 72884 28288
rect 72939 28328 72981 28337
rect 72939 28288 72940 28328
rect 72980 28288 72981 28328
rect 72939 28279 72981 28288
rect 73036 28328 73076 28783
rect 73036 28279 73076 28288
rect 72940 28194 72980 28279
rect 72651 27404 72693 27413
rect 72651 27364 72652 27404
rect 72692 27364 72693 27404
rect 72651 27355 72693 27364
rect 72364 26944 72500 26984
rect 72363 26816 72405 26825
rect 72363 26776 72364 26816
rect 72404 26776 72405 26816
rect 72363 26767 72405 26776
rect 72364 26682 72404 26767
rect 72268 26524 72404 26564
rect 71884 26144 71924 26524
rect 71884 26095 71924 26104
rect 71980 26144 72020 26153
rect 71595 26060 71637 26069
rect 71595 26020 71596 26060
rect 71636 26020 71637 26060
rect 71595 26011 71637 26020
rect 71980 25985 72020 26104
rect 72076 26144 72116 26153
rect 72076 26069 72116 26104
rect 72075 26060 72117 26069
rect 72075 26020 72076 26060
rect 72116 26020 72117 26060
rect 72075 26011 72117 26020
rect 71979 25976 72021 25985
rect 71979 25936 71980 25976
rect 72020 25936 72021 25976
rect 71979 25927 72021 25936
rect 71308 25600 71636 25640
rect 71500 25472 71540 25481
rect 71308 25432 71500 25472
rect 71116 25304 71156 25315
rect 71116 25229 71156 25264
rect 71211 25304 71253 25313
rect 71211 25264 71212 25304
rect 71252 25264 71253 25304
rect 71211 25255 71253 25264
rect 71115 25220 71157 25229
rect 71115 25180 71116 25220
rect 71156 25180 71157 25220
rect 71115 25171 71157 25180
rect 71212 25170 71252 25255
rect 71020 25083 71060 25092
rect 71308 24968 71348 25432
rect 71500 25423 71540 25432
rect 71596 25132 71636 25600
rect 71979 25304 72021 25313
rect 71979 25264 71980 25304
rect 72020 25264 72021 25304
rect 71979 25255 72021 25264
rect 72076 25304 72116 26011
rect 71980 25170 72020 25255
rect 71596 25092 71828 25132
rect 70828 24928 71348 24968
rect 71115 24464 71157 24473
rect 71115 24424 71116 24464
rect 71156 24424 71157 24464
rect 71115 24415 71157 24424
rect 70732 23020 70785 23060
rect 70539 22784 70581 22793
rect 70539 22744 70540 22784
rect 70580 22744 70581 22784
rect 70539 22735 70581 22744
rect 70745 22596 70785 23020
rect 70854 22784 70896 22793
rect 70854 22744 70855 22784
rect 70895 22744 70896 22784
rect 71116 22784 71156 24415
rect 71211 24128 71253 24137
rect 71211 24088 71212 24128
rect 71252 24088 71253 24128
rect 71211 24079 71253 24088
rect 71212 23792 71252 24079
rect 71212 23743 71252 23752
rect 71308 23792 71348 24928
rect 71692 24632 71732 24641
rect 71500 24380 71540 24389
rect 71540 24340 71636 24380
rect 71500 24331 71540 24340
rect 71499 23876 71541 23885
rect 71499 23836 71500 23876
rect 71540 23836 71541 23876
rect 71499 23827 71541 23836
rect 71308 23743 71348 23752
rect 71403 23792 71445 23801
rect 71403 23752 71404 23792
rect 71444 23752 71445 23792
rect 71403 23743 71445 23752
rect 71500 23792 71540 23827
rect 71404 23658 71444 23743
rect 71500 23741 71540 23752
rect 71596 23717 71636 24340
rect 71692 24137 71732 24592
rect 71691 24128 71733 24137
rect 71691 24088 71692 24128
rect 71732 24088 71733 24128
rect 71691 24079 71733 24088
rect 71595 23708 71637 23717
rect 71595 23668 71596 23708
rect 71636 23668 71637 23708
rect 71595 23659 71637 23668
rect 71307 23540 71349 23549
rect 71307 23500 71308 23540
rect 71348 23500 71349 23540
rect 71307 23491 71349 23500
rect 71308 23060 71348 23491
rect 71255 23020 71348 23060
rect 71116 22744 71185 22784
rect 70854 22735 70896 22744
rect 70855 22596 70895 22735
rect 71145 22596 71185 22744
rect 71255 22596 71295 23020
rect 71544 22868 71586 22877
rect 71544 22828 71545 22868
rect 71585 22828 71586 22868
rect 71544 22819 71586 22828
rect 71545 22596 71585 22819
rect 71788 22793 71828 25092
rect 71979 25052 72021 25061
rect 71979 25012 71980 25052
rect 72020 25012 72021 25052
rect 71979 25003 72021 25012
rect 71980 24632 72020 25003
rect 72076 24800 72116 25264
rect 72171 25304 72213 25313
rect 72171 25264 72172 25304
rect 72212 25264 72213 25304
rect 72171 25255 72213 25264
rect 72268 25304 72308 25313
rect 72172 25170 72212 25255
rect 72268 25229 72308 25264
rect 72267 25220 72309 25229
rect 72267 25180 72268 25220
rect 72308 25180 72309 25220
rect 72267 25171 72309 25180
rect 72268 24809 72308 25171
rect 72267 24800 72309 24809
rect 72076 24760 72212 24800
rect 72076 24632 72116 24641
rect 71980 24592 72076 24632
rect 72076 24583 72116 24592
rect 71883 24380 71925 24389
rect 71883 24340 71884 24380
rect 71924 24340 71925 24380
rect 71883 24331 71925 24340
rect 71884 23060 71924 24331
rect 72075 24044 72117 24053
rect 72075 24004 72076 24044
rect 72116 24004 72117 24044
rect 72075 23995 72117 24004
rect 71979 23960 72021 23969
rect 71979 23920 71980 23960
rect 72020 23920 72021 23960
rect 71979 23911 72021 23920
rect 71980 23826 72020 23911
rect 72076 23792 72116 23995
rect 72172 23885 72212 24760
rect 72267 24760 72268 24800
rect 72308 24760 72309 24800
rect 72267 24751 72309 24760
rect 72364 24632 72404 26524
rect 72460 25397 72500 26944
rect 72652 26312 72692 27355
rect 73132 27245 73172 29548
rect 73453 29168 73493 29177
rect 73708 29168 73748 30547
rect 74091 30512 74133 30521
rect 74091 30472 74092 30512
rect 74132 30472 74133 30512
rect 74091 30463 74133 30472
rect 73803 30260 73845 30269
rect 73803 30220 73804 30260
rect 73844 30220 73845 30260
rect 73803 30211 73845 30220
rect 73804 29924 73844 30211
rect 74092 30092 74132 30463
rect 74092 30043 74132 30052
rect 73804 29875 73844 29884
rect 73995 29840 74037 29849
rect 73995 29800 73996 29840
rect 74036 29800 74037 29840
rect 73995 29791 74037 29800
rect 73996 29706 74036 29791
rect 73493 29128 73748 29168
rect 74092 29672 74132 29681
rect 73453 29119 73493 29128
rect 73227 28328 73269 28337
rect 73227 28288 73228 28328
rect 73268 28288 73269 28328
rect 73227 28279 73269 28288
rect 73708 28328 73748 28339
rect 74092 28328 74132 29632
rect 73228 27665 73268 28279
rect 73708 28253 73748 28288
rect 73804 28288 74132 28328
rect 73707 28244 73749 28253
rect 73707 28204 73708 28244
rect 73748 28204 73749 28244
rect 73707 28195 73749 28204
rect 73611 28160 73653 28169
rect 73611 28120 73612 28160
rect 73652 28120 73653 28160
rect 73611 28111 73653 28120
rect 73612 28026 73652 28111
rect 73227 27656 73269 27665
rect 73227 27616 73228 27656
rect 73268 27616 73269 27656
rect 73227 27607 73269 27616
rect 73131 27236 73173 27245
rect 73131 27196 73132 27236
rect 73172 27196 73173 27236
rect 73131 27187 73173 27196
rect 72939 27152 72981 27161
rect 72939 27112 72940 27152
rect 72980 27112 72981 27152
rect 72939 27103 72981 27112
rect 72652 26263 72692 26272
rect 72748 26144 72788 26155
rect 72748 26069 72788 26104
rect 72843 26144 72885 26153
rect 72843 26104 72844 26144
rect 72884 26104 72885 26144
rect 72843 26095 72885 26104
rect 72940 26144 72980 27103
rect 73131 26816 73173 26825
rect 73131 26776 73132 26816
rect 73172 26776 73173 26816
rect 73131 26767 73173 26776
rect 73228 26816 73268 27607
rect 73228 26767 73268 26776
rect 72747 26060 72789 26069
rect 72747 26020 72748 26060
rect 72788 26020 72789 26060
rect 72747 26011 72789 26020
rect 72844 26010 72884 26095
rect 72459 25388 72501 25397
rect 72459 25348 72460 25388
rect 72500 25348 72501 25388
rect 72459 25339 72501 25348
rect 72843 25304 72885 25313
rect 72843 25264 72844 25304
rect 72884 25264 72885 25304
rect 72843 25255 72885 25264
rect 72268 24592 72404 24632
rect 72171 23876 72213 23885
rect 72171 23836 72172 23876
rect 72212 23836 72213 23876
rect 72171 23827 72213 23836
rect 72076 23549 72116 23752
rect 72268 23708 72308 24592
rect 72844 24557 72884 25255
rect 72940 24809 72980 26104
rect 73132 25145 73172 26767
rect 73323 26144 73365 26153
rect 73323 26104 73324 26144
rect 73364 26104 73365 26144
rect 73323 26095 73365 26104
rect 73707 26144 73749 26153
rect 73707 26104 73708 26144
rect 73748 26104 73749 26144
rect 73707 26095 73749 26104
rect 73324 26010 73364 26095
rect 73419 25976 73461 25985
rect 73419 25936 73420 25976
rect 73460 25936 73461 25976
rect 73419 25927 73461 25936
rect 73420 25842 73460 25927
rect 73612 25304 73652 25313
rect 73227 25220 73269 25229
rect 73227 25180 73228 25220
rect 73268 25180 73269 25220
rect 73227 25171 73269 25180
rect 73131 25136 73173 25145
rect 73131 25096 73132 25136
rect 73172 25096 73173 25136
rect 73131 25087 73173 25096
rect 73228 25086 73268 25171
rect 73612 25145 73652 25264
rect 73611 25136 73653 25145
rect 73611 25096 73612 25136
rect 73652 25096 73653 25136
rect 73611 25087 73653 25096
rect 72939 24800 72981 24809
rect 72939 24760 72940 24800
rect 72980 24760 72981 24800
rect 72939 24751 72981 24760
rect 72939 24632 72981 24641
rect 72939 24592 72940 24632
rect 72980 24592 72981 24632
rect 72939 24583 72981 24592
rect 72843 24548 72885 24557
rect 72843 24508 72844 24548
rect 72884 24508 72885 24548
rect 72843 24499 72885 24508
rect 72651 23960 72693 23969
rect 72651 23920 72652 23960
rect 72692 23920 72693 23960
rect 72651 23911 72693 23920
rect 72460 23792 72500 23803
rect 72460 23717 72500 23752
rect 72172 23668 72308 23708
rect 72459 23708 72501 23717
rect 72459 23668 72460 23708
rect 72500 23668 72501 23708
rect 72075 23540 72117 23549
rect 72075 23500 72076 23540
rect 72116 23500 72117 23540
rect 72075 23491 72117 23500
rect 72172 23060 72212 23668
rect 72459 23659 72501 23668
rect 72363 23624 72405 23633
rect 72363 23584 72364 23624
rect 72404 23584 72405 23624
rect 72363 23575 72405 23584
rect 72364 23490 72404 23575
rect 72459 23456 72501 23465
rect 72459 23416 72460 23456
rect 72500 23416 72501 23456
rect 72459 23407 72501 23416
rect 72363 23372 72405 23381
rect 72363 23332 72364 23372
rect 72404 23332 72405 23372
rect 72363 23323 72405 23332
rect 72364 23060 72404 23323
rect 72460 23060 72500 23407
rect 71884 23020 71985 23060
rect 71654 22784 71696 22793
rect 71654 22744 71655 22784
rect 71695 22744 71696 22784
rect 71654 22735 71696 22744
rect 71787 22784 71829 22793
rect 71787 22744 71788 22784
rect 71828 22744 71829 22784
rect 71787 22735 71829 22744
rect 71655 22596 71695 22735
rect 71945 22596 71985 23020
rect 72055 23020 72212 23060
rect 72345 23020 72404 23060
rect 72455 23020 72500 23060
rect 72652 23060 72692 23911
rect 72747 23792 72789 23801
rect 72747 23752 72748 23792
rect 72788 23752 72789 23792
rect 72747 23743 72789 23752
rect 72844 23792 72884 24499
rect 72940 24498 72980 24583
rect 73611 24548 73653 24557
rect 73611 24508 73612 24548
rect 73652 24508 73653 24548
rect 73611 24499 73653 24508
rect 72844 23743 72884 23752
rect 72748 23658 72788 23743
rect 73227 23708 73269 23717
rect 73227 23668 73228 23708
rect 73268 23668 73269 23708
rect 73227 23659 73269 23668
rect 73131 23624 73173 23633
rect 73131 23584 73132 23624
rect 73172 23584 73173 23624
rect 73131 23575 73173 23584
rect 72843 23540 72885 23549
rect 72843 23500 72844 23540
rect 72884 23500 72885 23540
rect 72843 23491 72885 23500
rect 72844 23060 72884 23491
rect 73132 23060 73172 23575
rect 73228 23060 73268 23659
rect 73515 23624 73557 23633
rect 73515 23584 73516 23624
rect 73556 23584 73557 23624
rect 73515 23575 73557 23584
rect 73323 23204 73365 23213
rect 73323 23164 73324 23204
rect 73364 23164 73471 23204
rect 73323 23155 73365 23164
rect 73324 23147 73364 23155
rect 72652 23020 72785 23060
rect 72844 23020 72895 23060
rect 73132 23020 73185 23060
rect 73228 23020 73295 23060
rect 72055 22596 72095 23020
rect 72345 22596 72385 23020
rect 72455 22596 72495 23020
rect 72745 22596 72785 23020
rect 72855 22596 72895 23020
rect 73145 22596 73185 23020
rect 73255 22596 73295 23020
rect 73431 22897 73471 23164
rect 73516 23060 73556 23575
rect 73612 23213 73652 24499
rect 73611 23204 73653 23213
rect 73611 23164 73612 23204
rect 73652 23164 73653 23204
rect 73611 23155 73653 23164
rect 73516 23020 73585 23060
rect 73420 22793 73471 22897
rect 73419 22784 73471 22793
rect 73419 22744 73420 22784
rect 73460 22744 73471 22784
rect 73419 22735 73461 22744
rect 73545 22596 73585 23020
rect 73708 22952 73748 26095
rect 73804 23549 73844 28288
rect 73995 28160 74037 28169
rect 73995 28120 73996 28160
rect 74036 28120 74037 28160
rect 73995 28111 74037 28120
rect 73899 25976 73941 25985
rect 73899 25936 73900 25976
rect 73940 25936 73941 25976
rect 73899 25927 73941 25936
rect 73803 23540 73845 23549
rect 73803 23500 73804 23540
rect 73844 23500 73845 23540
rect 73803 23491 73845 23500
rect 73900 22952 73940 25927
rect 73996 23060 74036 28111
rect 74091 24548 74133 24557
rect 74091 24508 74092 24548
rect 74132 24508 74133 24548
rect 74091 24499 74133 24508
rect 74092 24414 74132 24499
rect 74188 23717 74228 31639
rect 74380 31529 74420 35848
rect 74667 35839 74709 35848
rect 74475 35720 74517 35729
rect 74475 35680 74476 35720
rect 74516 35680 74517 35720
rect 74475 35671 74517 35680
rect 74860 35720 74900 35923
rect 74476 35586 74516 35671
rect 74860 35645 74900 35680
rect 74859 35636 74901 35645
rect 74859 35596 74860 35636
rect 74900 35596 74901 35636
rect 74859 35587 74901 35596
rect 74572 35216 74612 35225
rect 74956 35216 74996 37360
rect 75052 37351 75092 37360
rect 75340 37157 75380 37435
rect 76588 37400 76628 37411
rect 76107 37232 76149 37241
rect 76107 37192 76108 37232
rect 76148 37192 76149 37232
rect 76107 37183 76149 37192
rect 76204 37232 76244 37243
rect 76492 37241 76532 37326
rect 76588 37325 76628 37360
rect 76587 37316 76629 37325
rect 76587 37276 76588 37316
rect 76628 37276 76629 37316
rect 76587 37267 76629 37276
rect 76780 37316 76820 37325
rect 75339 37148 75381 37157
rect 75339 37108 75340 37148
rect 75380 37108 75381 37148
rect 75339 37099 75381 37108
rect 75340 36728 75380 37099
rect 75340 36679 75380 36688
rect 75628 36728 75668 36737
rect 75436 36485 75476 36570
rect 75435 36476 75477 36485
rect 75435 36436 75436 36476
rect 75476 36436 75477 36476
rect 75435 36427 75477 36436
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 75628 35645 75668 36688
rect 75724 36728 75764 36737
rect 75724 36140 75764 36688
rect 75820 36728 75860 36739
rect 75820 36653 75860 36688
rect 75915 36728 75957 36737
rect 75915 36688 75916 36728
rect 75956 36688 75957 36728
rect 75915 36679 75957 36688
rect 76108 36728 76148 37183
rect 76204 37157 76244 37192
rect 76491 37232 76533 37241
rect 76491 37192 76492 37232
rect 76532 37192 76533 37232
rect 76491 37183 76533 37192
rect 76203 37148 76245 37157
rect 76203 37108 76204 37148
rect 76244 37108 76245 37148
rect 76203 37099 76245 37108
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 76780 36896 76820 37276
rect 77068 36905 77108 38116
rect 77260 38107 77300 38116
rect 77452 37988 77492 37997
rect 77356 37948 77452 37988
rect 77164 37400 77204 37409
rect 77356 37400 77396 37948
rect 77452 37939 77492 37948
rect 77204 37360 77396 37400
rect 77164 37351 77204 37360
rect 75819 36644 75861 36653
rect 75819 36604 75820 36644
rect 75860 36604 75861 36644
rect 75819 36595 75861 36604
rect 75916 36594 75956 36679
rect 75724 36100 75860 36140
rect 75627 35636 75669 35645
rect 75627 35596 75628 35636
rect 75668 35596 75669 35636
rect 75627 35587 75669 35596
rect 75051 35384 75093 35393
rect 75051 35344 75052 35384
rect 75092 35344 75093 35384
rect 75051 35335 75093 35344
rect 75723 35384 75765 35393
rect 75723 35344 75724 35384
rect 75764 35344 75765 35384
rect 75723 35335 75765 35344
rect 74612 35176 74996 35216
rect 74572 34385 74612 35176
rect 75052 34964 75092 35335
rect 75724 35250 75764 35335
rect 75820 34973 75860 36100
rect 76108 36065 76148 36688
rect 76300 36856 76820 36896
rect 77067 36896 77109 36905
rect 77067 36856 77068 36896
rect 77108 36856 77109 36896
rect 76203 36644 76245 36653
rect 76203 36604 76204 36644
rect 76244 36604 76245 36644
rect 76203 36595 76245 36604
rect 76204 36510 76244 36595
rect 76300 36560 76340 36856
rect 77067 36847 77109 36856
rect 76492 36728 76532 36737
rect 76300 36511 76340 36520
rect 76396 36644 76436 36653
rect 76396 36149 76436 36604
rect 76492 36233 76532 36688
rect 76683 36728 76725 36737
rect 76683 36688 76684 36728
rect 76724 36688 76725 36728
rect 76683 36679 76725 36688
rect 77068 36728 77108 36737
rect 77108 36688 77204 36728
rect 76684 36594 76724 36679
rect 77068 36569 77108 36688
rect 77067 36560 77109 36569
rect 77067 36520 77068 36560
rect 77108 36520 77109 36560
rect 77067 36511 77109 36520
rect 76491 36224 76533 36233
rect 76491 36184 76492 36224
rect 76532 36184 76533 36224
rect 76491 36175 76533 36184
rect 76395 36140 76437 36149
rect 76395 36100 76396 36140
rect 76436 36100 76437 36140
rect 76395 36091 76437 36100
rect 76107 36056 76149 36065
rect 76107 36016 76108 36056
rect 76148 36016 76149 36056
rect 76107 36007 76149 36016
rect 76588 36016 77012 36056
rect 76491 35972 76533 35981
rect 76491 35932 76492 35972
rect 76532 35932 76533 35972
rect 76491 35923 76533 35932
rect 76300 35888 76340 35897
rect 76300 35729 76340 35848
rect 76396 35888 76436 35899
rect 76396 35813 76436 35848
rect 76492 35888 76532 35923
rect 76492 35837 76532 35848
rect 76588 35888 76628 36016
rect 76588 35839 76628 35848
rect 76779 35888 76821 35897
rect 76779 35848 76780 35888
rect 76820 35848 76821 35888
rect 76779 35839 76821 35848
rect 76876 35888 76916 35897
rect 76395 35804 76437 35813
rect 76395 35764 76396 35804
rect 76436 35764 76437 35804
rect 76395 35755 76437 35764
rect 76299 35720 76341 35729
rect 76299 35680 76300 35720
rect 76340 35680 76341 35720
rect 76299 35671 76341 35680
rect 76780 35716 76820 35839
rect 76876 35729 76916 35848
rect 76972 35888 77012 36016
rect 76972 35839 77012 35848
rect 77067 35804 77109 35813
rect 77067 35764 77068 35804
rect 77108 35764 77109 35804
rect 77067 35755 77109 35764
rect 76780 35667 76820 35676
rect 76875 35720 76917 35729
rect 76875 35680 76876 35720
rect 76916 35680 76917 35720
rect 76875 35671 76917 35680
rect 76203 35636 76245 35645
rect 76203 35596 76204 35636
rect 76244 35596 76245 35636
rect 76203 35587 76245 35596
rect 74860 34924 75092 34964
rect 75819 34964 75861 34973
rect 75819 34924 75820 34964
rect 75860 34924 75861 34964
rect 74571 34376 74613 34385
rect 74571 34336 74572 34376
rect 74612 34336 74613 34376
rect 74571 34327 74613 34336
rect 74764 34208 74804 34217
rect 74572 34168 74764 34208
rect 74572 33713 74612 34168
rect 74764 34159 74804 34168
rect 74571 33704 74613 33713
rect 74571 33664 74572 33704
rect 74612 33664 74613 33704
rect 74571 33655 74613 33664
rect 74764 33704 74804 33713
rect 74860 33704 74900 34924
rect 75819 34915 75861 34924
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 76107 34376 76149 34385
rect 76107 34336 76108 34376
rect 76148 34336 76149 34376
rect 76107 34327 76149 34336
rect 76108 34242 76148 34327
rect 74956 34208 74996 34217
rect 74956 33881 74996 34168
rect 76204 33965 76244 35587
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 76299 35384 76341 35393
rect 77068 35384 77108 35755
rect 76299 35344 76300 35384
rect 76340 35344 76341 35384
rect 76299 35335 76341 35344
rect 76876 35344 77108 35384
rect 76300 34889 76340 35335
rect 76876 35225 76916 35344
rect 77164 35300 77204 36688
rect 77259 36644 77301 36653
rect 77259 36604 77260 36644
rect 77300 36604 77301 36644
rect 77259 36595 77301 36604
rect 77260 36140 77300 36595
rect 77260 36091 77300 36100
rect 77164 35260 77205 35300
rect 76875 35216 76917 35225
rect 76875 35176 76876 35216
rect 76916 35176 76917 35216
rect 76875 35167 76917 35176
rect 77067 35216 77109 35225
rect 77067 35176 77068 35216
rect 77108 35176 77109 35216
rect 77067 35167 77109 35176
rect 76876 35082 76916 35167
rect 77068 35082 77108 35167
rect 77165 35132 77205 35260
rect 77259 35216 77301 35225
rect 77259 35176 77260 35216
rect 77300 35176 77301 35216
rect 77356 35216 77396 37360
rect 78028 37400 78068 37409
rect 77932 36728 77972 36737
rect 78028 36728 78068 37360
rect 79179 37316 79221 37325
rect 79179 37276 79180 37316
rect 79220 37276 79221 37316
rect 79179 37267 79221 37276
rect 79180 37232 79220 37267
rect 79180 37181 79220 37192
rect 77972 36688 78164 36728
rect 77932 36679 77972 36688
rect 77547 36224 77589 36233
rect 77547 36184 77548 36224
rect 77588 36184 77589 36224
rect 77547 36175 77589 36184
rect 77451 36140 77493 36149
rect 77451 36100 77452 36140
rect 77492 36100 77493 36140
rect 77451 36091 77493 36100
rect 77452 36006 77492 36091
rect 77452 35888 77492 35897
rect 77548 35888 77588 36175
rect 77492 35848 77588 35888
rect 77452 35839 77492 35848
rect 77452 35216 77492 35225
rect 77356 35176 77452 35216
rect 77259 35167 77301 35176
rect 77164 35092 77205 35132
rect 76779 34964 76821 34973
rect 76779 34924 76780 34964
rect 76820 34924 76821 34964
rect 76779 34915 76821 34924
rect 76299 34880 76341 34889
rect 76299 34840 76300 34880
rect 76340 34840 76341 34880
rect 76299 34831 76341 34840
rect 76780 34830 76820 34915
rect 76875 34880 76917 34889
rect 76875 34840 76876 34880
rect 76916 34840 76917 34880
rect 76875 34831 76917 34840
rect 76876 34208 76916 34831
rect 76972 34376 77012 34385
rect 77164 34376 77204 35092
rect 77012 34336 77204 34376
rect 76972 34327 77012 34336
rect 76876 34168 77012 34208
rect 76352 34040 76720 34049
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 76203 33956 76245 33965
rect 76203 33916 76204 33956
rect 76244 33916 76245 33956
rect 76203 33907 76245 33916
rect 76875 33956 76917 33965
rect 76875 33916 76876 33956
rect 76916 33916 76917 33956
rect 76875 33907 76917 33916
rect 74955 33872 74997 33881
rect 74955 33832 74956 33872
rect 74996 33832 74997 33872
rect 74955 33823 74997 33832
rect 76299 33872 76341 33881
rect 76299 33832 76300 33872
rect 76340 33832 76341 33872
rect 76299 33823 76341 33832
rect 76587 33872 76629 33881
rect 76587 33832 76588 33872
rect 76628 33832 76629 33872
rect 76587 33823 76629 33832
rect 76779 33872 76821 33881
rect 76779 33832 76780 33872
rect 76820 33832 76821 33872
rect 76779 33823 76821 33832
rect 76876 33872 76916 33907
rect 76300 33704 76340 33823
rect 74804 33664 74996 33704
rect 74764 33655 74804 33664
rect 74572 33140 74612 33655
rect 74859 33452 74901 33461
rect 74859 33412 74860 33452
rect 74900 33412 74901 33452
rect 74859 33403 74901 33412
rect 74860 33318 74900 33403
rect 74956 33140 74996 33664
rect 76300 33461 76340 33664
rect 76395 33704 76437 33713
rect 76395 33664 76396 33704
rect 76436 33664 76437 33704
rect 76395 33655 76437 33664
rect 76588 33704 76628 33823
rect 76588 33655 76628 33664
rect 76683 33704 76725 33713
rect 76683 33664 76684 33704
rect 76724 33664 76725 33704
rect 76683 33655 76725 33664
rect 76780 33704 76820 33823
rect 76876 33821 76916 33832
rect 76780 33655 76820 33664
rect 76396 33570 76436 33655
rect 76684 33570 76724 33655
rect 75723 33452 75765 33461
rect 75723 33412 75724 33452
rect 75764 33412 75765 33452
rect 75723 33403 75765 33412
rect 76299 33452 76341 33461
rect 76299 33412 76300 33452
rect 76340 33412 76341 33452
rect 76299 33403 76341 33412
rect 75112 33284 75480 33293
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75112 33235 75480 33244
rect 74572 33100 74708 33140
rect 74956 33100 75668 33140
rect 74379 31520 74421 31529
rect 74379 31480 74380 31520
rect 74420 31480 74421 31520
rect 74379 31471 74421 31480
rect 74475 31352 74517 31361
rect 74475 31312 74476 31352
rect 74516 31312 74517 31352
rect 74475 31303 74517 31312
rect 74476 31218 74516 31303
rect 74379 31184 74421 31193
rect 74379 31144 74380 31184
rect 74420 31144 74421 31184
rect 74379 31135 74421 31144
rect 74380 28001 74420 31135
rect 74572 28916 74612 28925
rect 74572 28253 74612 28876
rect 74476 28244 74516 28253
rect 74379 27992 74421 28001
rect 74379 27952 74380 27992
rect 74420 27952 74421 27992
rect 74379 27943 74421 27952
rect 74476 27497 74516 28204
rect 74571 28244 74613 28253
rect 74571 28204 74572 28244
rect 74612 28204 74613 28244
rect 74571 28195 74613 28204
rect 74475 27488 74517 27497
rect 74475 27448 74476 27488
rect 74516 27448 74517 27488
rect 74475 27439 74517 27448
rect 74572 27152 74612 28195
rect 74284 27112 74612 27152
rect 74284 24464 74324 27112
rect 74475 26816 74517 26825
rect 74475 26776 74476 26816
rect 74516 26776 74517 26816
rect 74475 26767 74517 26776
rect 74380 26648 74420 26657
rect 74380 26153 74420 26608
rect 74379 26144 74421 26153
rect 74379 26104 74380 26144
rect 74420 26104 74421 26144
rect 74379 26095 74421 26104
rect 74476 25304 74516 26767
rect 74572 26732 74612 26741
rect 74572 26237 74612 26692
rect 74571 26228 74613 26237
rect 74571 26188 74572 26228
rect 74612 26188 74613 26228
rect 74571 26179 74613 26188
rect 74571 26060 74613 26069
rect 74571 26020 74572 26060
rect 74612 26020 74613 26060
rect 74571 26011 74613 26020
rect 74476 24641 74516 25264
rect 74475 24632 74517 24641
rect 74475 24592 74476 24632
rect 74516 24592 74517 24632
rect 74475 24583 74517 24592
rect 74284 24424 74516 24464
rect 74187 23708 74229 23717
rect 74187 23668 74188 23708
rect 74228 23668 74229 23708
rect 74187 23659 74229 23668
rect 74187 23540 74229 23549
rect 74187 23500 74188 23540
rect 74228 23500 74229 23540
rect 74187 23491 74229 23500
rect 73996 23045 74132 23060
rect 73996 23036 74133 23045
rect 73996 23020 74092 23036
rect 74091 22996 74092 23020
rect 74132 22996 74133 23036
rect 74091 22987 74133 22996
rect 73708 22912 73844 22952
rect 73900 22912 73985 22952
rect 73804 22793 73844 22912
rect 73654 22784 73696 22793
rect 73654 22744 73655 22784
rect 73695 22744 73696 22784
rect 73654 22735 73696 22744
rect 73803 22784 73845 22793
rect 73803 22744 73804 22784
rect 73844 22744 73845 22784
rect 73803 22735 73845 22744
rect 73655 22596 73695 22735
rect 73945 22596 73985 22912
rect 74188 22793 74228 23491
rect 74476 23060 74516 24424
rect 74572 23549 74612 26011
rect 74668 24557 74708 33100
rect 75244 31940 75284 31949
rect 74956 31900 75244 31940
rect 74956 31361 74996 31900
rect 75244 31891 75284 31900
rect 75112 31772 75480 31781
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75112 31723 75480 31732
rect 74955 31352 74997 31361
rect 74955 31312 74956 31352
rect 74996 31312 74997 31352
rect 74955 31303 74997 31312
rect 74860 30848 74900 30857
rect 74860 30596 74900 30808
rect 74764 30556 74900 30596
rect 74764 29849 74804 30556
rect 74956 30269 74996 31303
rect 75052 30680 75092 30689
rect 75052 30521 75092 30640
rect 75435 30680 75477 30689
rect 75435 30640 75436 30680
rect 75476 30640 75477 30680
rect 75435 30631 75477 30640
rect 75436 30546 75476 30631
rect 75051 30512 75093 30521
rect 75051 30472 75052 30512
rect 75092 30472 75093 30512
rect 75051 30463 75093 30472
rect 75531 30428 75573 30437
rect 75531 30388 75532 30428
rect 75572 30388 75573 30428
rect 75531 30379 75573 30388
rect 74955 30260 74997 30269
rect 74955 30220 74956 30260
rect 74996 30220 74997 30260
rect 74955 30211 74997 30220
rect 75112 30260 75480 30269
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75112 30211 75480 30220
rect 75436 29924 75476 29933
rect 74763 29840 74805 29849
rect 74763 29800 74764 29840
rect 74804 29800 74805 29840
rect 74763 29791 74805 29800
rect 74764 28160 74804 29791
rect 75436 29597 75476 29884
rect 75435 29588 75477 29597
rect 75435 29548 75436 29588
rect 75476 29548 75477 29588
rect 75435 29539 75477 29548
rect 75112 28748 75480 28757
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75112 28699 75480 28708
rect 74860 28328 74900 28337
rect 74900 28288 74996 28328
rect 74860 28279 74900 28288
rect 74764 28120 74900 28160
rect 74763 27992 74805 28001
rect 74763 27952 74764 27992
rect 74804 27952 74805 27992
rect 74763 27943 74805 27952
rect 74764 26069 74804 27943
rect 74860 27161 74900 28120
rect 74859 27152 74901 27161
rect 74859 27112 74860 27152
rect 74900 27112 74901 27152
rect 74859 27103 74901 27112
rect 74956 26816 74996 28288
rect 75112 27236 75480 27245
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75112 27187 75480 27196
rect 74956 26741 74996 26776
rect 74955 26732 74997 26741
rect 74955 26692 74956 26732
rect 74996 26692 74997 26732
rect 74955 26683 74997 26692
rect 74859 26648 74901 26657
rect 74859 26608 74860 26648
rect 74900 26608 74901 26648
rect 74859 26599 74901 26608
rect 74763 26060 74805 26069
rect 74763 26020 74764 26060
rect 74804 26020 74805 26060
rect 74763 26011 74805 26020
rect 74860 24632 74900 26599
rect 75243 26480 75285 26489
rect 75243 26440 75244 26480
rect 75284 26440 75285 26480
rect 75243 26431 75285 26440
rect 75244 26060 75284 26431
rect 75244 26011 75284 26020
rect 75435 25976 75477 25985
rect 75435 25936 75436 25976
rect 75476 25936 75477 25976
rect 75435 25927 75477 25936
rect 75436 25842 75476 25927
rect 75112 25724 75480 25733
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75112 25675 75480 25684
rect 75051 25220 75093 25229
rect 75051 25180 75052 25220
rect 75092 25180 75093 25220
rect 75051 25171 75093 25180
rect 74764 24592 74860 24632
rect 74667 24548 74709 24557
rect 74667 24508 74668 24548
rect 74708 24508 74709 24548
rect 74667 24499 74709 24508
rect 74764 23792 74804 24592
rect 74860 24583 74900 24592
rect 74956 24548 74996 24557
rect 74860 24044 74900 24053
rect 74956 24044 74996 24508
rect 75052 24464 75092 25171
rect 75532 24977 75572 30379
rect 75628 30176 75668 33100
rect 75724 30437 75764 33403
rect 76780 32873 76820 32958
rect 76972 32873 77012 34168
rect 77067 34040 77109 34049
rect 77067 34000 77068 34040
rect 77108 34000 77109 34040
rect 77067 33991 77109 34000
rect 77068 33704 77108 33991
rect 77163 33872 77205 33881
rect 77163 33832 77164 33872
rect 77204 33832 77205 33872
rect 77163 33823 77205 33832
rect 77068 33655 77108 33664
rect 77164 33620 77204 33823
rect 77164 33571 77204 33580
rect 77260 33536 77300 35167
rect 77452 34889 77492 35176
rect 77451 34880 77493 34889
rect 77451 34840 77452 34880
rect 77492 34840 77493 34880
rect 77451 34831 77493 34840
rect 77548 34712 77588 35848
rect 77644 35888 77684 35897
rect 77644 35393 77684 35848
rect 77739 35888 77781 35897
rect 77739 35848 77740 35888
rect 77780 35848 77781 35888
rect 77739 35839 77781 35848
rect 78027 35888 78069 35897
rect 78027 35848 78028 35888
rect 78068 35848 78069 35888
rect 78027 35839 78069 35848
rect 77740 35754 77780 35839
rect 78028 35754 78068 35839
rect 77932 35720 77972 35729
rect 77643 35384 77685 35393
rect 77643 35344 77644 35384
rect 77684 35344 77685 35384
rect 77643 35335 77685 35344
rect 77548 34672 77684 34712
rect 77548 34544 77588 34553
rect 77452 34504 77548 34544
rect 77356 34292 77396 34301
rect 77356 33965 77396 34252
rect 77355 33956 77397 33965
rect 77355 33916 77356 33956
rect 77396 33916 77397 33956
rect 77355 33907 77397 33916
rect 77452 33881 77492 34504
rect 77548 34495 77588 34504
rect 77547 34376 77589 34385
rect 77547 34336 77548 34376
rect 77588 34336 77589 34376
rect 77547 34327 77589 34336
rect 77451 33872 77493 33881
rect 77451 33832 77452 33872
rect 77492 33832 77493 33872
rect 77451 33823 77493 33832
rect 77451 33704 77493 33713
rect 77451 33664 77452 33704
rect 77492 33664 77493 33704
rect 77451 33655 77493 33664
rect 77356 33620 77396 33631
rect 77356 33545 77396 33580
rect 77260 33487 77300 33496
rect 77355 33536 77397 33545
rect 77355 33496 77356 33536
rect 77396 33496 77397 33536
rect 77355 33487 77397 33496
rect 77452 33140 77492 33655
rect 77164 33100 77492 33140
rect 77548 33140 77588 34327
rect 77644 33713 77684 34672
rect 77932 34544 77972 35680
rect 78124 35216 78164 36688
rect 79084 36476 79124 36485
rect 79084 35813 79124 36436
rect 79467 35888 79509 35897
rect 79467 35848 79468 35888
rect 79508 35848 79509 35888
rect 79467 35839 79509 35848
rect 79083 35804 79125 35813
rect 79083 35764 79084 35804
rect 79124 35764 79125 35804
rect 79083 35755 79125 35764
rect 79468 35384 79508 35839
rect 79468 35335 79508 35344
rect 78316 35216 78356 35225
rect 78124 35176 78316 35216
rect 78316 34553 78356 35176
rect 78411 35132 78453 35141
rect 78411 35092 78412 35132
rect 78452 35092 78453 35132
rect 78411 35083 78453 35092
rect 78315 34544 78357 34553
rect 77932 34504 78068 34544
rect 78028 34460 78068 34504
rect 78315 34504 78316 34544
rect 78356 34504 78357 34544
rect 78315 34495 78357 34504
rect 78028 34420 78070 34460
rect 77835 34376 77877 34385
rect 77835 34336 77836 34376
rect 77876 34336 77877 34376
rect 77835 34327 77877 34336
rect 77932 34376 77972 34385
rect 77836 34242 77876 34327
rect 77932 34133 77972 34336
rect 78030 34292 78070 34420
rect 78028 34252 78070 34292
rect 78220 34376 78260 34385
rect 78028 34204 78068 34252
rect 77931 34124 77973 34133
rect 77931 34084 77932 34124
rect 77972 34084 77973 34124
rect 77931 34075 77973 34084
rect 78028 34049 78068 34164
rect 78220 34133 78260 34336
rect 78316 34376 78356 34387
rect 78316 34301 78356 34336
rect 78412 34376 78452 35083
rect 78315 34292 78357 34301
rect 78315 34252 78316 34292
rect 78356 34252 78357 34292
rect 78315 34243 78357 34252
rect 78219 34124 78261 34133
rect 78219 34084 78220 34124
rect 78260 34084 78261 34124
rect 78219 34075 78261 34084
rect 78027 34040 78069 34049
rect 78027 34000 78028 34040
rect 78068 34000 78069 34040
rect 78027 33991 78069 34000
rect 77643 33704 77685 33713
rect 77643 33664 77644 33704
rect 77684 33664 77685 33704
rect 77643 33655 77685 33664
rect 77836 33704 77876 33713
rect 77643 33536 77685 33545
rect 77643 33496 77644 33536
rect 77684 33496 77685 33536
rect 77643 33487 77685 33496
rect 77644 33402 77684 33487
rect 77548 33100 77684 33140
rect 76779 32864 76821 32873
rect 76779 32824 76780 32864
rect 76820 32824 76821 32864
rect 76779 32815 76821 32824
rect 76971 32864 77013 32873
rect 76971 32824 76972 32864
rect 77012 32824 77013 32864
rect 76971 32815 77013 32824
rect 76396 32780 76436 32789
rect 76396 32696 76436 32740
rect 76396 32656 76916 32696
rect 76352 32528 76720 32537
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76352 32479 76720 32488
rect 76779 32444 76821 32453
rect 76779 32395 76780 32444
rect 76820 32395 76821 32444
rect 76491 32360 76533 32369
rect 76491 32320 76492 32360
rect 76532 32320 76533 32360
rect 76491 32311 76533 32320
rect 75915 32192 75957 32201
rect 75915 32152 75916 32192
rect 75956 32152 75957 32192
rect 75915 32143 75957 32152
rect 75916 31184 75956 32143
rect 76300 31940 76340 31949
rect 76300 31529 76340 31900
rect 76299 31520 76341 31529
rect 76299 31480 76300 31520
rect 76340 31480 76341 31520
rect 76299 31471 76341 31480
rect 76012 31361 76052 31446
rect 76107 31436 76149 31445
rect 76107 31396 76108 31436
rect 76148 31396 76149 31436
rect 76107 31387 76149 31396
rect 76011 31352 76053 31361
rect 76011 31312 76012 31352
rect 76052 31312 76053 31352
rect 76011 31303 76053 31312
rect 76108 31352 76148 31387
rect 76108 31301 76148 31312
rect 76204 31352 76244 31361
rect 76300 31352 76340 31471
rect 76244 31312 76340 31352
rect 76492 31352 76532 32311
rect 76780 32309 76820 32378
rect 76683 32276 76725 32285
rect 76683 32236 76684 32276
rect 76724 32236 76725 32276
rect 76683 32227 76725 32236
rect 76588 32192 76628 32201
rect 76588 31697 76628 32152
rect 76684 32192 76724 32227
rect 76684 32141 76724 32152
rect 76876 32024 76916 32656
rect 76971 32192 77013 32201
rect 76971 32152 76972 32192
rect 77012 32152 77013 32192
rect 76971 32143 77013 32152
rect 76972 32058 77012 32143
rect 76684 31984 76916 32024
rect 76587 31688 76629 31697
rect 76587 31648 76588 31688
rect 76628 31648 76629 31688
rect 76587 31639 76629 31648
rect 76587 31520 76629 31529
rect 76587 31480 76588 31520
rect 76628 31480 76629 31520
rect 76587 31471 76629 31480
rect 76684 31520 76724 31984
rect 77068 31520 77108 31529
rect 76684 31471 76724 31480
rect 76780 31480 77068 31520
rect 76588 31436 76628 31471
rect 76588 31385 76628 31396
rect 76780 31436 76820 31480
rect 77068 31471 77108 31480
rect 76780 31387 76820 31396
rect 76204 31303 76244 31312
rect 76492 31303 76532 31312
rect 76876 31352 76916 31361
rect 77068 31352 77108 31361
rect 77164 31352 77204 33100
rect 77644 32873 77684 33100
rect 77355 32864 77397 32873
rect 77355 32824 77356 32864
rect 77396 32824 77397 32864
rect 77355 32815 77397 32824
rect 77643 32864 77685 32873
rect 77643 32824 77644 32864
rect 77684 32824 77685 32864
rect 77643 32815 77685 32824
rect 77356 32192 77396 32815
rect 77644 32730 77684 32815
rect 77396 32152 77492 32192
rect 77356 32143 77396 32152
rect 77259 31604 77301 31613
rect 77259 31564 77260 31604
rect 77300 31564 77301 31604
rect 77259 31555 77301 31564
rect 76916 31312 77068 31352
rect 77108 31312 77204 31352
rect 77260 31352 77300 31555
rect 76300 31184 76340 31193
rect 75916 31144 76300 31184
rect 76300 31135 76340 31144
rect 76352 31016 76720 31025
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76352 30967 76720 30976
rect 76299 30680 76341 30689
rect 76299 30640 76300 30680
rect 76340 30640 76341 30680
rect 76299 30631 76341 30640
rect 76300 30546 76340 30631
rect 76011 30512 76053 30521
rect 76011 30472 76012 30512
rect 76052 30472 76053 30512
rect 76011 30463 76053 30472
rect 75723 30428 75765 30437
rect 75723 30388 75724 30428
rect 75764 30388 75765 30428
rect 75723 30379 75765 30388
rect 75628 30136 75764 30176
rect 75627 30008 75669 30017
rect 75627 29968 75628 30008
rect 75668 29968 75669 30008
rect 75627 29959 75669 29968
rect 75628 29874 75668 29959
rect 75724 29084 75764 30136
rect 75819 30008 75861 30017
rect 75819 29968 75820 30008
rect 75860 29968 75861 30008
rect 75819 29959 75861 29968
rect 76012 30008 76052 30463
rect 76876 30017 76916 31312
rect 77068 31303 77108 31312
rect 77260 31268 77300 31312
rect 77145 31228 77300 31268
rect 77356 31352 77396 31361
rect 77145 31184 77185 31228
rect 76972 31144 77185 31184
rect 76396 30008 76436 30017
rect 76012 29959 76052 29968
rect 76108 29968 76396 30008
rect 75820 29840 75860 29959
rect 75820 29261 75860 29800
rect 75916 29924 75956 29933
rect 75916 29345 75956 29884
rect 76108 29924 76148 29968
rect 76396 29959 76436 29968
rect 76875 30008 76917 30017
rect 76875 29968 76876 30008
rect 76916 29968 76917 30008
rect 76875 29959 76917 29968
rect 75915 29336 75957 29345
rect 75915 29296 75916 29336
rect 75956 29296 75957 29336
rect 75915 29287 75957 29296
rect 75819 29252 75861 29261
rect 75819 29212 75820 29252
rect 75860 29212 75861 29252
rect 75819 29203 75861 29212
rect 76108 29177 76148 29884
rect 76779 29924 76821 29933
rect 76779 29884 76780 29924
rect 76820 29884 76821 29924
rect 76779 29875 76821 29884
rect 76204 29840 76244 29851
rect 76204 29765 76244 29800
rect 76683 29840 76725 29849
rect 76683 29800 76684 29840
rect 76724 29800 76725 29840
rect 76683 29791 76725 29800
rect 76780 29840 76820 29875
rect 76203 29756 76245 29765
rect 76203 29716 76204 29756
rect 76244 29716 76245 29756
rect 76203 29707 76245 29716
rect 76684 29706 76724 29791
rect 76780 29789 76820 29800
rect 76875 29756 76917 29765
rect 76875 29716 76876 29756
rect 76916 29716 76917 29756
rect 76875 29707 76917 29716
rect 76876 29668 76916 29707
rect 76876 29619 76916 29628
rect 76352 29504 76720 29513
rect 76972 29504 77012 31144
rect 77259 31100 77301 31109
rect 77259 31060 77260 31100
rect 77300 31060 77301 31100
rect 77259 31051 77301 31060
rect 77260 30605 77300 31051
rect 77356 30848 77396 31312
rect 77452 31109 77492 32152
rect 77547 31688 77589 31697
rect 77547 31648 77548 31688
rect 77588 31648 77589 31688
rect 77547 31639 77589 31648
rect 77548 31352 77588 31639
rect 77836 31613 77876 33664
rect 77932 33704 77972 33713
rect 78219 33704 78261 33713
rect 77972 33664 78220 33704
rect 78260 33664 78261 33704
rect 77932 33655 77972 33664
rect 78219 33655 78261 33664
rect 78220 33570 78260 33655
rect 78124 33452 78164 33461
rect 78124 32453 78164 33412
rect 78219 32864 78261 32873
rect 78219 32824 78220 32864
rect 78260 32824 78261 32864
rect 78219 32815 78261 32824
rect 78123 32444 78165 32453
rect 78123 32404 78124 32444
rect 78164 32404 78165 32444
rect 78123 32395 78165 32404
rect 77931 32276 77973 32285
rect 77931 32236 77932 32276
rect 77972 32236 77973 32276
rect 77931 32227 77973 32236
rect 77835 31604 77877 31613
rect 77835 31564 77836 31604
rect 77876 31564 77877 31604
rect 77835 31555 77877 31564
rect 77548 31303 77588 31312
rect 77643 31352 77685 31361
rect 77643 31312 77644 31352
rect 77684 31312 77685 31352
rect 77643 31303 77685 31312
rect 77740 31352 77780 31363
rect 77644 31218 77684 31303
rect 77740 31277 77780 31312
rect 77836 31352 77876 31361
rect 77932 31352 77972 32227
rect 78220 32192 78260 32815
rect 78123 31940 78165 31949
rect 78123 31900 78124 31940
rect 78164 31900 78165 31940
rect 78123 31891 78165 31900
rect 78027 31436 78069 31445
rect 78027 31396 78028 31436
rect 78068 31396 78069 31436
rect 78027 31387 78069 31396
rect 77876 31312 77972 31352
rect 77739 31268 77781 31277
rect 77739 31228 77740 31268
rect 77780 31228 77781 31268
rect 77739 31219 77781 31228
rect 77451 31100 77493 31109
rect 77451 31060 77452 31100
rect 77492 31060 77493 31100
rect 77451 31051 77493 31060
rect 77452 30848 77492 30857
rect 77356 30808 77452 30848
rect 77492 30808 77684 30848
rect 77452 30799 77492 30808
rect 77644 30680 77684 30808
rect 77644 30631 77684 30640
rect 77259 30596 77301 30605
rect 77259 30556 77260 30596
rect 77300 30556 77301 30596
rect 77259 30547 77301 30556
rect 77451 30596 77493 30605
rect 77451 30556 77452 30596
rect 77492 30556 77493 30596
rect 77451 30547 77493 30556
rect 77259 30260 77301 30269
rect 77259 30220 77260 30260
rect 77300 30220 77301 30260
rect 77259 30211 77301 30220
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76352 29455 76720 29464
rect 76780 29464 77012 29504
rect 77068 29756 77108 29765
rect 76587 29336 76629 29345
rect 76780 29336 76820 29464
rect 76587 29296 76588 29336
rect 76628 29296 76629 29336
rect 76587 29287 76629 29296
rect 76684 29296 76820 29336
rect 76491 29252 76533 29261
rect 76491 29212 76492 29252
rect 76532 29212 76533 29252
rect 76491 29203 76533 29212
rect 76107 29168 76149 29177
rect 76107 29128 76108 29168
rect 76148 29128 76149 29168
rect 76107 29119 76149 29128
rect 76492 29168 76532 29203
rect 76588 29202 76628 29287
rect 76492 29117 76532 29128
rect 76684 29168 76724 29296
rect 76972 29261 77012 29346
rect 77068 29345 77108 29716
rect 77067 29336 77109 29345
rect 77067 29296 77068 29336
rect 77108 29296 77109 29336
rect 77067 29287 77109 29296
rect 76971 29252 77013 29261
rect 76971 29212 76972 29252
rect 77012 29212 77013 29252
rect 76971 29203 77013 29212
rect 76684 29119 76724 29128
rect 76780 29168 76820 29177
rect 75724 29044 75860 29084
rect 75723 28328 75765 28337
rect 75723 28288 75724 28328
rect 75764 28288 75765 28328
rect 75723 28279 75765 28288
rect 75724 28194 75764 28279
rect 75723 27656 75765 27665
rect 75628 27616 75724 27656
rect 75764 27616 75765 27656
rect 75628 26144 75668 27616
rect 75723 27607 75765 27616
rect 75724 27522 75764 27607
rect 75723 27404 75765 27413
rect 75723 27364 75724 27404
rect 75764 27364 75765 27404
rect 75723 27355 75765 27364
rect 75724 27270 75764 27355
rect 75820 27236 75860 29044
rect 76780 28580 76820 29128
rect 77067 29168 77109 29177
rect 77067 29120 77068 29168
rect 77108 29120 77109 29168
rect 77260 29168 77300 30211
rect 77355 29840 77397 29849
rect 77355 29800 77356 29840
rect 77396 29800 77397 29840
rect 77355 29791 77397 29800
rect 77452 29840 77492 30547
rect 77452 29791 77492 29800
rect 77740 30428 77780 30437
rect 77356 29336 77396 29791
rect 77740 29765 77780 30388
rect 77836 29933 77876 31312
rect 78028 31184 78068 31387
rect 78124 31352 78164 31891
rect 78124 31277 78164 31312
rect 78123 31268 78165 31277
rect 78123 31228 78124 31268
rect 78164 31228 78165 31268
rect 78123 31219 78165 31228
rect 78028 30269 78068 31144
rect 78027 30260 78069 30269
rect 78027 30220 78028 30260
rect 78068 30220 78069 30260
rect 78027 30211 78069 30220
rect 77835 29924 77877 29933
rect 77835 29884 77836 29924
rect 77876 29884 77877 29924
rect 77835 29875 77877 29884
rect 77739 29756 77781 29765
rect 77739 29716 77740 29756
rect 77780 29716 77781 29756
rect 77739 29707 77781 29716
rect 77452 29336 77492 29345
rect 77356 29296 77452 29336
rect 77452 29287 77492 29296
rect 77548 29168 77588 29177
rect 77067 29119 77109 29120
rect 77164 29126 77204 29135
rect 77068 29033 77108 29119
rect 77300 29128 77548 29168
rect 77260 29119 77300 29128
rect 77548 29119 77588 29128
rect 77643 29168 77685 29177
rect 77643 29128 77644 29168
rect 77684 29128 77685 29168
rect 77643 29119 77685 29128
rect 77740 29168 77780 29177
rect 77836 29168 77876 29875
rect 77780 29128 77876 29168
rect 78027 29168 78069 29177
rect 78027 29128 78028 29168
rect 78068 29128 78069 29168
rect 77740 29119 77780 29128
rect 78027 29119 78069 29128
rect 77164 28925 77204 29086
rect 77644 29034 77684 29119
rect 78028 29034 78068 29119
rect 77163 28916 77205 28925
rect 77163 28876 77164 28916
rect 77204 28876 77205 28916
rect 77163 28867 77205 28876
rect 77931 28916 77973 28925
rect 78124 28916 78164 31219
rect 78220 30689 78260 32152
rect 78412 31361 78452 34336
rect 78507 34376 78549 34385
rect 78507 34336 78508 34376
rect 78548 34336 78549 34376
rect 78507 34327 78549 34336
rect 78508 34242 78548 34327
rect 78795 33704 78837 33713
rect 78795 33664 78796 33704
rect 78836 33664 78837 33704
rect 78795 33655 78837 33664
rect 78796 33116 78836 33655
rect 78796 33067 78836 33076
rect 79371 31940 79413 31949
rect 79371 31900 79372 31940
rect 79412 31900 79413 31940
rect 79371 31891 79413 31900
rect 79372 31806 79412 31891
rect 78411 31352 78453 31361
rect 78411 31312 78412 31352
rect 78452 31312 78453 31352
rect 78411 31303 78453 31312
rect 78219 30680 78261 30689
rect 78219 30640 78220 30680
rect 78260 30640 78261 30680
rect 78219 30631 78261 30640
rect 78220 29840 78260 30631
rect 78316 29840 78356 29849
rect 78220 29800 78316 29840
rect 78316 29791 78356 29800
rect 79468 29672 79508 29681
rect 79468 29177 79508 29632
rect 78699 29168 78741 29177
rect 78699 29128 78700 29168
rect 78740 29128 78741 29168
rect 78699 29119 78741 29128
rect 79467 29168 79509 29177
rect 79467 29128 79468 29168
rect 79508 29128 79509 29168
rect 79467 29119 79509 29128
rect 77931 28876 77932 28916
rect 77972 28876 77973 28916
rect 77931 28867 77973 28876
rect 78028 28876 78164 28916
rect 77932 28782 77972 28867
rect 76876 28580 76916 28589
rect 76780 28540 76876 28580
rect 76876 28337 76916 28540
rect 77068 28496 77108 28505
rect 77068 28412 77108 28456
rect 77068 28372 77300 28412
rect 76875 28328 76917 28337
rect 76875 28288 76876 28328
rect 76916 28288 76917 28328
rect 76875 28279 76917 28288
rect 76352 27992 76720 28001
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76352 27943 76720 27952
rect 76876 27749 76916 27780
rect 76011 27740 76053 27749
rect 76011 27700 76012 27740
rect 76052 27700 76053 27740
rect 76011 27691 76053 27700
rect 76875 27740 76917 27749
rect 76875 27700 76876 27740
rect 76916 27700 76917 27740
rect 76875 27691 76917 27700
rect 75916 27656 75956 27667
rect 75916 27581 75956 27616
rect 76012 27656 76052 27691
rect 76012 27605 76052 27616
rect 76203 27656 76245 27665
rect 76203 27616 76204 27656
rect 76244 27616 76245 27656
rect 76203 27607 76245 27616
rect 76587 27656 76629 27665
rect 76587 27616 76588 27656
rect 76628 27616 76629 27656
rect 76587 27607 76629 27616
rect 76876 27656 76916 27691
rect 75915 27572 75957 27581
rect 75915 27532 75916 27572
rect 75956 27532 75957 27572
rect 75915 27523 75957 27532
rect 76107 27572 76149 27581
rect 76107 27532 76108 27572
rect 76148 27532 76149 27572
rect 76107 27523 76149 27532
rect 76108 27320 76148 27523
rect 76204 27522 76244 27607
rect 76300 27572 76340 27581
rect 76300 27413 76340 27532
rect 76491 27572 76533 27581
rect 76491 27532 76492 27572
rect 76532 27532 76533 27572
rect 76491 27523 76533 27532
rect 76395 27488 76437 27497
rect 76395 27448 76396 27488
rect 76436 27448 76437 27488
rect 76395 27439 76437 27448
rect 76299 27404 76341 27413
rect 76299 27364 76300 27404
rect 76340 27364 76341 27404
rect 76299 27355 76341 27364
rect 76396 27354 76436 27439
rect 76492 27438 76532 27523
rect 76588 27522 76628 27607
rect 76780 27404 76820 27413
rect 76108 27280 76244 27320
rect 75820 27196 76148 27236
rect 75819 26816 75861 26825
rect 75819 26776 75820 26816
rect 75860 26776 75861 26816
rect 75819 26767 75861 26776
rect 75820 26682 75860 26767
rect 75819 26228 75861 26237
rect 75819 26188 75820 26228
rect 75860 26188 75861 26228
rect 75819 26179 75861 26188
rect 75628 25985 75668 26104
rect 75724 26060 75764 26069
rect 75627 25976 75669 25985
rect 75627 25936 75628 25976
rect 75668 25936 75669 25976
rect 75627 25927 75669 25936
rect 75628 25472 75668 25927
rect 75724 25556 75764 26020
rect 75820 25976 75860 26179
rect 76011 26144 76053 26153
rect 76011 26104 76012 26144
rect 76052 26104 76053 26144
rect 76011 26095 76053 26104
rect 75916 26060 75956 26071
rect 75916 25985 75956 26020
rect 76012 26010 76052 26095
rect 75820 25927 75860 25936
rect 75915 25976 75957 25985
rect 75915 25936 75916 25976
rect 75956 25936 75957 25976
rect 75915 25927 75957 25936
rect 76108 25724 76148 27196
rect 76204 26144 76244 27280
rect 76352 26480 76720 26489
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76352 26431 76720 26440
rect 76587 26312 76629 26321
rect 76587 26272 76588 26312
rect 76628 26272 76629 26312
rect 76587 26263 76629 26272
rect 76684 26316 76724 26325
rect 76780 26312 76820 27364
rect 76876 27068 76916 27616
rect 77068 27656 77108 27665
rect 76972 27068 77012 27077
rect 76876 27028 76972 27068
rect 76972 27019 77012 27028
rect 77068 26816 77108 27616
rect 77260 27581 77300 28372
rect 77356 28328 77396 28337
rect 77259 27572 77301 27581
rect 77259 27532 77260 27572
rect 77300 27532 77301 27572
rect 77259 27523 77301 27532
rect 77164 26816 77204 26825
rect 77068 26776 77164 26816
rect 77164 26767 77204 26776
rect 77260 26816 77300 27523
rect 77356 27488 77396 28288
rect 77452 28328 77492 28337
rect 77739 28328 77781 28337
rect 77492 28288 77684 28328
rect 77452 28279 77492 28288
rect 77548 28102 77588 28111
rect 77451 28076 77493 28085
rect 77451 28036 77452 28076
rect 77492 28036 77493 28076
rect 77451 28027 77493 28036
rect 77452 27656 77492 28027
rect 77548 27665 77588 28062
rect 77452 27607 77492 27616
rect 77547 27656 77589 27665
rect 77547 27616 77548 27656
rect 77588 27616 77589 27656
rect 77547 27607 77589 27616
rect 77644 27572 77684 28288
rect 77739 28288 77740 28328
rect 77780 28288 77781 28328
rect 77739 28279 77781 28288
rect 77740 28194 77780 28279
rect 77836 28160 77876 28169
rect 77836 27665 77876 28120
rect 77835 27656 77877 27665
rect 77835 27616 77836 27656
rect 77876 27616 77877 27656
rect 77835 27607 77877 27616
rect 77644 27532 77780 27572
rect 77356 27448 77684 27488
rect 77260 26767 77300 26776
rect 77355 26816 77397 26825
rect 77355 26776 77356 26816
rect 77396 26776 77397 26816
rect 77355 26767 77397 26776
rect 77452 26816 77492 26825
rect 77356 26682 77396 26767
rect 76724 26276 76820 26312
rect 76684 26272 76820 26276
rect 77452 26648 77492 26776
rect 77644 26816 77684 27448
rect 77740 27077 77780 27532
rect 77835 27404 77877 27413
rect 77835 27364 77836 27404
rect 77876 27364 77877 27404
rect 77835 27355 77877 27364
rect 77739 27068 77781 27077
rect 77739 27028 77740 27068
rect 77780 27028 77781 27068
rect 77739 27019 77781 27028
rect 77644 26767 77684 26776
rect 77740 26816 77780 26825
rect 77740 26648 77780 26776
rect 77836 26816 77876 27355
rect 77931 27068 77973 27077
rect 77931 27028 77932 27068
rect 77972 27028 77973 27068
rect 77931 27019 77973 27028
rect 77836 26767 77876 26776
rect 77932 26816 77972 27019
rect 77452 26608 77780 26648
rect 77835 26648 77877 26657
rect 77835 26608 77836 26648
rect 77876 26608 77877 26648
rect 76492 26144 76532 26153
rect 76204 26104 76340 26144
rect 76203 25976 76245 25985
rect 76203 25936 76204 25976
rect 76244 25936 76245 25976
rect 76203 25927 76245 25936
rect 76204 25842 76244 25927
rect 76108 25684 76244 25724
rect 76108 25556 76148 25565
rect 75724 25516 76108 25556
rect 76108 25507 76148 25516
rect 75628 25432 76052 25472
rect 75820 25304 75860 25313
rect 75628 25136 75668 25145
rect 75820 25136 75860 25264
rect 75915 25304 75957 25313
rect 75915 25264 75916 25304
rect 75956 25264 75957 25304
rect 76012 25304 76052 25432
rect 76108 25304 76148 25313
rect 76012 25264 76108 25304
rect 75915 25255 75957 25264
rect 76108 25255 76148 25264
rect 75916 25170 75956 25255
rect 76204 25136 76244 25684
rect 76300 25313 76340 26104
rect 76492 25313 76532 26104
rect 76588 26144 76628 26263
rect 76684 26153 76724 26272
rect 76588 26095 76628 26104
rect 76683 26144 76725 26153
rect 76876 26144 76916 26153
rect 76683 26104 76684 26144
rect 76724 26104 76725 26144
rect 76683 26095 76725 26104
rect 76780 26104 76876 26144
rect 76299 25304 76341 25313
rect 76299 25264 76300 25304
rect 76340 25264 76341 25304
rect 76299 25255 76341 25264
rect 76491 25304 76533 25313
rect 76491 25264 76492 25304
rect 76532 25264 76533 25304
rect 76491 25255 76533 25264
rect 76780 25304 76820 26104
rect 76876 26095 76916 26104
rect 77259 26144 77301 26153
rect 77259 26104 77260 26144
rect 77300 26104 77301 26144
rect 77259 26095 77301 26104
rect 77260 26010 77300 26095
rect 76875 25976 76917 25985
rect 76875 25936 76876 25976
rect 76916 25936 76917 25976
rect 76875 25927 76917 25936
rect 76780 25255 76820 25264
rect 76876 25304 76916 25927
rect 77452 25472 77492 26608
rect 77835 26599 77877 26608
rect 77739 26480 77781 26489
rect 77739 26440 77740 26480
rect 77780 26440 77781 26480
rect 77739 26431 77781 26440
rect 77643 26312 77685 26321
rect 77643 26272 77644 26312
rect 77684 26272 77685 26312
rect 77643 26263 77685 26272
rect 77260 25432 77492 25472
rect 76876 25255 76916 25264
rect 76972 25304 77012 25315
rect 76972 25229 77012 25264
rect 77068 25304 77108 25313
rect 77260 25304 77300 25432
rect 77108 25264 77300 25304
rect 77355 25304 77397 25313
rect 77355 25264 77356 25304
rect 77396 25264 77397 25304
rect 76971 25220 77013 25229
rect 76971 25180 76972 25220
rect 77012 25180 77013 25220
rect 76971 25171 77013 25180
rect 75668 25096 75860 25136
rect 76012 25096 76244 25136
rect 76875 25136 76917 25145
rect 76875 25096 76876 25136
rect 76916 25096 76917 25136
rect 75628 25087 75668 25096
rect 75531 24968 75573 24977
rect 75531 24928 75532 24968
rect 75572 24928 75573 24968
rect 75531 24919 75573 24928
rect 75436 24804 75476 24813
rect 75244 24725 75284 24756
rect 75436 24725 75476 24764
rect 75531 24800 75573 24809
rect 75531 24760 75532 24800
rect 75572 24760 75573 24800
rect 75531 24751 75573 24760
rect 75243 24716 75285 24725
rect 75243 24676 75244 24716
rect 75284 24676 75285 24716
rect 75243 24667 75285 24676
rect 75435 24716 75477 24725
rect 75435 24676 75436 24716
rect 75476 24676 75477 24716
rect 75435 24667 75477 24676
rect 75244 24632 75284 24667
rect 75147 24548 75189 24557
rect 75147 24508 75148 24548
rect 75188 24508 75189 24548
rect 75147 24499 75189 24508
rect 75052 24415 75092 24424
rect 75148 24414 75188 24499
rect 75244 24389 75284 24592
rect 75532 24632 75572 24751
rect 75532 24583 75572 24592
rect 75627 24632 75669 24641
rect 75627 24592 75628 24632
rect 75668 24592 75669 24632
rect 75627 24583 75669 24592
rect 75628 24498 75668 24583
rect 75435 24464 75477 24473
rect 75435 24424 75436 24464
rect 75476 24424 75477 24464
rect 75435 24415 75477 24424
rect 75243 24380 75285 24389
rect 75243 24340 75244 24380
rect 75284 24340 75285 24380
rect 75243 24331 75285 24340
rect 75051 24296 75093 24305
rect 75051 24256 75052 24296
rect 75092 24256 75093 24296
rect 75051 24247 75093 24256
rect 74900 24004 74996 24044
rect 74860 23995 74900 24004
rect 74860 23792 74900 23801
rect 74764 23752 74860 23792
rect 74860 23743 74900 23752
rect 75052 23792 75092 24247
rect 75148 23801 75188 23886
rect 75436 23876 75476 24415
rect 75531 24380 75573 24389
rect 75531 24340 75532 24380
rect 75572 24340 75573 24380
rect 75531 24331 75573 24340
rect 75532 24044 75572 24331
rect 75532 23995 75572 24004
rect 75436 23836 75572 23876
rect 75052 23743 75092 23752
rect 75147 23792 75189 23801
rect 75147 23752 75148 23792
rect 75188 23752 75189 23792
rect 75147 23743 75189 23752
rect 75435 23708 75477 23717
rect 75435 23668 75436 23708
rect 75476 23668 75477 23708
rect 75435 23659 75477 23668
rect 74859 23624 74901 23633
rect 74859 23584 74860 23624
rect 74900 23584 74901 23624
rect 74859 23575 74901 23584
rect 74571 23540 74613 23549
rect 74571 23500 74572 23540
rect 74612 23500 74613 23540
rect 74571 23491 74613 23500
rect 74344 23036 74386 23045
rect 74344 22996 74345 23036
rect 74385 22996 74386 23036
rect 74344 22987 74386 22996
rect 74455 23020 74516 23060
rect 74054 22784 74096 22793
rect 74054 22744 74055 22784
rect 74095 22744 74096 22784
rect 74054 22735 74096 22744
rect 74187 22784 74229 22793
rect 74187 22744 74188 22784
rect 74228 22744 74229 22784
rect 74187 22735 74229 22744
rect 74055 22596 74095 22735
rect 74345 22596 74385 22987
rect 74455 22596 74495 23020
rect 74860 22868 74900 23575
rect 75147 23540 75189 23549
rect 75147 23500 75148 23540
rect 75188 23500 75189 23540
rect 75147 23491 75189 23500
rect 75148 23060 75188 23491
rect 74855 22828 74900 22868
rect 75145 23020 75188 23060
rect 75254 23036 75296 23045
rect 74744 22784 74786 22793
rect 74744 22744 74745 22784
rect 74785 22744 74786 22784
rect 74744 22735 74786 22744
rect 74745 22596 74785 22735
rect 74855 22596 74895 22828
rect 75145 22596 75185 23020
rect 75254 22996 75255 23036
rect 75295 22996 75296 23036
rect 75254 22987 75296 22996
rect 75255 22596 75295 22987
rect 75436 22784 75476 23659
rect 75532 23060 75572 23836
rect 75628 23792 75668 23801
rect 75724 23792 75764 25096
rect 75819 24968 75861 24977
rect 75819 24928 75820 24968
rect 75860 24928 75861 24968
rect 75819 24919 75861 24928
rect 75820 24296 75860 24919
rect 75915 24548 75957 24557
rect 75915 24508 75916 24548
rect 75956 24508 75957 24548
rect 75915 24499 75957 24508
rect 75916 24464 75956 24499
rect 75916 24413 75956 24424
rect 75820 24256 75956 24296
rect 75819 24128 75861 24137
rect 75819 24088 75820 24128
rect 75860 24088 75861 24128
rect 75819 24079 75861 24088
rect 75668 23752 75764 23792
rect 75628 23743 75668 23752
rect 75532 23020 75695 23060
rect 75436 22744 75585 22784
rect 75545 22596 75585 22744
rect 75655 22596 75695 23020
rect 75820 22793 75860 24079
rect 75916 23060 75956 24256
rect 76012 24137 76052 25096
rect 76875 25087 76917 25096
rect 76352 24968 76720 24977
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76352 24919 76720 24928
rect 76203 24884 76245 24893
rect 76203 24844 76204 24884
rect 76244 24844 76245 24884
rect 76203 24835 76245 24844
rect 76107 24548 76149 24557
rect 76107 24508 76108 24548
rect 76148 24508 76149 24548
rect 76107 24499 76149 24508
rect 76204 24548 76244 24835
rect 76683 24800 76725 24809
rect 76683 24760 76684 24800
rect 76724 24760 76725 24800
rect 76683 24751 76725 24760
rect 76395 24716 76437 24725
rect 76395 24676 76396 24716
rect 76436 24676 76437 24716
rect 76395 24667 76437 24676
rect 76204 24499 76244 24508
rect 76011 24128 76053 24137
rect 76011 24088 76012 24128
rect 76052 24088 76053 24128
rect 76011 24079 76053 24088
rect 76108 23792 76148 24499
rect 76396 24380 76436 24667
rect 76588 24632 76628 24641
rect 76204 23792 76244 23801
rect 76108 23752 76204 23792
rect 76204 23743 76244 23752
rect 76300 23792 76340 23801
rect 76107 23624 76149 23633
rect 76107 23584 76108 23624
rect 76148 23584 76149 23624
rect 76107 23575 76149 23584
rect 76108 23490 76148 23575
rect 76300 23381 76340 23752
rect 76396 23792 76436 24340
rect 76396 23743 76436 23752
rect 76492 24592 76588 24632
rect 76492 23633 76532 24592
rect 76588 24583 76628 24592
rect 76684 24464 76724 24751
rect 76588 24424 76724 24464
rect 76588 23792 76628 24424
rect 76779 24044 76821 24053
rect 76779 24004 76780 24044
rect 76820 24004 76821 24044
rect 76779 23995 76821 24004
rect 76683 23960 76725 23969
rect 76683 23920 76684 23960
rect 76724 23920 76725 23960
rect 76683 23911 76725 23920
rect 76588 23743 76628 23752
rect 76684 23792 76724 23911
rect 76684 23743 76724 23752
rect 76780 23792 76820 23995
rect 76876 23792 76916 25087
rect 76971 25052 77013 25061
rect 76971 25012 76972 25052
rect 77012 25012 77013 25052
rect 76971 25003 77013 25012
rect 76972 24632 77012 25003
rect 77068 24809 77108 25264
rect 77355 25255 77397 25264
rect 77452 25304 77492 25313
rect 77356 25170 77396 25255
rect 77067 24800 77109 24809
rect 77067 24760 77068 24800
rect 77108 24760 77109 24800
rect 77067 24751 77109 24760
rect 76972 24583 77012 24592
rect 77067 24632 77109 24641
rect 77067 24592 77068 24632
rect 77108 24592 77109 24632
rect 77067 24583 77109 24592
rect 76876 23752 77012 23792
rect 76780 23743 76820 23752
rect 76491 23624 76533 23633
rect 76491 23584 76492 23624
rect 76532 23584 76533 23624
rect 76491 23575 76533 23584
rect 76875 23624 76917 23633
rect 76875 23584 76876 23624
rect 76916 23584 76917 23624
rect 76875 23575 76917 23584
rect 76395 23540 76437 23549
rect 76395 23500 76396 23540
rect 76436 23500 76437 23540
rect 76395 23491 76437 23500
rect 76299 23372 76341 23381
rect 76299 23332 76300 23372
rect 76340 23332 76341 23372
rect 76299 23323 76341 23332
rect 76299 23204 76341 23213
rect 76299 23164 76300 23204
rect 76340 23164 76341 23204
rect 76299 23155 76341 23164
rect 75916 23020 75985 23060
rect 75819 22784 75861 22793
rect 75819 22744 75820 22784
rect 75860 22744 75861 22784
rect 75819 22735 75861 22744
rect 75945 22596 75985 23020
rect 76054 22784 76096 22793
rect 76054 22744 76055 22784
rect 76095 22744 76096 22784
rect 76300 22784 76340 23155
rect 76396 22868 76436 23491
rect 76876 23490 76916 23575
rect 76972 23060 77012 23752
rect 77068 23633 77108 24583
rect 77452 24053 77492 25264
rect 77547 25304 77589 25313
rect 77547 25264 77548 25304
rect 77588 25264 77589 25304
rect 77547 25255 77589 25264
rect 77644 25304 77684 26263
rect 77644 25255 77684 25264
rect 77548 25170 77588 25255
rect 77451 24044 77493 24053
rect 77451 24004 77452 24044
rect 77492 24004 77493 24044
rect 77451 23995 77493 24004
rect 77259 23960 77301 23969
rect 77259 23920 77260 23960
rect 77300 23920 77301 23960
rect 77259 23911 77301 23920
rect 77260 23792 77300 23911
rect 77260 23743 77300 23752
rect 77067 23624 77109 23633
rect 77067 23584 77068 23624
rect 77108 23584 77109 23624
rect 77067 23575 77109 23584
rect 77164 23624 77204 23633
rect 77164 23381 77204 23584
rect 77259 23624 77301 23633
rect 77259 23584 77260 23624
rect 77300 23584 77301 23624
rect 77259 23575 77301 23584
rect 77163 23372 77205 23381
rect 77163 23332 77164 23372
rect 77204 23332 77205 23372
rect 77163 23323 77205 23332
rect 77260 23060 77300 23575
rect 77740 23060 77780 26431
rect 77836 26144 77876 26599
rect 77932 26321 77972 26776
rect 78028 26489 78068 28876
rect 78316 27656 78356 27665
rect 78220 27616 78316 27656
rect 78123 27068 78165 27077
rect 78123 27028 78124 27068
rect 78164 27028 78165 27068
rect 78123 27019 78165 27028
rect 78124 26934 78164 27019
rect 78220 26657 78260 27616
rect 78316 27607 78356 27616
rect 78603 27404 78645 27413
rect 78603 27364 78604 27404
rect 78644 27364 78645 27404
rect 78603 27355 78645 27364
rect 78315 27320 78357 27329
rect 78315 27280 78316 27320
rect 78356 27280 78357 27320
rect 78315 27271 78357 27280
rect 78316 26900 78356 27271
rect 78316 26851 78356 26860
rect 78507 26816 78549 26825
rect 78507 26776 78508 26816
rect 78548 26776 78549 26816
rect 78507 26767 78549 26776
rect 78604 26816 78644 27355
rect 78219 26648 78261 26657
rect 78219 26608 78220 26648
rect 78260 26608 78261 26648
rect 78219 26599 78261 26608
rect 78508 26648 78548 26767
rect 78027 26480 78069 26489
rect 78027 26440 78028 26480
rect 78068 26440 78069 26480
rect 78027 26431 78069 26440
rect 77931 26312 77973 26321
rect 77931 26272 77932 26312
rect 77972 26272 77973 26312
rect 77931 26263 77973 26272
rect 78124 26144 78164 26153
rect 77836 26104 78124 26144
rect 77836 24632 77876 26104
rect 78124 26095 78164 26104
rect 78508 25472 78548 26608
rect 78316 25432 78548 25472
rect 78219 25304 78261 25313
rect 78219 25264 78220 25304
rect 78260 25264 78261 25304
rect 78219 25255 78261 25264
rect 78123 25136 78165 25145
rect 78123 25096 78124 25136
rect 78164 25096 78165 25136
rect 78123 25087 78165 25096
rect 78124 25002 78164 25087
rect 77836 24583 77876 24592
rect 76745 23020 77012 23060
rect 77255 23020 77300 23060
rect 77544 23036 77586 23045
rect 76396 22828 76495 22868
rect 76300 22744 76385 22784
rect 76054 22735 76096 22744
rect 76055 22596 76095 22735
rect 76345 22596 76385 22744
rect 76455 22596 76495 22828
rect 76745 22596 76785 23020
rect 76854 22784 76896 22793
rect 76854 22744 76855 22784
rect 76895 22744 76896 22784
rect 76854 22735 76896 22744
rect 77144 22784 77186 22793
rect 77144 22744 77145 22784
rect 77185 22744 77186 22784
rect 77144 22735 77186 22744
rect 76855 22596 76895 22735
rect 77145 22596 77185 22735
rect 77255 22596 77295 23020
rect 77544 22996 77545 23036
rect 77585 22996 77586 23036
rect 77544 22987 77586 22996
rect 77655 23020 77780 23060
rect 77545 22596 77585 22987
rect 77655 22596 77695 23020
rect 78220 22961 78260 25255
rect 78316 23060 78356 25432
rect 78604 25388 78644 26776
rect 78508 25348 78644 25388
rect 78508 23060 78548 25348
rect 78700 25304 78740 29119
rect 79467 27404 79509 27413
rect 79467 27364 79468 27404
rect 79508 27364 79509 27404
rect 79467 27355 79509 27364
rect 79468 27270 79508 27355
rect 79276 25892 79316 25901
rect 79276 25313 79316 25852
rect 78316 23020 78385 23060
rect 78219 22952 78261 22961
rect 78219 22912 78220 22952
rect 78260 22912 78261 22952
rect 78219 22903 78261 22912
rect 77944 22784 77986 22793
rect 77944 22744 77945 22784
rect 77985 22744 77986 22784
rect 77944 22735 77986 22744
rect 78054 22784 78096 22793
rect 78054 22744 78055 22784
rect 78095 22744 78096 22784
rect 78054 22735 78096 22744
rect 77945 22596 77985 22735
rect 78055 22596 78095 22735
rect 78345 22596 78385 23020
rect 78455 23020 78548 23060
rect 78604 25264 78740 25304
rect 79275 25304 79317 25313
rect 79275 25264 79276 25304
rect 79316 25264 79317 25304
rect 78455 22596 78495 23020
rect 78604 22793 78644 25264
rect 79275 25255 79317 25264
rect 78891 25136 78933 25145
rect 78891 25096 78892 25136
rect 78932 25096 78933 25136
rect 78891 25087 78933 25096
rect 78796 23792 78836 23801
rect 78796 23633 78836 23752
rect 78700 23624 78740 23633
rect 78700 23213 78740 23584
rect 78795 23624 78837 23633
rect 78795 23584 78796 23624
rect 78836 23584 78837 23624
rect 78795 23575 78837 23584
rect 78699 23204 78741 23213
rect 78699 23164 78700 23204
rect 78740 23164 78741 23204
rect 78699 23155 78741 23164
rect 78892 23060 78932 25087
rect 78988 24548 79028 24557
rect 78988 23969 79028 24508
rect 78987 23960 79029 23969
rect 78987 23920 78988 23960
rect 79028 23920 79316 23960
rect 78987 23911 79029 23920
rect 78987 23792 79029 23801
rect 78987 23752 78988 23792
rect 79028 23752 79029 23792
rect 78987 23743 79029 23752
rect 78988 23658 79028 23743
rect 79083 23624 79125 23633
rect 79083 23584 79084 23624
rect 79124 23584 79125 23624
rect 79083 23575 79125 23584
rect 79084 23490 79124 23575
rect 79083 23372 79125 23381
rect 79083 23332 79084 23372
rect 79124 23332 79125 23372
rect 79083 23323 79125 23332
rect 78796 23020 78932 23060
rect 79084 23060 79124 23323
rect 79276 23060 79316 23920
rect 79563 23624 79605 23633
rect 79563 23584 79564 23624
rect 79604 23584 79605 23624
rect 79563 23575 79605 23584
rect 79564 23060 79604 23575
rect 79084 23020 79185 23060
rect 78796 22868 78836 23020
rect 78891 22952 78933 22961
rect 78891 22912 78892 22952
rect 78932 22912 78933 22952
rect 78891 22903 78933 22912
rect 78745 22828 78836 22868
rect 78603 22784 78645 22793
rect 78603 22744 78604 22784
rect 78644 22744 78645 22784
rect 78603 22735 78645 22744
rect 78745 22596 78785 22828
rect 78892 22784 78932 22903
rect 78855 22744 78932 22784
rect 78855 22596 78895 22744
rect 79145 22596 79185 23020
rect 79255 23020 79316 23060
rect 79545 23020 79604 23060
rect 79654 23036 79696 23045
rect 79255 22596 79295 23020
rect 79545 22596 79585 23020
rect 79654 22996 79655 23036
rect 79695 22996 79696 23036
rect 79654 22987 79696 22996
rect 79655 22596 79695 22987
rect 53067 21608 53109 21617
rect 53067 21568 53068 21608
rect 53108 21568 53109 21608
rect 53067 21559 53109 21568
rect 53067 18668 53109 18677
rect 53067 18628 53068 18668
rect 53108 18628 53109 18668
rect 53067 18619 53109 18628
rect 53068 17417 53108 18619
rect 53067 17408 53109 17417
rect 53067 17368 53068 17408
rect 53108 17368 53109 17408
rect 53067 17359 53109 17368
rect 52875 17240 52917 17249
rect 52875 17200 52876 17240
rect 52916 17200 53108 17240
rect 52875 17191 52917 17200
rect 52779 17072 52821 17081
rect 52779 17032 52780 17072
rect 52820 17032 52821 17072
rect 52779 17023 52821 17032
rect 52587 16988 52629 16997
rect 52587 16948 52588 16988
rect 52628 16948 52629 16988
rect 52587 16939 52629 16948
rect 52299 16904 52341 16913
rect 52299 16864 52300 16904
rect 52340 16864 52341 16904
rect 52299 16855 52341 16864
rect 52011 16820 52053 16829
rect 52011 16780 52012 16820
rect 52052 16780 52053 16820
rect 52011 16771 52053 16780
rect 52684 16820 52724 16831
rect 52684 16745 52724 16780
rect 52683 16736 52725 16745
rect 52683 16696 52684 16736
rect 52724 16696 52725 16736
rect 52683 16687 52725 16696
rect 52780 16577 52820 17023
rect 52587 16568 52629 16577
rect 52587 16528 52588 16568
rect 52628 16528 52629 16568
rect 52587 16519 52629 16528
rect 52779 16568 52821 16577
rect 52779 16528 52780 16568
rect 52820 16528 52821 16568
rect 52779 16519 52821 16528
rect 52203 16232 52245 16241
rect 52203 16192 52204 16232
rect 52244 16192 52245 16232
rect 52203 16183 52245 16192
rect 52204 16098 52244 16183
rect 52588 16157 52628 16519
rect 52876 16232 52916 16241
rect 52492 16148 52532 16157
rect 52299 16064 52341 16073
rect 52299 16024 52300 16064
rect 52340 16024 52341 16064
rect 52299 16015 52341 16024
rect 52300 15930 52340 16015
rect 51915 15812 51957 15821
rect 51915 15772 51916 15812
rect 51956 15772 51957 15812
rect 51915 15763 51957 15772
rect 52300 15728 52340 15737
rect 52492 15728 52532 16108
rect 52587 16148 52629 16157
rect 52587 16108 52588 16148
rect 52628 16108 52629 16148
rect 52587 16099 52629 16108
rect 52340 15688 52532 15728
rect 52587 15728 52629 15737
rect 52587 15688 52588 15728
rect 52628 15688 52629 15728
rect 52300 15679 52340 15688
rect 52587 15679 52629 15688
rect 52396 15560 52436 15569
rect 51819 15140 51861 15149
rect 51819 15100 51820 15140
rect 51860 15100 51861 15140
rect 51819 15091 51861 15100
rect 51723 14972 51765 14981
rect 52300 14972 52340 14981
rect 52396 14972 52436 15520
rect 52492 15560 52532 15569
rect 52492 14981 52532 15520
rect 52588 15560 52628 15679
rect 52588 15485 52628 15520
rect 52587 15476 52629 15485
rect 52587 15436 52588 15476
rect 52628 15436 52629 15476
rect 52587 15427 52629 15436
rect 52588 15396 52628 15427
rect 52876 15392 52916 16192
rect 53068 15560 53108 17200
rect 53545 17156 53585 17472
rect 53452 17116 53585 17156
rect 53452 16913 53492 17116
rect 53655 17072 53695 17472
rect 53945 17072 53985 17472
rect 54055 17072 54095 17472
rect 54345 17072 54385 17472
rect 54455 17249 54495 17472
rect 54745 17333 54785 17472
rect 54744 17324 54786 17333
rect 54744 17284 54745 17324
rect 54785 17284 54786 17324
rect 54744 17275 54786 17284
rect 54454 17240 54496 17249
rect 54454 17200 54455 17240
rect 54495 17200 54496 17240
rect 54454 17191 54496 17200
rect 54855 17072 54895 17472
rect 55145 17156 55185 17472
rect 53644 17032 53695 17072
rect 53932 17032 53985 17072
rect 54028 17032 54095 17072
rect 54316 17032 54385 17072
rect 54796 17032 54895 17072
rect 55084 17116 55185 17156
rect 53547 16988 53589 16997
rect 53644 16988 53684 17032
rect 53547 16948 53548 16988
rect 53588 16948 53684 16988
rect 53547 16939 53589 16948
rect 53451 16904 53493 16913
rect 53451 16864 53452 16904
rect 53492 16864 53493 16904
rect 53451 16855 53493 16864
rect 53932 16577 53972 17032
rect 54028 16829 54068 17032
rect 54027 16820 54069 16829
rect 54027 16780 54028 16820
rect 54068 16780 54069 16820
rect 54027 16771 54069 16780
rect 53931 16568 53973 16577
rect 53931 16528 53932 16568
rect 53972 16528 53973 16568
rect 53931 16519 53973 16528
rect 53355 16232 53397 16241
rect 53547 16232 53589 16241
rect 53355 16192 53356 16232
rect 53396 16192 53492 16232
rect 53355 16183 53397 16192
rect 53355 15896 53397 15905
rect 53355 15856 53356 15896
rect 53396 15856 53397 15896
rect 53355 15847 53397 15856
rect 53356 15653 53396 15847
rect 53355 15644 53397 15653
rect 53355 15604 53356 15644
rect 53396 15604 53397 15644
rect 53355 15595 53397 15604
rect 53068 15511 53108 15520
rect 52876 15352 53108 15392
rect 51723 14932 51724 14972
rect 51764 14932 51765 14972
rect 51723 14923 51765 14932
rect 52012 14932 52300 14972
rect 52340 14932 52436 14972
rect 52491 14972 52533 14981
rect 52491 14932 52492 14972
rect 52532 14932 52533 14972
rect 51627 14804 51669 14813
rect 51627 14764 51628 14804
rect 51668 14764 51669 14804
rect 51627 14755 51669 14764
rect 51724 14720 51764 14923
rect 51915 14888 51957 14897
rect 51915 14848 51916 14888
rect 51956 14848 51957 14888
rect 51915 14839 51957 14848
rect 51724 14132 51764 14680
rect 51532 14083 51572 14092
rect 51628 14092 51764 14132
rect 51820 14804 51860 14813
rect 51052 13796 51092 13805
rect 50956 13756 51052 13796
rect 50956 13217 50996 13756
rect 51052 13747 51092 13756
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 51435 13460 51477 13469
rect 51435 13420 51436 13460
rect 51476 13420 51477 13460
rect 51435 13411 51477 13420
rect 51436 13326 51476 13411
rect 51628 13376 51668 14092
rect 51723 13964 51765 13973
rect 51723 13924 51724 13964
rect 51764 13924 51765 13964
rect 51723 13915 51765 13924
rect 51532 13336 51668 13376
rect 50955 13208 50997 13217
rect 51148 13208 51188 13217
rect 50955 13168 50956 13208
rect 50996 13168 51148 13208
rect 50955 13159 50997 13168
rect 51148 13159 51188 13168
rect 51244 13208 51284 13217
rect 50956 13074 50996 13159
rect 51244 13049 51284 13168
rect 51436 13208 51476 13217
rect 51532 13208 51572 13336
rect 51476 13168 51572 13208
rect 51436 13159 51476 13168
rect 51243 13040 51285 13049
rect 51243 13000 51244 13040
rect 51284 13000 51285 13040
rect 51243 12991 51285 13000
rect 50476 12940 50612 12980
rect 50476 11864 50516 12940
rect 50860 12704 50900 12713
rect 50900 12664 51380 12704
rect 50860 12655 50900 12664
rect 51340 12620 51380 12664
rect 51340 12571 51380 12580
rect 50571 12536 50613 12545
rect 50571 12496 50572 12536
rect 50612 12496 50613 12536
rect 50571 12487 50613 12496
rect 50956 12536 50996 12545
rect 50572 11948 50612 12487
rect 50668 12284 50708 12293
rect 50708 12244 50900 12284
rect 50668 12235 50708 12244
rect 50668 11948 50708 11957
rect 50572 11908 50668 11948
rect 50668 11899 50708 11908
rect 50476 11824 50612 11864
rect 50188 11068 50324 11108
rect 50379 11108 50421 11117
rect 50379 11068 50380 11108
rect 50420 11068 50421 11108
rect 49900 10816 50132 10856
rect 49132 9976 49364 10016
rect 49420 10772 49460 10781
rect 49035 9512 49077 9521
rect 49035 9472 49036 9512
rect 49076 9472 49077 9512
rect 49035 9463 49077 9472
rect 48747 8756 48789 8765
rect 48747 8716 48748 8756
rect 48788 8716 48789 8756
rect 48747 8707 48789 8716
rect 48652 8672 48692 8681
rect 48652 8513 48692 8632
rect 48748 8672 48788 8707
rect 48748 8622 48788 8632
rect 48939 8672 48981 8681
rect 49036 8672 49076 9463
rect 49132 9092 49172 9976
rect 49420 9773 49460 10732
rect 49995 10100 50037 10109
rect 49995 10060 49996 10100
rect 50036 10060 50037 10100
rect 49995 10051 50037 10060
rect 49419 9764 49461 9773
rect 49419 9724 49420 9764
rect 49460 9724 49461 9764
rect 49419 9715 49461 9724
rect 49708 9680 49748 9691
rect 49708 9605 49748 9640
rect 49707 9596 49749 9605
rect 49420 9556 49652 9596
rect 49324 9512 49364 9521
rect 49420 9512 49460 9556
rect 49364 9472 49460 9512
rect 49324 9463 49364 9472
rect 49515 9428 49557 9437
rect 49515 9388 49516 9428
rect 49556 9388 49557 9428
rect 49515 9379 49557 9388
rect 49516 9294 49556 9379
rect 49228 9260 49268 9269
rect 49268 9220 49460 9260
rect 49228 9211 49268 9220
rect 49132 9052 49268 9092
rect 49131 8924 49173 8933
rect 49131 8884 49132 8924
rect 49172 8884 49173 8924
rect 49131 8875 49173 8884
rect 48939 8632 48940 8672
rect 48980 8632 49076 8672
rect 49132 8672 49172 8875
rect 48939 8623 48981 8632
rect 49132 8623 49172 8632
rect 49228 8672 49268 9052
rect 49323 8756 49365 8765
rect 49323 8716 49324 8756
rect 49364 8716 49365 8756
rect 49323 8707 49365 8716
rect 49228 8623 49268 8632
rect 49324 8672 49364 8707
rect 48843 8588 48885 8597
rect 48843 8548 48844 8588
rect 48884 8548 48885 8588
rect 48843 8539 48885 8548
rect 48651 8504 48693 8513
rect 48651 8464 48652 8504
rect 48692 8464 48693 8504
rect 48651 8455 48693 8464
rect 48844 8500 48884 8539
rect 48844 8451 48884 8460
rect 48940 8252 48980 8623
rect 49324 8621 49364 8632
rect 49420 8597 49460 9220
rect 49419 8588 49461 8597
rect 49419 8548 49420 8588
rect 49460 8548 49461 8588
rect 49419 8539 49461 8548
rect 49035 8504 49077 8513
rect 49035 8464 49036 8504
rect 49076 8464 49077 8504
rect 49035 8455 49077 8464
rect 49036 8370 49076 8455
rect 48940 8212 49172 8252
rect 48459 8000 48501 8009
rect 48459 7960 48460 8000
rect 48500 7960 48501 8000
rect 48459 7951 48501 7960
rect 49132 8000 49172 8212
rect 49612 8177 49652 9556
rect 49707 9556 49708 9596
rect 49748 9556 49749 9596
rect 49707 9547 49749 9556
rect 49900 9512 49940 9521
rect 49900 8849 49940 9472
rect 49899 8840 49941 8849
rect 49899 8800 49900 8840
rect 49940 8800 49941 8840
rect 49899 8791 49941 8800
rect 49707 8756 49749 8765
rect 49707 8716 49708 8756
rect 49748 8716 49749 8756
rect 49707 8707 49749 8716
rect 49708 8622 49748 8707
rect 49900 8504 49940 8513
rect 49996 8504 50036 10051
rect 50092 8756 50132 10816
rect 50188 8924 50228 11068
rect 50379 11059 50421 11068
rect 50283 10940 50325 10949
rect 50283 10900 50284 10940
rect 50324 10900 50325 10940
rect 50283 10891 50325 10900
rect 50284 10806 50324 10891
rect 50380 10436 50420 11059
rect 50380 10387 50420 10396
rect 50476 10772 50516 10781
rect 50476 10193 50516 10732
rect 50572 10268 50612 11824
rect 50860 11524 50900 12244
rect 50956 11948 50996 12496
rect 51051 12536 51093 12545
rect 51051 12496 51052 12536
rect 51092 12496 51093 12536
rect 51051 12487 51093 12496
rect 51148 12536 51188 12547
rect 51052 12402 51092 12487
rect 51148 12461 51188 12496
rect 51147 12452 51189 12461
rect 51147 12412 51148 12452
rect 51188 12412 51189 12452
rect 51147 12403 51189 12412
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 51340 11948 51380 11957
rect 51532 11948 51572 13168
rect 51627 13208 51669 13217
rect 51627 13168 51628 13208
rect 51668 13168 51669 13208
rect 51627 13159 51669 13168
rect 51724 13208 51764 13915
rect 51820 13469 51860 14764
rect 51916 14754 51956 14839
rect 52012 14804 52052 14932
rect 52300 14923 52340 14932
rect 52491 14923 52533 14932
rect 53068 14888 53108 15352
rect 53452 15233 53492 16192
rect 53547 16192 53548 16232
rect 53588 16192 53589 16232
rect 53547 16183 53589 16192
rect 53740 16232 53780 16241
rect 53451 15224 53493 15233
rect 53451 15184 53452 15224
rect 53492 15184 53493 15224
rect 53451 15175 53493 15184
rect 53451 14972 53493 14981
rect 53451 14932 53452 14972
rect 53492 14932 53493 14972
rect 53451 14923 53493 14932
rect 52012 14755 52052 14764
rect 52588 14848 53012 14888
rect 53068 14848 53396 14888
rect 52108 14720 52148 14729
rect 52011 14636 52053 14645
rect 52011 14596 52012 14636
rect 52052 14596 52053 14636
rect 52011 14587 52053 14596
rect 51916 14048 51956 14057
rect 51916 13889 51956 14008
rect 51915 13880 51957 13889
rect 51915 13840 51916 13880
rect 51956 13840 51957 13880
rect 51915 13831 51957 13840
rect 51819 13460 51861 13469
rect 51819 13420 51820 13460
rect 51860 13420 51861 13460
rect 51819 13411 51861 13420
rect 52012 13460 52052 14587
rect 52108 14561 52148 14680
rect 52588 14720 52628 14848
rect 52588 14671 52628 14680
rect 52684 14720 52724 14729
rect 52972 14720 53012 14848
rect 52724 14680 52916 14720
rect 52684 14671 52724 14680
rect 52107 14552 52149 14561
rect 52107 14512 52108 14552
rect 52148 14512 52149 14552
rect 52107 14503 52149 14512
rect 52779 14552 52821 14561
rect 52779 14508 52780 14552
rect 52820 14508 52821 14552
rect 52779 14503 52821 14508
rect 52780 14417 52820 14503
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 52876 14309 52916 14680
rect 52972 14671 53012 14680
rect 53068 14720 53108 14729
rect 53068 14477 53108 14680
rect 53163 14720 53205 14729
rect 53163 14680 53164 14720
rect 53204 14680 53205 14720
rect 53163 14671 53205 14680
rect 53260 14699 53300 14731
rect 53164 14586 53204 14671
rect 53260 14645 53300 14659
rect 53259 14636 53301 14645
rect 53259 14596 53260 14636
rect 53300 14596 53301 14636
rect 53259 14587 53301 14596
rect 53067 14468 53109 14477
rect 53067 14428 53068 14468
rect 53108 14428 53109 14468
rect 53067 14419 53109 14428
rect 52107 14300 52149 14309
rect 52107 14260 52108 14300
rect 52148 14260 52149 14300
rect 52107 14251 52149 14260
rect 52875 14300 52917 14309
rect 52875 14260 52876 14300
rect 52916 14260 52917 14300
rect 52875 14251 52917 14260
rect 53259 14300 53301 14309
rect 53259 14260 53260 14300
rect 53300 14260 53301 14300
rect 53259 14251 53301 14260
rect 52012 13411 52052 13420
rect 52108 13292 52148 14251
rect 53260 14141 53300 14251
rect 53259 14132 53301 14141
rect 53259 14092 53260 14132
rect 53300 14092 53301 14132
rect 53259 14083 53301 14092
rect 52779 14048 52821 14057
rect 52779 14008 52780 14048
rect 52820 14008 52821 14048
rect 52779 13999 52821 14008
rect 52203 13880 52245 13889
rect 52203 13840 52204 13880
rect 52244 13840 52245 13880
rect 52203 13831 52245 13840
rect 51628 12461 51668 13159
rect 51724 13133 51764 13168
rect 51820 13252 52148 13292
rect 51723 13124 51765 13133
rect 51723 13084 51724 13124
rect 51764 13084 51765 13124
rect 51723 13075 51765 13084
rect 51723 12956 51765 12965
rect 51723 12916 51724 12956
rect 51764 12916 51765 12956
rect 51723 12907 51765 12916
rect 51724 12536 51764 12907
rect 51724 12487 51764 12496
rect 51627 12452 51669 12461
rect 51627 12412 51628 12452
rect 51668 12412 51669 12452
rect 51627 12403 51669 12412
rect 50956 11908 51340 11948
rect 51340 11899 51380 11908
rect 51436 11908 51572 11948
rect 50955 11696 50997 11705
rect 50955 11656 50956 11696
rect 50996 11656 50997 11696
rect 50955 11647 50997 11656
rect 51052 11696 51092 11705
rect 50956 11562 50996 11647
rect 51052 11537 51092 11656
rect 51436 11612 51476 11908
rect 51628 11696 51668 12403
rect 51723 11948 51765 11957
rect 51723 11908 51724 11948
rect 51764 11908 51765 11948
rect 51723 11899 51765 11908
rect 51628 11647 51668 11656
rect 51724 11696 51764 11899
rect 51820 11705 51860 13252
rect 51915 13124 51957 13133
rect 51915 13084 51916 13124
rect 51956 13084 51957 13124
rect 51915 13075 51957 13084
rect 51724 11647 51764 11656
rect 51819 11696 51861 11705
rect 51819 11656 51820 11696
rect 51860 11656 51861 11696
rect 51819 11647 51861 11656
rect 51244 11570 51284 11579
rect 50860 11360 50900 11484
rect 51051 11528 51093 11537
rect 51051 11488 51052 11528
rect 51092 11488 51093 11528
rect 51051 11479 51093 11488
rect 50668 11320 50900 11360
rect 50668 11024 50708 11320
rect 51244 11276 51284 11530
rect 50668 10975 50708 10984
rect 50764 11236 51284 11276
rect 51340 11572 51476 11612
rect 51531 11612 51573 11621
rect 51531 11572 51532 11612
rect 51572 11572 51573 11612
rect 50764 10940 50804 11236
rect 51052 11024 51092 11033
rect 51340 11024 51380 11572
rect 51531 11563 51573 11572
rect 51532 11478 51572 11563
rect 51820 11562 51860 11647
rect 51627 11192 51669 11201
rect 51916 11192 51956 13075
rect 52204 12965 52244 13831
rect 52684 13208 52724 13217
rect 52780 13208 52820 13999
rect 53356 13889 53396 14848
rect 53452 14838 53492 14923
rect 53452 14729 53492 14748
rect 53451 14720 53493 14729
rect 53548 14720 53588 16183
rect 53451 14680 53452 14720
rect 53492 14680 53548 14720
rect 53451 14671 53493 14680
rect 53548 14671 53588 14680
rect 53643 14720 53685 14729
rect 53643 14680 53644 14720
rect 53684 14680 53685 14720
rect 53643 14671 53685 14680
rect 53547 14468 53589 14477
rect 53547 14428 53548 14468
rect 53588 14428 53589 14468
rect 53547 14419 53589 14428
rect 53355 13880 53397 13889
rect 53355 13840 53356 13880
rect 53396 13840 53397 13880
rect 53355 13831 53397 13840
rect 52724 13168 52820 13208
rect 52684 13159 52724 13168
rect 53548 12980 53588 14419
rect 53644 13133 53684 14671
rect 53740 14057 53780 16192
rect 53835 14804 53877 14813
rect 53835 14764 53836 14804
rect 53876 14764 53877 14804
rect 53835 14755 53877 14764
rect 53739 14048 53781 14057
rect 53739 14008 53740 14048
rect 53780 14008 53781 14048
rect 53739 13999 53781 14008
rect 53836 13217 53876 14755
rect 54028 14729 54068 14814
rect 53932 14720 53972 14729
rect 53932 14393 53972 14680
rect 54027 14720 54069 14729
rect 54027 14680 54028 14720
rect 54068 14680 54069 14720
rect 54027 14671 54069 14680
rect 54219 14720 54261 14729
rect 54219 14680 54220 14720
rect 54260 14680 54261 14720
rect 54219 14671 54261 14680
rect 54220 14586 54260 14671
rect 54124 14552 54164 14561
rect 54028 14512 54124 14552
rect 53931 14384 53973 14393
rect 53931 14344 53932 14384
rect 53972 14344 53973 14384
rect 53931 14335 53973 14344
rect 53932 14216 53972 14335
rect 53932 14167 53972 14176
rect 54028 13628 54068 14512
rect 54124 14503 54164 14512
rect 54316 14309 54356 17032
rect 54796 15821 54836 17032
rect 54891 16904 54933 16913
rect 54891 16864 54892 16904
rect 54932 16864 54933 16904
rect 54891 16855 54933 16864
rect 54892 16484 54932 16855
rect 55084 16745 55124 17116
rect 55255 17072 55295 17472
rect 55180 17032 55295 17072
rect 55545 17072 55585 17472
rect 55655 17072 55695 17472
rect 55945 17072 55985 17472
rect 56055 17072 56095 17472
rect 55545 17032 55604 17072
rect 55655 17032 55700 17072
rect 55945 17032 55988 17072
rect 55083 16736 55125 16745
rect 55083 16696 55084 16736
rect 55124 16696 55125 16736
rect 55083 16687 55125 16696
rect 55180 16661 55220 17032
rect 55179 16652 55221 16661
rect 55179 16612 55180 16652
rect 55220 16612 55221 16652
rect 55179 16603 55221 16612
rect 54892 16241 54932 16444
rect 55276 16241 55316 16326
rect 54891 16232 54933 16241
rect 55180 16232 55220 16241
rect 54891 16192 54892 16232
rect 54932 16192 54933 16232
rect 54891 16183 54933 16192
rect 54988 16192 55180 16232
rect 54795 15812 54837 15821
rect 54795 15772 54796 15812
rect 54836 15772 54837 15812
rect 54795 15763 54837 15772
rect 54603 15308 54645 15317
rect 54603 15268 54604 15308
rect 54644 15268 54645 15308
rect 54603 15259 54645 15268
rect 54604 15174 54644 15259
rect 54699 15224 54741 15233
rect 54699 15184 54700 15224
rect 54740 15184 54741 15224
rect 54699 15175 54741 15184
rect 54603 14888 54645 14897
rect 54603 14848 54604 14888
rect 54644 14848 54645 14888
rect 54603 14839 54645 14848
rect 54412 14720 54452 14729
rect 54412 14393 54452 14680
rect 54507 14552 54549 14561
rect 54507 14512 54508 14552
rect 54548 14512 54549 14552
rect 54507 14503 54549 14512
rect 54508 14418 54548 14503
rect 54411 14384 54453 14393
rect 54411 14344 54412 14384
rect 54452 14344 54453 14384
rect 54411 14335 54453 14344
rect 54315 14300 54357 14309
rect 54315 14260 54316 14300
rect 54356 14260 54357 14300
rect 54315 14251 54357 14260
rect 54124 14048 54164 14057
rect 54124 13712 54164 14008
rect 54508 14048 54548 14057
rect 54508 13889 54548 14008
rect 54507 13880 54549 13889
rect 54507 13840 54508 13880
rect 54548 13840 54549 13880
rect 54507 13831 54549 13840
rect 54124 13672 54548 13712
rect 54028 13588 54452 13628
rect 54412 13292 54452 13588
rect 54508 13376 54548 13672
rect 54508 13327 54548 13336
rect 54412 13243 54452 13252
rect 54604 13292 54644 14839
rect 54700 14477 54740 15175
rect 54988 14888 55028 16192
rect 55180 16183 55220 16192
rect 55275 16232 55317 16241
rect 55275 16192 55276 16232
rect 55316 16192 55317 16232
rect 55275 16183 55317 16192
rect 55372 16232 55412 16241
rect 55412 16192 55508 16232
rect 55372 16183 55412 16192
rect 55084 16064 55124 16073
rect 55124 16024 55412 16064
rect 55084 16015 55124 16024
rect 55372 15644 55412 16024
rect 55372 15595 55412 15604
rect 55468 15485 55508 16192
rect 55564 15989 55604 17032
rect 55660 16325 55700 17032
rect 55659 16316 55701 16325
rect 55659 16276 55660 16316
rect 55700 16276 55701 16316
rect 55659 16267 55701 16276
rect 55948 16157 55988 17032
rect 56044 17032 56095 17072
rect 56345 17072 56385 17472
rect 56455 17249 56495 17472
rect 56745 17333 56785 17472
rect 56744 17324 56786 17333
rect 56744 17284 56745 17324
rect 56785 17284 56786 17324
rect 56744 17275 56786 17284
rect 56855 17249 56895 17472
rect 57145 17333 57185 17472
rect 57255 17333 57295 17472
rect 57144 17324 57186 17333
rect 57144 17284 57145 17324
rect 57185 17284 57186 17324
rect 57144 17275 57186 17284
rect 57254 17324 57296 17333
rect 57254 17284 57255 17324
rect 57295 17284 57296 17324
rect 57254 17275 57296 17284
rect 57545 17249 57585 17472
rect 57655 17249 57695 17472
rect 56454 17240 56496 17249
rect 56454 17200 56455 17240
rect 56495 17200 56496 17240
rect 56454 17191 56496 17200
rect 56854 17240 56896 17249
rect 56854 17200 56855 17240
rect 56895 17200 56896 17240
rect 56854 17191 56896 17200
rect 57544 17240 57586 17249
rect 57544 17200 57545 17240
rect 57585 17200 57586 17240
rect 57544 17191 57586 17200
rect 57654 17240 57696 17249
rect 57654 17200 57655 17240
rect 57695 17200 57696 17240
rect 57654 17191 57696 17200
rect 57945 17165 57985 17472
rect 58055 17249 58095 17472
rect 58054 17240 58096 17249
rect 58054 17200 58055 17240
rect 58095 17200 58096 17240
rect 58054 17191 58096 17200
rect 57944 17156 57986 17165
rect 57944 17116 57945 17156
rect 57985 17116 57986 17156
rect 57944 17107 57986 17116
rect 58345 17072 58385 17472
rect 58455 17249 58495 17472
rect 58745 17333 58785 17472
rect 58855 17333 58895 17472
rect 58744 17324 58786 17333
rect 58744 17284 58745 17324
rect 58785 17284 58786 17324
rect 58744 17275 58786 17284
rect 58854 17324 58896 17333
rect 58854 17284 58855 17324
rect 58895 17284 58896 17324
rect 58854 17275 58896 17284
rect 58454 17240 58496 17249
rect 58454 17200 58455 17240
rect 58495 17200 58496 17240
rect 58454 17191 58496 17200
rect 59145 17072 59185 17472
rect 59255 17333 59295 17472
rect 59545 17333 59585 17472
rect 59655 17333 59695 17472
rect 59254 17324 59296 17333
rect 59254 17284 59255 17324
rect 59295 17284 59296 17324
rect 59254 17275 59296 17284
rect 59544 17324 59586 17333
rect 59544 17284 59545 17324
rect 59585 17284 59586 17324
rect 59544 17275 59586 17284
rect 59654 17324 59696 17333
rect 59654 17284 59655 17324
rect 59695 17284 59696 17324
rect 59654 17275 59696 17284
rect 59691 17156 59733 17165
rect 59691 17116 59692 17156
rect 59732 17116 59733 17156
rect 59691 17107 59733 17116
rect 56345 17032 56468 17072
rect 58345 17032 58388 17072
rect 56044 16493 56084 17032
rect 56043 16484 56085 16493
rect 56043 16444 56044 16484
rect 56084 16444 56085 16484
rect 56043 16435 56085 16444
rect 56331 16484 56373 16493
rect 56331 16444 56332 16484
rect 56372 16444 56373 16484
rect 56331 16435 56373 16444
rect 56332 16350 56372 16435
rect 56044 16316 56084 16325
rect 56084 16276 56180 16316
rect 56044 16267 56084 16276
rect 55947 16148 55989 16157
rect 55947 16108 55948 16148
rect 55988 16108 55989 16148
rect 55947 16099 55989 16108
rect 55852 16064 55892 16073
rect 55756 16024 55852 16064
rect 55563 15980 55605 15989
rect 55563 15940 55564 15980
rect 55604 15940 55605 15980
rect 55563 15931 55605 15940
rect 55756 15569 55796 16024
rect 55852 16015 55892 16024
rect 55947 15980 55989 15989
rect 55947 15940 55948 15980
rect 55988 15940 55989 15980
rect 55947 15931 55989 15940
rect 55755 15560 55797 15569
rect 55755 15520 55756 15560
rect 55796 15520 55797 15560
rect 55755 15511 55797 15520
rect 55467 15476 55509 15485
rect 55467 15436 55468 15476
rect 55508 15436 55509 15476
rect 55467 15427 55509 15436
rect 55756 15426 55796 15511
rect 55851 15476 55893 15485
rect 55851 15436 55852 15476
rect 55892 15436 55893 15476
rect 55851 15427 55893 15436
rect 55083 14888 55125 14897
rect 54988 14848 55084 14888
rect 55124 14848 55125 14888
rect 55083 14839 55125 14848
rect 55372 14848 55796 14888
rect 55084 14754 55124 14839
rect 55372 14720 55412 14848
rect 55372 14671 55412 14680
rect 55467 14720 55509 14729
rect 55467 14680 55468 14720
rect 55508 14680 55509 14720
rect 55467 14671 55509 14680
rect 55756 14720 55796 14848
rect 55756 14671 55796 14680
rect 55852 14720 55892 15427
rect 55468 14586 55508 14671
rect 55564 14494 55604 14503
rect 54699 14468 54741 14477
rect 54699 14428 54700 14468
rect 54740 14428 54741 14468
rect 54699 14419 54741 14428
rect 54795 14300 54837 14309
rect 54795 14260 54796 14300
rect 54836 14260 54837 14300
rect 54795 14251 54837 14260
rect 54699 13460 54741 13469
rect 54699 13420 54700 13460
rect 54740 13420 54741 13460
rect 54699 13411 54741 13420
rect 54604 13243 54644 13252
rect 53835 13208 53877 13217
rect 53835 13168 53836 13208
rect 53876 13168 53877 13208
rect 53835 13159 53877 13168
rect 54315 13208 54357 13217
rect 54315 13168 54316 13208
rect 54356 13168 54357 13208
rect 54315 13159 54357 13168
rect 54700 13208 54740 13411
rect 54700 13159 54740 13168
rect 53643 13124 53685 13133
rect 53643 13084 53644 13124
rect 53684 13084 53685 13124
rect 53643 13075 53685 13084
rect 54316 13074 54356 13159
rect 52203 12956 52245 12965
rect 52203 12916 52204 12956
rect 52244 12916 52245 12956
rect 53548 12940 53780 12980
rect 52203 12907 52245 12916
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 52779 12788 52821 12797
rect 52779 12748 52780 12788
rect 52820 12748 52821 12788
rect 52779 12739 52821 12748
rect 52587 12704 52629 12713
rect 52587 12664 52588 12704
rect 52628 12664 52629 12704
rect 52587 12655 52629 12664
rect 52588 12536 52628 12655
rect 52588 12487 52628 12496
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 52780 11201 52820 12739
rect 53740 12704 53780 12940
rect 53740 12655 53780 12664
rect 53740 12284 53780 12293
rect 53740 11957 53780 12244
rect 53739 11948 53781 11957
rect 53739 11908 53740 11948
rect 53780 11908 53781 11948
rect 53739 11899 53781 11908
rect 54796 11873 54836 14251
rect 55371 14048 55413 14057
rect 55371 14008 55372 14048
rect 55412 14008 55413 14048
rect 55371 13999 55413 14008
rect 55372 13914 55412 13999
rect 55564 13469 55604 14454
rect 55755 13796 55797 13805
rect 55755 13756 55756 13796
rect 55796 13756 55797 13796
rect 55755 13747 55797 13756
rect 55179 13460 55221 13469
rect 55179 13420 55180 13460
rect 55220 13420 55221 13460
rect 55179 13411 55221 13420
rect 55563 13460 55605 13469
rect 55563 13420 55564 13460
rect 55604 13420 55605 13460
rect 55563 13411 55605 13420
rect 55180 13326 55220 13411
rect 55275 13208 55317 13217
rect 55275 13168 55276 13208
rect 55316 13168 55317 13208
rect 55275 13159 55317 13168
rect 55468 13208 55508 13219
rect 55756 13217 55796 13747
rect 55276 13074 55316 13159
rect 55468 13133 55508 13168
rect 55660 13208 55700 13217
rect 55467 13124 55509 13133
rect 55467 13084 55468 13124
rect 55508 13084 55509 13124
rect 55467 13075 55509 13084
rect 55083 13040 55125 13049
rect 55083 13000 55084 13040
rect 55124 13000 55125 13040
rect 55083 12991 55125 13000
rect 55564 13040 55604 13049
rect 54795 11864 54837 11873
rect 54795 11824 54796 11864
rect 54836 11824 54837 11864
rect 54795 11815 54837 11824
rect 53355 11780 53397 11789
rect 53355 11740 53356 11780
rect 53396 11740 53397 11780
rect 53355 11731 53397 11740
rect 53356 11646 53396 11731
rect 54508 11696 54548 11705
rect 54548 11656 54740 11696
rect 54508 11647 54548 11656
rect 54123 11276 54165 11285
rect 54123 11236 54124 11276
rect 54164 11236 54165 11276
rect 54123 11227 54165 11236
rect 51627 11152 51628 11192
rect 51668 11152 51669 11192
rect 51627 11143 51669 11152
rect 51820 11152 51956 11192
rect 52779 11192 52821 11201
rect 52779 11152 52780 11192
rect 52820 11152 52821 11192
rect 51092 10984 51380 11024
rect 51436 11024 51476 11033
rect 51052 10975 51092 10984
rect 50764 10891 50804 10900
rect 50956 10940 50996 10949
rect 51436 10940 51476 10984
rect 50859 10856 50901 10865
rect 50859 10816 50860 10856
rect 50900 10816 50901 10856
rect 50859 10807 50901 10816
rect 50860 10722 50900 10807
rect 50956 10436 50996 10900
rect 51340 10900 51476 10940
rect 51532 11024 51572 11033
rect 51340 10781 51380 10900
rect 51339 10772 51381 10781
rect 51339 10732 51340 10772
rect 51380 10732 51381 10772
rect 51339 10723 51381 10732
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 51148 10436 51188 10445
rect 50956 10396 51148 10436
rect 51148 10387 51188 10396
rect 51243 10436 51285 10445
rect 51243 10396 51244 10436
rect 51284 10396 51285 10436
rect 51243 10387 51285 10396
rect 50764 10268 50804 10277
rect 50572 10228 50764 10268
rect 50475 10184 50517 10193
rect 50475 10144 50476 10184
rect 50516 10144 50517 10184
rect 50475 10135 50517 10144
rect 50283 9596 50325 9605
rect 50283 9556 50284 9596
rect 50324 9556 50325 9596
rect 50283 9547 50325 9556
rect 50284 9512 50324 9547
rect 50284 9461 50324 9472
rect 50284 8924 50324 8933
rect 50188 8884 50284 8924
rect 50188 8765 50228 8884
rect 50284 8875 50324 8884
rect 50092 8707 50132 8716
rect 50187 8756 50229 8765
rect 50187 8716 50188 8756
rect 50228 8716 50229 8756
rect 50187 8707 50229 8716
rect 50476 8672 50516 10135
rect 50764 9101 50804 10228
rect 50955 10268 50997 10277
rect 50955 10228 50956 10268
rect 50996 10228 50997 10268
rect 50955 10219 50997 10228
rect 50956 10016 50996 10219
rect 51147 10184 51189 10193
rect 51244 10184 51284 10387
rect 51532 10268 51572 10984
rect 51628 11024 51668 11143
rect 51628 10975 51668 10984
rect 51724 11024 51764 11035
rect 51724 10949 51764 10984
rect 51723 10940 51765 10949
rect 51723 10900 51724 10940
rect 51764 10900 51765 10940
rect 51723 10891 51765 10900
rect 51723 10772 51765 10781
rect 51723 10732 51724 10772
rect 51764 10732 51765 10772
rect 51723 10723 51765 10732
rect 51532 10228 51668 10268
rect 51147 10144 51148 10184
rect 51188 10144 51284 10184
rect 51340 10184 51380 10195
rect 51147 10135 51189 10144
rect 51148 10050 51188 10135
rect 51340 10109 51380 10144
rect 51435 10184 51477 10193
rect 51435 10144 51436 10184
rect 51476 10144 51477 10184
rect 51435 10135 51477 10144
rect 51339 10100 51381 10109
rect 51339 10060 51340 10100
rect 51380 10060 51381 10100
rect 51339 10051 51381 10060
rect 51436 10050 51476 10135
rect 51531 10100 51573 10109
rect 51531 10060 51532 10100
rect 51572 10060 51573 10100
rect 51531 10051 51573 10060
rect 50956 9967 50996 9976
rect 51147 9512 51189 9521
rect 51147 9472 51148 9512
rect 51188 9472 51189 9512
rect 51147 9463 51189 9472
rect 51148 9378 51188 9463
rect 50763 9092 50805 9101
rect 50763 9052 50764 9092
rect 50804 9052 50805 9092
rect 50763 9043 50805 9052
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 50763 8924 50805 8933
rect 50763 8884 50764 8924
rect 50804 8884 50805 8924
rect 50763 8875 50805 8884
rect 51243 8924 51285 8933
rect 51243 8884 51244 8924
rect 51284 8884 51285 8924
rect 51243 8875 51285 8884
rect 50667 8840 50709 8849
rect 50667 8800 50668 8840
rect 50708 8800 50709 8840
rect 50667 8791 50709 8800
rect 49940 8464 50228 8504
rect 49900 8455 49940 8464
rect 49611 8168 49653 8177
rect 49611 8128 49612 8168
rect 49652 8128 49653 8168
rect 49611 8119 49653 8128
rect 50091 8168 50133 8177
rect 50091 8128 50092 8168
rect 50132 8128 50133 8168
rect 50091 8119 50133 8128
rect 49132 7951 49172 7960
rect 48308 7120 48404 7160
rect 50092 7160 50132 8119
rect 48268 7111 48308 7120
rect 50092 7111 50132 7120
rect 50188 7160 50228 8464
rect 50283 8168 50325 8177
rect 50283 8128 50284 8168
rect 50324 8128 50325 8168
rect 50283 8119 50325 8128
rect 50284 8034 50324 8119
rect 50379 7412 50421 7421
rect 50379 7372 50380 7412
rect 50420 7372 50421 7412
rect 50379 7363 50421 7372
rect 50380 7278 50420 7363
rect 47884 7026 47924 7111
rect 50188 6749 50228 7120
rect 50380 7160 50420 7169
rect 50476 7160 50516 8632
rect 50572 8756 50612 8765
rect 50572 7421 50612 8716
rect 50668 8706 50708 8791
rect 50764 8756 50804 8875
rect 51244 8790 51284 8875
rect 50764 8707 50804 8716
rect 50859 8672 50901 8681
rect 50859 8632 50860 8672
rect 50900 8632 50901 8672
rect 50859 8623 50901 8632
rect 51532 8672 51572 10051
rect 51628 8933 51668 10228
rect 51724 10184 51764 10723
rect 51724 10135 51764 10144
rect 51627 8924 51669 8933
rect 51627 8884 51628 8924
rect 51668 8884 51669 8924
rect 51627 8875 51669 8884
rect 51627 8756 51669 8765
rect 51627 8716 51628 8756
rect 51668 8716 51669 8756
rect 51627 8707 51669 8716
rect 51532 8623 51572 8632
rect 51628 8672 51668 8707
rect 51820 8672 51860 11152
rect 52779 11143 52821 11152
rect 52204 11068 52628 11108
rect 51916 11024 51956 11033
rect 51916 10109 51956 10984
rect 52012 11024 52052 11033
rect 52012 10949 52052 10984
rect 52107 11024 52149 11033
rect 52107 10984 52108 11024
rect 52148 10984 52149 11024
rect 52107 10975 52149 10984
rect 52204 11024 52244 11068
rect 52204 10975 52244 10984
rect 52011 10940 52053 10949
rect 52011 10900 52012 10940
rect 52052 10900 52053 10940
rect 52011 10891 52053 10900
rect 52012 10697 52052 10891
rect 52108 10890 52148 10975
rect 52395 10940 52437 10949
rect 52395 10900 52396 10940
rect 52436 10900 52437 10940
rect 52395 10891 52437 10900
rect 52396 10806 52436 10891
rect 52588 10772 52628 11068
rect 52780 11058 52820 11143
rect 52875 11024 52917 11033
rect 52875 10984 52876 11024
rect 52916 10984 52917 11024
rect 52875 10975 52917 10984
rect 52628 10732 52820 10772
rect 52588 10723 52628 10732
rect 52011 10688 52053 10697
rect 52011 10648 52012 10688
rect 52052 10648 52053 10688
rect 52011 10639 52053 10648
rect 52012 10277 52052 10639
rect 52011 10268 52053 10277
rect 52011 10228 52012 10268
rect 52052 10228 52053 10268
rect 52011 10219 52053 10228
rect 52108 10184 52148 10193
rect 51915 10100 51957 10109
rect 51915 10060 51916 10100
rect 51956 10060 51957 10100
rect 51915 10051 51957 10060
rect 52108 9689 52148 10144
rect 52203 10184 52245 10193
rect 52203 10144 52204 10184
rect 52244 10144 52245 10184
rect 52203 10135 52245 10144
rect 52107 9680 52149 9689
rect 52107 9640 52108 9680
rect 52148 9640 52149 9680
rect 52204 9680 52244 10135
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 52300 9680 52340 9689
rect 52204 9640 52300 9680
rect 52340 9640 52532 9680
rect 52107 9631 52149 9640
rect 52300 9631 52340 9640
rect 52011 9512 52053 9521
rect 52011 9472 52012 9512
rect 52052 9472 52053 9512
rect 52011 9463 52053 9472
rect 52492 9512 52532 9640
rect 52492 9463 52532 9472
rect 52012 8840 52052 9463
rect 52588 9260 52628 9269
rect 52107 8840 52149 8849
rect 52012 8800 52108 8840
rect 52148 8800 52149 8840
rect 52107 8791 52149 8800
rect 52299 8840 52341 8849
rect 52299 8800 52300 8840
rect 52340 8800 52341 8840
rect 52299 8791 52341 8800
rect 52012 8672 52052 8681
rect 51820 8632 52012 8672
rect 50860 8538 50900 8623
rect 51628 8621 51668 8632
rect 52012 8623 52052 8632
rect 51724 8446 51764 8515
rect 51723 8380 51724 8429
rect 51764 8380 51765 8429
rect 52108 8420 52148 8791
rect 52300 8706 52340 8791
rect 52588 8681 52628 9220
rect 52780 8756 52820 10732
rect 52876 10529 52916 10975
rect 54124 10529 54164 11227
rect 52875 10520 52917 10529
rect 52875 10480 52876 10520
rect 52916 10480 52917 10520
rect 52875 10471 52917 10480
rect 54123 10520 54165 10529
rect 54123 10480 54124 10520
rect 54164 10480 54165 10520
rect 54123 10471 54165 10480
rect 54124 10436 54164 10471
rect 54124 10386 54164 10396
rect 53451 10352 53493 10361
rect 53451 10312 53452 10352
rect 53492 10312 53493 10352
rect 53451 10303 53493 10312
rect 52972 10184 53012 10193
rect 52972 10109 53012 10144
rect 52971 10100 53013 10109
rect 52971 10060 52972 10100
rect 53012 10060 53013 10100
rect 52971 10051 53013 10060
rect 52875 8756 52917 8765
rect 52780 8716 52876 8756
rect 52916 8716 52917 8756
rect 52875 8707 52917 8716
rect 52587 8672 52629 8681
rect 52587 8632 52588 8672
rect 52628 8632 52629 8672
rect 52587 8623 52629 8632
rect 51723 8371 51765 8380
rect 51916 8380 52148 8420
rect 50667 8000 50709 8009
rect 51052 8000 51092 8009
rect 50667 7960 50668 8000
rect 50708 7960 50709 8000
rect 50667 7951 50709 7960
rect 50956 7960 51052 8000
rect 50668 7866 50708 7951
rect 50571 7412 50613 7421
rect 50571 7372 50572 7412
rect 50612 7372 50613 7412
rect 50571 7363 50613 7372
rect 50420 7120 50516 7160
rect 50187 6740 50229 6749
rect 50187 6700 50188 6740
rect 50228 6700 50229 6740
rect 50187 6691 50229 6700
rect 50380 6413 50420 7120
rect 50956 7001 50996 7960
rect 51052 7951 51092 7960
rect 51916 8000 51956 8380
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 52587 8168 52629 8177
rect 52587 8128 52588 8168
rect 52628 8128 52629 8168
rect 52587 8119 52629 8128
rect 51916 7951 51956 7960
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 51724 7160 51764 7169
rect 50955 6992 50997 7001
rect 50955 6952 50956 6992
rect 50996 6952 50997 6992
rect 50955 6943 50997 6952
rect 51724 6581 51764 7120
rect 51819 7160 51861 7169
rect 51819 7120 51820 7160
rect 51860 7120 51861 7160
rect 51819 7111 51861 7120
rect 51916 7160 51956 7169
rect 51820 7026 51860 7111
rect 51723 6572 51765 6581
rect 51723 6532 51724 6572
rect 51764 6532 51765 6572
rect 51723 6523 51765 6532
rect 50379 6404 50421 6413
rect 50379 6364 50380 6404
rect 50420 6364 50421 6404
rect 50379 6355 50421 6364
rect 51916 6329 51956 7120
rect 52012 7160 52052 7169
rect 52204 7160 52244 7169
rect 52052 7120 52204 7160
rect 52012 7111 52052 7120
rect 52204 7111 52244 7120
rect 52588 7160 52628 8119
rect 52876 7421 52916 8707
rect 52972 8672 53012 10051
rect 53452 9596 53492 10303
rect 54700 10109 54740 11656
rect 55084 10949 55124 12991
rect 55564 12980 55604 13000
rect 55276 12940 55604 12980
rect 55660 12965 55700 13168
rect 55755 13208 55797 13217
rect 55755 13168 55756 13208
rect 55796 13168 55797 13208
rect 55755 13159 55797 13168
rect 55852 13133 55892 14680
rect 55948 14720 55988 15931
rect 56140 15905 56180 16276
rect 56236 16232 56276 16241
rect 56236 15980 56276 16192
rect 56236 15940 56372 15980
rect 56139 15896 56181 15905
rect 56139 15856 56140 15896
rect 56180 15856 56181 15896
rect 56139 15847 56181 15856
rect 56043 15644 56085 15653
rect 56043 15604 56044 15644
rect 56084 15604 56085 15644
rect 56043 15595 56085 15604
rect 56044 14729 56084 15595
rect 55948 14671 55988 14680
rect 56043 14720 56085 14729
rect 56043 14680 56044 14720
rect 56084 14680 56085 14720
rect 56043 14671 56085 14680
rect 56140 14552 56180 15847
rect 55948 14512 56180 14552
rect 55851 13124 55893 13133
rect 55948 13124 55988 14512
rect 56043 14384 56085 14393
rect 56043 14344 56044 14384
rect 56084 14344 56085 14384
rect 56043 14335 56085 14344
rect 56044 13124 56084 14335
rect 56332 13721 56372 15940
rect 56428 15737 56468 17032
rect 57291 16820 57333 16829
rect 57291 16780 57292 16820
rect 57332 16780 57333 16820
rect 57291 16771 57333 16780
rect 56619 16736 56661 16745
rect 56619 16696 56620 16736
rect 56660 16696 56661 16736
rect 56619 16687 56661 16696
rect 56620 16232 56660 16687
rect 57003 16484 57045 16493
rect 57003 16444 57004 16484
rect 57044 16444 57045 16484
rect 57003 16435 57045 16444
rect 57292 16484 57332 16771
rect 58348 16577 58388 17032
rect 59020 17032 59185 17072
rect 59595 17072 59637 17081
rect 59595 17032 59596 17072
rect 59636 17032 59637 17072
rect 58347 16568 58389 16577
rect 58347 16528 58348 16568
rect 58388 16528 58389 16568
rect 58347 16519 58389 16528
rect 57292 16435 57332 16444
rect 57004 16241 57044 16435
rect 58156 16241 58196 16326
rect 58731 16316 58773 16325
rect 58731 16276 58732 16316
rect 58772 16276 58773 16316
rect 58731 16267 58773 16276
rect 56620 15821 56660 16192
rect 56908 16232 56948 16241
rect 56716 16064 56756 16073
rect 56619 15812 56661 15821
rect 56619 15772 56620 15812
rect 56660 15772 56661 15812
rect 56619 15763 56661 15772
rect 56716 15737 56756 16024
rect 56908 15989 56948 16192
rect 57003 16232 57045 16241
rect 57003 16192 57004 16232
rect 57044 16192 57045 16232
rect 57003 16183 57045 16192
rect 57196 16232 57236 16241
rect 56907 15980 56949 15989
rect 56907 15940 56908 15980
rect 56948 15940 56949 15980
rect 56907 15931 56949 15940
rect 56427 15728 56469 15737
rect 56427 15688 56428 15728
rect 56468 15688 56469 15728
rect 56427 15679 56469 15688
rect 56715 15728 56757 15737
rect 56715 15688 56716 15728
rect 56756 15688 56757 15728
rect 56715 15679 56757 15688
rect 56620 15560 56660 15569
rect 56620 14057 56660 15520
rect 56716 14813 56756 15679
rect 57099 15560 57141 15569
rect 57099 15520 57100 15560
rect 57140 15520 57141 15560
rect 57099 15511 57141 15520
rect 56907 15140 56949 15149
rect 56907 15100 56908 15140
rect 56948 15100 56949 15140
rect 56907 15091 56949 15100
rect 56715 14804 56757 14813
rect 56715 14764 56716 14804
rect 56756 14764 56757 14804
rect 56715 14755 56757 14764
rect 56908 14729 56948 15091
rect 56907 14720 56949 14729
rect 56907 14680 56908 14720
rect 56948 14680 56949 14720
rect 56907 14671 56949 14680
rect 56619 14048 56661 14057
rect 56619 14008 56620 14048
rect 56660 14008 56661 14048
rect 56619 13999 56661 14008
rect 56523 13796 56565 13805
rect 56523 13756 56524 13796
rect 56564 13756 56565 13796
rect 56523 13747 56565 13756
rect 56331 13712 56373 13721
rect 56331 13672 56332 13712
rect 56372 13672 56373 13712
rect 56331 13663 56373 13672
rect 56524 13662 56564 13747
rect 56236 13336 56756 13376
rect 56236 13208 56276 13336
rect 56236 13159 56276 13168
rect 56332 13208 56372 13217
rect 55851 13084 55852 13124
rect 55892 13084 55893 13124
rect 55851 13075 55893 13084
rect 55945 13084 55988 13124
rect 56043 13084 56084 13124
rect 55755 13040 55797 13049
rect 55755 13000 55756 13040
rect 55796 13000 55797 13040
rect 55945 13040 55985 13084
rect 55945 13000 55988 13040
rect 55755 12991 55797 13000
rect 55659 12956 55701 12965
rect 55180 12536 55220 12545
rect 55180 11201 55220 12496
rect 55276 12452 55316 12940
rect 55659 12916 55660 12956
rect 55700 12916 55701 12956
rect 55659 12907 55701 12916
rect 55563 12704 55605 12713
rect 55563 12664 55564 12704
rect 55604 12664 55605 12704
rect 55563 12655 55605 12664
rect 55564 12536 55604 12655
rect 55564 12487 55604 12496
rect 55276 12403 55316 12412
rect 55468 12452 55508 12461
rect 55372 12368 55412 12377
rect 55468 12368 55508 12412
rect 55756 12368 55796 12991
rect 55948 12704 55988 13000
rect 56043 12980 56083 13084
rect 56332 13049 56372 13168
rect 56427 13208 56469 13217
rect 56427 13168 56428 13208
rect 56468 13168 56469 13208
rect 56427 13159 56469 13168
rect 56524 13208 56564 13219
rect 56428 13074 56468 13159
rect 56524 13133 56564 13168
rect 56716 13208 56756 13336
rect 56716 13159 56756 13168
rect 56523 13124 56565 13133
rect 56523 13084 56524 13124
rect 56564 13084 56565 13124
rect 56523 13075 56565 13084
rect 56331 13040 56373 13049
rect 56331 13000 56332 13040
rect 56372 13000 56373 13040
rect 56331 12991 56373 13000
rect 56043 12940 56084 12980
rect 56044 12788 56084 12940
rect 56044 12748 56180 12788
rect 55945 12664 55988 12704
rect 55945 12620 55985 12664
rect 56043 12620 56085 12629
rect 55945 12580 55988 12620
rect 55468 12328 55756 12368
rect 55372 12032 55412 12328
rect 55756 12319 55796 12328
rect 55372 11992 55796 12032
rect 55275 11864 55317 11873
rect 55275 11824 55276 11864
rect 55316 11824 55317 11864
rect 55275 11815 55317 11824
rect 55276 11696 55316 11815
rect 55467 11780 55509 11789
rect 55467 11740 55468 11780
rect 55508 11740 55509 11780
rect 55467 11731 55509 11740
rect 55756 11738 55796 11992
rect 55372 11696 55412 11705
rect 55276 11656 55372 11696
rect 55372 11647 55412 11656
rect 55179 11192 55221 11201
rect 55179 11152 55180 11192
rect 55220 11152 55221 11192
rect 55179 11143 55221 11152
rect 55180 11033 55220 11143
rect 55179 11024 55221 11033
rect 55372 11024 55412 11033
rect 55179 10984 55180 11024
rect 55220 10984 55221 11024
rect 55179 10975 55221 10984
rect 55276 10984 55372 11024
rect 54795 10940 54837 10949
rect 54795 10900 54796 10940
rect 54836 10900 54837 10940
rect 54795 10891 54837 10900
rect 55083 10940 55125 10949
rect 55083 10900 55084 10940
rect 55124 10900 55125 10940
rect 55083 10891 55125 10900
rect 54796 10781 54836 10891
rect 55180 10890 55220 10975
rect 54795 10772 54837 10781
rect 55180 10772 55220 10781
rect 54795 10732 54796 10772
rect 54836 10732 54837 10772
rect 54795 10723 54837 10732
rect 54892 10732 55180 10772
rect 54892 10268 54932 10732
rect 55180 10723 55220 10732
rect 54987 10352 55029 10361
rect 54987 10312 54988 10352
rect 55028 10312 55029 10352
rect 54987 10303 55029 10312
rect 54892 10219 54932 10228
rect 54988 10218 55028 10303
rect 55083 10268 55125 10277
rect 55083 10228 55084 10268
rect 55124 10228 55125 10268
rect 55083 10219 55125 10228
rect 54796 10184 54836 10193
rect 54699 10100 54741 10109
rect 54699 10060 54700 10100
rect 54740 10060 54741 10100
rect 54699 10051 54741 10060
rect 53835 9680 53877 9689
rect 53835 9640 53836 9680
rect 53876 9640 53877 9680
rect 53835 9631 53877 9640
rect 53452 9547 53492 9556
rect 53836 9512 53876 9631
rect 53355 9344 53397 9353
rect 53355 9304 53356 9344
rect 53396 9304 53397 9344
rect 53355 9295 53397 9304
rect 53164 8672 53204 8681
rect 53012 8632 53164 8672
rect 52972 8623 53012 8632
rect 53067 7916 53109 7925
rect 53067 7876 53068 7916
rect 53108 7876 53109 7916
rect 53067 7867 53109 7876
rect 53068 7782 53108 7867
rect 52875 7412 52917 7421
rect 52875 7372 52876 7412
rect 52916 7372 52917 7412
rect 52875 7363 52917 7372
rect 52588 7001 52628 7120
rect 52107 6992 52149 7001
rect 52107 6952 52108 6992
rect 52148 6952 52149 6992
rect 52107 6943 52149 6952
rect 52587 6992 52629 7001
rect 52587 6952 52588 6992
rect 52628 6952 52629 6992
rect 52587 6943 52629 6952
rect 51915 6320 51957 6329
rect 51915 6280 51916 6320
rect 51956 6280 51957 6320
rect 51915 6271 51957 6280
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 52108 5648 52148 6943
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 52683 6656 52725 6665
rect 52683 6616 52684 6656
rect 52724 6616 52725 6656
rect 52683 6607 52725 6616
rect 52780 6660 52820 6669
rect 52876 6665 52916 7363
rect 53164 7220 53204 8632
rect 53356 8168 53396 9295
rect 53836 8177 53876 9472
rect 54700 9512 54740 10051
rect 54796 10025 54836 10144
rect 55084 10134 55124 10219
rect 55180 10184 55220 10195
rect 55180 10109 55220 10144
rect 55179 10100 55221 10109
rect 55179 10060 55180 10100
rect 55220 10060 55221 10100
rect 55179 10051 55221 10060
rect 54795 10016 54837 10025
rect 54795 9976 54796 10016
rect 54836 9976 54837 10016
rect 54795 9967 54837 9976
rect 54700 9463 54740 9472
rect 54507 8672 54549 8681
rect 54507 8632 54508 8672
rect 54548 8632 54549 8672
rect 54796 8672 54836 9967
rect 55276 9764 55316 10984
rect 55372 10975 55412 10984
rect 55468 11024 55508 11731
rect 55948 11705 55988 12580
rect 56043 12580 56044 12620
rect 56084 12580 56085 12620
rect 56043 12571 56085 12580
rect 56044 12536 56084 12571
rect 56140 12545 56180 12748
rect 56236 12713 56276 12798
rect 56235 12708 56277 12713
rect 56235 12664 56236 12708
rect 56276 12664 56277 12708
rect 56235 12655 56277 12664
rect 56044 12485 56084 12496
rect 56139 12536 56181 12545
rect 56139 12496 56140 12536
rect 56180 12496 56181 12536
rect 56139 12487 56181 12496
rect 56140 12402 56180 12487
rect 56139 12032 56181 12041
rect 56139 11992 56140 12032
rect 56180 11992 56181 12032
rect 56139 11983 56181 11992
rect 56043 11948 56085 11957
rect 56043 11908 56044 11948
rect 56084 11908 56085 11948
rect 56043 11899 56085 11908
rect 55756 11689 55796 11698
rect 55947 11696 55989 11705
rect 55947 11656 55948 11696
rect 55988 11656 55989 11696
rect 55947 11647 55989 11656
rect 56044 11696 56084 11899
rect 56140 11738 56180 11983
rect 56236 11957 56276 12655
rect 56428 12629 56468 12714
rect 56427 12620 56469 12629
rect 56427 12580 56428 12620
rect 56468 12580 56469 12620
rect 56427 12571 56469 12580
rect 56524 12536 56564 13075
rect 56619 12620 56661 12629
rect 56619 12580 56620 12620
rect 56660 12580 56661 12620
rect 56619 12571 56661 12580
rect 56524 12200 56564 12496
rect 56620 12536 56660 12571
rect 56620 12485 56660 12496
rect 56715 12536 56757 12545
rect 56715 12496 56716 12536
rect 56756 12496 56757 12536
rect 56715 12487 56757 12496
rect 56716 12402 56756 12487
rect 56811 12452 56853 12461
rect 56811 12412 56812 12452
rect 56852 12412 56853 12452
rect 56811 12403 56853 12412
rect 56332 12160 56564 12200
rect 56235 11948 56277 11957
rect 56235 11908 56236 11948
rect 56276 11908 56277 11948
rect 56235 11899 56277 11908
rect 56332 11705 56372 12160
rect 56523 11948 56565 11957
rect 56523 11908 56524 11948
rect 56564 11908 56565 11948
rect 56523 11899 56565 11908
rect 56524 11814 56564 11899
rect 56619 11864 56661 11873
rect 56619 11824 56620 11864
rect 56660 11824 56661 11864
rect 56619 11815 56661 11824
rect 56427 11780 56469 11789
rect 56427 11740 56428 11780
rect 56468 11740 56469 11780
rect 56427 11731 56469 11740
rect 56140 11689 56180 11698
rect 56331 11696 56373 11705
rect 56044 11647 56084 11656
rect 56236 11675 56276 11684
rect 56331 11656 56332 11696
rect 56372 11656 56373 11696
rect 56331 11647 56373 11656
rect 56428 11696 56468 11731
rect 56428 11645 56468 11656
rect 55948 11528 55988 11537
rect 55948 11369 55988 11488
rect 56043 11528 56085 11537
rect 56043 11488 56044 11528
rect 56084 11488 56085 11528
rect 56043 11479 56085 11488
rect 55563 11360 55605 11369
rect 55563 11320 55564 11360
rect 55604 11320 55605 11360
rect 55563 11311 55605 11320
rect 55947 11360 55989 11369
rect 55947 11320 55948 11360
rect 55988 11320 55989 11360
rect 55947 11311 55989 11320
rect 55468 10975 55508 10984
rect 55467 10184 55509 10193
rect 55467 10144 55468 10184
rect 55508 10144 55509 10184
rect 55467 10135 55509 10144
rect 55564 10184 55604 11311
rect 55755 11024 55797 11033
rect 55755 10984 55756 11024
rect 55796 10984 55797 11024
rect 55755 10975 55797 10984
rect 55852 11024 55892 11033
rect 55756 10890 55796 10975
rect 55852 10352 55892 10984
rect 55948 11024 55988 11033
rect 55948 10865 55988 10984
rect 56044 11024 56084 11479
rect 56139 11360 56181 11369
rect 56139 11320 56140 11360
rect 56180 11320 56181 11360
rect 56139 11311 56181 11320
rect 56044 10975 56084 10984
rect 55947 10856 55989 10865
rect 55947 10816 55948 10856
rect 55988 10816 55989 10856
rect 55947 10807 55989 10816
rect 55947 10688 55989 10697
rect 55947 10648 55948 10688
rect 55988 10648 55989 10688
rect 55947 10639 55989 10648
rect 55852 10277 55892 10312
rect 55851 10268 55893 10277
rect 55851 10228 55852 10268
rect 55892 10228 55893 10268
rect 55851 10219 55893 10228
rect 55564 10135 55604 10144
rect 55371 10100 55413 10109
rect 55371 10060 55372 10100
rect 55412 10060 55413 10100
rect 55371 10051 55413 10060
rect 55084 9724 55316 9764
rect 55372 9958 55412 10051
rect 55468 10050 55508 10135
rect 54891 8672 54933 8681
rect 54796 8632 54892 8672
rect 54932 8632 54933 8672
rect 54507 8623 54549 8632
rect 54891 8623 54933 8632
rect 55084 8672 55124 9724
rect 55372 8924 55412 9918
rect 55852 9260 55892 9269
rect 55372 8875 55412 8884
rect 55468 9220 55852 9260
rect 53356 8119 53396 8128
rect 53835 8168 53877 8177
rect 53835 8128 53836 8168
rect 53876 8128 53877 8168
rect 53835 8119 53877 8128
rect 54123 8168 54165 8177
rect 54123 8128 54124 8168
rect 54164 8128 54165 8168
rect 54123 8119 54165 8128
rect 53452 8000 53492 8009
rect 53356 7748 53396 7757
rect 53356 7337 53396 7708
rect 53452 7505 53492 7960
rect 53836 8000 53876 8009
rect 53547 7916 53589 7925
rect 53547 7876 53548 7916
rect 53588 7876 53589 7916
rect 53547 7867 53589 7876
rect 53548 7664 53588 7867
rect 53836 7664 53876 7960
rect 53932 8000 53972 8009
rect 54124 8000 54164 8119
rect 53972 7960 54124 8000
rect 53932 7951 53972 7960
rect 54124 7951 54164 7960
rect 54315 8000 54357 8009
rect 54315 7960 54316 8000
rect 54356 7960 54357 8000
rect 54315 7951 54357 7960
rect 54508 8000 54548 8623
rect 54892 8538 54932 8623
rect 54988 8504 55028 8513
rect 54700 8177 54740 8181
rect 54699 8172 54741 8177
rect 54699 8128 54700 8172
rect 54740 8128 54741 8172
rect 54699 8119 54741 8128
rect 54700 8037 54740 8119
rect 54795 8084 54837 8093
rect 54795 8044 54796 8084
rect 54836 8044 54837 8084
rect 54795 8035 54837 8044
rect 54220 7916 54260 7925
rect 54220 7757 54260 7876
rect 54316 7832 54356 7951
rect 54411 7916 54453 7925
rect 54411 7876 54412 7916
rect 54452 7876 54453 7916
rect 54411 7867 54453 7876
rect 54316 7783 54356 7792
rect 54412 7782 54452 7867
rect 54219 7748 54261 7757
rect 54219 7708 54220 7748
rect 54260 7708 54261 7748
rect 54219 7699 54261 7708
rect 53548 7624 53876 7664
rect 53451 7496 53493 7505
rect 53451 7456 53452 7496
rect 53492 7456 53493 7496
rect 53451 7447 53493 7456
rect 53355 7328 53397 7337
rect 53355 7288 53356 7328
rect 53396 7288 53397 7328
rect 53355 7279 53397 7288
rect 53068 7180 53396 7220
rect 52587 6488 52629 6497
rect 52587 6448 52588 6488
rect 52628 6448 52629 6488
rect 52587 6439 52629 6448
rect 52684 6488 52724 6607
rect 52684 6439 52724 6448
rect 52588 6354 52628 6439
rect 52299 6320 52341 6329
rect 52780 6320 52820 6620
rect 52875 6656 52917 6665
rect 52875 6616 52876 6656
rect 52916 6616 52917 6656
rect 52875 6607 52917 6616
rect 52972 6488 53012 6499
rect 52972 6413 53012 6448
rect 52971 6404 53013 6413
rect 52971 6364 52972 6404
rect 53012 6364 53013 6404
rect 52971 6355 53013 6364
rect 51724 5564 51764 5573
rect 45771 4976 45813 4985
rect 45771 4936 45772 4976
rect 45812 4936 45813 4976
rect 45771 4927 45813 4936
rect 51724 4817 51764 5524
rect 51723 4808 51765 4817
rect 51723 4768 51724 4808
rect 51764 4768 51765 4808
rect 51723 4759 51765 4768
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 52108 3977 52148 5608
rect 52204 6280 52300 6320
rect 52340 6280 52341 6320
rect 52204 5144 52244 6280
rect 52299 6271 52341 6280
rect 52684 6280 52820 6320
rect 52300 6186 52340 6271
rect 52684 5741 52724 6280
rect 52972 6236 53012 6245
rect 52780 6196 52972 6236
rect 52683 5732 52725 5741
rect 52683 5692 52684 5732
rect 52724 5692 52725 5732
rect 52683 5683 52725 5692
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 52780 5144 52820 6196
rect 52972 6187 53012 6196
rect 52875 5732 52917 5741
rect 52875 5692 52876 5732
rect 52916 5692 52917 5732
rect 52875 5683 52917 5692
rect 52204 5104 52340 5144
rect 52204 4976 52244 4987
rect 52204 4901 52244 4936
rect 52203 4892 52245 4901
rect 52203 4852 52204 4892
rect 52244 4852 52245 4892
rect 52203 4843 52245 4852
rect 52300 4892 52340 5104
rect 52300 4843 52340 4852
rect 52492 5104 52820 5144
rect 52492 4892 52532 5104
rect 52492 4843 52532 4852
rect 52588 4976 52628 4985
rect 52588 4817 52628 4936
rect 52876 4901 52916 5683
rect 52972 5648 53012 5657
rect 53068 5648 53108 7180
rect 53356 7160 53396 7180
rect 53452 7160 53492 7169
rect 53356 7120 53452 7160
rect 53452 7111 53492 7120
rect 53548 6824 53588 7624
rect 53643 7496 53685 7505
rect 53643 7456 53644 7496
rect 53684 7456 53685 7496
rect 53643 7447 53685 7456
rect 53278 6784 53588 6824
rect 53163 6656 53205 6665
rect 53163 6616 53164 6656
rect 53204 6616 53205 6656
rect 53163 6607 53205 6616
rect 53164 6488 53204 6607
rect 53164 6439 53204 6448
rect 53278 6495 53318 6784
rect 53548 6581 53588 6612
rect 53547 6572 53589 6581
rect 53547 6532 53548 6572
rect 53588 6532 53589 6572
rect 53547 6523 53589 6532
rect 53278 6446 53318 6455
rect 53451 6488 53493 6497
rect 53451 6448 53452 6488
rect 53492 6448 53493 6488
rect 53451 6439 53493 6448
rect 53548 6488 53588 6523
rect 53452 6354 53492 6439
rect 53548 6329 53588 6448
rect 53644 6488 53684 7447
rect 53739 7412 53781 7421
rect 53739 7372 53740 7412
rect 53780 7372 53781 7412
rect 53739 7363 53781 7372
rect 53644 6439 53684 6448
rect 53740 6488 53780 7363
rect 54508 7220 54548 7960
rect 54796 8000 54836 8035
rect 54603 7496 54645 7505
rect 54603 7456 54604 7496
rect 54644 7456 54645 7496
rect 54603 7447 54645 7456
rect 54604 7412 54644 7447
rect 54796 7421 54836 7960
rect 54891 8000 54933 8009
rect 54891 7960 54892 8000
rect 54932 7960 54933 8000
rect 54891 7951 54933 7960
rect 54892 7866 54932 7951
rect 54988 7925 55028 8464
rect 54987 7916 55029 7925
rect 54987 7876 54988 7916
rect 55028 7876 55029 7916
rect 54987 7867 55029 7876
rect 54604 7361 54644 7372
rect 54795 7412 54837 7421
rect 54795 7372 54796 7412
rect 54836 7372 54837 7412
rect 54795 7363 54837 7372
rect 54412 7180 54548 7220
rect 54219 6656 54261 6665
rect 54219 6616 54220 6656
rect 54260 6616 54261 6656
rect 54219 6607 54261 6616
rect 53740 6439 53780 6448
rect 53163 6320 53205 6329
rect 53163 6280 53164 6320
rect 53204 6280 53205 6320
rect 53163 6271 53205 6280
rect 53547 6320 53589 6329
rect 53547 6280 53548 6320
rect 53588 6280 53589 6320
rect 53547 6271 53589 6280
rect 53012 5608 53108 5648
rect 52972 5599 53012 5608
rect 52875 4892 52917 4901
rect 52875 4852 52876 4892
rect 52916 4852 52917 4892
rect 52875 4843 52917 4852
rect 52395 4808 52437 4817
rect 52395 4768 52396 4808
rect 52436 4768 52437 4808
rect 52395 4759 52437 4768
rect 52587 4808 52629 4817
rect 52587 4768 52588 4808
rect 52628 4768 52629 4808
rect 52587 4759 52629 4768
rect 52396 4674 52436 4759
rect 53068 4313 53108 5608
rect 53164 4817 53204 6271
rect 54220 5825 54260 6607
rect 54219 5816 54261 5825
rect 54219 5776 54220 5816
rect 54260 5776 54261 5816
rect 54219 5767 54261 5776
rect 54124 5480 54164 5489
rect 53932 5440 54124 5480
rect 53452 4976 53492 4985
rect 53932 4976 53972 5440
rect 54124 5431 54164 5440
rect 54220 5312 54260 5767
rect 53492 4936 53932 4976
rect 53452 4927 53492 4936
rect 53932 4927 53972 4936
rect 54028 5272 54260 5312
rect 54028 4976 54068 5272
rect 54220 4976 54260 4985
rect 54028 4927 54068 4936
rect 54124 4936 54220 4976
rect 53355 4892 53397 4901
rect 53355 4852 53356 4892
rect 53396 4852 53397 4892
rect 53355 4843 53397 4852
rect 53163 4808 53205 4817
rect 53163 4768 53164 4808
rect 53204 4768 53205 4808
rect 53163 4759 53205 4768
rect 53356 4758 53396 4843
rect 54124 4817 54164 4936
rect 54220 4927 54260 4936
rect 54412 4976 54452 7180
rect 55084 6824 55124 8632
rect 55180 8672 55220 8681
rect 55468 8672 55508 9220
rect 55852 9211 55892 9220
rect 55220 8632 55468 8672
rect 55180 8623 55220 8632
rect 55468 8623 55508 8632
rect 55755 8672 55797 8681
rect 55755 8632 55756 8672
rect 55796 8632 55797 8672
rect 55755 8623 55797 8632
rect 55660 8588 55700 8597
rect 55564 8548 55660 8588
rect 55372 8168 55412 8177
rect 55564 8168 55604 8548
rect 55660 8539 55700 8548
rect 55659 8420 55701 8429
rect 55659 8380 55660 8420
rect 55700 8380 55701 8420
rect 55659 8371 55701 8380
rect 55412 8128 55604 8168
rect 55372 8119 55412 8128
rect 55468 8000 55508 8009
rect 55468 7757 55508 7960
rect 55564 8000 55604 8009
rect 55564 7841 55604 7960
rect 55660 8000 55700 8371
rect 55563 7832 55605 7841
rect 55563 7792 55564 7832
rect 55604 7792 55605 7832
rect 55563 7783 55605 7792
rect 55179 7748 55221 7757
rect 55179 7708 55180 7748
rect 55220 7708 55221 7748
rect 55179 7699 55221 7708
rect 55467 7748 55509 7757
rect 55467 7708 55468 7748
rect 55508 7708 55509 7748
rect 55467 7699 55509 7708
rect 55180 7614 55220 7699
rect 55275 7076 55317 7085
rect 55275 7036 55276 7076
rect 55316 7036 55317 7076
rect 55275 7027 55317 7036
rect 54988 6784 55124 6824
rect 54988 6665 55028 6784
rect 54987 6656 55029 6665
rect 54987 6616 54988 6656
rect 55028 6616 55029 6656
rect 54987 6607 55029 6616
rect 55083 6572 55125 6581
rect 55083 6532 55084 6572
rect 55124 6532 55125 6572
rect 55083 6523 55125 6532
rect 55084 6438 55124 6523
rect 55180 6488 55220 6497
rect 55180 5816 55220 6448
rect 55276 6488 55316 7027
rect 55563 6572 55605 6581
rect 55563 6532 55564 6572
rect 55604 6532 55605 6572
rect 55563 6523 55605 6532
rect 55276 6439 55316 6448
rect 55371 6488 55413 6497
rect 55371 6448 55372 6488
rect 55412 6448 55413 6488
rect 55371 6439 55413 6448
rect 55372 6354 55412 6439
rect 55564 6438 55604 6523
rect 55660 6497 55700 7960
rect 55756 6581 55796 8623
rect 55851 8000 55893 8009
rect 55851 7960 55852 8000
rect 55892 7960 55893 8000
rect 55851 7951 55893 7960
rect 55948 8000 55988 10639
rect 56043 10016 56085 10025
rect 56043 9976 56044 10016
rect 56084 9976 56085 10016
rect 56043 9967 56085 9976
rect 56044 9882 56084 9967
rect 56140 9437 56180 11311
rect 56236 11192 56276 11635
rect 56236 11152 56372 11192
rect 56235 11024 56277 11033
rect 56235 10984 56236 11024
rect 56276 10984 56277 11024
rect 56235 10975 56277 10984
rect 56236 10890 56276 10975
rect 56235 10436 56277 10445
rect 56235 10396 56236 10436
rect 56276 10396 56277 10436
rect 56235 10387 56277 10396
rect 56236 10277 56276 10387
rect 56235 10268 56277 10277
rect 56235 10228 56236 10268
rect 56276 10228 56277 10268
rect 56235 10219 56277 10228
rect 56236 10134 56276 10219
rect 56332 10193 56372 11152
rect 56620 11024 56660 11815
rect 56620 10975 56660 10984
rect 56523 10352 56565 10361
rect 56523 10312 56524 10352
rect 56564 10312 56565 10352
rect 56523 10303 56565 10312
rect 56331 10184 56373 10193
rect 56331 10144 56332 10184
rect 56372 10144 56373 10184
rect 56331 10135 56373 10144
rect 56139 9428 56181 9437
rect 56332 9428 56372 10135
rect 56139 9388 56140 9428
rect 56180 9388 56181 9428
rect 56139 9379 56181 9388
rect 56236 9388 56372 9428
rect 56140 9294 56180 9379
rect 56043 8672 56085 8681
rect 56043 8632 56044 8672
rect 56084 8632 56085 8672
rect 56043 8623 56085 8632
rect 56044 8538 56084 8623
rect 56236 8588 56276 9388
rect 56331 9260 56373 9269
rect 56331 9220 56332 9260
rect 56372 9220 56373 9260
rect 56331 9211 56373 9220
rect 56332 8681 56372 9211
rect 56331 8672 56373 8681
rect 56331 8632 56332 8672
rect 56372 8632 56373 8672
rect 56331 8623 56373 8632
rect 56140 8548 56276 8588
rect 56140 8093 56180 8548
rect 56139 8084 56181 8093
rect 56139 8044 56140 8084
rect 56180 8044 56181 8084
rect 56139 8035 56181 8044
rect 55852 7866 55892 7951
rect 55948 6824 55988 7960
rect 56043 8000 56085 8009
rect 56043 7960 56044 8000
rect 56084 7960 56085 8000
rect 56043 7951 56085 7960
rect 56140 8000 56180 8035
rect 56140 7951 56180 7960
rect 56044 7866 56084 7951
rect 56236 7244 56276 7253
rect 56524 7244 56564 10303
rect 56812 7505 56852 12403
rect 56908 10781 56948 14671
rect 57100 13208 57140 15511
rect 57196 13469 57236 16192
rect 58060 16232 58100 16241
rect 58060 16148 58100 16192
rect 58155 16232 58197 16241
rect 58155 16192 58156 16232
rect 58196 16192 58197 16232
rect 58155 16183 58197 16192
rect 58252 16232 58292 16241
rect 58636 16232 58676 16241
rect 57868 16108 58100 16148
rect 57292 16064 57332 16073
rect 57195 13460 57237 13469
rect 57195 13420 57196 13460
rect 57236 13420 57237 13460
rect 57195 13411 57237 13420
rect 57100 12545 57140 13168
rect 57196 12629 57236 13411
rect 57292 13217 57332 16024
rect 57771 15980 57813 15989
rect 57771 15940 57772 15980
rect 57812 15940 57813 15980
rect 57771 15931 57813 15940
rect 57772 15728 57812 15931
rect 57772 15679 57812 15688
rect 57868 15485 57908 16108
rect 57963 15812 58005 15821
rect 57963 15772 57964 15812
rect 58004 15772 58005 15812
rect 57963 15763 58005 15772
rect 57964 15644 58004 15763
rect 57964 15595 58004 15604
rect 57867 15476 57909 15485
rect 57867 15436 57868 15476
rect 57908 15436 57909 15476
rect 57867 15427 57909 15436
rect 58252 14972 58292 16192
rect 58444 16192 58636 16232
rect 58348 16064 58388 16073
rect 58348 15821 58388 16024
rect 58347 15812 58389 15821
rect 58347 15772 58348 15812
rect 58388 15772 58389 15812
rect 58347 15763 58389 15772
rect 58444 15653 58484 16192
rect 58636 16183 58676 16192
rect 58732 16232 58772 16267
rect 58732 16181 58772 16192
rect 58828 16232 58868 16241
rect 58539 15812 58581 15821
rect 58539 15772 58540 15812
rect 58580 15772 58581 15812
rect 58539 15763 58581 15772
rect 58443 15644 58485 15653
rect 58443 15604 58444 15644
rect 58484 15604 58485 15644
rect 58443 15595 58485 15604
rect 58347 15560 58389 15569
rect 58347 15520 58348 15560
rect 58388 15520 58389 15560
rect 58347 15511 58389 15520
rect 58348 15426 58388 15511
rect 58443 15140 58485 15149
rect 58443 15100 58444 15140
rect 58484 15100 58485 15140
rect 58443 15091 58485 15100
rect 58156 14932 58252 14972
rect 57579 14804 57621 14813
rect 57579 14764 57580 14804
rect 57620 14764 57621 14804
rect 57579 14755 57621 14764
rect 57387 14132 57429 14141
rect 57387 14092 57388 14132
rect 57428 14092 57429 14132
rect 57387 14083 57429 14092
rect 57388 13973 57428 14083
rect 57387 13964 57429 13973
rect 57387 13924 57388 13964
rect 57428 13924 57429 13964
rect 57387 13915 57429 13924
rect 57580 13301 57620 14755
rect 57963 14048 58005 14057
rect 57963 14008 57964 14048
rect 58004 14008 58005 14048
rect 57963 13999 58005 14008
rect 58060 14048 58100 14059
rect 57675 13880 57717 13889
rect 57675 13840 57676 13880
rect 57716 13840 57717 13880
rect 57675 13831 57717 13840
rect 57579 13292 57621 13301
rect 57579 13252 57580 13292
rect 57620 13252 57621 13292
rect 57579 13243 57621 13252
rect 57291 13208 57333 13217
rect 57291 13168 57292 13208
rect 57332 13168 57333 13208
rect 57291 13159 57333 13168
rect 57195 12620 57237 12629
rect 57195 12580 57196 12620
rect 57236 12580 57237 12620
rect 57195 12571 57237 12580
rect 57676 12620 57716 13831
rect 57964 13217 58004 13999
rect 58060 13973 58100 14008
rect 58059 13964 58101 13973
rect 58059 13924 58060 13964
rect 58100 13924 58101 13964
rect 58059 13915 58101 13924
rect 58156 13964 58196 14932
rect 58252 14923 58292 14932
rect 58444 14216 58484 15091
rect 58540 14720 58580 15763
rect 58635 15560 58677 15569
rect 58635 15520 58636 15560
rect 58676 15520 58677 15560
rect 58635 15511 58677 15520
rect 58636 15233 58676 15511
rect 58828 15485 58868 16192
rect 58924 16064 58964 16073
rect 58924 15821 58964 16024
rect 58923 15812 58965 15821
rect 58923 15772 58924 15812
rect 58964 15772 58965 15812
rect 58923 15763 58965 15772
rect 58827 15476 58869 15485
rect 58827 15436 58828 15476
rect 58868 15436 58869 15476
rect 58827 15427 58869 15436
rect 58635 15224 58677 15233
rect 58635 15184 58636 15224
rect 58676 15184 58677 15224
rect 58635 15175 58677 15184
rect 58828 14972 58868 15427
rect 59020 15401 59060 17032
rect 59595 17023 59637 17032
rect 59596 16484 59636 17023
rect 59116 16316 59156 16325
rect 59116 15905 59156 16276
rect 59499 16316 59541 16325
rect 59499 16276 59500 16316
rect 59540 16276 59541 16316
rect 59499 16267 59541 16276
rect 59500 16232 59540 16267
rect 59596 16241 59636 16444
rect 59500 16181 59540 16192
rect 59595 16232 59637 16241
rect 59595 16192 59596 16232
rect 59636 16192 59637 16232
rect 59595 16183 59637 16192
rect 59308 16064 59348 16073
rect 59348 16024 59444 16064
rect 59308 16015 59348 16024
rect 59115 15896 59157 15905
rect 59115 15856 59116 15896
rect 59156 15856 59157 15896
rect 59115 15847 59157 15856
rect 59404 15821 59444 16024
rect 59403 15812 59445 15821
rect 59403 15772 59404 15812
rect 59444 15772 59445 15812
rect 59403 15763 59445 15772
rect 59115 15728 59157 15737
rect 59115 15688 59116 15728
rect 59156 15688 59157 15728
rect 59115 15679 59157 15688
rect 59019 15392 59061 15401
rect 59019 15352 59020 15392
rect 59060 15352 59061 15392
rect 59019 15343 59061 15352
rect 58924 14972 58964 14981
rect 58828 14932 58924 14972
rect 58924 14923 58964 14932
rect 59116 14804 59156 15679
rect 59116 14755 59156 14764
rect 59212 15560 59252 15569
rect 58540 14671 58580 14680
rect 58635 14720 58677 14729
rect 58635 14680 58636 14720
rect 58676 14680 58677 14720
rect 58635 14671 58677 14680
rect 58636 14586 58676 14671
rect 58923 14552 58965 14561
rect 58923 14512 58924 14552
rect 58964 14512 58965 14552
rect 58923 14503 58965 14512
rect 59115 14552 59157 14561
rect 59115 14512 59116 14552
rect 59156 14512 59157 14552
rect 59115 14503 59157 14512
rect 58732 14494 58772 14503
rect 58444 14176 58580 14216
rect 58444 14048 58484 14057
rect 58156 13915 58196 13924
rect 58348 13964 58388 13973
rect 58251 13880 58293 13889
rect 58251 13840 58252 13880
rect 58292 13840 58293 13880
rect 58251 13831 58293 13840
rect 58252 13746 58292 13831
rect 58059 13712 58101 13721
rect 58059 13672 58060 13712
rect 58100 13672 58101 13712
rect 58059 13663 58101 13672
rect 57963 13208 58005 13217
rect 57676 12571 57716 12580
rect 57772 13168 57964 13208
rect 58004 13168 58005 13208
rect 57099 12536 57141 12545
rect 57099 12496 57100 12536
rect 57140 12496 57141 12536
rect 57099 12487 57141 12496
rect 57100 11873 57140 12487
rect 57099 11864 57141 11873
rect 57099 11824 57100 11864
rect 57140 11824 57141 11864
rect 57099 11815 57141 11824
rect 57772 11033 57812 13168
rect 57963 13159 58005 13168
rect 57964 13074 58004 13159
rect 58060 12980 58100 13663
rect 57964 12940 58100 12980
rect 57483 11024 57525 11033
rect 57483 10984 57484 11024
rect 57524 10984 57525 11024
rect 57483 10975 57525 10984
rect 57771 11024 57813 11033
rect 57771 10984 57772 11024
rect 57812 10984 57813 11024
rect 57771 10975 57813 10984
rect 57484 10890 57524 10975
rect 56907 10772 56949 10781
rect 56907 10732 56908 10772
rect 56948 10732 56949 10772
rect 56907 10723 56949 10732
rect 56908 10361 56948 10723
rect 56907 10352 56949 10361
rect 56907 10312 56908 10352
rect 56948 10312 56949 10352
rect 56907 10303 56949 10312
rect 57099 9512 57141 9521
rect 57099 9472 57100 9512
rect 57140 9472 57141 9512
rect 57099 9463 57141 9472
rect 57484 9512 57524 9521
rect 57100 9378 57140 9463
rect 57484 9269 57524 9472
rect 57483 9260 57525 9269
rect 57483 9220 57484 9260
rect 57524 9220 57525 9260
rect 57483 9211 57525 9220
rect 57867 9092 57909 9101
rect 57867 9052 57868 9092
rect 57908 9052 57909 9092
rect 57867 9043 57909 9052
rect 56907 8672 56949 8681
rect 56907 8632 56908 8672
rect 56948 8632 56949 8672
rect 56907 8623 56949 8632
rect 56908 8538 56948 8623
rect 56811 7496 56853 7505
rect 56811 7456 56812 7496
rect 56852 7456 56853 7496
rect 56811 7447 56853 7456
rect 56276 7204 56564 7244
rect 56236 7195 56276 7204
rect 56620 7160 56660 7169
rect 56044 6992 56084 7001
rect 56084 6952 56276 6992
rect 56044 6943 56084 6952
rect 55948 6784 56084 6824
rect 55755 6572 55797 6581
rect 55755 6532 55756 6572
rect 55796 6532 55797 6572
rect 55755 6523 55797 6532
rect 55947 6572 55989 6581
rect 55947 6532 55948 6572
rect 55988 6532 55989 6572
rect 55947 6523 55989 6532
rect 55659 6488 55701 6497
rect 55659 6448 55660 6488
rect 55700 6448 55701 6488
rect 55659 6439 55701 6448
rect 55948 6488 55988 6523
rect 55948 6437 55988 6448
rect 56044 6329 56084 6784
rect 56043 6320 56085 6329
rect 56043 6280 56044 6320
rect 56084 6280 56085 6320
rect 56043 6271 56085 6280
rect 54795 5144 54837 5153
rect 54795 5104 54796 5144
rect 54836 5104 54837 5144
rect 54795 5095 54837 5104
rect 54123 4808 54165 4817
rect 54123 4768 54124 4808
rect 54164 4768 54165 4808
rect 54123 4759 54165 4768
rect 54219 4724 54261 4733
rect 54219 4684 54220 4724
rect 54260 4684 54261 4724
rect 54219 4675 54261 4684
rect 54220 4590 54260 4675
rect 53067 4304 53109 4313
rect 53067 4264 53068 4304
rect 53108 4264 53109 4304
rect 53067 4255 53109 4264
rect 53835 4220 53877 4229
rect 53835 4180 53836 4220
rect 53876 4180 53877 4220
rect 53835 4171 53877 4180
rect 53836 4136 53876 4171
rect 54412 4145 54452 4936
rect 54796 4976 54836 5095
rect 54796 4927 54836 4936
rect 55180 4901 55220 5776
rect 55468 5776 55988 5816
rect 55468 5648 55508 5776
rect 55468 5599 55508 5608
rect 55563 5648 55605 5657
rect 55563 5608 55564 5648
rect 55604 5608 55605 5648
rect 55563 5599 55605 5608
rect 55948 5648 55988 5776
rect 55948 5599 55988 5608
rect 56044 5648 56084 6271
rect 56236 5657 56276 6952
rect 56620 6917 56660 7120
rect 57099 7160 57141 7169
rect 57099 7120 57100 7160
rect 57140 7120 57141 7160
rect 57099 7111 57141 7120
rect 57484 7160 57524 7169
rect 57524 7120 57620 7160
rect 57484 7111 57524 7120
rect 56715 7076 56757 7085
rect 56715 7036 56716 7076
rect 56756 7036 56757 7076
rect 56715 7027 56757 7036
rect 56716 6942 56756 7027
rect 57100 7026 57140 7111
rect 56331 6908 56373 6917
rect 56331 6868 56332 6908
rect 56372 6868 56373 6908
rect 56331 6859 56373 6868
rect 56619 6908 56661 6917
rect 56619 6868 56620 6908
rect 56660 6868 56661 6908
rect 56619 6859 56661 6868
rect 55564 5514 55604 5599
rect 55660 5422 55700 5431
rect 55660 5144 55700 5382
rect 55755 5144 55797 5153
rect 55660 5104 55756 5144
rect 55796 5104 55797 5144
rect 55755 5095 55797 5104
rect 55756 5010 55796 5095
rect 55851 4976 55893 4985
rect 55851 4936 55852 4976
rect 55892 4936 55893 4976
rect 55851 4927 55893 4936
rect 54508 4892 54548 4901
rect 54508 4733 54548 4852
rect 54699 4892 54741 4901
rect 54699 4852 54700 4892
rect 54740 4852 54741 4892
rect 54699 4843 54741 4852
rect 55179 4892 55221 4901
rect 55179 4852 55180 4892
rect 55220 4852 55221 4892
rect 55179 4843 55221 4852
rect 54604 4808 54644 4817
rect 54507 4724 54549 4733
rect 54507 4684 54508 4724
rect 54548 4684 54549 4724
rect 54507 4675 54549 4684
rect 54604 4229 54644 4768
rect 54700 4758 54740 4843
rect 55852 4842 55892 4927
rect 56044 4817 56084 5608
rect 56140 5648 56180 5657
rect 56140 5396 56180 5608
rect 56235 5648 56277 5657
rect 56235 5608 56236 5648
rect 56276 5608 56277 5648
rect 56235 5599 56277 5608
rect 56236 5514 56276 5599
rect 56332 5396 56372 6859
rect 57580 6581 57620 7120
rect 57868 7085 57908 9043
rect 57964 8924 58004 12940
rect 58059 12536 58101 12545
rect 58059 12496 58060 12536
rect 58100 12496 58101 12536
rect 58059 12487 58101 12496
rect 58060 12402 58100 12487
rect 58059 12116 58101 12125
rect 58059 12076 58060 12116
rect 58100 12076 58101 12116
rect 58059 12067 58101 12076
rect 58060 9092 58100 12067
rect 58251 11192 58293 11201
rect 58251 11152 58252 11192
rect 58292 11152 58293 11192
rect 58251 11143 58293 11152
rect 58252 10352 58292 11143
rect 58348 10436 58388 13924
rect 58444 11201 58484 14008
rect 58443 11192 58485 11201
rect 58443 11152 58444 11192
rect 58484 11152 58485 11192
rect 58443 11143 58485 11152
rect 58444 10436 58484 10445
rect 58348 10396 58444 10436
rect 58444 10387 58484 10396
rect 58252 10312 58388 10352
rect 58251 10184 58293 10193
rect 58251 10144 58252 10184
rect 58292 10144 58293 10184
rect 58251 10135 58293 10144
rect 58252 10050 58292 10135
rect 58155 10016 58197 10025
rect 58155 9976 58156 10016
rect 58196 9976 58197 10016
rect 58348 10016 58388 10312
rect 58443 10268 58485 10277
rect 58443 10228 58444 10268
rect 58484 10228 58485 10268
rect 58443 10219 58485 10228
rect 58444 10184 58484 10219
rect 58444 10133 58484 10144
rect 58348 9976 58484 10016
rect 58155 9967 58197 9976
rect 58156 9882 58196 9967
rect 58348 9512 58388 9521
rect 58252 9472 58348 9512
rect 58060 9052 58196 9092
rect 58060 8924 58100 8933
rect 57964 8884 58060 8924
rect 57964 8009 58004 8884
rect 58060 8875 58100 8884
rect 57963 8000 58005 8009
rect 57963 7960 57964 8000
rect 58004 7960 58005 8000
rect 57963 7951 58005 7960
rect 57867 7076 57909 7085
rect 57867 7036 57868 7076
rect 57908 7036 57909 7076
rect 57867 7027 57909 7036
rect 57963 6908 58005 6917
rect 57963 6868 57964 6908
rect 58004 6868 58005 6908
rect 57963 6859 58005 6868
rect 57964 6656 58004 6859
rect 57964 6607 58004 6616
rect 57579 6572 57621 6581
rect 57579 6532 57580 6572
rect 57620 6532 57621 6572
rect 57579 6523 57621 6532
rect 56811 6488 56853 6497
rect 56811 6448 56812 6488
rect 56852 6448 56853 6488
rect 56811 6439 56853 6448
rect 56812 6354 56852 6439
rect 56907 6404 56949 6413
rect 56907 6364 56908 6404
rect 56948 6364 56949 6404
rect 56907 6355 56949 6364
rect 56523 5816 56565 5825
rect 56523 5776 56524 5816
rect 56564 5776 56565 5816
rect 56523 5767 56565 5776
rect 56140 5356 56372 5396
rect 56235 4976 56277 4985
rect 56235 4936 56236 4976
rect 56276 4936 56277 4976
rect 56235 4927 56277 4936
rect 56043 4808 56085 4817
rect 56043 4768 56044 4808
rect 56084 4768 56085 4808
rect 56043 4759 56085 4768
rect 55083 4304 55125 4313
rect 55083 4264 55084 4304
rect 55124 4264 55125 4304
rect 55083 4255 55125 4264
rect 56236 4304 56276 4927
rect 56276 4264 56468 4304
rect 56236 4255 56276 4264
rect 54603 4220 54645 4229
rect 54603 4180 54604 4220
rect 54644 4180 54645 4220
rect 54603 4171 54645 4180
rect 53836 4085 53876 4096
rect 54220 4136 54260 4145
rect 54220 3977 54260 4096
rect 54411 4136 54453 4145
rect 54411 4096 54412 4136
rect 54452 4096 54453 4136
rect 54411 4087 54453 4096
rect 55084 4136 55124 4255
rect 52107 3968 52149 3977
rect 52107 3928 52108 3968
rect 52148 3928 52149 3968
rect 52107 3919 52149 3928
rect 54219 3968 54261 3977
rect 54219 3928 54220 3968
rect 54260 3928 54261 3968
rect 54219 3919 54261 3928
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 5163 3632 5205 3641
rect 5163 3592 5164 3632
rect 5204 3592 5205 3632
rect 5163 3583 5205 3592
rect 7371 3632 7413 3641
rect 7371 3592 7372 3632
rect 7412 3592 7413 3632
rect 7371 3583 7413 3592
rect 5164 3498 5204 3583
rect 55084 3473 55124 4096
rect 56331 4136 56373 4145
rect 56331 4096 56332 4136
rect 56372 4096 56373 4136
rect 56331 4087 56373 4096
rect 56428 4136 56468 4264
rect 56524 4229 56564 5767
rect 56908 4976 56948 6355
rect 57483 5648 57525 5657
rect 57483 5608 57484 5648
rect 57524 5608 57525 5648
rect 57483 5599 57525 5608
rect 56908 4927 56948 4936
rect 57003 4976 57045 4985
rect 57003 4936 57004 4976
rect 57044 4936 57045 4976
rect 57003 4927 57045 4936
rect 57100 4976 57140 4985
rect 57004 4842 57044 4927
rect 57004 4304 57044 4313
rect 57100 4304 57140 4936
rect 57196 4976 57236 4985
rect 57388 4976 57428 4985
rect 57236 4936 57388 4976
rect 57196 4927 57236 4936
rect 57388 4927 57428 4936
rect 57484 4808 57524 5599
rect 57580 4976 57620 6523
rect 58060 5732 58100 5741
rect 58156 5732 58196 9052
rect 58252 8681 58292 9472
rect 58348 9463 58388 9472
rect 58251 8672 58293 8681
rect 58251 8632 58252 8672
rect 58292 8632 58293 8672
rect 58444 8672 58484 9976
rect 58540 9101 58580 14176
rect 58732 13889 58772 14454
rect 58924 14418 58964 14503
rect 58827 14384 58869 14393
rect 58827 14344 58828 14384
rect 58868 14344 58869 14384
rect 58827 14335 58869 14344
rect 58731 13880 58773 13889
rect 58731 13840 58732 13880
rect 58772 13840 58773 13880
rect 58731 13831 58773 13840
rect 58828 13721 58868 14335
rect 58827 13712 58869 13721
rect 58827 13672 58828 13712
rect 58868 13672 58869 13712
rect 58827 13663 58869 13672
rect 59116 13628 59156 14503
rect 59212 14057 59252 15520
rect 59692 14813 59732 17107
rect 59945 17072 59985 17472
rect 60055 17165 60095 17472
rect 60054 17156 60096 17165
rect 60054 17116 60055 17156
rect 60095 17116 60096 17156
rect 60054 17107 60096 17116
rect 60345 17072 60385 17472
rect 60455 17249 60495 17472
rect 60454 17240 60496 17249
rect 60454 17200 60455 17240
rect 60495 17200 60496 17240
rect 60454 17191 60496 17200
rect 59788 17032 59985 17072
rect 60268 17032 60385 17072
rect 60745 17072 60785 17472
rect 60855 17249 60895 17472
rect 60854 17240 60896 17249
rect 60854 17200 60855 17240
rect 60895 17200 60896 17240
rect 60854 17191 60896 17200
rect 61035 17156 61077 17165
rect 61035 17116 61036 17156
rect 61076 17116 61077 17156
rect 61035 17107 61077 17116
rect 60745 17032 60788 17072
rect 59691 14804 59733 14813
rect 59691 14764 59692 14804
rect 59732 14764 59733 14804
rect 59691 14755 59733 14764
rect 59788 14225 59828 17032
rect 60075 16988 60117 16997
rect 60075 16948 60076 16988
rect 60116 16948 60117 16988
rect 60075 16939 60117 16948
rect 60076 16232 60116 16939
rect 59884 16192 60076 16232
rect 59787 14216 59829 14225
rect 59787 14176 59788 14216
rect 59828 14176 59829 14216
rect 59787 14167 59829 14176
rect 59211 14048 59253 14057
rect 59211 14008 59212 14048
rect 59252 14008 59253 14048
rect 59211 13999 59253 14008
rect 59308 14048 59348 14057
rect 59500 14048 59540 14057
rect 59348 14008 59500 14048
rect 59308 13999 59348 14008
rect 59211 13880 59253 13889
rect 59211 13840 59212 13880
rect 59252 13840 59253 13880
rect 59211 13831 59253 13840
rect 59212 13746 59252 13831
rect 59116 13588 59252 13628
rect 59115 13460 59157 13469
rect 59115 13420 59116 13460
rect 59156 13420 59157 13460
rect 59115 13411 59157 13420
rect 58923 13208 58965 13217
rect 58923 13168 58924 13208
rect 58964 13168 58965 13208
rect 58923 13159 58965 13168
rect 58924 12536 58964 13159
rect 59116 13133 59156 13411
rect 59115 13124 59157 13133
rect 59115 13084 59116 13124
rect 59156 13084 59157 13124
rect 59115 13075 59157 13084
rect 58924 12487 58964 12496
rect 58635 12032 58677 12041
rect 58635 11992 58636 12032
rect 58676 11992 58677 12032
rect 58635 11983 58677 11992
rect 58636 11192 58676 11983
rect 59020 11696 59060 11705
rect 58636 11143 58676 11152
rect 58924 11528 58964 11537
rect 58924 11108 58964 11488
rect 58924 11059 58964 11068
rect 58635 10940 58677 10949
rect 58635 10900 58636 10940
rect 58676 10900 58677 10940
rect 58635 10891 58677 10900
rect 58636 10184 58676 10891
rect 58924 10352 58964 10361
rect 59020 10352 59060 11656
rect 59115 11696 59157 11705
rect 59115 11656 59116 11696
rect 59156 11656 59157 11696
rect 59115 11647 59157 11656
rect 59212 11696 59252 13588
rect 59500 12713 59540 14008
rect 59596 14048 59636 14057
rect 59788 14048 59828 14057
rect 59596 13217 59636 14008
rect 59692 14008 59788 14048
rect 59692 13469 59732 14008
rect 59788 13999 59828 14008
rect 59787 13796 59829 13805
rect 59787 13756 59788 13796
rect 59828 13756 59829 13796
rect 59787 13747 59829 13756
rect 59788 13662 59828 13747
rect 59691 13460 59733 13469
rect 59691 13420 59692 13460
rect 59732 13420 59733 13460
rect 59691 13411 59733 13420
rect 59884 13376 59924 16192
rect 60076 16183 60116 16192
rect 60172 16064 60212 16073
rect 60075 15812 60117 15821
rect 60075 15772 60076 15812
rect 60116 15772 60117 15812
rect 60075 15763 60117 15772
rect 59980 14048 60020 14059
rect 59980 13973 60020 14008
rect 59979 13964 60021 13973
rect 59979 13924 59980 13964
rect 60020 13924 60021 13964
rect 59979 13915 60021 13924
rect 59979 13544 60021 13553
rect 59979 13504 59980 13544
rect 60020 13504 60021 13544
rect 59979 13495 60021 13504
rect 59788 13336 59924 13376
rect 59595 13208 59637 13217
rect 59595 13168 59596 13208
rect 59636 13168 59637 13208
rect 59595 13159 59637 13168
rect 59788 12980 59828 13336
rect 59980 13292 60020 13495
rect 59692 12940 59828 12980
rect 59884 13252 59980 13292
rect 59499 12704 59541 12713
rect 59499 12664 59500 12704
rect 59540 12664 59541 12704
rect 59499 12655 59541 12664
rect 59307 12536 59349 12545
rect 59307 12496 59308 12536
rect 59348 12496 59349 12536
rect 59307 12487 59349 12496
rect 59212 11647 59252 11656
rect 59116 11562 59156 11647
rect 59308 11024 59348 12487
rect 59596 11696 59636 11705
rect 59500 11528 59540 11537
rect 59308 10975 59348 10984
rect 59404 11488 59500 11528
rect 59404 10856 59444 11488
rect 59500 11479 59540 11488
rect 58828 10312 58924 10352
rect 58964 10312 59060 10352
rect 59212 10816 59444 10856
rect 58636 10109 58676 10144
rect 58731 10184 58773 10193
rect 58731 10144 58732 10184
rect 58772 10144 58773 10184
rect 58731 10135 58773 10144
rect 58635 10100 58677 10109
rect 58635 10060 58636 10100
rect 58676 10060 58677 10100
rect 58635 10051 58677 10060
rect 58636 10020 58676 10051
rect 58732 10050 58772 10135
rect 58731 9512 58773 9521
rect 58731 9472 58732 9512
rect 58772 9472 58773 9512
rect 58731 9463 58773 9472
rect 58539 9092 58581 9101
rect 58539 9052 58540 9092
rect 58580 9052 58581 9092
rect 58539 9043 58581 9052
rect 58635 8840 58677 8849
rect 58635 8800 58636 8840
rect 58676 8800 58677 8840
rect 58635 8791 58677 8800
rect 58732 8840 58772 9463
rect 58732 8791 58772 8800
rect 58636 8756 58676 8791
rect 58636 8705 58676 8716
rect 58828 8756 58868 10312
rect 58924 10303 58964 10312
rect 59212 10184 59252 10816
rect 59596 10613 59636 11656
rect 59692 11696 59732 12940
rect 59692 11201 59732 11656
rect 59788 11696 59828 11705
rect 59691 11192 59733 11201
rect 59691 11152 59692 11192
rect 59732 11152 59733 11192
rect 59691 11143 59733 11152
rect 59788 10856 59828 11656
rect 59692 10816 59828 10856
rect 59595 10604 59637 10613
rect 59595 10564 59596 10604
rect 59636 10564 59637 10604
rect 59595 10555 59637 10564
rect 59596 10436 59636 10445
rect 59692 10436 59732 10816
rect 59787 10688 59829 10697
rect 59787 10648 59788 10688
rect 59828 10648 59829 10688
rect 59787 10639 59829 10648
rect 59636 10396 59732 10436
rect 59596 10387 59636 10396
rect 59788 10268 59828 10639
rect 59788 10219 59828 10228
rect 59212 10135 59252 10144
rect 59308 10184 59348 10195
rect 59308 10109 59348 10144
rect 59499 10184 59541 10193
rect 59499 10144 59500 10184
rect 59540 10144 59541 10184
rect 59499 10135 59541 10144
rect 59115 10100 59157 10109
rect 59115 10060 59116 10100
rect 59156 10060 59157 10100
rect 59115 10051 59157 10060
rect 59307 10100 59349 10109
rect 59307 10060 59308 10100
rect 59348 10060 59349 10100
rect 59307 10051 59349 10060
rect 58923 10016 58965 10025
rect 58923 9976 58924 10016
rect 58964 9976 58965 10016
rect 58923 9967 58965 9976
rect 58828 8707 58868 8716
rect 58540 8672 58580 8681
rect 58444 8632 58540 8672
rect 58251 8623 58293 8632
rect 58540 8623 58580 8632
rect 58924 8672 58964 9967
rect 59019 9932 59061 9941
rect 59019 9892 59020 9932
rect 59060 9892 59061 9932
rect 59019 9883 59061 9892
rect 59020 8715 59060 9883
rect 59116 9101 59156 10051
rect 59403 10016 59445 10025
rect 59403 9972 59404 10016
rect 59444 9972 59445 10016
rect 59403 9967 59445 9972
rect 59404 9881 59444 9967
rect 59500 9680 59540 10135
rect 59595 10016 59637 10025
rect 59595 9976 59596 10016
rect 59636 9976 59637 10016
rect 59595 9967 59637 9976
rect 59596 9882 59636 9967
rect 59500 9631 59540 9640
rect 59884 9512 59924 13252
rect 59980 13243 60020 13252
rect 60076 13124 60116 15763
rect 60172 15401 60212 16024
rect 60171 15392 60213 15401
rect 60171 15352 60172 15392
rect 60212 15352 60213 15392
rect 60171 15343 60213 15352
rect 60172 14813 60212 15343
rect 60171 14804 60213 14813
rect 60171 14764 60172 14804
rect 60212 14764 60213 14804
rect 60171 14755 60213 14764
rect 60172 14552 60212 14561
rect 60172 13637 60212 14512
rect 60268 14309 60308 17032
rect 60748 16661 60788 17032
rect 60747 16652 60789 16661
rect 60747 16612 60748 16652
rect 60788 16612 60789 16652
rect 60747 16603 60789 16612
rect 60748 16409 60788 16422
rect 60747 16400 60789 16409
rect 60747 16360 60748 16400
rect 60788 16360 60789 16400
rect 60747 16351 60789 16360
rect 60748 16327 60788 16351
rect 60363 16316 60405 16325
rect 60363 16276 60364 16316
rect 60404 16276 60405 16316
rect 60748 16278 60788 16287
rect 60363 16267 60405 16276
rect 60364 15728 60404 16267
rect 60459 16232 60501 16241
rect 60459 16192 60460 16232
rect 60500 16192 60501 16232
rect 60459 16183 60501 16192
rect 60556 16232 60596 16243
rect 60460 16098 60500 16183
rect 60556 16157 60596 16192
rect 61036 16157 61076 17107
rect 61145 17072 61185 17472
rect 61255 17333 61295 17472
rect 61254 17324 61296 17333
rect 61254 17284 61255 17324
rect 61295 17284 61296 17324
rect 61254 17275 61296 17284
rect 61545 17072 61585 17472
rect 61132 17032 61185 17072
rect 61420 17032 61585 17072
rect 61655 17072 61695 17472
rect 61945 17072 61985 17472
rect 62055 17333 62095 17472
rect 62054 17324 62096 17333
rect 62054 17284 62055 17324
rect 62095 17284 62096 17324
rect 62054 17275 62096 17284
rect 62345 17072 62385 17472
rect 62455 17249 62495 17472
rect 62454 17240 62496 17249
rect 62454 17200 62455 17240
rect 62495 17200 62496 17240
rect 62454 17191 62496 17200
rect 61655 17032 61748 17072
rect 61132 16409 61172 17032
rect 61131 16400 61173 16409
rect 61131 16360 61132 16400
rect 61172 16360 61173 16400
rect 61131 16351 61173 16360
rect 60555 16148 60597 16157
rect 60555 16108 60556 16148
rect 60596 16108 60597 16148
rect 60555 16099 60597 16108
rect 61035 16148 61077 16157
rect 61035 16108 61036 16148
rect 61076 16108 61077 16148
rect 61035 16099 61077 16108
rect 61132 16148 61172 16157
rect 60940 16064 60980 16073
rect 60940 15905 60980 16024
rect 60939 15896 60981 15905
rect 60939 15856 60940 15896
rect 60980 15856 60981 15896
rect 60939 15847 60981 15856
rect 60364 15679 60404 15688
rect 60940 15728 60980 15737
rect 61132 15728 61172 16108
rect 61420 16073 61460 17032
rect 61516 16232 61556 16241
rect 61556 16192 61652 16232
rect 61516 16183 61556 16192
rect 61419 16064 61461 16073
rect 61419 16024 61420 16064
rect 61460 16024 61461 16064
rect 61419 16015 61461 16024
rect 61419 15896 61461 15905
rect 61419 15856 61420 15896
rect 61460 15856 61461 15896
rect 61419 15847 61461 15856
rect 60980 15688 61172 15728
rect 60940 15679 60980 15688
rect 60939 15560 60981 15569
rect 60939 15520 60940 15560
rect 60980 15520 60981 15560
rect 60939 15511 60981 15520
rect 61036 15560 61076 15569
rect 60459 15056 60501 15065
rect 60459 15016 60460 15056
rect 60500 15016 60501 15056
rect 60459 15007 60501 15016
rect 60363 14804 60405 14813
rect 60363 14764 60364 14804
rect 60404 14764 60405 14804
rect 60363 14755 60405 14764
rect 60364 14670 60404 14755
rect 60267 14300 60309 14309
rect 60267 14260 60268 14300
rect 60308 14260 60309 14300
rect 60267 14251 60309 14260
rect 60364 14048 60404 14057
rect 60460 14048 60500 15007
rect 60651 14888 60693 14897
rect 60651 14848 60652 14888
rect 60692 14848 60693 14888
rect 60651 14839 60693 14848
rect 60404 14008 60500 14048
rect 60364 13999 60404 14008
rect 60555 13964 60597 13973
rect 60555 13924 60556 13964
rect 60596 13924 60597 13964
rect 60555 13915 60597 13924
rect 60459 13796 60501 13805
rect 60459 13756 60460 13796
rect 60500 13756 60501 13796
rect 60459 13747 60501 13756
rect 60171 13628 60213 13637
rect 60171 13588 60172 13628
rect 60212 13588 60213 13628
rect 60171 13579 60213 13588
rect 60171 13460 60213 13469
rect 60171 13420 60172 13460
rect 60212 13420 60213 13460
rect 60171 13411 60213 13420
rect 60363 13460 60405 13469
rect 60363 13420 60364 13460
rect 60404 13420 60405 13460
rect 60363 13411 60405 13420
rect 60172 13326 60212 13411
rect 60267 13376 60309 13385
rect 60267 13336 60268 13376
rect 60308 13336 60309 13376
rect 60267 13327 60309 13336
rect 59980 13084 60116 13124
rect 59980 11780 60020 13084
rect 60075 12704 60117 12713
rect 60075 12664 60076 12704
rect 60116 12664 60117 12704
rect 60075 12655 60117 12664
rect 60076 12570 60116 12655
rect 60268 12620 60308 13327
rect 60364 13208 60404 13411
rect 60460 13292 60500 13747
rect 60556 13376 60596 13915
rect 60556 13327 60596 13336
rect 60460 13243 60500 13252
rect 60652 13292 60692 14839
rect 60843 14636 60885 14645
rect 60843 14596 60844 14636
rect 60884 14596 60885 14636
rect 60843 14587 60885 14596
rect 60747 13880 60789 13889
rect 60747 13840 60748 13880
rect 60788 13840 60789 13880
rect 60747 13831 60789 13840
rect 60652 13243 60692 13252
rect 60364 13159 60404 13168
rect 60748 13208 60788 13831
rect 60748 13159 60788 13168
rect 60363 12956 60405 12965
rect 60363 12916 60364 12956
rect 60404 12916 60405 12956
rect 60363 12907 60405 12916
rect 60651 12956 60693 12965
rect 60651 12916 60652 12956
rect 60692 12916 60693 12956
rect 60651 12907 60693 12916
rect 60268 12571 60308 12580
rect 59980 11731 60020 11740
rect 60172 11528 60212 11537
rect 60076 11488 60172 11528
rect 59979 10604 60021 10613
rect 59979 10564 59980 10604
rect 60020 10564 60021 10604
rect 59979 10555 60021 10564
rect 59980 10436 60020 10555
rect 59980 10387 60020 10396
rect 60076 10268 60116 11488
rect 60172 11479 60212 11488
rect 60171 11024 60213 11033
rect 60171 10984 60172 11024
rect 60212 10984 60213 11024
rect 60171 10975 60213 10984
rect 60172 10890 60212 10975
rect 60171 10268 60213 10277
rect 60076 10228 60172 10268
rect 60212 10228 60213 10268
rect 60171 10219 60213 10228
rect 60172 10134 60212 10219
rect 60267 10016 60309 10025
rect 60267 9976 60268 10016
rect 60308 9976 60309 10016
rect 60267 9967 60309 9976
rect 59212 9472 59924 9512
rect 59115 9092 59157 9101
rect 59115 9052 59116 9092
rect 59156 9052 59157 9092
rect 59115 9043 59157 9052
rect 59116 8849 59156 8934
rect 59115 8840 59157 8849
rect 59115 8800 59116 8840
rect 59156 8800 59157 8840
rect 59115 8791 59157 8800
rect 59020 8675 59156 8715
rect 58924 8623 58964 8632
rect 59116 8672 59156 8675
rect 59116 8623 59156 8632
rect 58252 7160 58292 8623
rect 59019 8588 59061 8597
rect 59019 8548 59020 8588
rect 59060 8548 59061 8588
rect 59019 8539 59061 8548
rect 58347 8168 58389 8177
rect 59020 8168 59060 8539
rect 58347 8128 58348 8168
rect 58388 8128 58389 8168
rect 58347 8119 58389 8128
rect 58636 8128 59020 8168
rect 58348 8034 58388 8119
rect 58443 8000 58485 8009
rect 58443 7960 58444 8000
rect 58484 7960 58485 8000
rect 58443 7951 58485 7960
rect 58444 7866 58484 7951
rect 58636 7916 58676 8128
rect 59020 8119 59060 8128
rect 58636 7867 58676 7876
rect 59212 7916 59252 9472
rect 60171 9428 60213 9437
rect 60171 9388 60172 9428
rect 60212 9388 60213 9428
rect 60171 9379 60213 9388
rect 60268 9428 60308 9967
rect 60268 9379 60308 9388
rect 60076 9260 60116 9269
rect 59500 9220 60076 9260
rect 59307 9092 59349 9101
rect 59307 9052 59308 9092
rect 59348 9052 59349 9092
rect 59307 9043 59349 9052
rect 59308 8672 59348 9043
rect 59308 8623 59348 8632
rect 59404 8672 59444 8681
rect 59404 8420 59444 8632
rect 59308 8380 59444 8420
rect 59308 8009 59348 8380
rect 59404 8177 59444 8263
rect 59403 8172 59445 8177
rect 59403 8128 59404 8172
rect 59444 8128 59445 8172
rect 59403 8119 59445 8128
rect 59500 8093 59540 9220
rect 60076 9211 60116 9220
rect 60172 8672 60212 9379
rect 60364 9260 60404 12907
rect 60652 12545 60692 12907
rect 60651 12536 60693 12545
rect 60651 12496 60652 12536
rect 60692 12496 60693 12536
rect 60651 12487 60693 12496
rect 60652 12402 60692 12487
rect 60651 10856 60693 10865
rect 60651 10816 60652 10856
rect 60692 10816 60693 10856
rect 60651 10807 60693 10816
rect 60555 10604 60597 10613
rect 60555 10564 60556 10604
rect 60596 10564 60597 10604
rect 60555 10555 60597 10564
rect 60459 10268 60501 10277
rect 60459 10228 60460 10268
rect 60500 10228 60501 10268
rect 60459 10219 60501 10228
rect 60460 10109 60500 10219
rect 60459 10100 60501 10109
rect 60459 10060 60460 10100
rect 60500 10060 60501 10100
rect 60459 10051 60501 10060
rect 60172 8623 60212 8632
rect 60268 9220 60404 9260
rect 59788 8588 59828 8597
rect 59828 8548 60116 8588
rect 59788 8539 59828 8548
rect 59691 8168 59733 8177
rect 59691 8128 59692 8168
rect 59732 8128 59733 8168
rect 59691 8119 59733 8128
rect 60076 8168 60116 8548
rect 60076 8119 60116 8128
rect 59499 8084 59541 8093
rect 59499 8044 59500 8084
rect 59540 8044 59541 8084
rect 59499 8035 59541 8044
rect 59307 8000 59349 8009
rect 59307 7960 59308 8000
rect 59348 7960 59349 8000
rect 59307 7951 59349 7960
rect 59500 8000 59540 8035
rect 59212 7867 59252 7876
rect 58828 7748 58868 7757
rect 58348 7160 58388 7169
rect 58252 7120 58348 7160
rect 58348 6497 58388 7120
rect 58828 7001 58868 7708
rect 59308 7412 59348 7951
rect 59500 7950 59540 7960
rect 59595 8000 59637 8009
rect 59595 7960 59596 8000
rect 59636 7960 59637 8000
rect 59595 7951 59637 7960
rect 59596 7866 59636 7951
rect 59500 7412 59540 7421
rect 59308 7372 59500 7412
rect 59500 7363 59540 7372
rect 59692 7160 59732 8119
rect 60172 8000 60212 8009
rect 59884 7748 59924 7757
rect 60172 7748 60212 7960
rect 60268 8000 60308 9220
rect 60268 7951 60308 7960
rect 60364 8000 60404 8009
rect 60460 8000 60500 10051
rect 60556 8168 60596 10555
rect 60652 10184 60692 10807
rect 60652 10135 60692 10144
rect 60844 9353 60884 14587
rect 60940 11117 60980 15511
rect 61036 14897 61076 15520
rect 61131 15560 61173 15569
rect 61131 15520 61132 15560
rect 61172 15520 61173 15560
rect 61131 15511 61173 15520
rect 61228 15560 61268 15571
rect 61132 15426 61172 15511
rect 61228 15485 61268 15520
rect 61227 15476 61269 15485
rect 61420 15476 61460 15847
rect 61612 15728 61652 16192
rect 61612 15679 61652 15688
rect 61227 15436 61228 15476
rect 61268 15436 61269 15476
rect 61227 15427 61269 15436
rect 61324 15436 61420 15476
rect 61324 15056 61364 15436
rect 61420 15427 61460 15436
rect 61612 15308 61652 15317
rect 61612 15065 61652 15268
rect 61228 15016 61364 15056
rect 61611 15056 61653 15065
rect 61611 15016 61612 15056
rect 61652 15016 61653 15056
rect 61035 14888 61077 14897
rect 61035 14848 61036 14888
rect 61076 14848 61077 14888
rect 61035 14839 61077 14848
rect 61036 14754 61076 14839
rect 61228 14384 61268 15016
rect 61611 15007 61653 15016
rect 61323 14888 61365 14897
rect 61323 14848 61324 14888
rect 61364 14848 61365 14888
rect 61323 14839 61365 14848
rect 61324 14720 61364 14839
rect 61324 14671 61364 14680
rect 61419 14720 61461 14729
rect 61419 14680 61420 14720
rect 61460 14680 61461 14720
rect 61419 14671 61461 14680
rect 61420 14586 61460 14671
rect 61516 14494 61556 14503
rect 61228 14344 61460 14384
rect 61323 14216 61365 14225
rect 61323 14176 61324 14216
rect 61364 14176 61365 14216
rect 61323 14167 61365 14176
rect 61035 14132 61077 14141
rect 61035 14092 61036 14132
rect 61076 14092 61077 14132
rect 61035 14083 61077 14092
rect 61036 12980 61076 14083
rect 61227 14048 61269 14057
rect 61227 14008 61228 14048
rect 61268 14008 61269 14048
rect 61227 13999 61269 14008
rect 61228 13049 61268 13999
rect 61227 13040 61269 13049
rect 61227 13000 61228 13040
rect 61268 13000 61269 13040
rect 61227 12991 61269 13000
rect 61036 12940 61172 12980
rect 61035 11864 61077 11873
rect 61035 11824 61036 11864
rect 61076 11824 61077 11864
rect 61035 11815 61077 11824
rect 60939 11108 60981 11117
rect 60939 11068 60940 11108
rect 60980 11068 60981 11108
rect 60939 11059 60981 11068
rect 61036 10940 61076 11815
rect 61132 11285 61172 12940
rect 61324 12797 61364 14167
rect 61323 12788 61365 12797
rect 61323 12748 61324 12788
rect 61364 12748 61365 12788
rect 61323 12739 61365 12748
rect 61228 11864 61268 11873
rect 61131 11276 61173 11285
rect 61131 11236 61132 11276
rect 61172 11236 61173 11276
rect 61131 11227 61173 11236
rect 60940 10900 61076 10940
rect 60843 9344 60885 9353
rect 60843 9304 60844 9344
rect 60884 9304 60885 9344
rect 60843 9295 60885 9304
rect 60747 8924 60789 8933
rect 60747 8884 60748 8924
rect 60788 8884 60789 8924
rect 60747 8875 60789 8884
rect 60556 8128 60692 8168
rect 60404 7960 60500 8000
rect 60555 8000 60597 8009
rect 60555 7960 60556 8000
rect 60596 7960 60597 8000
rect 60364 7951 60404 7960
rect 60555 7951 60597 7960
rect 60652 8000 60692 8128
rect 60556 7866 60596 7951
rect 59788 7708 59884 7748
rect 59924 7708 60212 7748
rect 59788 7244 59828 7708
rect 59884 7699 59924 7708
rect 59788 7195 59828 7204
rect 59884 7328 59924 7337
rect 59884 7169 59924 7288
rect 59980 7244 60020 7253
rect 59692 7111 59732 7120
rect 59883 7160 59925 7169
rect 59883 7120 59884 7160
rect 59924 7120 59925 7160
rect 59883 7111 59925 7120
rect 58827 6992 58869 7001
rect 58827 6952 58828 6992
rect 58868 6952 58869 6992
rect 58827 6943 58869 6952
rect 59980 6656 60020 7204
rect 60076 7160 60116 7169
rect 60076 7001 60116 7120
rect 60652 7085 60692 7960
rect 60748 8000 60788 8875
rect 60843 8084 60885 8093
rect 60843 8044 60844 8084
rect 60884 8044 60885 8084
rect 60843 8035 60885 8044
rect 60748 7951 60788 7960
rect 60844 8000 60884 8035
rect 60844 7949 60884 7960
rect 60651 7076 60693 7085
rect 60651 7036 60652 7076
rect 60692 7036 60693 7076
rect 60651 7027 60693 7036
rect 60075 6992 60117 7001
rect 60075 6952 60076 6992
rect 60116 6952 60117 6992
rect 60075 6943 60117 6952
rect 59980 6607 60020 6616
rect 58347 6488 58389 6497
rect 58347 6448 58348 6488
rect 58388 6448 58389 6488
rect 58347 6439 58389 6448
rect 59788 6488 59828 6497
rect 58348 5825 58388 6439
rect 58347 5816 58389 5825
rect 58347 5776 58348 5816
rect 58388 5776 58389 5816
rect 58347 5767 58389 5776
rect 58100 5692 58196 5732
rect 59403 5732 59445 5741
rect 59403 5692 59404 5732
rect 59444 5692 59445 5732
rect 57964 5648 58004 5659
rect 57964 5573 58004 5608
rect 57963 5564 58005 5573
rect 57868 5524 57964 5564
rect 58004 5524 58005 5564
rect 57772 4976 57812 4985
rect 57580 4936 57772 4976
rect 57772 4927 57812 4936
rect 57044 4264 57140 4304
rect 57388 4768 57524 4808
rect 57771 4808 57813 4817
rect 57771 4768 57772 4808
rect 57812 4768 57813 4808
rect 56523 4220 56565 4229
rect 56523 4180 56524 4220
rect 56564 4180 56565 4220
rect 56523 4171 56565 4180
rect 56428 4087 56468 4096
rect 56524 4136 56564 4171
rect 5068 3415 5108 3424
rect 55083 3464 55125 3473
rect 55083 3424 55084 3464
rect 55124 3424 55125 3464
rect 55083 3415 55125 3424
rect 56044 3464 56084 3473
rect 843 3380 885 3389
rect 843 3340 844 3380
rect 884 3340 885 3380
rect 843 3331 885 3340
rect 2475 3380 2517 3389
rect 2475 3340 2476 3380
rect 2516 3340 2517 3380
rect 2475 3331 2517 3340
rect 844 3246 884 3331
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 56044 2801 56084 3424
rect 56043 2792 56085 2801
rect 56043 2752 56044 2792
rect 56084 2752 56085 2792
rect 56043 2743 56085 2752
rect 844 2708 884 2717
rect 556 2668 844 2708
rect 844 2659 884 2668
rect 56332 2624 56372 4087
rect 56524 4085 56564 4096
rect 56715 4136 56757 4145
rect 56715 4096 56716 4136
rect 56756 4096 56757 4136
rect 56715 4087 56757 4096
rect 56716 4002 56756 4087
rect 56427 3968 56469 3977
rect 56620 3968 56660 3977
rect 56427 3928 56428 3968
rect 56468 3928 56469 3968
rect 56427 3919 56469 3928
rect 56524 3928 56620 3968
rect 56428 3464 56468 3919
rect 56428 3415 56468 3424
rect 56524 2900 56564 3928
rect 56620 3919 56660 3928
rect 56428 2860 56564 2900
rect 57004 2876 57044 4264
rect 57388 4229 57428 4768
rect 57771 4759 57813 4768
rect 57387 4220 57429 4229
rect 57387 4180 57388 4220
rect 57428 4180 57429 4220
rect 57387 4171 57429 4180
rect 57099 4136 57141 4145
rect 57099 4096 57100 4136
rect 57140 4096 57141 4136
rect 57099 4087 57141 4096
rect 57291 4136 57333 4145
rect 57291 4096 57292 4136
rect 57332 4096 57333 4136
rect 57291 4087 57333 4096
rect 57388 4136 57428 4171
rect 56428 2708 56468 2860
rect 56620 2836 57044 2876
rect 56523 2792 56565 2801
rect 56523 2752 56524 2792
rect 56564 2752 56565 2792
rect 56523 2743 56565 2752
rect 56428 2659 56468 2668
rect 56524 2658 56564 2743
rect 56620 2708 56660 2836
rect 57100 2801 57140 4087
rect 57292 4002 57332 4087
rect 57388 4086 57428 4096
rect 57675 4136 57717 4145
rect 57675 4096 57676 4136
rect 57716 4096 57717 4136
rect 57675 4087 57717 4096
rect 57772 4136 57812 4759
rect 57772 4087 57812 4096
rect 57868 4136 57908 5524
rect 57963 5515 58005 5524
rect 58060 4985 58100 5692
rect 59403 5683 59445 5692
rect 59404 5648 59444 5683
rect 59404 5597 59444 5608
rect 59788 5489 59828 6448
rect 59884 6488 59924 6497
rect 59884 5993 59924 6448
rect 60076 6488 60116 6943
rect 60652 6488 60692 7027
rect 60940 6992 60980 10900
rect 61131 10436 61173 10445
rect 61228 10436 61268 11824
rect 61420 11780 61460 14344
rect 61516 13889 61556 14454
rect 61708 14225 61748 17032
rect 61900 17032 61985 17072
rect 62284 17032 62385 17072
rect 62745 17072 62785 17472
rect 62855 17072 62895 17472
rect 62955 17156 62997 17165
rect 62955 17116 62956 17156
rect 62996 17116 62997 17156
rect 62955 17107 62997 17116
rect 62745 17032 62804 17072
rect 62855 17032 62900 17072
rect 61900 15737 61940 17032
rect 62284 16157 62324 17032
rect 62764 16913 62804 17032
rect 62763 16904 62805 16913
rect 62763 16864 62764 16904
rect 62804 16864 62805 16904
rect 62763 16855 62805 16864
rect 62571 16568 62613 16577
rect 62571 16528 62572 16568
rect 62612 16528 62613 16568
rect 62571 16519 62613 16528
rect 62380 16232 62420 16241
rect 62283 16148 62325 16157
rect 62283 16108 62284 16148
rect 62324 16108 62325 16148
rect 62283 16099 62325 16108
rect 61995 16064 62037 16073
rect 61995 16024 61996 16064
rect 62036 16024 62037 16064
rect 61995 16015 62037 16024
rect 61899 15728 61941 15737
rect 61899 15688 61900 15728
rect 61940 15688 61941 15728
rect 61899 15679 61941 15688
rect 61996 15581 62036 16015
rect 61804 15560 61844 15569
rect 61804 14897 61844 15520
rect 61900 15560 61940 15570
rect 61996 15532 62036 15541
rect 62092 15560 62132 15569
rect 61900 15485 61940 15520
rect 61899 15476 61941 15485
rect 61899 15436 61900 15476
rect 61940 15465 61941 15476
rect 61940 15436 62036 15465
rect 61899 15427 62036 15436
rect 61900 15425 62036 15427
rect 61899 15308 61941 15317
rect 61899 15268 61900 15308
rect 61940 15268 61941 15308
rect 61899 15259 61941 15268
rect 61803 14888 61845 14897
rect 61803 14848 61804 14888
rect 61844 14848 61845 14888
rect 61803 14839 61845 14848
rect 61900 14804 61940 15259
rect 61900 14755 61940 14764
rect 61996 14561 62036 15425
rect 62092 14729 62132 15520
rect 62283 15476 62325 15485
rect 62283 15436 62284 15476
rect 62324 15436 62325 15476
rect 62283 15427 62325 15436
rect 62284 15342 62324 15427
rect 62380 14888 62420 16192
rect 62475 15308 62517 15317
rect 62475 15268 62476 15308
rect 62516 15268 62517 15308
rect 62475 15259 62517 15268
rect 62476 15174 62516 15259
rect 62572 15056 62612 16519
rect 62284 14848 62420 14888
rect 62476 15016 62612 15056
rect 62091 14720 62133 14729
rect 62091 14680 62092 14720
rect 62132 14680 62133 14720
rect 62091 14671 62133 14680
rect 61995 14552 62037 14561
rect 61995 14512 61996 14552
rect 62036 14512 62037 14552
rect 61995 14503 62037 14512
rect 62092 14552 62132 14671
rect 61707 14216 61749 14225
rect 61707 14176 61708 14216
rect 61748 14176 61749 14216
rect 61707 14167 61749 14176
rect 62092 14141 62132 14512
rect 62091 14132 62133 14141
rect 62091 14092 62092 14132
rect 62132 14092 62133 14132
rect 62091 14083 62133 14092
rect 62284 14057 62324 14848
rect 62380 14720 62420 14729
rect 62380 14561 62420 14680
rect 62476 14720 62516 15016
rect 62860 14981 62900 17032
rect 62859 14972 62901 14981
rect 62859 14932 62860 14972
rect 62900 14932 62901 14972
rect 62859 14923 62901 14932
rect 62476 14671 62516 14680
rect 62572 14720 62612 14729
rect 62379 14552 62421 14561
rect 62379 14512 62380 14552
rect 62420 14512 62421 14552
rect 62379 14503 62421 14512
rect 62283 14048 62325 14057
rect 62283 14008 62284 14048
rect 62324 14008 62325 14048
rect 62283 13999 62325 14008
rect 62380 13973 62420 14503
rect 62572 14216 62612 14680
rect 62668 14636 62708 14645
rect 62860 14636 62900 14645
rect 62708 14596 62860 14636
rect 62668 14587 62708 14596
rect 62860 14587 62900 14596
rect 62956 14468 62996 17107
rect 63145 17072 63185 17472
rect 63255 17072 63295 17472
rect 63545 17072 63585 17472
rect 63655 17072 63695 17472
rect 63819 17240 63861 17249
rect 63819 17200 63820 17240
rect 63860 17200 63861 17240
rect 63819 17191 63861 17200
rect 63145 17032 63188 17072
rect 63148 15989 63188 17032
rect 63244 17032 63295 17072
rect 63532 17032 63585 17072
rect 63628 17032 63695 17072
rect 63244 16493 63284 17032
rect 63243 16484 63285 16493
rect 63243 16444 63244 16484
rect 63284 16444 63285 16484
rect 63243 16435 63285 16444
rect 63532 16232 63572 17032
rect 63628 16829 63668 17032
rect 63627 16820 63669 16829
rect 63627 16780 63628 16820
rect 63668 16780 63669 16820
rect 63627 16771 63669 16780
rect 63820 16400 63860 17191
rect 63945 17072 63985 17472
rect 63916 17032 63985 17072
rect 64055 17072 64095 17472
rect 64345 17249 64385 17472
rect 64455 17333 64495 17472
rect 64454 17324 64496 17333
rect 64454 17284 64455 17324
rect 64495 17284 64496 17324
rect 64454 17275 64496 17284
rect 64344 17240 64386 17249
rect 64344 17200 64345 17240
rect 64385 17200 64386 17240
rect 64344 17191 64386 17200
rect 64745 17072 64785 17472
rect 64855 17300 64895 17472
rect 64855 17260 64916 17300
rect 64055 17032 64148 17072
rect 63916 16745 63956 17032
rect 63915 16736 63957 16745
rect 63915 16696 63916 16736
rect 63956 16696 63957 16736
rect 63915 16687 63957 16696
rect 63915 16484 63957 16493
rect 63915 16444 63916 16484
rect 63956 16444 63957 16484
rect 63915 16435 63957 16444
rect 63724 16360 63860 16400
rect 63532 16192 63668 16232
rect 63435 16148 63477 16157
rect 63435 16108 63436 16148
rect 63476 16108 63477 16148
rect 63435 16099 63477 16108
rect 63147 15980 63189 15989
rect 63147 15940 63148 15980
rect 63188 15940 63189 15980
rect 63147 15931 63189 15940
rect 63436 15308 63476 16099
rect 63531 16064 63573 16073
rect 63531 16024 63532 16064
rect 63572 16024 63573 16064
rect 63531 16015 63573 16024
rect 63532 15930 63572 16015
rect 63436 15268 63572 15308
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 63243 14972 63285 14981
rect 63243 14932 63244 14972
rect 63284 14932 63285 14972
rect 63243 14923 63285 14932
rect 63244 14720 63284 14923
rect 63244 14477 63284 14680
rect 63532 14636 63572 15268
rect 63436 14596 63572 14636
rect 62476 14176 62612 14216
rect 62764 14428 62996 14468
rect 63243 14468 63285 14477
rect 63436 14468 63476 14596
rect 63243 14428 63244 14468
rect 63284 14428 63285 14468
rect 62379 13964 62421 13973
rect 62379 13924 62380 13964
rect 62420 13924 62421 13964
rect 62379 13915 62421 13924
rect 61515 13880 61557 13889
rect 61515 13840 61516 13880
rect 61556 13840 61557 13880
rect 61515 13831 61557 13840
rect 61803 13796 61845 13805
rect 61803 13756 61804 13796
rect 61844 13756 61845 13796
rect 61803 13747 61845 13756
rect 62379 13796 62421 13805
rect 62379 13756 62380 13796
rect 62420 13756 62421 13796
rect 62379 13747 62421 13756
rect 61515 13460 61557 13469
rect 61515 13420 61516 13460
rect 61556 13420 61557 13460
rect 61515 13411 61557 13420
rect 61516 13208 61556 13411
rect 61611 13292 61653 13301
rect 61611 13252 61612 13292
rect 61652 13252 61653 13292
rect 61611 13243 61653 13252
rect 61516 13159 61556 13168
rect 61612 13124 61652 13243
rect 61707 13208 61749 13217
rect 61707 13168 61708 13208
rect 61748 13168 61749 13208
rect 61707 13159 61749 13168
rect 61804 13208 61844 13747
rect 62380 13662 62420 13747
rect 61995 13460 62037 13469
rect 62476 13460 62516 14176
rect 62572 14048 62612 14057
rect 62572 13805 62612 14008
rect 62668 13889 62708 13974
rect 62667 13880 62709 13889
rect 62667 13840 62668 13880
rect 62708 13840 62709 13880
rect 62667 13831 62709 13840
rect 62571 13796 62613 13805
rect 62571 13756 62572 13796
rect 62612 13756 62613 13796
rect 62571 13747 62613 13756
rect 62667 13712 62709 13721
rect 62667 13672 62668 13712
rect 62708 13672 62709 13712
rect 62667 13663 62709 13672
rect 62572 13460 62612 13469
rect 61995 13420 61996 13460
rect 62036 13420 62037 13460
rect 61995 13411 62037 13420
rect 62284 13420 62572 13460
rect 61804 13159 61844 13168
rect 61996 13208 62036 13411
rect 62187 13376 62229 13385
rect 62187 13336 62188 13376
rect 62228 13336 62229 13376
rect 62187 13327 62229 13336
rect 62091 13292 62133 13301
rect 62091 13252 62092 13292
rect 62132 13252 62133 13292
rect 62091 13243 62133 13252
rect 61612 13075 61652 13084
rect 61515 13040 61557 13049
rect 61515 13000 61516 13040
rect 61556 13000 61557 13040
rect 61515 12991 61557 13000
rect 61516 12536 61556 12991
rect 61516 12487 61556 12496
rect 61708 11957 61748 13159
rect 61899 12620 61941 12629
rect 61899 12580 61900 12620
rect 61940 12580 61941 12620
rect 61899 12571 61941 12580
rect 61707 11948 61749 11957
rect 61707 11908 61708 11948
rect 61748 11908 61749 11948
rect 61707 11899 61749 11908
rect 61420 11705 61460 11740
rect 61707 11780 61749 11789
rect 61707 11740 61708 11780
rect 61748 11740 61749 11780
rect 61707 11731 61749 11740
rect 61419 11696 61461 11705
rect 61419 11656 61420 11696
rect 61460 11656 61461 11696
rect 61419 11647 61461 11656
rect 61420 11616 61460 11647
rect 61323 11192 61365 11201
rect 61323 11152 61324 11192
rect 61364 11152 61365 11192
rect 61323 11143 61365 11152
rect 61324 11058 61364 11143
rect 61708 11024 61748 11731
rect 61803 11612 61845 11621
rect 61803 11572 61804 11612
rect 61844 11572 61845 11612
rect 61803 11563 61845 11572
rect 61708 10975 61748 10984
rect 61804 10982 61844 11563
rect 61900 11117 61940 12571
rect 61996 11789 62036 13168
rect 62092 13158 62132 13243
rect 62188 13242 62228 13327
rect 62284 13292 62324 13420
rect 62572 13411 62612 13420
rect 62284 13243 62324 13252
rect 62380 13208 62420 13217
rect 62091 13040 62133 13049
rect 62091 13000 62092 13040
rect 62132 13000 62133 13040
rect 62091 12991 62133 13000
rect 62092 12629 62132 12991
rect 62380 12881 62420 13168
rect 62668 13049 62708 13663
rect 62667 13040 62709 13049
rect 62667 13000 62668 13040
rect 62708 13000 62709 13040
rect 62667 12991 62709 13000
rect 62379 12872 62421 12881
rect 62379 12832 62380 12872
rect 62420 12832 62421 12872
rect 62379 12823 62421 12832
rect 62091 12620 62133 12629
rect 62091 12580 62092 12620
rect 62132 12580 62133 12620
rect 62091 12571 62133 12580
rect 62764 12452 62804 14428
rect 63243 14419 63285 14428
rect 63340 14428 63476 14468
rect 63531 14468 63573 14477
rect 63531 14428 63532 14468
rect 63572 14428 63573 14468
rect 63340 14069 63380 14428
rect 63531 14419 63573 14428
rect 63436 14141 63476 14172
rect 63435 14132 63477 14141
rect 63435 14092 63436 14132
rect 63476 14092 63477 14132
rect 63435 14083 63477 14092
rect 63148 14048 63188 14057
rect 62860 14008 63148 14048
rect 62860 13208 62900 14008
rect 63148 13999 63188 14008
rect 63244 14048 63284 14057
rect 63340 14020 63380 14029
rect 63436 14048 63476 14083
rect 63244 13889 63284 14008
rect 63436 13973 63476 14008
rect 63435 13964 63477 13973
rect 63435 13924 63436 13964
rect 63476 13924 63477 13964
rect 63435 13915 63477 13924
rect 63243 13880 63285 13889
rect 63243 13840 63244 13880
rect 63284 13840 63285 13880
rect 63243 13831 63285 13840
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 62860 13159 62900 13168
rect 62955 13208 62997 13217
rect 62955 13168 62956 13208
rect 62996 13168 62997 13208
rect 62955 13159 62997 13168
rect 62956 13074 62996 13159
rect 63052 12982 63092 12991
rect 62956 12942 63052 12980
rect 63532 12965 63572 14419
rect 63628 13133 63668 16192
rect 63724 14309 63764 16360
rect 63916 16350 63956 16435
rect 63820 16232 63860 16243
rect 63820 16157 63860 16192
rect 63819 16148 63861 16157
rect 63819 16108 63820 16148
rect 63860 16108 63861 16148
rect 63819 16099 63861 16108
rect 64108 15737 64148 17032
rect 64204 17032 64785 17072
rect 64107 15728 64149 15737
rect 64107 15688 64108 15728
rect 64148 15688 64149 15728
rect 64107 15679 64149 15688
rect 64108 14720 64148 14729
rect 63723 14300 63765 14309
rect 63723 14260 63724 14300
rect 63764 14260 63765 14300
rect 63723 14251 63765 14260
rect 64108 14057 64148 14680
rect 64107 14048 64149 14057
rect 64107 14008 64108 14048
rect 64148 14008 64149 14048
rect 64107 13999 64149 14008
rect 63819 13964 63861 13973
rect 63819 13924 63820 13964
rect 63860 13924 63861 13964
rect 63819 13915 63861 13924
rect 63820 13385 63860 13915
rect 63819 13376 63861 13385
rect 63819 13336 63820 13376
rect 63860 13336 63861 13376
rect 63819 13327 63861 13336
rect 63820 13217 63860 13327
rect 63819 13208 63861 13217
rect 63819 13168 63820 13208
rect 63860 13168 63861 13208
rect 63819 13159 63861 13168
rect 63627 13124 63669 13133
rect 63627 13084 63628 13124
rect 63668 13084 63669 13124
rect 63627 13075 63669 13084
rect 62956 12940 63092 12942
rect 62956 12881 62996 12940
rect 63052 12933 63092 12940
rect 63531 12956 63573 12965
rect 63531 12916 63532 12956
rect 63572 12916 63573 12956
rect 63531 12907 63573 12916
rect 62955 12872 62997 12881
rect 62955 12832 62956 12872
rect 62996 12832 62997 12872
rect 62955 12823 62997 12832
rect 62956 12704 62996 12823
rect 63723 12788 63765 12797
rect 63723 12748 63724 12788
rect 63764 12748 63765 12788
rect 63723 12739 63765 12748
rect 62956 12655 62996 12664
rect 63724 12704 63764 12739
rect 63724 12653 63764 12664
rect 62092 12412 62804 12452
rect 62860 12536 62900 12545
rect 61995 11780 62037 11789
rect 61995 11740 61996 11780
rect 62036 11740 62037 11780
rect 61995 11731 62037 11740
rect 62092 11360 62132 12412
rect 62668 12284 62708 12293
rect 62860 12284 62900 12496
rect 63627 12536 63669 12545
rect 63627 12496 63628 12536
rect 63668 12496 63669 12536
rect 63627 12487 63669 12496
rect 62708 12244 62900 12284
rect 62379 11864 62421 11873
rect 62379 11824 62380 11864
rect 62420 11824 62421 11864
rect 62379 11815 62421 11824
rect 62187 11780 62229 11789
rect 62187 11740 62188 11780
rect 62228 11740 62229 11780
rect 62187 11731 62229 11740
rect 62188 11696 62228 11731
rect 62188 11645 62228 11656
rect 62380 11696 62420 11815
rect 62380 11647 62420 11656
rect 62476 11696 62516 11705
rect 62668 11696 62708 12244
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 63148 11705 63188 11790
rect 62516 11656 62708 11696
rect 63147 11696 63189 11705
rect 63147 11656 63148 11696
rect 63188 11656 63189 11696
rect 62476 11647 62516 11656
rect 63147 11647 63189 11656
rect 62283 11612 62325 11621
rect 62283 11572 62284 11612
rect 62324 11572 62325 11612
rect 62283 11563 62325 11572
rect 62764 11612 62804 11621
rect 63339 11612 63381 11621
rect 62804 11572 62996 11612
rect 62764 11563 62804 11572
rect 62284 11478 62324 11563
rect 62092 11320 62228 11360
rect 62091 11192 62133 11201
rect 62091 11152 62092 11192
rect 62132 11152 62133 11192
rect 62091 11143 62133 11152
rect 61899 11108 61941 11117
rect 61899 11068 61900 11108
rect 61940 11068 61941 11108
rect 61899 11059 61941 11068
rect 62092 11024 62132 11143
rect 61804 10933 61844 10942
rect 61900 10865 61940 10950
rect 62092 10949 62132 10984
rect 61996 10940 62036 10949
rect 61899 10856 61941 10865
rect 61899 10816 61900 10856
rect 61940 10816 61941 10856
rect 61899 10807 61941 10816
rect 61996 10781 62036 10900
rect 62091 10940 62133 10949
rect 62091 10900 62092 10940
rect 62132 10900 62133 10940
rect 62091 10891 62133 10900
rect 61995 10772 62037 10781
rect 61995 10732 61996 10772
rect 62036 10732 62037 10772
rect 61995 10723 62037 10732
rect 61131 10396 61132 10436
rect 61172 10396 61268 10436
rect 61131 10387 61173 10396
rect 61036 10184 61076 10193
rect 61036 9176 61076 10144
rect 61132 9437 61172 10387
rect 61899 10184 61941 10193
rect 61899 10144 61900 10184
rect 61940 10144 61941 10184
rect 61899 10135 61941 10144
rect 61900 10050 61940 10135
rect 61131 9428 61173 9437
rect 61131 9388 61132 9428
rect 61172 9388 61173 9428
rect 61131 9379 61173 9388
rect 61419 9428 61461 9437
rect 61419 9388 61420 9428
rect 61460 9388 61461 9428
rect 61419 9379 61461 9388
rect 61132 9294 61172 9379
rect 61324 9260 61364 9269
rect 61324 9176 61364 9220
rect 61036 9136 61364 9176
rect 61036 8672 61076 8681
rect 61036 7169 61076 8632
rect 61324 8009 61364 9136
rect 61323 8000 61365 8009
rect 61323 7960 61324 8000
rect 61364 7960 61365 8000
rect 61323 7951 61365 7960
rect 61035 7160 61077 7169
rect 61035 7120 61036 7160
rect 61076 7120 61077 7160
rect 61035 7111 61077 7120
rect 60940 6952 61076 6992
rect 60747 6572 60789 6581
rect 60747 6532 60748 6572
rect 60788 6532 60789 6572
rect 60747 6523 60789 6532
rect 59883 5984 59925 5993
rect 59883 5944 59884 5984
rect 59924 5944 59925 5984
rect 59883 5935 59925 5944
rect 60076 5909 60116 6448
rect 60460 6448 60652 6488
rect 60075 5900 60117 5909
rect 60075 5860 60076 5900
rect 60116 5860 60117 5900
rect 60075 5851 60117 5860
rect 60268 5648 60308 5657
rect 60076 5608 60268 5648
rect 59883 5564 59925 5573
rect 59883 5524 59884 5564
rect 59924 5524 59925 5564
rect 59883 5515 59925 5524
rect 58251 5480 58293 5489
rect 58251 5440 58252 5480
rect 58292 5440 58293 5480
rect 58251 5431 58293 5440
rect 59787 5480 59829 5489
rect 59787 5440 59788 5480
rect 59828 5440 59829 5480
rect 59787 5431 59829 5440
rect 58252 5346 58292 5431
rect 59788 4985 59828 5431
rect 58059 4976 58101 4985
rect 58059 4936 58060 4976
rect 58100 4936 58101 4976
rect 58059 4927 58101 4936
rect 58636 4976 58676 4985
rect 57963 4220 58005 4229
rect 57963 4180 57964 4220
rect 58004 4180 58005 4220
rect 57963 4171 58005 4180
rect 57868 4087 57908 4096
rect 57964 4136 58004 4171
rect 57676 4002 57716 4087
rect 57964 4085 58004 4096
rect 57484 3910 57524 3919
rect 57291 3464 57333 3473
rect 57291 3424 57292 3464
rect 57332 3424 57333 3464
rect 57291 3415 57333 3424
rect 57292 3330 57332 3415
rect 57484 2885 57524 3870
rect 58636 3473 58676 4936
rect 59787 4976 59829 4985
rect 59787 4936 59788 4976
rect 59828 4936 59829 4976
rect 59787 4927 59829 4936
rect 59788 4808 59828 4817
rect 59884 4808 59924 5515
rect 59828 4768 59924 4808
rect 59788 4759 59828 4768
rect 60076 3977 60116 5608
rect 60268 5599 60308 5608
rect 60460 5144 60500 6448
rect 60652 6439 60692 6448
rect 60748 6488 60788 6523
rect 60748 6437 60788 6448
rect 60844 6488 60884 6497
rect 60844 5816 60884 6448
rect 60939 6488 60981 6497
rect 60939 6448 60940 6488
rect 60980 6448 60981 6488
rect 60939 6439 60981 6448
rect 60940 6354 60980 6439
rect 60940 5816 60980 5825
rect 60844 5776 60940 5816
rect 60364 5104 60500 5144
rect 60652 5564 60692 5573
rect 60364 4724 60404 5104
rect 60555 5060 60597 5069
rect 60555 5020 60556 5060
rect 60596 5020 60597 5060
rect 60555 5011 60597 5020
rect 60459 4976 60501 4985
rect 60459 4936 60460 4976
rect 60500 4936 60501 4976
rect 60459 4927 60501 4936
rect 60460 4842 60500 4927
rect 60556 4926 60596 5011
rect 60652 4724 60692 5524
rect 60747 5060 60789 5069
rect 60747 5020 60748 5060
rect 60788 5020 60789 5060
rect 60747 5011 60789 5020
rect 60748 4976 60788 5011
rect 60748 4925 60788 4936
rect 60844 4892 60884 5776
rect 60940 5767 60980 5776
rect 61036 5489 61076 6952
rect 61131 6488 61173 6497
rect 61131 6448 61132 6488
rect 61172 6448 61173 6488
rect 61420 6488 61460 9379
rect 62188 8933 62228 11320
rect 62764 11201 62804 11287
rect 62763 11196 62805 11201
rect 62763 11152 62764 11196
rect 62804 11152 62805 11196
rect 62763 11143 62805 11152
rect 62956 11192 62996 11572
rect 63244 11572 63340 11612
rect 63380 11572 63381 11612
rect 63244 11528 63284 11572
rect 63339 11563 63381 11572
rect 63340 11544 63380 11563
rect 62956 11143 62996 11152
rect 63148 11488 63284 11528
rect 62475 11108 62517 11117
rect 62475 11068 62476 11108
rect 62516 11068 62517 11108
rect 62475 11059 62517 11068
rect 62283 10772 62325 10781
rect 62283 10732 62284 10772
rect 62324 10732 62325 10772
rect 62283 10723 62325 10732
rect 62284 10638 62324 10723
rect 62187 8924 62229 8933
rect 62187 8884 62188 8924
rect 62228 8884 62229 8924
rect 62187 8875 62229 8884
rect 62188 8790 62228 8875
rect 62091 8252 62133 8261
rect 62091 8212 62092 8252
rect 62132 8212 62133 8252
rect 62091 8203 62133 8212
rect 61803 8084 61845 8093
rect 61803 8044 61804 8084
rect 61844 8044 61845 8084
rect 61803 8035 61845 8044
rect 61612 7160 61652 7171
rect 61612 7085 61652 7120
rect 61708 7160 61748 7169
rect 61611 7076 61653 7085
rect 61611 7036 61612 7076
rect 61652 7036 61653 7076
rect 61611 7027 61653 7036
rect 61516 6992 61556 7001
rect 61516 6656 61556 6952
rect 61708 6749 61748 7120
rect 61804 7160 61844 8035
rect 62092 7328 62132 8203
rect 62187 8084 62229 8093
rect 62187 8044 62188 8084
rect 62228 8044 62229 8084
rect 62187 8035 62229 8044
rect 62188 7950 62228 8035
rect 62283 7748 62325 7757
rect 62283 7708 62284 7748
rect 62324 7708 62325 7748
rect 62283 7699 62325 7708
rect 62092 7288 62228 7328
rect 61707 6740 61749 6749
rect 61707 6700 61708 6740
rect 61748 6700 61749 6740
rect 61707 6691 61749 6700
rect 61516 6616 61652 6656
rect 61516 6488 61556 6497
rect 61420 6448 61516 6488
rect 61131 6439 61173 6448
rect 61516 6439 61556 6448
rect 61132 6354 61172 6439
rect 61612 6320 61652 6616
rect 61228 6280 61652 6320
rect 61131 5900 61173 5909
rect 61131 5860 61132 5900
rect 61172 5860 61173 5900
rect 61131 5851 61173 5860
rect 61035 5480 61077 5489
rect 61035 5440 61036 5480
rect 61076 5440 61077 5480
rect 61035 5431 61077 5440
rect 61132 4976 61172 5851
rect 61228 5648 61268 6280
rect 61804 6068 61844 7120
rect 62092 7160 62132 7169
rect 62092 6749 62132 7120
rect 62188 7160 62228 7288
rect 62091 6740 62133 6749
rect 62091 6700 62092 6740
rect 62132 6700 62133 6740
rect 62091 6691 62133 6700
rect 62188 6581 62228 7120
rect 62187 6572 62229 6581
rect 62187 6532 62188 6572
rect 62228 6532 62229 6572
rect 62187 6523 62229 6532
rect 61899 6488 61941 6497
rect 61899 6448 61900 6488
rect 61940 6448 61941 6488
rect 61899 6439 61941 6448
rect 61228 5599 61268 5608
rect 61324 6028 61844 6068
rect 61324 5648 61364 6028
rect 61324 5599 61364 5608
rect 61323 5480 61365 5489
rect 61323 5440 61324 5480
rect 61364 5440 61365 5480
rect 61323 5431 61365 5440
rect 61172 4936 61268 4976
rect 61132 4927 61172 4936
rect 60844 4843 60884 4852
rect 61036 4892 61076 4901
rect 60940 4808 60980 4817
rect 60940 4724 60980 4768
rect 60364 4684 60500 4724
rect 60652 4684 60980 4724
rect 60268 4136 60308 4145
rect 60171 4052 60213 4061
rect 60171 4012 60172 4052
rect 60212 4012 60213 4052
rect 60171 4003 60213 4012
rect 60075 3968 60117 3977
rect 60075 3928 60076 3968
rect 60116 3928 60117 3968
rect 60075 3919 60117 3928
rect 60172 3918 60212 4003
rect 60268 3800 60308 4096
rect 60363 4136 60405 4145
rect 60363 4096 60364 4136
rect 60404 4096 60405 4136
rect 60363 4087 60405 4096
rect 60460 4136 60500 4684
rect 61036 4397 61076 4852
rect 61035 4388 61077 4397
rect 61035 4348 61036 4388
rect 61076 4348 61077 4388
rect 61035 4339 61077 4348
rect 60747 4304 60789 4313
rect 60747 4264 60748 4304
rect 60788 4264 60789 4304
rect 60747 4255 60789 4264
rect 60500 4096 60596 4136
rect 60460 4087 60500 4096
rect 60364 4002 60404 4087
rect 59788 3760 60308 3800
rect 60556 3800 60596 4096
rect 60651 4052 60693 4061
rect 60651 4012 60652 4052
rect 60692 4012 60693 4052
rect 60651 4003 60693 4012
rect 60652 3918 60692 4003
rect 60556 3760 60692 3800
rect 58635 3464 58677 3473
rect 58635 3424 58636 3464
rect 58676 3424 58677 3464
rect 58635 3415 58677 3424
rect 59788 3296 59828 3760
rect 60268 3636 60308 3645
rect 60171 3548 60213 3557
rect 60171 3508 60172 3548
rect 60212 3508 60213 3548
rect 60171 3499 60213 3508
rect 60075 3464 60117 3473
rect 60075 3424 60076 3464
rect 60116 3424 60117 3464
rect 60075 3415 60117 3424
rect 60172 3464 60212 3499
rect 60076 3330 60116 3415
rect 60172 3413 60212 3424
rect 59212 3256 59788 3296
rect 58444 3212 58484 3221
rect 57483 2876 57525 2885
rect 57483 2836 57484 2876
rect 57524 2836 57525 2876
rect 57483 2827 57525 2836
rect 57867 2876 57909 2885
rect 57867 2836 57868 2876
rect 57908 2836 57909 2876
rect 57867 2827 57909 2836
rect 57099 2792 57141 2801
rect 57099 2752 57100 2792
rect 57140 2752 57141 2792
rect 57099 2743 57141 2752
rect 57868 2742 57908 2827
rect 56620 2659 56660 2668
rect 56332 2549 56372 2584
rect 56715 2624 56757 2633
rect 56715 2584 56716 2624
rect 56756 2584 56757 2624
rect 56715 2575 56757 2584
rect 57964 2624 58004 2633
rect 58444 2624 58484 3172
rect 58539 2792 58581 2801
rect 58539 2752 58540 2792
rect 58580 2752 58581 2792
rect 58539 2743 58581 2752
rect 58732 2792 58772 2801
rect 59116 2792 59156 2801
rect 58772 2752 59060 2792
rect 58732 2743 58772 2752
rect 58004 2584 58444 2624
rect 57964 2575 58004 2584
rect 58444 2575 58484 2584
rect 58540 2624 58580 2743
rect 59020 2708 59060 2752
rect 59020 2659 59060 2668
rect 58540 2575 58580 2584
rect 58731 2624 58773 2633
rect 58731 2584 58732 2624
rect 58772 2584 58773 2624
rect 58731 2575 58773 2584
rect 58923 2624 58965 2633
rect 58923 2584 58924 2624
rect 58964 2584 58965 2624
rect 58923 2575 58965 2584
rect 56331 2540 56373 2549
rect 56331 2500 56332 2540
rect 56372 2500 56373 2540
rect 56331 2491 56373 2500
rect 652 2456 692 2465
rect 56332 2460 56372 2491
rect 56716 2490 56756 2575
rect 58732 2490 58772 2575
rect 58924 2490 58964 2575
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 59116 2045 59156 2752
rect 59212 2708 59252 3256
rect 59788 3247 59828 3256
rect 60172 2876 60212 2885
rect 60268 2876 60308 3596
rect 60555 3464 60597 3473
rect 60555 3424 60556 3464
rect 60596 3424 60597 3464
rect 60555 3415 60597 3424
rect 60652 3464 60692 3760
rect 60556 3330 60596 3415
rect 60652 2885 60692 3424
rect 60748 3464 60788 4255
rect 61036 4136 61076 4145
rect 61036 3977 61076 4096
rect 61035 3968 61077 3977
rect 61035 3928 61036 3968
rect 61076 3928 61077 3968
rect 61035 3919 61077 3928
rect 60843 3716 60885 3725
rect 60843 3676 60844 3716
rect 60884 3676 60885 3716
rect 60843 3667 60885 3676
rect 60844 3557 60884 3667
rect 60843 3548 60885 3557
rect 60843 3508 60844 3548
rect 60884 3508 60885 3548
rect 60843 3499 60885 3508
rect 60748 3415 60788 3424
rect 60844 3464 60884 3499
rect 60844 3414 60884 3424
rect 61036 2969 61076 3919
rect 61228 3464 61268 4936
rect 61324 4892 61364 5431
rect 61420 5422 61460 5431
rect 61420 5069 61460 5382
rect 61419 5060 61461 5069
rect 61419 5020 61420 5060
rect 61460 5020 61461 5060
rect 61419 5011 61461 5020
rect 61420 4892 61460 4901
rect 61324 4852 61420 4892
rect 61420 4649 61460 4852
rect 61419 4640 61461 4649
rect 61419 4600 61420 4640
rect 61460 4600 61461 4640
rect 61419 4591 61461 4600
rect 61419 4388 61461 4397
rect 61419 4348 61420 4388
rect 61460 4348 61461 4388
rect 61419 4339 61461 4348
rect 61420 3632 61460 4339
rect 61516 3725 61556 6028
rect 61611 5900 61653 5909
rect 61611 5860 61612 5900
rect 61652 5860 61653 5900
rect 61611 5851 61653 5860
rect 61612 5144 61652 5851
rect 61900 5825 61940 6439
rect 61899 5816 61941 5825
rect 61899 5776 61900 5816
rect 61940 5776 61941 5816
rect 61899 5767 61941 5776
rect 61612 5095 61652 5104
rect 61803 4892 61845 4901
rect 61803 4852 61804 4892
rect 61844 4852 61845 4892
rect 61803 4843 61845 4852
rect 61804 4758 61844 4843
rect 61612 4724 61652 4733
rect 61515 3716 61557 3725
rect 61515 3676 61516 3716
rect 61556 3676 61557 3716
rect 61515 3667 61557 3676
rect 61420 3583 61460 3592
rect 61612 3548 61652 4684
rect 61803 4640 61845 4649
rect 61803 4600 61804 4640
rect 61844 4600 61845 4640
rect 61803 4591 61845 4600
rect 61804 3632 61844 4591
rect 61804 3583 61844 3592
rect 61900 4136 61940 5767
rect 62284 5144 62324 7699
rect 62379 7160 62421 7169
rect 62379 7120 62380 7160
rect 62420 7120 62421 7160
rect 62379 7111 62421 7120
rect 62380 6497 62420 7111
rect 62379 6488 62421 6497
rect 62379 6448 62380 6488
rect 62420 6448 62421 6488
rect 62379 6439 62421 6448
rect 62380 6354 62420 6439
rect 62284 5095 62324 5104
rect 62188 4976 62228 4985
rect 62476 4976 62516 11059
rect 62571 11024 62613 11033
rect 62571 10984 62572 11024
rect 62612 10984 62613 11024
rect 62571 10975 62613 10984
rect 62668 11024 62708 11033
rect 62572 10890 62612 10975
rect 62668 10940 62708 10984
rect 63052 11024 63092 11033
rect 62668 10900 62900 10940
rect 62763 10352 62805 10361
rect 62763 10312 62764 10352
rect 62804 10312 62805 10352
rect 62763 10303 62805 10312
rect 62764 10109 62804 10303
rect 62763 10100 62805 10109
rect 62763 10060 62764 10100
rect 62804 10060 62805 10100
rect 62763 10051 62805 10060
rect 62860 10025 62900 10900
rect 63052 10781 63092 10984
rect 63148 11024 63188 11488
rect 63531 11192 63573 11201
rect 63148 10975 63188 10984
rect 63244 11152 63532 11192
rect 63572 11152 63573 11192
rect 63244 11024 63284 11152
rect 63531 11143 63573 11152
rect 63244 10975 63284 10984
rect 63435 11024 63477 11033
rect 63435 10984 63436 11024
rect 63476 10984 63477 11024
rect 63435 10975 63477 10984
rect 63532 11024 63572 11143
rect 63532 10975 63572 10984
rect 63628 11024 63668 12487
rect 63724 12284 63764 12293
rect 63724 11621 63764 12244
rect 63723 11612 63765 11621
rect 63723 11572 63724 11612
rect 63764 11572 63765 11612
rect 63723 11563 63765 11572
rect 63628 10975 63668 10984
rect 63724 11024 63764 11033
rect 63820 11024 63860 13159
rect 64204 12461 64244 17032
rect 64876 16241 64916 17260
rect 65145 17165 65185 17472
rect 65144 17156 65186 17165
rect 65144 17116 65145 17156
rect 65185 17116 65186 17156
rect 65144 17107 65186 17116
rect 65255 17072 65295 17472
rect 65545 17249 65585 17472
rect 65655 17333 65695 17472
rect 65654 17324 65696 17333
rect 65654 17284 65655 17324
rect 65695 17284 65696 17324
rect 65654 17275 65696 17284
rect 65544 17240 65586 17249
rect 65544 17200 65545 17240
rect 65585 17200 65586 17240
rect 65544 17191 65586 17200
rect 65945 17072 65985 17472
rect 66055 17333 66095 17472
rect 66054 17324 66096 17333
rect 66054 17284 66055 17324
rect 66095 17284 66096 17324
rect 66054 17275 66096 17284
rect 66345 17081 66385 17472
rect 66455 17165 66495 17472
rect 66745 17165 66785 17472
rect 66855 17249 66895 17472
rect 66854 17240 66896 17249
rect 66854 17200 66855 17240
rect 66895 17200 66896 17240
rect 66854 17191 66896 17200
rect 66454 17156 66496 17165
rect 66454 17116 66455 17156
rect 66495 17116 66496 17156
rect 66454 17107 66496 17116
rect 66744 17156 66786 17165
rect 66744 17116 66745 17156
rect 66785 17116 66786 17156
rect 66744 17107 66786 17116
rect 65255 17032 65300 17072
rect 64875 16232 64917 16241
rect 64875 16192 64876 16232
rect 64916 16192 64917 16232
rect 64875 16183 64917 16192
rect 64876 14645 64916 16183
rect 64971 15980 65013 15989
rect 64971 15940 64972 15980
rect 65012 15940 65013 15980
rect 64971 15931 65013 15940
rect 64875 14636 64917 14645
rect 64875 14596 64876 14636
rect 64916 14596 64917 14636
rect 64875 14587 64917 14596
rect 64779 14552 64821 14561
rect 64779 14512 64780 14552
rect 64820 14512 64821 14552
rect 64779 14503 64821 14512
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 64780 14216 64820 14503
rect 64588 14176 64820 14216
rect 64588 14132 64628 14176
rect 64588 14083 64628 14092
rect 64972 14048 65012 15931
rect 65067 15812 65109 15821
rect 65067 15772 65068 15812
rect 65108 15772 65109 15812
rect 65067 15763 65109 15772
rect 65068 15476 65108 15763
rect 65260 15476 65300 17032
rect 65932 17032 65985 17072
rect 66315 17072 66385 17081
rect 66315 17032 66316 17072
rect 66356 17032 66385 17072
rect 67145 17081 67185 17472
rect 67255 17333 67295 17472
rect 67254 17324 67296 17333
rect 67254 17284 67255 17324
rect 67295 17284 67296 17324
rect 67254 17275 67296 17284
rect 67371 17240 67413 17249
rect 67371 17200 67372 17240
rect 67412 17200 67413 17240
rect 67371 17191 67413 17200
rect 67145 17072 67221 17081
rect 67145 17032 67180 17072
rect 67220 17032 67221 17072
rect 65739 16568 65781 16577
rect 65739 16528 65740 16568
rect 65780 16528 65781 16568
rect 65739 16519 65781 16528
rect 65740 16484 65780 16519
rect 65740 16433 65780 16444
rect 65643 16400 65685 16409
rect 65643 16360 65644 16400
rect 65684 16360 65685 16400
rect 65643 16351 65685 16360
rect 65644 16232 65684 16351
rect 65548 16192 65644 16232
rect 65451 16148 65493 16157
rect 65451 16108 65452 16148
rect 65492 16108 65493 16148
rect 65451 16099 65493 16108
rect 65355 15560 65397 15569
rect 65355 15520 65356 15560
rect 65396 15520 65397 15560
rect 65355 15511 65397 15520
rect 65068 15427 65108 15436
rect 65164 15436 65300 15476
rect 65067 15308 65109 15317
rect 65067 15268 65068 15308
rect 65108 15268 65109 15308
rect 65067 15259 65109 15268
rect 65068 14645 65108 15259
rect 65164 15233 65204 15436
rect 65260 15308 65300 15317
rect 65356 15308 65396 15511
rect 65300 15268 65396 15308
rect 65260 15259 65300 15268
rect 65163 15224 65205 15233
rect 65163 15184 65164 15224
rect 65204 15184 65205 15224
rect 65163 15175 65205 15184
rect 65452 15140 65492 16099
rect 65548 15485 65588 16192
rect 65644 16183 65684 16192
rect 65643 15896 65685 15905
rect 65643 15856 65644 15896
rect 65684 15856 65685 15896
rect 65643 15847 65685 15856
rect 65547 15476 65589 15485
rect 65547 15436 65548 15476
rect 65588 15436 65589 15476
rect 65547 15427 65589 15436
rect 65260 15100 65492 15140
rect 65163 14972 65205 14981
rect 65163 14932 65164 14972
rect 65204 14932 65205 14972
rect 65163 14923 65205 14932
rect 65260 14972 65300 15100
rect 65260 14923 65300 14932
rect 65067 14636 65109 14645
rect 65067 14596 65068 14636
rect 65108 14596 65109 14636
rect 65067 14587 65109 14596
rect 65067 14384 65109 14393
rect 65067 14344 65068 14384
rect 65108 14344 65109 14384
rect 65067 14335 65109 14344
rect 64972 13999 65012 14008
rect 64875 13544 64917 13553
rect 64875 13504 64876 13544
rect 64916 13504 64917 13544
rect 64875 13495 64917 13504
rect 64779 12956 64821 12965
rect 64779 12916 64780 12956
rect 64820 12916 64821 12956
rect 64779 12907 64821 12916
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 64396 12536 64436 12545
rect 64203 12452 64245 12461
rect 64203 12412 64204 12452
rect 64244 12412 64245 12452
rect 64203 12403 64245 12412
rect 64396 11873 64436 12496
rect 64780 12536 64820 12907
rect 64780 12461 64820 12496
rect 64779 12452 64821 12461
rect 64779 12412 64780 12452
rect 64820 12412 64821 12452
rect 64779 12403 64821 12412
rect 64395 11864 64437 11873
rect 64395 11824 64396 11864
rect 64436 11824 64437 11864
rect 64395 11815 64437 11824
rect 64876 11705 64916 13495
rect 64012 11696 64052 11705
rect 64012 11033 64052 11656
rect 64875 11696 64917 11705
rect 64875 11656 64876 11696
rect 64916 11656 64917 11696
rect 64875 11647 64917 11656
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 64779 11192 64821 11201
rect 64779 11152 64780 11192
rect 64820 11152 64821 11192
rect 64779 11143 64821 11152
rect 64780 11058 64820 11143
rect 63764 10984 63860 11024
rect 64011 11024 64053 11033
rect 64011 10984 64012 11024
rect 64052 10984 64053 11024
rect 63724 10975 63764 10984
rect 64011 10975 64053 10984
rect 63436 10890 63476 10975
rect 63531 10856 63573 10865
rect 63531 10816 63532 10856
rect 63572 10816 63573 10856
rect 63531 10807 63573 10816
rect 63051 10772 63093 10781
rect 63051 10732 63052 10772
rect 63092 10732 63093 10772
rect 63051 10723 63093 10732
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 63340 10436 63380 10445
rect 63532 10436 63572 10807
rect 63380 10396 63572 10436
rect 63340 10387 63380 10396
rect 63052 10268 63092 10277
rect 62956 10228 63052 10268
rect 63092 10228 63284 10268
rect 62859 10016 62901 10025
rect 62859 9976 62860 10016
rect 62900 9976 62901 10016
rect 62859 9967 62901 9976
rect 62668 9512 62708 9521
rect 62860 9512 62900 9521
rect 62572 9472 62668 9512
rect 62572 8168 62612 9472
rect 62668 9463 62708 9472
rect 62764 9472 62860 9512
rect 62668 9260 62708 9269
rect 62668 8765 62708 9220
rect 62667 8756 62709 8765
rect 62667 8716 62668 8756
rect 62708 8716 62709 8756
rect 62667 8707 62709 8716
rect 62572 8128 62708 8168
rect 62571 8000 62613 8009
rect 62571 7960 62572 8000
rect 62612 7960 62613 8000
rect 62571 7951 62613 7960
rect 62228 4936 62516 4976
rect 62188 4927 62228 4936
rect 61516 3508 61652 3548
rect 61324 3464 61364 3473
rect 61228 3424 61324 3464
rect 61035 2960 61077 2969
rect 61035 2920 61036 2960
rect 61076 2920 61077 2960
rect 61035 2911 61077 2920
rect 61324 2900 61364 3424
rect 61516 3464 61556 3508
rect 59212 2659 59252 2668
rect 59308 2836 60172 2876
rect 60212 2836 60308 2876
rect 60651 2876 60693 2885
rect 60651 2836 60652 2876
rect 60692 2836 60693 2876
rect 61324 2860 61460 2900
rect 59308 2624 59348 2836
rect 60172 2827 60212 2836
rect 60651 2827 60693 2836
rect 60748 2792 60788 2801
rect 61132 2792 61172 2801
rect 60788 2752 61076 2792
rect 60748 2743 60788 2752
rect 60555 2708 60597 2717
rect 60555 2668 60556 2708
rect 60596 2668 60597 2708
rect 60555 2659 60597 2668
rect 61036 2708 61076 2752
rect 61036 2659 61076 2668
rect 59308 2575 59348 2584
rect 60268 2624 60308 2633
rect 60460 2624 60500 2633
rect 60308 2584 60460 2624
rect 60268 2575 60308 2584
rect 60460 2120 60500 2584
rect 60556 2624 60596 2659
rect 60556 2573 60596 2584
rect 60747 2624 60789 2633
rect 60747 2584 60748 2624
rect 60788 2584 60789 2624
rect 60747 2575 60789 2584
rect 60939 2624 60981 2633
rect 60939 2584 60940 2624
rect 60980 2584 60981 2624
rect 60939 2575 60981 2584
rect 60748 2490 60788 2575
rect 60940 2490 60980 2575
rect 60748 2120 60788 2129
rect 61132 2120 61172 2752
rect 61227 2792 61269 2801
rect 61227 2752 61228 2792
rect 61268 2752 61269 2792
rect 61227 2743 61269 2752
rect 61228 2708 61268 2743
rect 61228 2657 61268 2668
rect 61420 2633 61460 2860
rect 61516 2717 61556 3424
rect 61612 3445 61652 3454
rect 61515 2708 61557 2717
rect 61515 2668 61516 2708
rect 61556 2668 61557 2708
rect 61515 2659 61557 2668
rect 61612 2633 61652 3405
rect 61707 2792 61749 2801
rect 61707 2752 61708 2792
rect 61748 2752 61749 2792
rect 61707 2743 61749 2752
rect 61708 2658 61748 2743
rect 61324 2624 61364 2633
rect 61324 2465 61364 2584
rect 61419 2624 61461 2633
rect 61419 2584 61420 2624
rect 61460 2584 61461 2624
rect 61419 2575 61461 2584
rect 61611 2624 61653 2633
rect 61611 2584 61612 2624
rect 61652 2584 61653 2624
rect 61611 2575 61653 2584
rect 61323 2456 61365 2465
rect 61323 2416 61324 2456
rect 61364 2416 61365 2456
rect 61323 2407 61365 2416
rect 60460 2080 60748 2120
rect 60748 2071 60788 2080
rect 61036 2080 61172 2120
rect 58347 2036 58389 2045
rect 58347 1996 58348 2036
rect 58388 1996 58389 2036
rect 58347 1987 58389 1996
rect 59115 2036 59157 2045
rect 59115 1996 59116 2036
rect 59156 1996 59157 2036
rect 59115 1987 59157 1996
rect 60267 2036 60309 2045
rect 60267 1996 60268 2036
rect 60308 1996 60309 2036
rect 60267 1987 60309 1996
rect 58348 1902 58388 1987
rect 58732 1952 58772 1961
rect 58732 1541 58772 1912
rect 59595 1952 59637 1961
rect 59595 1912 59596 1952
rect 59636 1912 59637 1952
rect 59595 1903 59637 1912
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 58731 1532 58773 1541
rect 58731 1492 58732 1532
rect 58772 1492 58773 1532
rect 58731 1483 58773 1492
rect 59596 1112 59636 1903
rect 60268 1541 60308 1987
rect 60267 1532 60309 1541
rect 60267 1492 60268 1532
rect 60308 1492 60309 1532
rect 60267 1483 60309 1492
rect 59596 1063 59636 1072
rect 59883 1112 59925 1121
rect 59883 1072 59884 1112
rect 59924 1072 59925 1112
rect 59883 1063 59925 1072
rect 60268 1112 60308 1483
rect 61036 1121 61076 2080
rect 61131 1952 61173 1961
rect 61131 1912 61132 1952
rect 61172 1912 61173 1952
rect 61131 1903 61173 1912
rect 61324 1952 61364 1963
rect 61900 1961 61940 4096
rect 61996 4724 62036 4733
rect 61996 3389 62036 4684
rect 62284 4724 62324 4733
rect 62284 4145 62324 4684
rect 62476 4313 62516 4936
rect 62475 4304 62517 4313
rect 62475 4264 62476 4304
rect 62516 4264 62517 4304
rect 62475 4255 62517 4264
rect 62283 4136 62325 4145
rect 62283 4096 62284 4136
rect 62324 4096 62325 4136
rect 62283 4087 62325 4096
rect 62572 3977 62612 7951
rect 62668 7001 62708 8128
rect 62764 7085 62804 9472
rect 62860 9463 62900 9472
rect 62956 9512 62996 10228
rect 63052 10219 63092 10228
rect 63244 10184 63284 10228
rect 64012 10193 64052 10975
rect 64971 10604 65013 10613
rect 64971 10564 64972 10604
rect 65012 10564 65013 10604
rect 64971 10555 65013 10564
rect 64683 10436 64725 10445
rect 64683 10396 64684 10436
rect 64724 10396 64725 10436
rect 64972 10436 65012 10555
rect 64972 10396 65022 10436
rect 64683 10387 64725 10396
rect 64684 10277 64724 10387
rect 64982 10277 65022 10396
rect 65068 10352 65108 14335
rect 65164 12545 65204 14923
rect 65548 14720 65588 14729
rect 65356 14680 65548 14720
rect 65260 13460 65300 13469
rect 65356 13460 65396 14680
rect 65548 14671 65588 14680
rect 65644 14720 65684 15847
rect 65739 15560 65781 15569
rect 65739 15520 65740 15560
rect 65780 15520 65781 15560
rect 65739 15511 65781 15520
rect 65644 14671 65684 14680
rect 65740 14720 65780 15511
rect 65451 14552 65493 14561
rect 65451 14512 65452 14552
rect 65492 14512 65493 14552
rect 65451 14503 65493 14512
rect 65643 14552 65685 14561
rect 65643 14512 65644 14552
rect 65684 14512 65685 14552
rect 65643 14503 65685 14512
rect 65452 14418 65492 14503
rect 65300 13420 65492 13460
rect 65260 13411 65300 13420
rect 65259 13208 65301 13217
rect 65259 13168 65260 13208
rect 65300 13168 65301 13208
rect 65259 13159 65301 13168
rect 65163 12536 65205 12545
rect 65163 12496 65164 12536
rect 65204 12496 65205 12536
rect 65163 12487 65205 12496
rect 65164 11948 65204 12487
rect 65164 11899 65204 11908
rect 65068 10312 65204 10352
rect 64683 10268 64725 10277
rect 64683 10228 64684 10268
rect 64724 10228 64725 10268
rect 64683 10219 64725 10228
rect 64972 10268 65022 10277
rect 65012 10228 65022 10268
rect 63244 10135 63284 10144
rect 64011 10184 64053 10193
rect 64011 10144 64012 10184
rect 64052 10144 64053 10184
rect 64011 10135 64053 10144
rect 64684 10134 64724 10219
rect 64875 10184 64917 10193
rect 64780 10144 64876 10184
rect 64916 10144 64917 10184
rect 63147 10100 63189 10109
rect 63147 10060 63148 10100
rect 63188 10060 63189 10100
rect 63147 10051 63189 10060
rect 62956 9463 62996 9472
rect 63148 9428 63188 10051
rect 64203 10016 64245 10025
rect 64203 9976 64204 10016
rect 64244 9976 64245 10016
rect 64203 9967 64245 9976
rect 64395 10016 64437 10025
rect 64492 10016 64532 10025
rect 64395 9976 64396 10016
rect 64436 9976 64492 10016
rect 64395 9967 64437 9976
rect 64492 9967 64532 9976
rect 63532 9689 63572 9774
rect 63531 9680 63573 9689
rect 63531 9640 63532 9680
rect 63572 9640 63573 9680
rect 63531 9631 63573 9640
rect 64011 9680 64053 9689
rect 64011 9640 64012 9680
rect 64052 9640 64053 9680
rect 64011 9631 64053 9640
rect 64012 9596 64052 9631
rect 64012 9545 64052 9556
rect 63628 9512 63668 9521
rect 63148 9379 63188 9388
rect 63532 9472 63628 9512
rect 63339 9344 63381 9353
rect 63339 9304 63340 9344
rect 63380 9304 63381 9344
rect 63339 9295 63381 9304
rect 63340 9210 63380 9295
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 63052 8840 63092 8849
rect 62955 8756 62997 8765
rect 62955 8716 62956 8756
rect 62996 8716 62997 8756
rect 62955 8707 62997 8716
rect 62859 8672 62901 8681
rect 62859 8632 62860 8672
rect 62900 8632 62901 8672
rect 62859 8623 62901 8632
rect 62860 8538 62900 8623
rect 62956 8622 62996 8707
rect 63052 8093 63092 8800
rect 63532 8840 63572 9472
rect 63628 9463 63668 9472
rect 63723 9512 63765 9521
rect 63723 9472 63724 9512
rect 63764 9472 63765 9512
rect 63723 9463 63765 9472
rect 63820 9512 63860 9521
rect 63724 9378 63764 9463
rect 63820 9353 63860 9472
rect 63819 9344 63861 9353
rect 63819 9304 63820 9344
rect 63860 9304 63861 9344
rect 63819 9295 63861 9304
rect 63820 8933 63860 9295
rect 64204 9260 64244 9967
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 64395 9680 64437 9689
rect 64395 9640 64396 9680
rect 64436 9640 64437 9680
rect 64395 9631 64437 9640
rect 64396 9512 64436 9631
rect 64396 9463 64436 9472
rect 64204 9220 64532 9260
rect 64395 9092 64437 9101
rect 64395 9052 64396 9092
rect 64436 9052 64437 9092
rect 64395 9043 64437 9052
rect 63819 8924 63861 8933
rect 63819 8884 63820 8924
rect 63860 8884 63861 8924
rect 63819 8875 63861 8884
rect 64299 8924 64341 8933
rect 64299 8884 64300 8924
rect 64340 8884 64341 8924
rect 64299 8875 64341 8884
rect 63532 8765 63572 8800
rect 63627 8840 63669 8849
rect 63627 8800 63628 8840
rect 63668 8800 63669 8840
rect 63627 8791 63669 8800
rect 63147 8756 63189 8765
rect 63147 8716 63148 8756
rect 63188 8716 63189 8756
rect 63147 8707 63189 8716
rect 63531 8756 63573 8765
rect 63531 8716 63532 8756
rect 63572 8716 63573 8756
rect 63531 8707 63573 8716
rect 63148 8622 63188 8707
rect 63244 8672 63284 8681
rect 63244 8513 63284 8632
rect 63243 8504 63285 8513
rect 63243 8464 63244 8504
rect 63284 8464 63285 8504
rect 63243 8455 63285 8464
rect 63147 8420 63189 8429
rect 63147 8380 63148 8420
rect 63188 8380 63189 8420
rect 63147 8371 63189 8380
rect 63051 8084 63093 8093
rect 63051 8044 63052 8084
rect 63092 8044 63093 8084
rect 63051 8035 63093 8044
rect 63148 7757 63188 8371
rect 63436 8000 63476 8009
rect 63476 7960 63572 8000
rect 63436 7951 63476 7960
rect 63147 7748 63189 7757
rect 63147 7708 63148 7748
rect 63188 7708 63189 7748
rect 63147 7699 63189 7708
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 63532 7169 63572 7960
rect 63531 7160 63573 7169
rect 63531 7120 63532 7160
rect 63572 7120 63573 7160
rect 63531 7111 63573 7120
rect 62763 7076 62805 7085
rect 62763 7036 62764 7076
rect 62804 7036 62805 7076
rect 62763 7027 62805 7036
rect 62667 6992 62709 7001
rect 62667 6952 62668 6992
rect 62708 6952 62709 6992
rect 62667 6943 62709 6952
rect 62764 5909 62804 7027
rect 63531 6740 63573 6749
rect 63531 6700 63532 6740
rect 63572 6700 63573 6740
rect 63531 6691 63573 6700
rect 63532 6656 63572 6691
rect 63532 6605 63572 6616
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 62763 5900 62805 5909
rect 62763 5860 62764 5900
rect 62804 5860 62805 5900
rect 62763 5851 62805 5860
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 63051 4304 63093 4313
rect 63628 4304 63668 8791
rect 63820 8716 64244 8756
rect 63820 8672 63860 8716
rect 64204 8672 64244 8716
rect 63820 8623 63860 8632
rect 63916 8662 63956 8671
rect 64204 8623 64244 8632
rect 64300 8672 64340 8875
rect 63916 8597 63956 8622
rect 63915 8588 63957 8597
rect 63915 8548 63916 8588
rect 63956 8548 63957 8588
rect 63915 8539 63957 8548
rect 63916 8527 63956 8539
rect 64012 8513 64052 8570
rect 64300 8513 64340 8632
rect 64396 8672 64436 9043
rect 64492 8765 64532 9220
rect 64780 9101 64820 10144
rect 64875 10135 64917 10144
rect 64876 10050 64916 10135
rect 64972 9521 65012 10228
rect 65164 10184 65204 10312
rect 65068 10144 65204 10184
rect 65068 10100 65108 10144
rect 65068 10060 65204 10100
rect 65067 9680 65109 9689
rect 65067 9640 65068 9680
rect 65108 9640 65109 9680
rect 65067 9631 65109 9640
rect 64971 9512 65013 9521
rect 64971 9472 64972 9512
rect 65012 9472 65013 9512
rect 64971 9463 65013 9472
rect 64779 9092 64821 9101
rect 64779 9052 64780 9092
rect 64820 9052 64821 9092
rect 64779 9043 64821 9052
rect 64491 8756 64533 8765
rect 64491 8716 64492 8756
rect 64532 8716 64533 8756
rect 64491 8707 64533 8716
rect 64396 8623 64436 8632
rect 64492 8672 64532 8707
rect 64492 8597 64532 8632
rect 64971 8672 65013 8681
rect 64971 8632 64972 8672
rect 65012 8632 65013 8672
rect 64971 8623 65013 8632
rect 64491 8588 64533 8597
rect 64491 8548 64492 8588
rect 64532 8548 64533 8588
rect 64491 8539 64533 8548
rect 64011 8504 64053 8513
rect 64011 8464 64012 8504
rect 64052 8464 64053 8504
rect 64011 8455 64053 8464
rect 64299 8504 64341 8513
rect 64492 8508 64532 8539
rect 64299 8464 64300 8504
rect 64340 8464 64341 8504
rect 64299 8455 64341 8464
rect 64012 8446 64052 8455
rect 64012 7412 64052 8406
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 64972 7916 65012 8623
rect 65068 8597 65108 9631
rect 65067 8588 65109 8597
rect 65067 8548 65068 8588
rect 65108 8548 65109 8588
rect 65067 8539 65109 8548
rect 64972 7867 65012 7876
rect 64588 7748 64628 7757
rect 64780 7748 64820 7757
rect 64012 7363 64052 7372
rect 64300 7708 64588 7748
rect 64108 7160 64148 7169
rect 64300 7160 64340 7708
rect 64588 7699 64628 7708
rect 64684 7708 64780 7748
rect 64588 7337 64628 7422
rect 64587 7328 64629 7337
rect 64587 7288 64588 7328
rect 64628 7288 64629 7328
rect 64587 7279 64629 7288
rect 64148 7120 64300 7160
rect 64108 7111 64148 7120
rect 64300 7111 64340 7120
rect 64396 7160 64436 7171
rect 64396 7085 64436 7120
rect 64588 7160 64628 7169
rect 64684 7160 64724 7708
rect 64780 7699 64820 7708
rect 64628 7120 64724 7160
rect 64779 7160 64821 7169
rect 64779 7120 64780 7160
rect 64820 7120 64821 7160
rect 64011 7076 64053 7085
rect 64011 7036 64012 7076
rect 64052 7036 64053 7076
rect 64011 7027 64053 7036
rect 64395 7076 64437 7085
rect 64395 7036 64396 7076
rect 64436 7036 64437 7076
rect 64395 7027 64437 7036
rect 63723 6656 63765 6665
rect 63723 6616 63724 6656
rect 63764 6616 63765 6656
rect 63723 6607 63765 6616
rect 63724 6522 63764 6607
rect 63051 4264 63052 4304
rect 63092 4264 63093 4304
rect 63051 4255 63093 4264
rect 63532 4264 63668 4304
rect 64012 4892 64052 7027
rect 64588 7001 64628 7120
rect 64779 7111 64821 7120
rect 64876 7160 64916 7169
rect 64203 6992 64245 7001
rect 64203 6952 64204 6992
rect 64244 6952 64245 6992
rect 64203 6943 64245 6952
rect 64587 6992 64629 7001
rect 64587 6952 64588 6992
rect 64628 6952 64629 6992
rect 64587 6943 64629 6952
rect 64107 6656 64149 6665
rect 64107 6616 64108 6656
rect 64148 6616 64149 6656
rect 64107 6607 64149 6616
rect 64108 4991 64148 6607
rect 64204 5732 64244 6943
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 64780 6488 64820 7111
rect 64876 6665 64916 7120
rect 65068 7085 65108 8539
rect 65067 7076 65109 7085
rect 65067 7036 65068 7076
rect 65108 7036 65109 7076
rect 65164 7076 65204 10060
rect 65260 9680 65300 13159
rect 65355 13124 65397 13133
rect 65355 13084 65356 13124
rect 65396 13084 65397 13124
rect 65355 13075 65397 13084
rect 65356 11696 65396 13075
rect 65452 11780 65492 13420
rect 65548 13208 65588 13217
rect 65548 12965 65588 13168
rect 65644 13208 65684 14503
rect 65740 13544 65780 14680
rect 65835 14048 65877 14057
rect 65835 14008 65836 14048
rect 65876 14008 65877 14048
rect 65835 13999 65877 14008
rect 65836 13914 65876 13999
rect 65932 13721 65972 17032
rect 66315 17023 66357 17032
rect 67179 17023 67221 17032
rect 66219 16904 66261 16913
rect 66219 16864 66220 16904
rect 66260 16864 66261 16904
rect 66219 16855 66261 16864
rect 66220 16745 66260 16855
rect 66219 16736 66261 16745
rect 66219 16696 66220 16736
rect 66260 16696 66261 16736
rect 66219 16687 66261 16696
rect 66603 16736 66645 16745
rect 66603 16696 66604 16736
rect 66644 16696 66645 16736
rect 66603 16687 66645 16696
rect 66123 16568 66165 16577
rect 66123 16528 66124 16568
rect 66164 16528 66165 16568
rect 66123 16519 66165 16528
rect 66124 16484 66164 16519
rect 66124 16433 66164 16444
rect 66028 16232 66068 16241
rect 66028 14225 66068 16192
rect 66315 16232 66357 16241
rect 66315 16192 66316 16232
rect 66356 16192 66357 16232
rect 66315 16183 66357 16192
rect 66604 16232 66644 16687
rect 66699 16652 66741 16661
rect 66699 16612 66700 16652
rect 66740 16612 66741 16652
rect 66699 16603 66741 16612
rect 66700 16484 66740 16603
rect 66700 16435 66740 16444
rect 67372 16409 67412 17191
rect 67545 17072 67585 17472
rect 67655 17324 67695 17472
rect 67655 17284 67700 17324
rect 67545 17032 67604 17072
rect 67564 16913 67604 17032
rect 67563 16904 67605 16913
rect 67563 16864 67564 16904
rect 67604 16864 67605 16904
rect 67563 16855 67605 16864
rect 67371 16400 67413 16409
rect 67371 16360 67372 16400
rect 67412 16360 67413 16400
rect 67371 16351 67413 16360
rect 67563 16400 67605 16409
rect 67563 16360 67564 16400
rect 67604 16360 67605 16400
rect 67563 16351 67605 16360
rect 66604 16183 66644 16192
rect 67276 16232 67316 16241
rect 66316 16098 66356 16183
rect 66892 16148 66932 16157
rect 66124 16064 66164 16073
rect 66124 15905 66164 16024
rect 66700 16064 66740 16075
rect 66700 15989 66740 16024
rect 66699 15980 66741 15989
rect 66699 15940 66700 15980
rect 66740 15940 66741 15980
rect 66699 15931 66741 15940
rect 66123 15896 66165 15905
rect 66123 15856 66124 15896
rect 66164 15856 66165 15896
rect 66123 15847 66165 15856
rect 66892 15728 66932 16108
rect 67083 15980 67125 15989
rect 67083 15940 67084 15980
rect 67124 15940 67125 15980
rect 67083 15931 67125 15940
rect 66892 15679 66932 15688
rect 66988 15560 67028 15569
rect 66988 14888 67028 15520
rect 67084 15560 67124 15931
rect 67276 15905 67316 16192
rect 67564 16073 67604 16351
rect 67563 16064 67605 16073
rect 67563 16024 67564 16064
rect 67604 16024 67605 16064
rect 67563 16015 67605 16024
rect 67275 15896 67317 15905
rect 67275 15856 67276 15896
rect 67316 15856 67317 15896
rect 67275 15847 67317 15856
rect 67467 15644 67509 15653
rect 67467 15604 67468 15644
rect 67508 15604 67509 15644
rect 67467 15595 67509 15604
rect 67084 15511 67124 15520
rect 67179 15560 67221 15569
rect 67179 15520 67180 15560
rect 67220 15520 67221 15560
rect 67179 15511 67221 15520
rect 67180 15426 67220 15511
rect 67468 15510 67508 15595
rect 67564 15560 67604 16015
rect 67564 15511 67604 15520
rect 67660 15401 67700 17284
rect 67945 17072 67985 17472
rect 68055 17072 68095 17472
rect 68345 17072 68385 17472
rect 68455 17072 68495 17472
rect 68745 17324 68785 17472
rect 67945 17032 67988 17072
rect 67948 16325 67988 17032
rect 68044 17032 68095 17072
rect 68332 17032 68385 17072
rect 68428 17032 68495 17072
rect 68620 17284 68785 17324
rect 68044 16829 68084 17032
rect 68043 16820 68085 16829
rect 68043 16780 68044 16820
rect 68084 16780 68085 16820
rect 68043 16771 68085 16780
rect 68332 16409 68372 17032
rect 68331 16400 68373 16409
rect 68331 16360 68332 16400
rect 68372 16360 68373 16400
rect 68331 16351 68373 16360
rect 67947 16316 67989 16325
rect 67947 16276 67948 16316
rect 67988 16276 67989 16316
rect 67947 16267 67989 16276
rect 67755 16232 67797 16241
rect 67755 16192 67756 16232
rect 67796 16192 67797 16232
rect 67755 16183 67797 16192
rect 68140 16232 68180 16241
rect 68180 16192 68372 16232
rect 68140 16183 68180 16192
rect 67659 15392 67701 15401
rect 67659 15352 67660 15392
rect 67700 15352 67701 15392
rect 67659 15343 67701 15352
rect 67371 15308 67413 15317
rect 67371 15268 67372 15308
rect 67412 15268 67413 15308
rect 67371 15259 67413 15268
rect 67180 14888 67220 14897
rect 66988 14848 67180 14888
rect 67220 14848 67316 14888
rect 67180 14839 67220 14848
rect 66315 14384 66357 14393
rect 66315 14344 66316 14384
rect 66356 14344 66357 14384
rect 66315 14335 66357 14344
rect 66027 14216 66069 14225
rect 66027 14176 66028 14216
rect 66068 14176 66164 14216
rect 66027 14167 66069 14176
rect 65931 13712 65973 13721
rect 65931 13672 65932 13712
rect 65972 13672 65973 13712
rect 65931 13663 65973 13672
rect 65740 13504 66068 13544
rect 65547 12956 65589 12965
rect 65547 12916 65548 12956
rect 65588 12916 65589 12956
rect 65547 12907 65589 12916
rect 65644 12704 65684 13168
rect 66028 13208 66068 13504
rect 65739 13124 65781 13133
rect 65739 13084 65740 13124
rect 65780 13084 65781 13124
rect 65739 13075 65781 13084
rect 65740 13036 65780 13075
rect 65932 13049 65972 13134
rect 65740 12987 65780 12996
rect 65931 13040 65973 13049
rect 65931 13000 65932 13040
rect 65972 13000 65973 13040
rect 65931 12991 65973 13000
rect 66028 12980 66068 13168
rect 66124 13208 66164 14176
rect 66219 13376 66261 13385
rect 66219 13336 66220 13376
rect 66260 13336 66261 13376
rect 66219 13327 66261 13336
rect 66124 13159 66164 13168
rect 66220 13208 66260 13327
rect 66220 13159 66260 13168
rect 66028 12940 66260 12980
rect 65644 12664 66068 12704
rect 65643 12536 65685 12545
rect 65643 12496 65644 12536
rect 65684 12496 65685 12536
rect 65643 12487 65685 12496
rect 65644 12402 65684 12487
rect 65547 11864 65589 11873
rect 65932 11864 65972 11873
rect 65547 11824 65548 11864
rect 65588 11824 65589 11864
rect 65547 11815 65589 11824
rect 65644 11824 65932 11864
rect 65452 11731 65492 11740
rect 65548 11730 65588 11815
rect 65644 11780 65684 11824
rect 65932 11815 65972 11824
rect 65644 11731 65684 11740
rect 65356 11647 65396 11656
rect 65739 11696 65781 11705
rect 65739 11656 65740 11696
rect 65780 11656 65781 11696
rect 65739 11647 65781 11656
rect 65931 11696 65973 11705
rect 65931 11656 65932 11696
rect 65972 11656 65973 11696
rect 65931 11647 65973 11656
rect 65740 11562 65780 11647
rect 65932 11562 65972 11647
rect 66028 11444 66068 12664
rect 66220 12629 66260 12940
rect 66219 12620 66261 12629
rect 66219 12580 66220 12620
rect 66260 12580 66261 12620
rect 66219 12571 66261 12580
rect 66123 12032 66165 12041
rect 66123 11992 66124 12032
rect 66164 11992 66165 12032
rect 66123 11983 66165 11992
rect 66124 11696 66164 11983
rect 66124 11621 66164 11656
rect 66220 11696 66260 11705
rect 66123 11612 66165 11621
rect 66123 11572 66124 11612
rect 66164 11572 66165 11612
rect 66123 11563 66165 11572
rect 66220 11537 66260 11656
rect 66219 11528 66261 11537
rect 66219 11488 66220 11528
rect 66260 11488 66261 11528
rect 66219 11479 66261 11488
rect 66028 11404 66164 11444
rect 65931 11024 65973 11033
rect 65931 10984 65932 11024
rect 65972 10984 65973 11024
rect 65931 10975 65973 10984
rect 65260 9640 65492 9680
rect 65259 9512 65301 9521
rect 65259 9472 65260 9512
rect 65300 9472 65301 9512
rect 65259 9463 65301 9472
rect 65260 9378 65300 9463
rect 65259 8756 65301 8765
rect 65259 8716 65260 8756
rect 65300 8716 65301 8756
rect 65259 8707 65301 8716
rect 65260 7203 65300 8707
rect 65355 8336 65397 8345
rect 65355 8296 65356 8336
rect 65396 8296 65397 8336
rect 65355 8287 65397 8296
rect 65260 7154 65300 7163
rect 65356 7160 65396 8287
rect 65356 7111 65396 7120
rect 65164 7036 65300 7076
rect 65067 7027 65109 7036
rect 64972 6992 65012 7001
rect 64972 6908 65012 6952
rect 65164 6934 65204 6943
rect 64972 6894 65164 6908
rect 65260 6917 65300 7036
rect 64972 6868 65204 6894
rect 65259 6908 65301 6917
rect 65259 6868 65260 6908
rect 65300 6868 65301 6908
rect 64875 6656 64917 6665
rect 64875 6616 64876 6656
rect 64916 6616 64917 6656
rect 64875 6607 64917 6616
rect 64875 6488 64917 6497
rect 64780 6448 64876 6488
rect 64916 6448 64917 6488
rect 64875 6439 64917 6448
rect 64876 6354 64916 6439
rect 64972 6236 65012 6868
rect 65259 6859 65301 6868
rect 64876 6196 65012 6236
rect 64587 5900 64629 5909
rect 64587 5860 64588 5900
rect 64628 5860 64629 5900
rect 64587 5851 64629 5860
rect 64588 5732 64628 5851
rect 64683 5816 64725 5825
rect 64683 5776 64684 5816
rect 64724 5776 64725 5816
rect 64683 5767 64725 5776
rect 64204 5692 64532 5732
rect 64204 5144 64244 5692
rect 64492 5648 64532 5692
rect 64588 5683 64628 5692
rect 64684 5682 64724 5767
rect 64779 5732 64821 5741
rect 64779 5692 64780 5732
rect 64820 5692 64821 5732
rect 64779 5683 64821 5692
rect 64492 5599 64532 5608
rect 64780 5598 64820 5683
rect 64876 5648 64916 6196
rect 65355 5900 65397 5909
rect 65355 5860 65356 5900
rect 65396 5860 65397 5900
rect 65355 5851 65397 5860
rect 65260 5657 65300 5742
rect 65164 5648 65204 5657
rect 64876 5599 64916 5608
rect 64972 5608 65164 5648
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 64972 5153 65012 5608
rect 65164 5599 65204 5608
rect 65259 5648 65301 5657
rect 65259 5608 65260 5648
rect 65300 5608 65301 5648
rect 65259 5599 65301 5608
rect 65356 5648 65396 5851
rect 65356 5599 65396 5608
rect 65452 5573 65492 9640
rect 65932 9521 65972 10975
rect 66124 10697 66164 11404
rect 66220 11201 66260 11479
rect 66219 11192 66261 11201
rect 66219 11152 66220 11192
rect 66260 11152 66261 11192
rect 66219 11143 66261 11152
rect 66123 10688 66165 10697
rect 66123 10648 66124 10688
rect 66164 10648 66165 10688
rect 66123 10639 66165 10648
rect 65931 9512 65973 9521
rect 65931 9472 65932 9512
rect 65972 9472 65973 9512
rect 65931 9463 65973 9472
rect 65931 8924 65973 8933
rect 65931 8884 65932 8924
rect 65972 8884 65973 8924
rect 65931 8875 65973 8884
rect 65932 8790 65972 8875
rect 66027 8504 66069 8513
rect 66027 8464 66028 8504
rect 66068 8464 66069 8504
rect 66027 8455 66069 8464
rect 65931 8168 65973 8177
rect 65644 8128 65876 8168
rect 65644 7328 65684 8128
rect 65740 8000 65780 8009
rect 65740 7421 65780 7960
rect 65836 8000 65876 8128
rect 65931 8128 65932 8168
rect 65972 8128 65973 8168
rect 65931 8119 65973 8128
rect 65836 7951 65876 7960
rect 65932 8000 65972 8119
rect 66028 8009 66068 8455
rect 65932 7951 65972 7960
rect 66027 8000 66069 8009
rect 66027 7960 66028 8000
rect 66068 7960 66069 8000
rect 66027 7951 66069 7960
rect 66124 7832 66164 10639
rect 66316 8849 66356 14335
rect 66988 14225 67028 14310
rect 66987 14216 67029 14225
rect 66987 14176 66988 14216
rect 67028 14176 67029 14216
rect 66987 14167 67029 14176
rect 67180 14048 67220 14057
rect 66892 14008 67180 14048
rect 66699 13544 66741 13553
rect 66699 13504 66700 13544
rect 66740 13504 66741 13544
rect 66699 13495 66741 13504
rect 66508 13301 66548 13316
rect 66507 13292 66549 13301
rect 66507 13252 66508 13292
rect 66548 13252 66549 13292
rect 66507 13243 66549 13252
rect 66508 13221 66548 13243
rect 66508 13172 66548 13181
rect 66700 13208 66740 13495
rect 66795 13376 66837 13385
rect 66795 13336 66796 13376
rect 66836 13336 66837 13376
rect 66795 13327 66837 13336
rect 66892 13376 66932 14008
rect 67180 13999 67220 14008
rect 67276 13628 67316 14848
rect 67372 13712 67412 15259
rect 67467 14720 67509 14729
rect 67467 14680 67468 14720
rect 67508 14680 67509 14720
rect 67467 14671 67509 14680
rect 67564 14720 67604 14731
rect 67468 14586 67508 14671
rect 67564 14645 67604 14680
rect 67563 14636 67605 14645
rect 67563 14596 67564 14636
rect 67604 14596 67605 14636
rect 67563 14587 67605 14596
rect 67660 14494 67700 14503
rect 67564 14048 67604 14057
rect 67372 13672 67508 13712
rect 66892 13327 66932 13336
rect 66988 13588 67316 13628
rect 66796 13292 66836 13327
rect 66796 13241 66836 13252
rect 66988 13292 67028 13588
rect 67371 13544 67413 13553
rect 67371 13504 67372 13544
rect 67412 13504 67413 13544
rect 67371 13495 67413 13504
rect 67179 13460 67221 13469
rect 67179 13420 67180 13460
rect 67220 13420 67221 13460
rect 67179 13411 67221 13420
rect 66988 13243 67028 13252
rect 66700 13159 66740 13168
rect 67083 13208 67125 13217
rect 67083 13168 67084 13208
rect 67124 13168 67125 13208
rect 67083 13159 67125 13168
rect 66411 13124 66453 13133
rect 66411 13084 66412 13124
rect 66452 13084 66453 13124
rect 66411 13075 66453 13084
rect 66795 13124 66837 13133
rect 66795 13084 66796 13124
rect 66836 13084 66837 13124
rect 66795 13075 66837 13084
rect 66987 13124 67029 13133
rect 66987 13084 66988 13124
rect 67028 13084 67029 13124
rect 66987 13075 67029 13084
rect 66412 12990 66452 13075
rect 66796 12980 66836 13075
rect 66603 12956 66645 12965
rect 66603 12916 66604 12956
rect 66644 12916 66645 12956
rect 66603 12907 66645 12916
rect 66700 12940 66836 12980
rect 66604 12461 66644 12907
rect 66603 12452 66645 12461
rect 66603 12412 66604 12452
rect 66644 12412 66645 12452
rect 66603 12403 66645 12412
rect 66604 11024 66644 12403
rect 66700 11192 66740 12940
rect 66796 12704 66836 12713
rect 66988 12704 67028 13075
rect 67084 13074 67124 13159
rect 67180 12980 67220 13411
rect 67276 13385 67316 13470
rect 67275 13376 67317 13385
rect 67275 13336 67276 13376
rect 67316 13336 67317 13376
rect 67275 13327 67317 13336
rect 67276 13208 67316 13217
rect 67372 13208 67412 13495
rect 67468 13469 67508 13672
rect 67467 13460 67509 13469
rect 67467 13420 67468 13460
rect 67508 13420 67509 13460
rect 67467 13411 67509 13420
rect 67564 13385 67604 14008
rect 67563 13376 67605 13385
rect 67563 13336 67564 13376
rect 67604 13336 67605 13376
rect 67563 13327 67605 13336
rect 67660 13217 67700 14454
rect 67316 13168 67412 13208
rect 67468 13208 67508 13217
rect 67276 13159 67316 13168
rect 67180 12940 67316 12980
rect 66836 12664 67028 12704
rect 66796 12655 66836 12664
rect 67179 12620 67221 12629
rect 67179 12580 67180 12620
rect 67220 12580 67221 12620
rect 67179 12571 67221 12580
rect 66892 11696 66932 11705
rect 66892 11537 66932 11656
rect 67083 11696 67125 11705
rect 67083 11656 67084 11696
rect 67124 11656 67125 11696
rect 67083 11647 67125 11656
rect 67180 11696 67220 12571
rect 67180 11647 67220 11656
rect 67276 11696 67316 12940
rect 67468 11789 67508 13168
rect 67564 13208 67604 13217
rect 67564 13133 67604 13168
rect 67659 13208 67701 13217
rect 67659 13168 67660 13208
rect 67700 13168 67701 13208
rect 67659 13159 67701 13168
rect 67562 13124 67604 13133
rect 67562 13084 67563 13124
rect 67603 13084 67604 13124
rect 67562 13075 67604 13084
rect 67756 12713 67796 16183
rect 68139 16064 68181 16073
rect 68139 16024 68140 16064
rect 68180 16024 68181 16064
rect 68139 16015 68181 16024
rect 67948 15560 67988 15569
rect 67948 14729 67988 15520
rect 68043 15560 68085 15569
rect 68043 15520 68044 15560
rect 68084 15520 68085 15560
rect 68043 15511 68085 15520
rect 68140 15560 68180 16015
rect 68140 15511 68180 15520
rect 68236 15560 68276 15569
rect 68044 15426 68084 15511
rect 68139 15392 68181 15401
rect 68139 15352 68140 15392
rect 68180 15352 68181 15392
rect 68139 15343 68181 15352
rect 67947 14720 67989 14729
rect 67947 14680 67948 14720
rect 67988 14680 67989 14720
rect 67947 14671 67989 14680
rect 68140 13637 68180 15343
rect 68236 14645 68276 15520
rect 68235 14636 68277 14645
rect 68235 14596 68236 14636
rect 68276 14596 68277 14636
rect 68235 14587 68277 14596
rect 68332 14048 68372 16192
rect 68428 15737 68468 17032
rect 68620 16157 68660 17284
rect 68855 17072 68895 17472
rect 69145 17156 69185 17472
rect 68812 17032 68895 17072
rect 69100 17116 69185 17156
rect 68715 16736 68757 16745
rect 68715 16696 68716 16736
rect 68756 16696 68757 16736
rect 68715 16687 68757 16696
rect 68619 16148 68661 16157
rect 68619 16108 68620 16148
rect 68660 16108 68661 16148
rect 68619 16099 68661 16108
rect 68619 15896 68661 15905
rect 68619 15856 68620 15896
rect 68660 15856 68661 15896
rect 68619 15847 68661 15856
rect 68427 15728 68469 15737
rect 68427 15688 68428 15728
rect 68468 15688 68469 15728
rect 68427 15679 68469 15688
rect 68427 15560 68469 15569
rect 68427 15520 68428 15560
rect 68468 15520 68469 15560
rect 68427 15511 68469 15520
rect 68428 15426 68468 15511
rect 68523 15476 68565 15485
rect 68523 15436 68524 15476
rect 68564 15436 68565 15476
rect 68523 15427 68565 15436
rect 68524 15342 68564 15427
rect 68620 15140 68660 15847
rect 68524 15100 68660 15140
rect 68428 14804 68468 14813
rect 68428 14561 68468 14764
rect 68427 14552 68469 14561
rect 68427 14512 68428 14552
rect 68468 14512 68469 14552
rect 68427 14503 68469 14512
rect 68428 14048 68468 14057
rect 68332 14008 68428 14048
rect 68235 13796 68277 13805
rect 68235 13756 68236 13796
rect 68276 13756 68277 13796
rect 68235 13747 68277 13756
rect 68139 13628 68181 13637
rect 68139 13588 68140 13628
rect 68180 13588 68181 13628
rect 68139 13579 68181 13588
rect 68043 13292 68085 13301
rect 68043 13252 68044 13292
rect 68084 13252 68085 13292
rect 68043 13243 68085 13252
rect 68044 12980 68084 13243
rect 68139 13208 68181 13217
rect 68139 13168 68140 13208
rect 68180 13168 68181 13208
rect 68139 13159 68181 13168
rect 68236 13208 68276 13747
rect 68331 13292 68373 13301
rect 68331 13252 68332 13292
rect 68372 13252 68373 13292
rect 68331 13243 68373 13252
rect 68236 13159 68276 13168
rect 68140 13074 68180 13159
rect 68235 13040 68277 13049
rect 68235 13000 68236 13040
rect 68276 13000 68277 13040
rect 68235 12991 68277 13000
rect 68044 12940 68180 12980
rect 67755 12704 67797 12713
rect 67755 12664 67756 12704
rect 67796 12664 67797 12704
rect 67755 12655 67797 12664
rect 67947 12620 67989 12629
rect 67947 12580 67948 12620
rect 67988 12580 67989 12620
rect 67947 12571 67989 12580
rect 67852 12536 67892 12545
rect 67756 12496 67852 12536
rect 67467 11780 67509 11789
rect 67467 11740 67468 11780
rect 67508 11740 67509 11780
rect 67467 11731 67509 11740
rect 67276 11647 67316 11656
rect 67372 11696 67412 11705
rect 66891 11528 66933 11537
rect 66891 11488 66892 11528
rect 66932 11488 66933 11528
rect 66891 11479 66933 11488
rect 66988 11528 67028 11537
rect 66988 11285 67028 11488
rect 66987 11276 67029 11285
rect 66987 11236 66988 11276
rect 67028 11236 67029 11276
rect 66987 11227 67029 11236
rect 66700 11152 66932 11192
rect 66796 11024 66836 11033
rect 66604 10984 66796 11024
rect 66796 10975 66836 10984
rect 66795 10856 66837 10865
rect 66795 10816 66796 10856
rect 66836 10816 66837 10856
rect 66795 10807 66837 10816
rect 66411 10520 66453 10529
rect 66411 10480 66412 10520
rect 66452 10480 66453 10520
rect 66411 10471 66453 10480
rect 66412 10193 66452 10471
rect 66603 10268 66645 10277
rect 66603 10228 66604 10268
rect 66644 10228 66645 10268
rect 66603 10219 66645 10228
rect 66411 10184 66453 10193
rect 66411 10144 66412 10184
rect 66452 10144 66453 10184
rect 66411 10135 66453 10144
rect 66412 9680 66452 10135
rect 66507 10100 66549 10109
rect 66507 10060 66508 10100
rect 66548 10060 66549 10100
rect 66507 10051 66549 10060
rect 66412 9631 66452 9640
rect 66508 8924 66548 10051
rect 66412 8884 66548 8924
rect 66315 8840 66357 8849
rect 66315 8800 66316 8840
rect 66356 8800 66357 8840
rect 66315 8791 66357 8800
rect 66219 8336 66261 8345
rect 66219 8296 66220 8336
rect 66260 8296 66261 8336
rect 66219 8287 66261 8296
rect 66220 8168 66260 8287
rect 66412 8261 66452 8884
rect 66507 8756 66549 8765
rect 66507 8716 66508 8756
rect 66548 8716 66549 8756
rect 66507 8707 66549 8716
rect 66411 8252 66453 8261
rect 66411 8212 66412 8252
rect 66452 8212 66453 8252
rect 66411 8203 66453 8212
rect 66220 8119 66260 8128
rect 66411 8000 66453 8009
rect 66316 7958 66356 7967
rect 66315 7918 66316 7925
rect 66411 7960 66412 8000
rect 66452 7960 66453 8000
rect 66411 7951 66453 7960
rect 66508 8000 66548 8707
rect 66508 7951 66548 7960
rect 66356 7918 66357 7925
rect 66315 7916 66357 7918
rect 66315 7876 66316 7916
rect 66356 7876 66357 7916
rect 66315 7867 66357 7876
rect 66028 7792 66164 7832
rect 65739 7412 65781 7421
rect 65739 7372 65740 7412
rect 65780 7372 65781 7412
rect 65739 7363 65781 7372
rect 65548 7288 65644 7328
rect 65548 5741 65588 7288
rect 65644 7279 65684 7288
rect 65739 7076 65781 7085
rect 65739 7036 65740 7076
rect 65780 7036 65781 7076
rect 65739 7027 65781 7036
rect 65740 6488 65780 7027
rect 65740 6161 65780 6448
rect 65739 6152 65781 6161
rect 65739 6112 65740 6152
rect 65780 6112 65781 6152
rect 65739 6103 65781 6112
rect 65739 5984 65781 5993
rect 65739 5944 65740 5984
rect 65780 5944 65781 5984
rect 65739 5935 65781 5944
rect 65643 5900 65685 5909
rect 65643 5860 65644 5900
rect 65684 5860 65685 5900
rect 65643 5851 65685 5860
rect 65547 5732 65589 5741
rect 65547 5692 65548 5732
rect 65588 5692 65589 5732
rect 65547 5683 65589 5692
rect 65644 5657 65684 5851
rect 65643 5648 65685 5657
rect 65643 5608 65644 5648
rect 65684 5608 65685 5648
rect 65643 5599 65685 5608
rect 65740 5648 65780 5935
rect 65451 5564 65493 5573
rect 65451 5524 65452 5564
rect 65492 5524 65493 5564
rect 65451 5515 65493 5524
rect 65068 5480 65108 5489
rect 65548 5480 65588 5489
rect 65108 5440 65396 5480
rect 65068 5431 65108 5440
rect 64587 5144 64629 5153
rect 64204 5104 64436 5144
rect 64108 4942 64148 4951
rect 64204 4962 64244 4971
rect 64204 4892 64244 4922
rect 64012 4852 64244 4892
rect 63052 4170 63092 4255
rect 63244 4052 63284 4061
rect 62571 3968 62613 3977
rect 62571 3928 62572 3968
rect 62612 3928 62613 3968
rect 62571 3919 62613 3928
rect 62091 3716 62133 3725
rect 62091 3676 62092 3716
rect 62132 3676 62133 3716
rect 62091 3667 62133 3676
rect 61995 3380 62037 3389
rect 61995 3340 61996 3380
rect 62036 3340 62037 3380
rect 61995 3331 62037 3340
rect 61996 3246 62036 3331
rect 62092 2969 62132 3667
rect 63244 3305 63284 4012
rect 63243 3296 63285 3305
rect 63243 3256 63244 3296
rect 63284 3256 63285 3296
rect 63243 3247 63285 3256
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 62091 2960 62133 2969
rect 62091 2920 62092 2960
rect 62132 2920 62133 2960
rect 62091 2911 62133 2920
rect 62763 2960 62805 2969
rect 62763 2920 62764 2960
rect 62804 2920 62805 2960
rect 62763 2911 62805 2920
rect 61996 2624 62036 2633
rect 60268 1063 60308 1072
rect 61035 1112 61077 1121
rect 61035 1072 61036 1112
rect 61076 1072 61077 1112
rect 61035 1063 61077 1072
rect 61132 1112 61172 1903
rect 61324 1877 61364 1912
rect 61899 1952 61941 1961
rect 61899 1912 61900 1952
rect 61940 1912 61941 1952
rect 61899 1903 61941 1912
rect 61323 1868 61365 1877
rect 61323 1828 61324 1868
rect 61364 1828 61365 1868
rect 61323 1819 61365 1828
rect 61900 1784 61940 1903
rect 61900 1735 61940 1744
rect 61996 1196 62036 2584
rect 62092 2624 62132 2911
rect 62667 2876 62709 2885
rect 62667 2836 62668 2876
rect 62708 2836 62709 2876
rect 62667 2827 62709 2836
rect 62475 2792 62517 2801
rect 62475 2752 62476 2792
rect 62516 2752 62517 2792
rect 62475 2743 62517 2752
rect 62092 2575 62132 2584
rect 62283 2624 62325 2633
rect 62283 2584 62284 2624
rect 62324 2584 62325 2624
rect 62283 2575 62325 2584
rect 62476 2624 62516 2743
rect 62571 2708 62613 2717
rect 62571 2668 62572 2708
rect 62612 2668 62613 2708
rect 62571 2659 62613 2668
rect 62476 2575 62516 2584
rect 62572 2624 62612 2659
rect 62187 2456 62229 2465
rect 62187 2412 62188 2456
rect 62228 2412 62229 2456
rect 62187 2407 62229 2412
rect 62188 2321 62228 2407
rect 62284 1364 62324 2575
rect 62572 2573 62612 2584
rect 62668 2624 62708 2827
rect 62380 2456 62420 2465
rect 62380 2036 62420 2416
rect 62380 1987 62420 1996
rect 62284 1315 62324 1324
rect 61996 1156 62612 1196
rect 61132 1063 61172 1072
rect 62572 1112 62612 1156
rect 62572 1063 62612 1072
rect 62668 1112 62708 2584
rect 62764 2372 62804 2911
rect 63532 2900 63572 4264
rect 63628 4136 63668 4145
rect 63628 3977 63668 4096
rect 63627 3968 63669 3977
rect 63627 3928 63628 3968
rect 63668 3928 63669 3968
rect 63627 3919 63669 3928
rect 63340 2876 63572 2900
rect 63380 2860 63572 2876
rect 63340 2717 63380 2836
rect 63339 2708 63381 2717
rect 63339 2668 63340 2708
rect 63380 2668 63381 2708
rect 63339 2659 63381 2668
rect 62859 2624 62901 2633
rect 62859 2584 62860 2624
rect 62900 2584 62901 2624
rect 62859 2575 62901 2584
rect 63244 2624 63284 2633
rect 62860 2490 62900 2575
rect 62955 2456 62997 2465
rect 62955 2416 62956 2456
rect 62996 2416 62997 2456
rect 62955 2407 62997 2416
rect 62764 2332 62900 2372
rect 62763 2036 62805 2045
rect 62763 1996 62764 2036
rect 62804 1996 62805 2036
rect 62763 1987 62805 1996
rect 62764 1952 62804 1987
rect 62764 1901 62804 1912
rect 62763 1700 62805 1709
rect 62763 1660 62764 1700
rect 62804 1660 62805 1700
rect 62763 1651 62805 1660
rect 62668 1063 62708 1072
rect 62764 1112 62804 1651
rect 62764 1063 62804 1072
rect 62860 1112 62900 2332
rect 62956 2322 62996 2407
rect 63244 2129 63284 2584
rect 64012 2465 64052 4852
rect 64300 4808 64340 5104
rect 64396 4976 64436 5104
rect 64587 5104 64588 5144
rect 64628 5104 64629 5144
rect 64587 5095 64629 5104
rect 64971 5144 65013 5153
rect 64971 5104 64972 5144
rect 65012 5104 65013 5144
rect 64971 5095 65013 5104
rect 65068 5148 65108 5157
rect 64396 4927 64436 4936
rect 64108 4768 64340 4808
rect 64588 4808 64628 5095
rect 64875 4976 64917 4985
rect 64875 4936 64876 4976
rect 64916 4936 64917 4976
rect 64875 4927 64917 4936
rect 64972 4976 65012 4987
rect 64876 4842 64916 4927
rect 64972 4901 65012 4936
rect 64971 4892 65013 4901
rect 64971 4852 64972 4892
rect 65012 4852 65013 4892
rect 64971 4843 65013 4852
rect 64108 3464 64148 4768
rect 64588 4759 64628 4768
rect 64396 4724 64436 4733
rect 64204 4684 64396 4724
rect 64204 3632 64244 4684
rect 64396 4675 64436 4684
rect 64491 4304 64533 4313
rect 64491 4264 64492 4304
rect 64532 4264 64533 4304
rect 64491 4255 64533 4264
rect 64492 4136 64532 4255
rect 64492 4087 64532 4096
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 64876 3632 64916 3641
rect 65068 3632 65108 5108
rect 65356 5060 65396 5440
rect 65356 5011 65396 5020
rect 65548 4985 65588 5440
rect 65547 4976 65589 4985
rect 65547 4936 65548 4976
rect 65588 4936 65589 4976
rect 65547 4927 65589 4936
rect 65451 4892 65493 4901
rect 65451 4852 65452 4892
rect 65492 4852 65493 4892
rect 65451 4843 65493 4852
rect 65163 3968 65205 3977
rect 65163 3928 65164 3968
rect 65204 3928 65205 3968
rect 65163 3919 65205 3928
rect 64204 3592 64436 3632
rect 64300 3464 64340 3473
rect 64108 3424 64300 3464
rect 64300 2624 64340 3424
rect 64396 3380 64436 3592
rect 64684 3592 64876 3632
rect 64916 3592 65108 3632
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 64684 3464 64724 3592
rect 64876 3583 64916 3592
rect 64684 3415 64724 3424
rect 64972 3464 65012 3473
rect 65164 3464 65204 3919
rect 65012 3424 65204 3464
rect 65452 3464 65492 4843
rect 65644 4136 65684 5599
rect 65740 5153 65780 5608
rect 65836 5648 65876 5657
rect 65739 5144 65781 5153
rect 65739 5104 65740 5144
rect 65780 5104 65781 5144
rect 65739 5095 65781 5104
rect 65739 4976 65781 4985
rect 65739 4936 65740 4976
rect 65780 4936 65781 4976
rect 65739 4927 65781 4936
rect 65740 4842 65780 4927
rect 65836 4901 65876 5608
rect 65835 4892 65877 4901
rect 65835 4852 65836 4892
rect 65876 4852 65877 4892
rect 65835 4843 65877 4852
rect 65836 4388 65876 4843
rect 65836 4339 65876 4348
rect 66028 4220 66068 7792
rect 66123 7412 66165 7421
rect 66123 7372 66124 7412
rect 66164 7372 66165 7412
rect 66123 7363 66165 7372
rect 66124 7160 66164 7363
rect 66124 7111 66164 7120
rect 66124 6488 66164 6497
rect 66124 5825 66164 6448
rect 66123 5816 66165 5825
rect 66123 5776 66124 5816
rect 66164 5776 66165 5816
rect 66123 5767 66165 5776
rect 66316 5657 66356 7867
rect 66412 7866 66452 7951
rect 66508 7160 66548 7169
rect 66604 7160 66644 10219
rect 66699 8168 66741 8177
rect 66699 8128 66700 8168
rect 66740 8128 66741 8168
rect 66796 8168 66836 10807
rect 66892 8504 66932 11152
rect 67084 11108 67124 11647
rect 66988 11068 67124 11108
rect 66988 10184 67028 11068
rect 67180 11024 67220 11033
rect 67180 10352 67220 10984
rect 67372 10856 67412 11656
rect 67468 11612 67508 11621
rect 67660 11612 67700 11621
rect 67508 11572 67660 11612
rect 67468 11563 67508 11572
rect 67660 11563 67700 11572
rect 67563 11444 67605 11453
rect 67756 11444 67796 12496
rect 67852 12487 67892 12496
rect 67948 12536 67988 12571
rect 67948 12485 67988 12496
rect 68044 12536 68084 12547
rect 68044 12461 68084 12496
rect 68140 12536 68180 12940
rect 68043 12452 68085 12461
rect 68043 12412 68044 12452
rect 68084 12412 68085 12452
rect 68043 12403 68085 12412
rect 68140 12200 68180 12496
rect 67563 11404 67564 11444
rect 67604 11404 67605 11444
rect 67563 11395 67605 11404
rect 67660 11404 67796 11444
rect 67948 12160 68180 12200
rect 67467 11276 67509 11285
rect 67467 11236 67468 11276
rect 67508 11236 67509 11276
rect 67467 11227 67509 11236
rect 67180 10303 67220 10312
rect 67276 10816 67372 10856
rect 66988 10135 67028 10144
rect 67084 10268 67124 10277
rect 67084 9764 67124 10228
rect 67276 10268 67316 10816
rect 67372 10807 67412 10816
rect 67276 10219 67316 10228
rect 67372 10184 67412 10193
rect 67468 10184 67508 11227
rect 67564 10856 67604 11395
rect 67660 11024 67700 11404
rect 67851 11276 67893 11285
rect 67851 11227 67852 11276
rect 67892 11227 67893 11276
rect 67852 11141 67892 11210
rect 67660 10975 67700 10984
rect 67756 11024 67796 11033
rect 67948 11024 67988 12160
rect 68043 11696 68085 11705
rect 68043 11656 68044 11696
rect 68084 11656 68085 11696
rect 68043 11647 68085 11656
rect 68044 11562 68084 11647
rect 67796 10984 67988 11024
rect 67756 10975 67796 10984
rect 67564 10816 67700 10856
rect 67412 10144 67508 10184
rect 67372 10135 67412 10144
rect 67084 9724 67604 9764
rect 67564 9680 67604 9724
rect 67564 9631 67604 9640
rect 67371 9512 67413 9521
rect 67371 9472 67372 9512
rect 67412 9472 67413 9512
rect 67371 9463 67413 9472
rect 67468 9512 67508 9521
rect 67084 8672 67124 8681
rect 67372 8672 67412 9463
rect 67468 8681 67508 9472
rect 67660 9512 67700 10816
rect 68236 10520 68276 12991
rect 68332 11705 68372 13243
rect 68428 13217 68468 14008
rect 68427 13208 68469 13217
rect 68427 13168 68428 13208
rect 68468 13168 68469 13208
rect 68427 13159 68469 13168
rect 68428 12545 68468 13159
rect 68524 13133 68564 15100
rect 68619 14720 68661 14729
rect 68619 14680 68620 14720
rect 68660 14680 68661 14720
rect 68619 14671 68661 14680
rect 68620 14552 68660 14671
rect 68620 14503 68660 14512
rect 68619 13880 68661 13889
rect 68619 13840 68620 13880
rect 68660 13840 68661 13880
rect 68619 13831 68661 13840
rect 68620 13208 68660 13831
rect 68620 13159 68660 13168
rect 68523 13124 68565 13133
rect 68523 13084 68524 13124
rect 68564 13084 68565 13124
rect 68523 13075 68565 13084
rect 68716 12980 68756 16687
rect 68812 16493 68852 17032
rect 68811 16484 68853 16493
rect 68811 16444 68812 16484
rect 68852 16444 68853 16484
rect 68811 16435 68853 16444
rect 69100 14981 69140 17116
rect 69255 17072 69295 17472
rect 69545 17072 69585 17472
rect 69196 17032 69295 17072
rect 69388 17032 69585 17072
rect 69655 17072 69695 17472
rect 69945 17165 69985 17472
rect 70055 17165 70095 17472
rect 70345 17249 70385 17472
rect 70455 17333 70495 17472
rect 70454 17324 70496 17333
rect 70454 17284 70455 17324
rect 70495 17284 70496 17324
rect 70745 17300 70785 17472
rect 70855 17300 70895 17472
rect 70454 17275 70496 17284
rect 70732 17260 70785 17300
rect 70828 17260 70895 17300
rect 70344 17240 70386 17249
rect 70344 17200 70345 17240
rect 70385 17200 70386 17240
rect 70344 17191 70386 17200
rect 69944 17156 69986 17165
rect 69944 17116 69945 17156
rect 69985 17116 69986 17156
rect 69944 17107 69986 17116
rect 70054 17156 70096 17165
rect 70054 17116 70055 17156
rect 70095 17116 70096 17156
rect 70054 17107 70096 17116
rect 69655 17032 69812 17072
rect 69099 14972 69141 14981
rect 69099 14932 69100 14972
rect 69140 14932 69141 14972
rect 69099 14923 69141 14932
rect 69100 14729 69140 14814
rect 68812 14720 68852 14729
rect 68812 13805 68852 14680
rect 68908 14720 68948 14729
rect 68811 13796 68853 13805
rect 68811 13756 68812 13796
rect 68852 13756 68853 13796
rect 68811 13747 68853 13756
rect 68811 13628 68853 13637
rect 68811 13588 68812 13628
rect 68852 13588 68853 13628
rect 68811 13579 68853 13588
rect 68524 12940 68756 12980
rect 68427 12536 68469 12545
rect 68427 12496 68428 12536
rect 68468 12496 68469 12536
rect 68427 12487 68469 12496
rect 68331 11696 68373 11705
rect 68331 11656 68332 11696
rect 68372 11656 68373 11696
rect 68331 11647 68373 11656
rect 68140 10480 68276 10520
rect 67935 9523 67975 9532
rect 67660 9463 67700 9472
rect 67756 9512 67796 9521
rect 67796 9483 67935 9512
rect 67796 9472 67975 9483
rect 67659 9344 67701 9353
rect 67659 9304 67660 9344
rect 67700 9304 67701 9344
rect 67659 9295 67701 9304
rect 67124 8632 67412 8672
rect 67084 8623 67124 8632
rect 66892 8464 67124 8504
rect 66796 8128 66932 8168
rect 66699 8119 66741 8128
rect 66700 8034 66740 8119
rect 66795 8000 66837 8009
rect 66795 7960 66796 8000
rect 66836 7960 66837 8000
rect 66795 7951 66837 7960
rect 66796 7866 66836 7951
rect 66548 7120 66644 7160
rect 66508 7111 66548 7120
rect 66892 6749 66932 8128
rect 66891 6740 66933 6749
rect 66891 6700 66892 6740
rect 66932 6700 66933 6740
rect 66891 6691 66933 6700
rect 66603 6488 66645 6497
rect 66603 6448 66604 6488
rect 66644 6448 66645 6488
rect 66603 6439 66645 6448
rect 66315 5648 66357 5657
rect 66315 5608 66316 5648
rect 66356 5608 66357 5648
rect 66315 5599 66357 5608
rect 66604 4976 66644 6439
rect 66604 4313 66644 4936
rect 66795 4976 66837 4985
rect 66795 4936 66796 4976
rect 66836 4936 66837 4976
rect 66795 4927 66837 4936
rect 66603 4304 66645 4313
rect 66603 4264 66604 4304
rect 66644 4264 66645 4304
rect 66603 4255 66645 4264
rect 66028 4171 66068 4180
rect 66123 4220 66165 4229
rect 66123 4180 66124 4220
rect 66164 4180 66165 4220
rect 66123 4171 66165 4180
rect 65644 4096 65780 4136
rect 65643 3968 65685 3977
rect 65643 3928 65644 3968
rect 65684 3928 65685 3968
rect 65643 3919 65685 3928
rect 65644 3834 65684 3919
rect 65740 3716 65780 4096
rect 65644 3676 65780 3716
rect 65547 3632 65589 3641
rect 65547 3592 65548 3632
rect 65588 3592 65589 3632
rect 65547 3583 65589 3592
rect 64396 3331 64436 3340
rect 64588 3380 64628 3415
rect 64588 3329 64628 3340
rect 64491 3296 64533 3305
rect 64491 3256 64492 3296
rect 64532 3256 64533 3296
rect 64491 3247 64533 3256
rect 64492 3162 64532 3247
rect 64972 2900 65012 3424
rect 64780 2860 65012 2900
rect 65452 2900 65492 3424
rect 65548 3464 65588 3583
rect 65644 3557 65684 3676
rect 65643 3548 65685 3557
rect 65643 3508 65644 3548
rect 65684 3508 65685 3548
rect 65643 3499 65685 3508
rect 65548 3415 65588 3424
rect 65644 3464 65684 3499
rect 65644 3414 65684 3424
rect 65740 3464 65780 3473
rect 65452 2860 65684 2900
rect 64491 2708 64533 2717
rect 64491 2668 64492 2708
rect 64532 2668 64533 2708
rect 64491 2659 64533 2668
rect 64395 2624 64437 2633
rect 64300 2584 64396 2624
rect 64436 2584 64437 2624
rect 64395 2575 64437 2584
rect 64396 2490 64436 2575
rect 64492 2540 64532 2659
rect 64492 2491 64532 2500
rect 64588 2624 64628 2633
rect 64588 2465 64628 2584
rect 64684 2624 64724 2633
rect 64780 2624 64820 2860
rect 65068 2792 65108 2801
rect 64971 2708 65013 2717
rect 64971 2668 64972 2708
rect 65012 2668 65013 2708
rect 64971 2659 65013 2668
rect 64724 2584 64820 2624
rect 64875 2624 64917 2633
rect 64875 2584 64876 2624
rect 64916 2584 64917 2624
rect 64684 2575 64724 2584
rect 64875 2575 64917 2584
rect 64876 2490 64916 2575
rect 64972 2574 65012 2659
rect 64011 2456 64053 2465
rect 64011 2416 64012 2456
rect 64052 2416 64053 2456
rect 64011 2407 64053 2416
rect 64587 2456 64629 2465
rect 64587 2416 64588 2456
rect 64628 2416 64629 2456
rect 64587 2407 64629 2416
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 63243 2120 63285 2129
rect 63243 2080 63244 2120
rect 63284 2080 63285 2120
rect 63243 2071 63285 2080
rect 64779 2120 64821 2129
rect 64779 2080 64780 2120
rect 64820 2080 64821 2120
rect 64779 2071 64821 2080
rect 63244 1709 63284 2071
rect 64780 1986 64820 2071
rect 64972 2036 65012 2045
rect 65068 2036 65108 2752
rect 65163 2708 65205 2717
rect 65163 2668 65164 2708
rect 65204 2668 65205 2708
rect 65163 2659 65205 2668
rect 65164 2574 65204 2659
rect 65260 2624 65300 2633
rect 65644 2624 65684 2860
rect 65300 2584 65588 2624
rect 65260 2575 65300 2584
rect 65012 1996 65108 2036
rect 65548 2398 65588 2584
rect 65644 2575 65684 2584
rect 65740 2624 65780 3424
rect 65931 3464 65973 3473
rect 65931 3424 65932 3464
rect 65972 3424 65973 3464
rect 65931 3415 65973 3424
rect 66028 3464 66068 3473
rect 65932 3330 65972 3415
rect 66028 2792 66068 3424
rect 66124 3464 66164 4171
rect 66219 3548 66261 3557
rect 66219 3508 66220 3548
rect 66260 3508 66261 3548
rect 66219 3499 66261 3508
rect 66124 3415 66164 3424
rect 66220 3464 66260 3499
rect 66220 3413 66260 3424
rect 66411 3464 66453 3473
rect 66411 3424 66412 3464
rect 66452 3424 66453 3464
rect 66411 3415 66453 3424
rect 66796 3464 66836 4927
rect 66796 3415 66836 3424
rect 66412 3330 66452 3415
rect 67084 2900 67124 8464
rect 67372 7160 67412 8632
rect 67467 8672 67509 8681
rect 67467 8632 67468 8672
rect 67508 8632 67509 8672
rect 67467 8623 67509 8632
rect 67372 7111 67412 7120
rect 67660 3641 67700 9295
rect 67756 8933 67796 9472
rect 68140 9428 68180 10480
rect 68331 10436 68373 10445
rect 68331 10396 68332 10436
rect 68372 10396 68373 10436
rect 68331 10387 68373 10396
rect 68235 10352 68277 10361
rect 68235 10312 68236 10352
rect 68276 10312 68277 10352
rect 68235 10303 68277 10312
rect 68236 10184 68276 10303
rect 68236 10135 68276 10144
rect 68332 10184 68372 10387
rect 68524 10361 68564 12940
rect 68619 12704 68661 12713
rect 68619 12664 68620 12704
rect 68660 12664 68661 12704
rect 68619 12655 68661 12664
rect 68620 10604 68660 12655
rect 68812 12461 68852 13579
rect 68908 13133 68948 14680
rect 69099 14720 69141 14729
rect 69099 14680 69100 14720
rect 69140 14680 69141 14720
rect 69099 14671 69141 14680
rect 69004 14552 69044 14561
rect 69004 13973 69044 14512
rect 69003 13964 69045 13973
rect 69003 13924 69004 13964
rect 69044 13924 69045 13964
rect 69003 13915 69045 13924
rect 69003 13292 69045 13301
rect 69003 13252 69004 13292
rect 69044 13252 69045 13292
rect 69003 13243 69045 13252
rect 69004 13208 69044 13243
rect 69004 13157 69044 13168
rect 68907 13124 68949 13133
rect 68907 13084 68908 13124
rect 68948 13084 68949 13124
rect 68907 13075 68949 13084
rect 69196 12797 69236 17032
rect 69291 16484 69333 16493
rect 69291 16444 69292 16484
rect 69332 16444 69333 16484
rect 69291 16435 69333 16444
rect 69292 16350 69332 16435
rect 69291 16064 69333 16073
rect 69291 16024 69292 16064
rect 69332 16024 69333 16064
rect 69291 16015 69333 16024
rect 69292 15930 69332 16015
rect 69291 14804 69333 14813
rect 69291 14764 69292 14804
rect 69332 14764 69333 14804
rect 69291 14755 69333 14764
rect 69292 14670 69332 14755
rect 69388 12980 69428 17032
rect 69580 16232 69620 16243
rect 69580 16157 69620 16192
rect 69675 16232 69717 16241
rect 69675 16192 69676 16232
rect 69716 16192 69717 16232
rect 69675 16183 69717 16192
rect 69579 16148 69621 16157
rect 69579 16108 69580 16148
rect 69620 16108 69621 16148
rect 69579 16099 69621 16108
rect 69676 16098 69716 16183
rect 69484 15476 69524 15485
rect 69484 14981 69524 15436
rect 69676 15317 69716 15402
rect 69675 15308 69717 15317
rect 69675 15268 69676 15308
rect 69716 15268 69717 15308
rect 69675 15259 69717 15268
rect 69772 15056 69812 17032
rect 69963 16988 70005 16997
rect 69963 16948 69964 16988
rect 70004 16948 70005 16988
rect 69963 16939 70005 16948
rect 69964 16484 70004 16939
rect 70732 16829 70772 17260
rect 70731 16820 70773 16829
rect 70731 16780 70732 16820
rect 70772 16780 70773 16820
rect 70731 16771 70773 16780
rect 70828 16661 70868 17260
rect 71145 17072 71185 17472
rect 71255 17165 71295 17472
rect 71545 17333 71585 17472
rect 71545 17324 71589 17333
rect 71545 17284 71548 17324
rect 71588 17284 71589 17324
rect 71547 17275 71589 17284
rect 71254 17156 71296 17165
rect 71254 17116 71255 17156
rect 71295 17116 71296 17156
rect 71254 17107 71296 17116
rect 71655 17072 71695 17472
rect 71945 17072 71985 17472
rect 72055 17165 72095 17472
rect 72054 17156 72096 17165
rect 72054 17116 72055 17156
rect 72095 17116 72096 17156
rect 72054 17107 72096 17116
rect 71116 17032 71185 17072
rect 71596 17032 71695 17072
rect 71884 17032 71985 17072
rect 72345 17072 72385 17472
rect 72455 17240 72495 17472
rect 72745 17300 72785 17472
rect 72855 17300 72895 17472
rect 73145 17300 73185 17472
rect 72652 17260 72785 17300
rect 72844 17260 72895 17300
rect 73132 17260 73185 17300
rect 72455 17200 72596 17240
rect 72345 17032 72404 17072
rect 70827 16652 70869 16661
rect 70827 16612 70828 16652
rect 70868 16612 70869 16652
rect 70827 16603 70869 16612
rect 69964 16435 70004 16444
rect 70348 16316 70388 16325
rect 69867 16232 69909 16241
rect 69867 16192 69868 16232
rect 69908 16192 69909 16232
rect 69867 16183 69909 16192
rect 69868 16098 69908 16183
rect 69964 16064 70004 16073
rect 69964 15905 70004 16024
rect 70156 16064 70196 16073
rect 69963 15896 70005 15905
rect 69963 15856 69964 15896
rect 70004 15856 70005 15896
rect 69963 15847 70005 15856
rect 69867 15728 69909 15737
rect 69867 15688 69868 15728
rect 69908 15688 69909 15728
rect 69867 15679 69909 15688
rect 69868 15594 69908 15679
rect 69676 15016 69812 15056
rect 69964 15560 70004 15569
rect 69483 14972 69525 14981
rect 69483 14932 69484 14972
rect 69524 14932 69525 14972
rect 69483 14923 69525 14932
rect 69483 14552 69525 14561
rect 69483 14512 69484 14552
rect 69524 14512 69525 14552
rect 69483 14503 69525 14512
rect 69292 12940 69428 12980
rect 69484 12956 69524 14503
rect 69579 13796 69621 13805
rect 69579 13756 69580 13796
rect 69620 13756 69621 13796
rect 69579 13747 69621 13756
rect 69580 13662 69620 13747
rect 69195 12788 69237 12797
rect 69195 12748 69196 12788
rect 69236 12748 69237 12788
rect 69195 12739 69237 12748
rect 68907 12536 68949 12545
rect 68907 12496 68908 12536
rect 68948 12496 68949 12536
rect 68907 12487 68949 12496
rect 68811 12452 68853 12461
rect 68811 12412 68812 12452
rect 68852 12412 68853 12452
rect 68811 12403 68853 12412
rect 68908 11696 68948 12487
rect 68908 11647 68948 11656
rect 68907 10940 68949 10949
rect 68907 10900 68908 10940
rect 68948 10900 68949 10940
rect 68907 10891 68949 10900
rect 68908 10806 68948 10891
rect 68716 10772 68756 10781
rect 68756 10732 68852 10772
rect 68716 10723 68756 10732
rect 68620 10564 68756 10604
rect 68523 10352 68565 10361
rect 68523 10312 68524 10352
rect 68564 10312 68565 10352
rect 68523 10303 68565 10312
rect 68428 10226 68468 10235
rect 68468 10186 68660 10226
rect 68428 10177 68468 10186
rect 68332 10135 68372 10144
rect 68427 10100 68469 10109
rect 68427 10060 68428 10100
rect 68468 10060 68469 10100
rect 68427 10051 68469 10060
rect 68235 10016 68277 10025
rect 68235 9976 68236 10016
rect 68276 9976 68277 10016
rect 68235 9967 68277 9976
rect 68236 9596 68276 9967
rect 68236 9547 68276 9556
rect 67852 9388 68180 9428
rect 67755 8924 67797 8933
rect 67755 8884 67756 8924
rect 67796 8884 67797 8924
rect 67755 8875 67797 8884
rect 67755 5144 67797 5153
rect 67755 5104 67756 5144
rect 67796 5104 67797 5144
rect 67755 5095 67797 5104
rect 67756 5010 67796 5095
rect 67659 3632 67701 3641
rect 67659 3592 67660 3632
rect 67700 3592 67701 3632
rect 67659 3583 67701 3592
rect 66892 2876 67124 2900
rect 66028 2717 66068 2752
rect 66796 2860 67124 2876
rect 67660 3464 67700 3473
rect 67660 2900 67700 3424
rect 67852 2900 67892 9388
rect 68044 9260 68084 9269
rect 67948 8672 67988 8683
rect 67948 8597 67988 8632
rect 67947 8588 67989 8597
rect 67947 8548 67948 8588
rect 67988 8548 67989 8588
rect 67947 8539 67989 8548
rect 68044 8345 68084 9220
rect 68332 8588 68372 8597
rect 68140 8548 68332 8588
rect 68043 8336 68085 8345
rect 67948 8296 68044 8336
rect 68084 8296 68085 8336
rect 67948 8000 67988 8296
rect 68043 8287 68085 8296
rect 68044 8202 68084 8287
rect 67948 7951 67988 7960
rect 68043 7916 68085 7925
rect 68043 7876 68044 7916
rect 68084 7876 68085 7916
rect 68043 7867 68085 7876
rect 68044 7782 68084 7867
rect 68140 7832 68180 8548
rect 68332 8539 68372 8548
rect 68428 8009 68468 10051
rect 68523 10016 68565 10025
rect 68523 9976 68524 10016
rect 68564 9976 68565 10016
rect 68523 9967 68565 9976
rect 68524 9882 68564 9967
rect 68620 9764 68660 10186
rect 68524 9724 68660 9764
rect 68524 8924 68564 9724
rect 68619 9596 68661 9605
rect 68619 9556 68620 9596
rect 68660 9556 68661 9596
rect 68619 9547 68661 9556
rect 68620 9512 68660 9547
rect 68620 9461 68660 9472
rect 68716 9344 68756 10564
rect 68812 9605 68852 10732
rect 69292 10529 69332 12940
rect 69474 12916 69524 12956
rect 69387 12872 69429 12881
rect 69474 12872 69514 12916
rect 69387 12832 69388 12872
rect 69428 12832 69514 12872
rect 69387 12823 69429 12832
rect 69291 10520 69333 10529
rect 69291 10480 69292 10520
rect 69332 10480 69333 10520
rect 69291 10471 69333 10480
rect 68907 10352 68949 10361
rect 68907 10312 68908 10352
rect 68948 10312 68949 10352
rect 68907 10303 68949 10312
rect 69291 10352 69333 10361
rect 69291 10312 69292 10352
rect 69332 10312 69333 10352
rect 69291 10303 69333 10312
rect 68811 9596 68853 9605
rect 68811 9556 68812 9596
rect 68852 9556 68853 9596
rect 68811 9547 68853 9556
rect 68332 8000 68372 8009
rect 68140 7783 68180 7792
rect 68236 7916 68276 7925
rect 68139 7664 68181 7673
rect 68139 7624 68140 7664
rect 68180 7624 68181 7664
rect 68139 7615 68181 7624
rect 68140 6509 68180 7615
rect 68236 6656 68276 7876
rect 68332 7757 68372 7960
rect 68427 8000 68469 8009
rect 68427 7960 68428 8000
rect 68468 7960 68469 8000
rect 68427 7951 68469 7960
rect 68331 7748 68373 7757
rect 68331 7708 68332 7748
rect 68372 7708 68373 7748
rect 68331 7699 68373 7708
rect 68428 7412 68468 7951
rect 68524 7925 68564 8884
rect 68620 9304 68756 9344
rect 68523 7916 68565 7925
rect 68523 7876 68524 7916
rect 68564 7876 68565 7916
rect 68523 7867 68565 7876
rect 68620 7673 68660 9304
rect 68811 9008 68853 9017
rect 68811 8968 68812 9008
rect 68852 8968 68853 9008
rect 68811 8959 68853 8968
rect 68812 8672 68852 8959
rect 68908 8681 68948 10303
rect 69099 10268 69141 10277
rect 69099 10228 69100 10268
rect 69140 10228 69141 10268
rect 69099 10219 69141 10228
rect 69100 10184 69140 10219
rect 69004 10016 69044 10025
rect 69004 9017 69044 9976
rect 69003 9008 69045 9017
rect 69003 8968 69004 9008
rect 69044 8968 69045 9008
rect 69003 8959 69045 8968
rect 68812 8623 68852 8632
rect 68907 8672 68949 8681
rect 68907 8632 68908 8672
rect 68948 8632 68949 8672
rect 69100 8672 69140 10144
rect 69195 10184 69237 10193
rect 69195 10144 69196 10184
rect 69236 10144 69237 10184
rect 69195 10135 69237 10144
rect 69292 10184 69332 10303
rect 69292 10135 69332 10144
rect 69196 10050 69236 10135
rect 69388 8756 69428 12823
rect 69483 12620 69525 12629
rect 69483 12580 69484 12620
rect 69524 12580 69525 12620
rect 69483 12571 69525 12580
rect 69484 12486 69524 12571
rect 69483 11612 69525 11621
rect 69483 11572 69484 11612
rect 69524 11572 69525 11612
rect 69483 11563 69525 11572
rect 69484 10268 69524 11563
rect 69676 10613 69716 15016
rect 69964 14888 70004 15520
rect 70059 15560 70101 15569
rect 70059 15520 70060 15560
rect 70100 15520 70101 15560
rect 70059 15511 70101 15520
rect 70156 15560 70196 16024
rect 70348 15905 70388 16276
rect 70732 16316 70772 16325
rect 70540 16064 70580 16073
rect 70732 16064 70772 16276
rect 70923 16316 70965 16325
rect 70923 16276 70924 16316
rect 70964 16276 70965 16316
rect 70923 16267 70965 16276
rect 70924 16182 70964 16267
rect 71116 16241 71156 17032
rect 71596 16409 71636 17032
rect 71595 16400 71637 16409
rect 71595 16360 71596 16400
rect 71636 16360 71637 16400
rect 71595 16351 71637 16360
rect 71787 16400 71829 16409
rect 71787 16360 71788 16400
rect 71828 16360 71829 16400
rect 71787 16351 71829 16360
rect 71788 16266 71828 16351
rect 71115 16232 71157 16241
rect 71115 16192 71116 16232
rect 71156 16192 71157 16232
rect 71115 16183 71157 16192
rect 71116 16064 71156 16073
rect 70732 16024 71116 16064
rect 70347 15896 70389 15905
rect 70347 15856 70348 15896
rect 70388 15856 70389 15896
rect 70347 15847 70389 15856
rect 70251 15812 70293 15821
rect 70251 15772 70252 15812
rect 70292 15772 70293 15812
rect 70251 15763 70293 15772
rect 70060 15426 70100 15511
rect 70156 14897 70196 15520
rect 70060 14888 70100 14897
rect 69964 14848 70060 14888
rect 69771 14720 69813 14729
rect 69771 14680 69772 14720
rect 69812 14680 69813 14720
rect 69771 14671 69813 14680
rect 69772 14141 69812 14671
rect 69771 14132 69813 14141
rect 69771 14092 69772 14132
rect 69812 14092 69813 14132
rect 69771 14083 69813 14092
rect 69772 14048 69812 14083
rect 69772 13997 69812 14008
rect 69867 13964 69909 13973
rect 69867 13924 69868 13964
rect 69908 13924 69909 13964
rect 69867 13915 69909 13924
rect 70060 13964 70100 14848
rect 70155 14888 70197 14897
rect 70155 14848 70156 14888
rect 70196 14848 70197 14888
rect 70155 14839 70197 14848
rect 70155 14048 70197 14057
rect 70155 14008 70156 14048
rect 70196 14008 70197 14048
rect 70155 13999 70197 14008
rect 70060 13915 70100 13924
rect 69868 13830 69908 13915
rect 70156 13914 70196 13999
rect 69963 13880 70005 13889
rect 69963 13840 69964 13880
rect 70004 13840 70005 13880
rect 69963 13831 70005 13840
rect 69964 13746 70004 13831
rect 70155 13796 70197 13805
rect 70155 13756 70156 13796
rect 70196 13756 70197 13796
rect 70155 13747 70197 13756
rect 69963 13292 70005 13301
rect 69963 13252 69964 13292
rect 70004 13252 70005 13292
rect 69963 13243 70005 13252
rect 69867 13208 69909 13217
rect 69867 13168 69868 13208
rect 69908 13168 69909 13208
rect 69867 13159 69909 13168
rect 69868 13074 69908 13159
rect 69964 12980 70004 13243
rect 69868 12940 70004 12980
rect 69868 12536 69908 12940
rect 69868 12487 69908 12496
rect 70059 12452 70101 12461
rect 70059 12412 70060 12452
rect 70100 12412 70101 12452
rect 70059 12403 70101 12412
rect 70060 11948 70100 12403
rect 70060 11899 70100 11908
rect 69963 11024 70005 11033
rect 69963 10984 69964 11024
rect 70004 10984 70005 11024
rect 69963 10975 70005 10984
rect 69964 10890 70004 10975
rect 69675 10604 69717 10613
rect 69675 10564 69676 10604
rect 69716 10564 69717 10604
rect 69675 10555 69717 10564
rect 70059 10520 70101 10529
rect 70059 10480 70060 10520
rect 70100 10480 70101 10520
rect 70059 10471 70101 10480
rect 70060 10436 70100 10471
rect 70060 10277 70100 10396
rect 69484 10219 69524 10228
rect 69868 10268 69908 10277
rect 69676 10016 69716 10025
rect 69868 10016 69908 10228
rect 70059 10268 70101 10277
rect 70059 10228 70060 10268
rect 70100 10228 70101 10268
rect 70059 10219 70101 10228
rect 69716 9976 69908 10016
rect 69676 9967 69716 9976
rect 69483 9512 69525 9521
rect 69483 9472 69484 9512
rect 69524 9472 69525 9512
rect 69483 9463 69525 9472
rect 69484 9378 69524 9463
rect 69868 8849 69908 9976
rect 69867 8840 69909 8849
rect 69867 8800 69868 8840
rect 69908 8800 69909 8840
rect 69867 8791 69909 8800
rect 69388 8707 69428 8716
rect 69675 8756 69717 8765
rect 69675 8716 69676 8756
rect 69716 8716 69717 8756
rect 69675 8707 69717 8716
rect 69100 8632 69332 8672
rect 68907 8623 68949 8632
rect 68908 8538 68948 8623
rect 69196 8504 69236 8513
rect 69100 8464 69196 8504
rect 69004 8446 69044 8455
rect 69004 8345 69044 8406
rect 69003 8336 69045 8345
rect 69003 8296 69004 8336
rect 69044 8296 69045 8336
rect 69003 8287 69045 8296
rect 68907 8252 68949 8261
rect 68907 8212 68908 8252
rect 68948 8212 68949 8252
rect 68907 8203 68949 8212
rect 68908 7916 68948 8203
rect 68908 7867 68948 7876
rect 69100 7916 69140 8464
rect 69196 8455 69236 8464
rect 69292 7916 69332 8632
rect 69676 8622 69716 8707
rect 70156 8177 70196 13747
rect 70252 11621 70292 15763
rect 70347 15728 70389 15737
rect 70347 15688 70348 15728
rect 70388 15688 70389 15728
rect 70347 15679 70389 15688
rect 70348 15644 70388 15679
rect 70540 15644 70580 16024
rect 70540 15604 70676 15644
rect 70348 15593 70388 15604
rect 70636 15560 70676 15604
rect 70732 15560 70772 15569
rect 70636 15520 70732 15560
rect 70443 15308 70485 15317
rect 70443 15268 70444 15308
rect 70484 15268 70485 15308
rect 70443 15259 70485 15268
rect 70347 14720 70389 14729
rect 70347 14680 70348 14720
rect 70388 14680 70389 14720
rect 70347 14671 70389 14680
rect 70444 14720 70484 15259
rect 70348 14586 70388 14671
rect 70444 14645 70484 14680
rect 70443 14636 70485 14645
rect 70443 14596 70444 14636
rect 70484 14596 70485 14636
rect 70443 14587 70485 14596
rect 70540 14494 70580 14503
rect 70347 14384 70389 14393
rect 70347 14344 70348 14384
rect 70388 14344 70389 14384
rect 70347 14335 70389 14344
rect 70348 13301 70388 14335
rect 70540 14216 70580 14454
rect 70636 14393 70676 15520
rect 70732 15511 70772 15520
rect 70827 15224 70869 15233
rect 70827 15184 70828 15224
rect 70868 15184 70869 15224
rect 70827 15175 70869 15184
rect 70731 14804 70773 14813
rect 70731 14764 70732 14804
rect 70772 14764 70773 14804
rect 70731 14755 70773 14764
rect 70732 14670 70772 14755
rect 70635 14384 70677 14393
rect 70635 14344 70636 14384
rect 70676 14344 70677 14384
rect 70635 14335 70677 14344
rect 70540 14057 70580 14176
rect 70539 14048 70581 14057
rect 70539 14008 70540 14048
rect 70580 14008 70581 14048
rect 70539 13999 70581 14008
rect 70636 14048 70676 14057
rect 70539 13880 70581 13889
rect 70539 13840 70540 13880
rect 70580 13840 70581 13880
rect 70539 13831 70581 13840
rect 70347 13292 70389 13301
rect 70347 13252 70348 13292
rect 70388 13252 70389 13292
rect 70347 13243 70389 13252
rect 70251 11612 70293 11621
rect 70251 11572 70252 11612
rect 70292 11572 70293 11612
rect 70251 11563 70293 11572
rect 70348 11024 70388 13243
rect 70443 11360 70485 11369
rect 70443 11320 70444 11360
rect 70484 11320 70485 11360
rect 70443 11311 70485 11320
rect 70348 10975 70388 10984
rect 70347 10436 70389 10445
rect 70444 10436 70484 11311
rect 70347 10396 70348 10436
rect 70388 10396 70484 10436
rect 70347 10387 70389 10396
rect 70348 10302 70388 10387
rect 70251 10184 70293 10193
rect 70540 10184 70580 13831
rect 70636 13637 70676 14008
rect 70828 13889 70868 15175
rect 71116 14981 71156 16024
rect 71307 15728 71349 15737
rect 71307 15688 71308 15728
rect 71348 15688 71349 15728
rect 71307 15679 71349 15688
rect 70923 14972 70965 14981
rect 70923 14932 70924 14972
rect 70964 14932 70965 14972
rect 70923 14923 70965 14932
rect 71115 14972 71157 14981
rect 71115 14932 71116 14972
rect 71156 14932 71157 14972
rect 71115 14923 71157 14932
rect 70924 14838 70964 14923
rect 71211 14888 71253 14897
rect 71211 14848 71212 14888
rect 71252 14848 71253 14888
rect 71211 14839 71253 14848
rect 71115 14720 71157 14729
rect 71115 14680 71116 14720
rect 71156 14680 71157 14720
rect 71115 14671 71157 14680
rect 71212 14720 71252 14839
rect 71212 14671 71252 14680
rect 71308 14720 71348 15679
rect 71596 15560 71636 15569
rect 71308 14671 71348 14680
rect 71404 14720 71444 14731
rect 71116 14586 71156 14671
rect 71404 14645 71444 14680
rect 71403 14636 71445 14645
rect 71403 14596 71404 14636
rect 71444 14596 71445 14636
rect 71403 14587 71445 14596
rect 70923 14552 70965 14561
rect 70923 14512 70924 14552
rect 70964 14512 70965 14552
rect 70923 14503 70965 14512
rect 70924 14418 70964 14503
rect 71020 14176 71540 14216
rect 70923 14132 70965 14141
rect 70923 14092 70924 14132
rect 70964 14092 70965 14132
rect 70923 14083 70965 14092
rect 70924 14048 70964 14083
rect 70924 13997 70964 14008
rect 71020 13964 71060 14176
rect 71308 14048 71348 14057
rect 71020 13915 71060 13924
rect 71211 13964 71253 13973
rect 71211 13924 71212 13964
rect 71252 13924 71253 13964
rect 71211 13915 71253 13924
rect 70827 13880 70869 13889
rect 70827 13840 70828 13880
rect 70868 13840 70869 13880
rect 70827 13831 70869 13840
rect 71116 13880 71156 13889
rect 70923 13796 70965 13805
rect 70923 13756 70924 13796
rect 70964 13756 70965 13796
rect 70923 13747 70965 13756
rect 70635 13628 70677 13637
rect 70635 13588 70636 13628
rect 70676 13588 70677 13628
rect 70635 13579 70677 13588
rect 70635 13376 70677 13385
rect 70635 13336 70636 13376
rect 70676 13336 70677 13376
rect 70635 13327 70677 13336
rect 70636 12629 70676 13327
rect 70731 13208 70773 13217
rect 70731 13168 70732 13208
rect 70772 13168 70773 13208
rect 70731 13159 70773 13168
rect 70635 12620 70677 12629
rect 70635 12580 70636 12620
rect 70676 12580 70677 12620
rect 70635 12571 70677 12580
rect 70732 12536 70772 13159
rect 70732 12487 70772 12496
rect 70251 10144 70252 10184
rect 70292 10144 70580 10184
rect 70251 10135 70293 10144
rect 70252 10050 70292 10135
rect 70540 9680 70580 10144
rect 70636 9680 70676 9689
rect 70540 9640 70636 9680
rect 70636 9631 70676 9640
rect 70443 9596 70485 9605
rect 70443 9556 70444 9596
rect 70484 9556 70485 9596
rect 70443 9547 70485 9556
rect 70444 8933 70484 9547
rect 70539 9512 70581 9521
rect 70539 9472 70540 9512
rect 70580 9472 70581 9512
rect 70539 9463 70581 9472
rect 70443 8924 70485 8933
rect 70443 8884 70444 8924
rect 70484 8884 70485 8924
rect 70443 8875 70485 8884
rect 70155 8168 70197 8177
rect 70155 8128 70156 8168
rect 70196 8128 70197 8168
rect 70155 8119 70197 8128
rect 69100 7841 69140 7876
rect 69196 7876 69332 7916
rect 69099 7832 69141 7841
rect 69004 7792 69100 7832
rect 69140 7792 69141 7832
rect 68716 7748 68756 7757
rect 68619 7664 68661 7673
rect 68619 7624 68620 7664
rect 68660 7624 68661 7664
rect 68619 7615 68661 7624
rect 68716 7589 68756 7708
rect 68715 7580 68757 7589
rect 68715 7540 68716 7580
rect 68756 7540 68757 7580
rect 68715 7531 68757 7540
rect 68524 7412 68564 7421
rect 68428 7372 68524 7412
rect 68524 7363 68564 7372
rect 68908 7244 68948 7253
rect 69004 7244 69044 7792
rect 69099 7783 69141 7792
rect 69196 7664 69236 7876
rect 69291 7748 69333 7757
rect 69291 7708 69292 7748
rect 69332 7708 69333 7748
rect 69291 7699 69333 7708
rect 68948 7204 69044 7244
rect 69100 7624 69236 7664
rect 68908 7195 68948 7204
rect 68716 6992 68756 7001
rect 68236 6616 68372 6656
rect 67947 6488 67989 6497
rect 67947 6448 67948 6488
rect 67988 6448 67989 6488
rect 67947 6439 67989 6448
rect 68044 6488 68084 6497
rect 68140 6460 68180 6469
rect 68236 6488 68276 6497
rect 67948 6354 67988 6439
rect 68044 5396 68084 6448
rect 68139 6320 68181 6329
rect 68236 6320 68276 6448
rect 68139 6280 68140 6320
rect 68180 6280 68276 6320
rect 68139 6271 68181 6280
rect 68332 5900 68372 6616
rect 68427 6488 68469 6497
rect 68427 6448 68428 6488
rect 68468 6448 68469 6488
rect 68427 6439 68469 6448
rect 68428 6354 68468 6439
rect 68236 5860 68372 5900
rect 68139 5732 68181 5741
rect 68139 5692 68140 5732
rect 68180 5692 68181 5732
rect 68139 5683 68181 5692
rect 68140 5648 68180 5683
rect 68140 5597 68180 5608
rect 68236 5564 68276 5860
rect 68620 5816 68660 5825
rect 68332 5648 68372 5659
rect 68332 5573 68372 5608
rect 68427 5648 68469 5657
rect 68427 5608 68428 5648
rect 68468 5608 68469 5648
rect 68427 5599 68469 5608
rect 68236 5515 68276 5524
rect 68331 5564 68373 5573
rect 68331 5524 68332 5564
rect 68372 5524 68373 5564
rect 68331 5515 68373 5524
rect 68428 5514 68468 5599
rect 68620 5396 68660 5776
rect 68716 5741 68756 6952
rect 68812 6488 68852 6499
rect 68812 6413 68852 6448
rect 68811 6404 68853 6413
rect 68811 6364 68812 6404
rect 68852 6364 68853 6404
rect 68811 6355 68853 6364
rect 69100 6329 69140 7624
rect 69292 7614 69332 7699
rect 70444 7160 70484 8875
rect 70060 7076 70100 7085
rect 69579 6656 69621 6665
rect 69579 6616 69580 6656
rect 69620 6616 69621 6656
rect 69579 6607 69621 6616
rect 69099 6320 69141 6329
rect 69099 6280 69100 6320
rect 69140 6280 69141 6320
rect 69099 6271 69141 6280
rect 69100 5984 69140 6271
rect 69100 5944 69524 5984
rect 68907 5816 68949 5825
rect 68907 5776 68908 5816
rect 68948 5776 68949 5816
rect 68907 5767 68949 5776
rect 69387 5816 69429 5825
rect 69387 5776 69388 5816
rect 69428 5776 69429 5816
rect 69387 5767 69429 5776
rect 68715 5732 68757 5741
rect 68715 5692 68716 5732
rect 68756 5692 68757 5732
rect 68715 5683 68757 5692
rect 68044 5356 68660 5396
rect 67948 4976 67988 4985
rect 67948 4640 67988 4936
rect 68331 4976 68373 4985
rect 68331 4936 68332 4976
rect 68372 4936 68373 4976
rect 68331 4927 68373 4936
rect 68332 4842 68372 4927
rect 67948 4600 68564 4640
rect 68427 4472 68469 4481
rect 68427 4432 68428 4472
rect 68468 4432 68469 4472
rect 68427 4423 68469 4432
rect 68428 4220 68468 4423
rect 68524 4304 68564 4600
rect 68620 4481 68660 5356
rect 68619 4472 68661 4481
rect 68619 4432 68620 4472
rect 68660 4432 68661 4472
rect 68619 4423 68661 4432
rect 68524 4255 68564 4264
rect 68428 4171 68468 4180
rect 68620 4220 68660 4229
rect 68331 4136 68373 4145
rect 68331 4096 68332 4136
rect 68372 4096 68373 4136
rect 68331 4087 68373 4096
rect 68332 4002 68372 4087
rect 67660 2860 67796 2900
rect 67852 2860 68372 2900
rect 66796 2836 66932 2860
rect 66796 2717 66836 2836
rect 66027 2708 66069 2717
rect 66027 2668 66028 2708
rect 66068 2668 66069 2708
rect 66027 2659 66069 2668
rect 66219 2708 66261 2717
rect 66219 2668 66220 2708
rect 66260 2668 66261 2708
rect 66219 2659 66261 2668
rect 66795 2708 66837 2717
rect 66795 2668 66796 2708
rect 66836 2668 66837 2708
rect 66795 2659 66837 2668
rect 65740 2575 65780 2584
rect 64972 1987 65012 1996
rect 63627 1952 63669 1961
rect 63627 1912 63628 1952
rect 63668 1912 63669 1952
rect 63627 1903 63669 1912
rect 65355 1952 65397 1961
rect 65355 1912 65356 1952
rect 65396 1912 65397 1952
rect 65355 1903 65397 1912
rect 63628 1818 63668 1903
rect 65356 1818 65396 1903
rect 63243 1700 63285 1709
rect 63243 1660 63244 1700
rect 63284 1660 63285 1700
rect 63243 1651 63285 1660
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 65548 1364 65588 2358
rect 66220 2129 66260 2659
rect 66604 2624 66644 2633
rect 66219 2120 66261 2129
rect 66219 2080 66220 2120
rect 66260 2080 66261 2120
rect 66219 2071 66261 2080
rect 66219 1952 66261 1961
rect 66219 1912 66220 1952
rect 66260 1912 66261 1952
rect 66219 1903 66261 1912
rect 66220 1818 66260 1903
rect 66604 1709 66644 2584
rect 66700 2624 66740 2633
rect 66700 2465 66740 2584
rect 66891 2624 66933 2633
rect 66891 2584 66892 2624
rect 66932 2584 66933 2624
rect 66891 2575 66933 2584
rect 67563 2624 67605 2633
rect 67563 2584 67564 2624
rect 67604 2584 67605 2624
rect 67563 2575 67605 2584
rect 66892 2490 66932 2575
rect 66699 2456 66741 2465
rect 66699 2416 66700 2456
rect 66740 2416 66741 2456
rect 66699 2407 66741 2416
rect 66796 2456 66836 2465
rect 66796 2045 66836 2416
rect 66795 2036 66837 2045
rect 66795 1996 66796 2036
rect 66836 1996 66837 2036
rect 66795 1987 66837 1996
rect 67564 1952 67604 2575
rect 67659 2036 67701 2045
rect 67659 1996 67660 2036
rect 67700 1996 67701 2036
rect 67659 1987 67701 1996
rect 67564 1903 67604 1912
rect 67660 1910 67700 1987
rect 67756 1961 67796 2860
rect 68236 2624 68276 2633
rect 68139 2456 68181 2465
rect 68139 2416 68140 2456
rect 68180 2416 68181 2456
rect 68139 2407 68181 2416
rect 68140 2322 68180 2407
rect 68236 2120 68276 2584
rect 68332 2624 68372 2860
rect 68620 2876 68660 4180
rect 68716 4136 68756 5683
rect 68908 5648 68948 5767
rect 68908 5599 68948 5608
rect 69004 5648 69044 5659
rect 69004 5573 69044 5608
rect 69291 5648 69333 5657
rect 69291 5608 69292 5648
rect 69332 5608 69333 5648
rect 69291 5599 69333 5608
rect 69388 5648 69428 5767
rect 69388 5599 69428 5608
rect 69484 5648 69524 5944
rect 68811 5564 68853 5573
rect 68811 5524 68812 5564
rect 68852 5524 68853 5564
rect 68811 5515 68853 5524
rect 69003 5564 69045 5573
rect 69003 5524 69004 5564
rect 69044 5524 69045 5564
rect 69003 5515 69045 5524
rect 68812 4304 68852 5515
rect 69100 5422 69140 5431
rect 69100 4388 69140 5382
rect 69195 4976 69237 4985
rect 69195 4936 69196 4976
rect 69236 4936 69237 4976
rect 69195 4927 69237 4936
rect 69196 4842 69236 4927
rect 69292 4808 69332 5599
rect 69292 4768 69428 4808
rect 69292 4388 69332 4397
rect 69100 4348 69292 4388
rect 68907 4304 68949 4313
rect 68812 4264 68908 4304
rect 68948 4264 68949 4304
rect 68907 4255 68949 4264
rect 68716 4061 68756 4096
rect 68715 4052 68757 4061
rect 68715 4012 68716 4052
rect 68756 4012 68757 4052
rect 68715 4003 68757 4012
rect 68620 2827 68660 2836
rect 68332 2575 68372 2584
rect 68427 2624 68469 2633
rect 68427 2584 68428 2624
rect 68468 2584 68469 2624
rect 68427 2575 68469 2584
rect 68620 2624 68660 2633
rect 68716 2624 68756 4003
rect 68811 3632 68853 3641
rect 68811 3592 68812 3632
rect 68852 3592 68853 3632
rect 68811 3583 68853 3592
rect 68812 3498 68852 3583
rect 68908 2900 68948 4255
rect 69100 4220 69140 4229
rect 69004 4180 69100 4220
rect 69004 3725 69044 4180
rect 69100 4171 69140 4180
rect 69196 4145 69236 4348
rect 69292 4339 69332 4348
rect 69195 4136 69237 4145
rect 69195 4096 69196 4136
rect 69236 4096 69237 4136
rect 69195 4087 69237 4096
rect 69388 4136 69428 4768
rect 69388 4087 69428 4096
rect 69003 3716 69045 3725
rect 69003 3676 69004 3716
rect 69044 3676 69045 3716
rect 69003 3667 69045 3676
rect 69004 3632 69044 3667
rect 69004 3581 69044 3592
rect 69195 3380 69237 3389
rect 69195 3340 69196 3380
rect 69236 3340 69237 3380
rect 69195 3331 69237 3340
rect 69196 3246 69236 3331
rect 68660 2584 68756 2624
rect 68812 2860 68948 2900
rect 68812 2624 68852 2860
rect 69484 2633 69524 5608
rect 69580 5648 69620 6607
rect 69675 6488 69717 6497
rect 69675 6448 69676 6488
rect 69716 6448 69717 6488
rect 69675 6439 69717 6448
rect 69676 6354 69716 6439
rect 70060 6329 70100 7036
rect 70444 6413 70484 7120
rect 70540 8672 70580 9463
rect 70827 8672 70869 8681
rect 70540 8632 70828 8672
rect 70868 8632 70869 8672
rect 70540 6497 70580 8632
rect 70827 8623 70869 8632
rect 70828 8538 70868 8623
rect 70827 6656 70869 6665
rect 70827 6616 70828 6656
rect 70868 6616 70869 6656
rect 70827 6607 70869 6616
rect 70828 6522 70868 6607
rect 70539 6488 70581 6497
rect 70539 6448 70540 6488
rect 70580 6448 70581 6488
rect 70539 6439 70581 6448
rect 70731 6488 70773 6497
rect 70731 6448 70732 6488
rect 70772 6448 70773 6488
rect 70731 6439 70773 6448
rect 70155 6404 70197 6413
rect 70155 6364 70156 6404
rect 70196 6364 70197 6404
rect 70155 6355 70197 6364
rect 70443 6404 70485 6413
rect 70443 6364 70444 6404
rect 70484 6364 70485 6404
rect 70443 6355 70485 6364
rect 70059 6320 70101 6329
rect 70059 6280 70060 6320
rect 70100 6280 70101 6320
rect 70059 6271 70101 6280
rect 69771 5732 69813 5741
rect 69771 5692 69772 5732
rect 69812 5692 69813 5732
rect 69771 5683 69813 5692
rect 69580 5599 69620 5608
rect 69676 5648 69716 5657
rect 69676 5573 69716 5608
rect 69675 5564 69717 5573
rect 69772 5564 69812 5683
rect 69675 5524 69676 5564
rect 69716 5524 69812 5564
rect 69675 5515 69717 5524
rect 69676 5430 69716 5515
rect 69675 4304 69717 4313
rect 69675 4264 69676 4304
rect 69716 4264 69717 4304
rect 69675 4255 69717 4264
rect 69676 3548 69716 4255
rect 69676 3499 69716 3508
rect 68620 2575 68660 2584
rect 68812 2575 68852 2584
rect 68908 2624 68948 2633
rect 69196 2624 69236 2633
rect 69483 2624 69525 2633
rect 68948 2584 69196 2624
rect 69236 2584 69332 2624
rect 68908 2575 68948 2584
rect 69196 2575 69236 2584
rect 68428 2490 68468 2575
rect 68811 2456 68853 2465
rect 68811 2416 68812 2456
rect 68852 2416 68853 2456
rect 68811 2407 68853 2416
rect 69100 2456 69140 2465
rect 68619 2204 68661 2213
rect 68619 2155 68620 2204
rect 67852 2080 68276 2120
rect 67755 1952 67797 1961
rect 67755 1912 67756 1952
rect 67796 1912 67797 1952
rect 67755 1903 67797 1912
rect 67660 1861 67700 1870
rect 67852 1868 67892 2080
rect 67852 1819 67892 1828
rect 67948 1952 67988 1961
rect 67948 1793 67988 1912
rect 68043 1952 68085 1961
rect 68043 1912 68044 1952
rect 68084 1912 68085 1952
rect 68043 1903 68085 1912
rect 67756 1784 67796 1793
rect 66219 1700 66261 1709
rect 66219 1660 66220 1700
rect 66260 1660 66261 1700
rect 66219 1651 66261 1660
rect 66603 1700 66645 1709
rect 66603 1660 66604 1700
rect 66644 1660 66645 1700
rect 66603 1651 66645 1660
rect 67371 1700 67413 1709
rect 67371 1660 67372 1700
rect 67412 1660 67413 1700
rect 67371 1651 67413 1660
rect 66124 1364 66164 1373
rect 65548 1324 66124 1364
rect 66124 1315 66164 1324
rect 62860 1063 62900 1072
rect 66220 1112 66260 1651
rect 67372 1566 67412 1651
rect 67179 1196 67221 1205
rect 67179 1156 67180 1196
rect 67220 1156 67221 1196
rect 67179 1147 67221 1156
rect 66220 1063 66260 1072
rect 66795 1112 66837 1121
rect 66795 1072 66796 1112
rect 66836 1072 66837 1112
rect 66795 1063 66837 1072
rect 67180 1112 67220 1147
rect 67756 1121 67796 1744
rect 67947 1784 67989 1793
rect 67947 1744 67948 1784
rect 67988 1744 67989 1784
rect 67947 1735 67989 1744
rect 59884 978 59924 1063
rect 66796 978 66836 1063
rect 67180 1061 67220 1072
rect 67755 1112 67797 1121
rect 67755 1072 67756 1112
rect 67796 1072 67797 1112
rect 67755 1063 67797 1072
rect 68044 1112 68084 1903
rect 68140 1784 68180 1793
rect 68236 1784 68276 2080
rect 68660 2155 68661 2204
rect 68180 1744 68276 1784
rect 68428 1952 68468 1961
rect 68140 1735 68180 1744
rect 68428 1121 68468 1912
rect 68524 1952 68564 1961
rect 68524 1709 68564 1912
rect 68620 1793 68660 2138
rect 68812 2036 68852 2407
rect 69100 2213 69140 2416
rect 69099 2204 69141 2213
rect 69099 2164 69100 2204
rect 69140 2164 69141 2204
rect 69099 2155 69141 2164
rect 68812 1987 68852 1996
rect 69195 2036 69237 2045
rect 69195 1996 69196 2036
rect 69236 1996 69237 2036
rect 69195 1987 69237 1996
rect 69196 1952 69236 1987
rect 69196 1901 69236 1912
rect 68619 1784 68661 1793
rect 68619 1744 68620 1784
rect 68660 1744 68661 1784
rect 68619 1735 68661 1744
rect 68523 1700 68565 1709
rect 68523 1660 68524 1700
rect 68564 1660 68565 1700
rect 68523 1651 68565 1660
rect 69196 1364 69236 1373
rect 69292 1364 69332 2584
rect 69483 2584 69484 2624
rect 69524 2584 69620 2624
rect 69483 2575 69525 2584
rect 69580 1541 69620 2584
rect 69772 1709 69812 5524
rect 70156 5153 70196 6355
rect 70347 5648 70389 5657
rect 70347 5608 70348 5648
rect 70388 5608 70389 5648
rect 70347 5599 70389 5608
rect 70155 5144 70197 5153
rect 70155 5104 70156 5144
rect 70196 5104 70197 5144
rect 70155 5095 70197 5104
rect 70348 5144 70388 5599
rect 70348 5095 70388 5104
rect 70060 3464 70100 3473
rect 70156 3464 70196 5095
rect 70539 5060 70581 5069
rect 70539 5020 70540 5060
rect 70580 5020 70581 5060
rect 70539 5011 70581 5020
rect 70540 4926 70580 5011
rect 70100 3424 70196 3464
rect 70060 3415 70100 3424
rect 70059 2876 70101 2885
rect 70059 2836 70060 2876
rect 70100 2836 70101 2876
rect 70059 2827 70101 2836
rect 70060 1961 70100 2827
rect 70156 2045 70196 3424
rect 70155 2036 70197 2045
rect 70155 1996 70156 2036
rect 70196 1996 70197 2036
rect 70155 1987 70197 1996
rect 70059 1952 70101 1961
rect 70059 1912 70060 1952
rect 70100 1912 70101 1952
rect 70059 1903 70101 1912
rect 70060 1818 70100 1903
rect 69771 1700 69813 1709
rect 69771 1660 69772 1700
rect 69812 1660 69813 1700
rect 69771 1651 69813 1660
rect 69579 1532 69621 1541
rect 69579 1492 69580 1532
rect 69620 1492 69621 1532
rect 69579 1483 69621 1492
rect 69236 1324 69332 1364
rect 69196 1315 69236 1324
rect 68044 1063 68084 1072
rect 68427 1112 68469 1121
rect 68427 1072 68428 1112
rect 68468 1072 68469 1112
rect 68427 1063 68469 1072
rect 69483 1112 69525 1121
rect 69483 1072 69484 1112
rect 69524 1072 69525 1112
rect 69483 1063 69525 1072
rect 69580 1112 69620 1483
rect 69675 1196 69717 1205
rect 69675 1156 69676 1196
rect 69716 1156 69717 1196
rect 69675 1147 69717 1156
rect 69580 1063 69620 1072
rect 69676 1112 69716 1147
rect 69484 978 69524 1063
rect 69676 1061 69716 1072
rect 69772 1112 69812 1651
rect 70732 1364 70772 6439
rect 70924 6068 70964 13747
rect 71019 13628 71061 13637
rect 71019 13588 71020 13628
rect 71060 13588 71061 13628
rect 71019 13579 71061 13588
rect 71020 13460 71060 13579
rect 71116 13553 71156 13840
rect 71212 13830 71252 13915
rect 71115 13544 71157 13553
rect 71115 13504 71116 13544
rect 71156 13504 71157 13544
rect 71115 13495 71157 13504
rect 71020 13376 71060 13420
rect 71308 13385 71348 14008
rect 71403 14048 71445 14057
rect 71403 14008 71404 14048
rect 71444 14008 71445 14048
rect 71403 13999 71445 14008
rect 71307 13376 71349 13385
rect 71020 13336 71252 13376
rect 71115 13208 71157 13217
rect 71115 13168 71116 13208
rect 71156 13168 71157 13208
rect 71115 13159 71157 13168
rect 71212 13208 71252 13336
rect 71307 13336 71308 13376
rect 71348 13336 71349 13376
rect 71307 13327 71349 13336
rect 71404 13292 71444 13999
rect 71500 13460 71540 14176
rect 71596 14057 71636 15520
rect 71884 15233 71924 17032
rect 72075 16232 72117 16241
rect 72075 16192 72076 16232
rect 72116 16192 72117 16232
rect 72075 16183 72117 16192
rect 72172 16232 72212 16241
rect 71979 16064 72021 16073
rect 71979 16024 71980 16064
rect 72020 16024 72021 16064
rect 71979 16015 72021 16024
rect 71883 15224 71925 15233
rect 71883 15184 71884 15224
rect 71924 15184 71925 15224
rect 71883 15175 71925 15184
rect 71884 14720 71924 14729
rect 71692 14680 71884 14720
rect 71595 14048 71637 14057
rect 71595 14008 71596 14048
rect 71636 14008 71637 14048
rect 71595 13999 71637 14008
rect 71500 13411 71540 13420
rect 71404 13252 71540 13292
rect 71212 13159 71252 13168
rect 71308 13208 71348 13217
rect 71116 11024 71156 13159
rect 71308 13124 71348 13168
rect 71500 13208 71540 13252
rect 71596 13217 71636 13999
rect 71692 13973 71732 14680
rect 71884 14671 71924 14680
rect 71980 14720 72020 16015
rect 72076 15560 72116 16183
rect 72172 15737 72212 16192
rect 72268 16064 72308 16073
rect 72268 15821 72308 16024
rect 72267 15812 72309 15821
rect 72267 15772 72268 15812
rect 72308 15772 72309 15812
rect 72267 15763 72309 15772
rect 72171 15728 72213 15737
rect 72171 15688 72172 15728
rect 72212 15688 72213 15728
rect 72171 15679 72213 15688
rect 72268 15569 72308 15763
rect 72364 15653 72404 17032
rect 72459 16652 72501 16661
rect 72459 16612 72460 16652
rect 72500 16612 72501 16652
rect 72459 16603 72501 16612
rect 72460 16493 72500 16603
rect 72459 16484 72501 16493
rect 72459 16444 72460 16484
rect 72500 16444 72501 16484
rect 72459 16435 72501 16444
rect 72460 16232 72500 16435
rect 72556 16325 72596 17200
rect 72555 16316 72597 16325
rect 72555 16276 72556 16316
rect 72596 16276 72597 16316
rect 72555 16267 72597 16276
rect 72460 16183 72500 16192
rect 72556 16064 72596 16073
rect 72556 15989 72596 16024
rect 72555 15980 72597 15989
rect 72555 15940 72556 15980
rect 72596 15940 72597 15980
rect 72555 15931 72597 15940
rect 72556 15929 72596 15931
rect 72363 15644 72405 15653
rect 72363 15604 72364 15644
rect 72404 15604 72405 15644
rect 72363 15595 72405 15604
rect 72267 15560 72309 15569
rect 72076 15520 72212 15560
rect 72075 14888 72117 14897
rect 72075 14848 72076 14888
rect 72116 14848 72117 14888
rect 72075 14839 72117 14848
rect 71980 14671 72020 14680
rect 72076 14720 72116 14839
rect 72076 14671 72116 14680
rect 72172 14561 72212 15520
rect 72267 15520 72268 15560
rect 72308 15520 72309 15560
rect 72267 15511 72309 15520
rect 72459 14636 72501 14645
rect 72459 14596 72460 14636
rect 72500 14596 72501 14636
rect 72459 14587 72501 14596
rect 71788 14552 71828 14561
rect 71788 14132 71828 14512
rect 72171 14552 72213 14561
rect 72171 14512 72172 14552
rect 72212 14512 72213 14552
rect 72171 14503 72213 14512
rect 71884 14132 71924 14141
rect 71788 14092 71884 14132
rect 71884 14083 71924 14092
rect 71691 13964 71733 13973
rect 71691 13924 71692 13964
rect 71732 13924 71733 13964
rect 71691 13915 71733 13924
rect 71692 13460 71732 13915
rect 72172 13796 72212 14503
rect 72267 14384 72309 14393
rect 72267 14344 72268 14384
rect 72308 14344 72309 14384
rect 72267 14335 72309 14344
rect 72268 14048 72308 14335
rect 72268 13973 72308 14008
rect 72267 13964 72309 13973
rect 72267 13924 72268 13964
rect 72308 13924 72309 13964
rect 72267 13915 72309 13924
rect 72172 13756 72308 13796
rect 71692 13411 71732 13420
rect 72171 13376 72213 13385
rect 72171 13336 72172 13376
rect 72212 13336 72213 13376
rect 72171 13327 72213 13336
rect 71403 13124 71445 13133
rect 71308 13084 71404 13124
rect 71444 13084 71445 13124
rect 71403 13075 71445 13084
rect 71500 11696 71540 13168
rect 71595 13208 71637 13217
rect 71595 13168 71596 13208
rect 71636 13168 71637 13208
rect 71595 13159 71637 13168
rect 71979 13208 72021 13217
rect 71979 13168 71980 13208
rect 72020 13168 72021 13208
rect 71979 13159 72021 13168
rect 72076 13208 72116 13217
rect 71787 13124 71829 13133
rect 71787 13084 71788 13124
rect 71828 13084 71829 13124
rect 71787 13075 71829 13084
rect 71596 11696 71636 11705
rect 71500 11656 71596 11696
rect 71212 11024 71252 11033
rect 71116 10984 71212 11024
rect 71019 10100 71061 10109
rect 71019 10060 71020 10100
rect 71060 10060 71061 10100
rect 71212 10100 71252 10984
rect 71596 10184 71636 11656
rect 71788 11696 71828 13075
rect 71980 13074 72020 13159
rect 72076 12965 72116 13168
rect 72172 13036 72212 13327
rect 72075 12956 72117 12965
rect 72075 12916 72076 12956
rect 72116 12916 72117 12956
rect 72075 12907 72117 12916
rect 72172 12704 72212 12996
rect 72172 12655 72212 12664
rect 72076 12536 72116 12545
rect 71788 11647 71828 11656
rect 71884 12452 71924 12461
rect 72076 12452 72116 12496
rect 71924 12412 72116 12452
rect 71884 11696 71924 12412
rect 71979 11864 72021 11873
rect 71979 11824 71980 11864
rect 72020 11824 72021 11864
rect 71979 11815 72021 11824
rect 71884 11647 71924 11656
rect 71692 11528 71732 11537
rect 71732 11488 71828 11528
rect 71692 11479 71732 11488
rect 71788 10268 71828 11488
rect 71883 11024 71925 11033
rect 71883 10984 71884 11024
rect 71924 10984 71925 11024
rect 71883 10975 71925 10984
rect 71884 10352 71924 10975
rect 71884 10303 71924 10312
rect 71788 10219 71828 10228
rect 71980 10268 72020 11815
rect 72172 11696 72212 11705
rect 72075 11528 72117 11537
rect 72075 11488 72076 11528
rect 72116 11488 72117 11528
rect 72075 11479 72117 11488
rect 71980 10219 72020 10228
rect 72076 10226 72116 11479
rect 72172 11192 72212 11656
rect 72268 11453 72308 13756
rect 72460 12965 72500 14587
rect 72555 14384 72597 14393
rect 72555 14344 72556 14384
rect 72596 14344 72597 14384
rect 72555 14335 72597 14344
rect 72459 12956 72501 12965
rect 72459 12916 72460 12956
rect 72500 12916 72501 12956
rect 72459 12907 72501 12916
rect 72460 11696 72500 12907
rect 72556 12284 72596 14335
rect 72652 14225 72692 17260
rect 72844 16577 72884 17260
rect 73132 16661 73172 17260
rect 73255 17072 73295 17472
rect 73545 17072 73585 17472
rect 73228 17032 73295 17072
rect 73516 17032 73585 17072
rect 73655 17072 73695 17472
rect 73945 17156 73985 17472
rect 73900 17116 73985 17156
rect 73655 17032 73748 17072
rect 73131 16652 73173 16661
rect 73131 16612 73132 16652
rect 73172 16612 73173 16652
rect 73131 16603 73173 16612
rect 72843 16568 72885 16577
rect 72843 16528 72844 16568
rect 72884 16528 72885 16568
rect 72843 16519 72885 16528
rect 73131 16400 73173 16409
rect 73131 16360 73132 16400
rect 73172 16360 73173 16400
rect 73131 16351 73173 16360
rect 72843 16316 72885 16325
rect 72843 16276 72844 16316
rect 72884 16276 72885 16316
rect 72843 16267 72885 16276
rect 72747 15728 72789 15737
rect 72747 15688 72748 15728
rect 72788 15688 72789 15728
rect 72747 15679 72789 15688
rect 72748 15594 72788 15679
rect 72844 15485 72884 16267
rect 72939 16148 72981 16157
rect 72939 16108 72940 16148
rect 72980 16108 72981 16148
rect 72939 16099 72981 16108
rect 72940 15728 72980 16099
rect 73132 15737 73172 16351
rect 73228 15989 73268 17032
rect 73420 16493 73460 16578
rect 73419 16484 73461 16493
rect 73419 16444 73420 16484
rect 73460 16444 73461 16484
rect 73419 16435 73461 16444
rect 73516 16409 73556 17032
rect 73515 16400 73557 16409
rect 73515 16360 73516 16400
rect 73556 16360 73557 16400
rect 73515 16351 73557 16360
rect 73419 16316 73461 16325
rect 73324 16276 73420 16316
rect 73460 16276 73461 16316
rect 73324 16232 73364 16276
rect 73419 16267 73461 16276
rect 73324 16183 73364 16192
rect 73419 16064 73461 16073
rect 73419 16024 73420 16064
rect 73460 16024 73461 16064
rect 73419 16015 73461 16024
rect 73611 16064 73653 16073
rect 73611 16024 73612 16064
rect 73652 16024 73653 16064
rect 73611 16015 73653 16024
rect 73227 15980 73269 15989
rect 73227 15940 73228 15980
rect 73268 15940 73269 15980
rect 73227 15931 73269 15940
rect 73420 15930 73460 16015
rect 72940 15679 72980 15688
rect 73131 15728 73173 15737
rect 73131 15688 73132 15728
rect 73172 15688 73173 15728
rect 73131 15679 73173 15688
rect 72843 15476 72885 15485
rect 72843 15436 72844 15476
rect 72884 15436 72885 15476
rect 72843 15427 72885 15436
rect 73438 14972 73480 14981
rect 73438 14932 73439 14972
rect 73479 14932 73480 14972
rect 73438 14923 73480 14932
rect 72747 14888 72789 14897
rect 72747 14848 72748 14888
rect 72788 14848 72789 14888
rect 72747 14839 72789 14848
rect 72651 14216 72693 14225
rect 72651 14176 72652 14216
rect 72692 14176 72693 14216
rect 72651 14167 72693 14176
rect 72651 13208 72693 13217
rect 72651 13168 72652 13208
rect 72692 13168 72693 13208
rect 72651 13159 72693 13168
rect 72748 13208 72788 14839
rect 73439 14799 73479 14923
rect 73439 14729 73479 14759
rect 73438 14720 73480 14729
rect 73612 14720 73652 16015
rect 73708 15821 73748 17032
rect 73900 16325 73940 17116
rect 74055 17072 74095 17472
rect 74187 17240 74229 17249
rect 74187 17200 74188 17240
rect 74228 17200 74229 17240
rect 74187 17191 74229 17200
rect 73996 17032 74095 17072
rect 73996 16493 74036 17032
rect 73995 16484 74037 16493
rect 73995 16444 73996 16484
rect 74036 16444 74037 16484
rect 73995 16435 74037 16444
rect 74188 16484 74228 17191
rect 74345 17072 74385 17472
rect 74188 16435 74228 16444
rect 74284 17032 74385 17072
rect 74455 17072 74495 17472
rect 74745 17240 74785 17472
rect 74855 17249 74895 17472
rect 74854 17240 74896 17249
rect 74745 17200 74804 17240
rect 74667 17156 74709 17165
rect 74667 17116 74668 17156
rect 74708 17116 74709 17156
rect 74667 17107 74709 17116
rect 74455 17032 74516 17072
rect 73899 16316 73941 16325
rect 73804 16276 73900 16316
rect 73940 16276 73941 16316
rect 73707 15812 73749 15821
rect 73707 15772 73708 15812
rect 73748 15772 73749 15812
rect 73707 15763 73749 15772
rect 73707 15476 73749 15485
rect 73707 15436 73708 15476
rect 73748 15436 73749 15476
rect 73707 15427 73749 15436
rect 73438 14680 73439 14720
rect 73479 14680 73480 14720
rect 73438 14671 73480 14680
rect 73545 14680 73652 14720
rect 73545 14636 73585 14680
rect 73516 14596 73585 14636
rect 73035 14552 73077 14561
rect 73035 14512 73036 14552
rect 73076 14512 73077 14552
rect 73035 14503 73077 14512
rect 72843 14216 72885 14225
rect 72843 14176 72844 14216
rect 72884 14176 72885 14216
rect 72843 14167 72885 14176
rect 72652 13074 72692 13159
rect 72748 12713 72788 13168
rect 72844 13208 72884 14167
rect 72844 13159 72884 13168
rect 72940 13208 72980 13217
rect 72940 12965 72980 13168
rect 72939 12956 72981 12965
rect 72939 12916 72940 12956
rect 72980 12916 72981 12956
rect 72939 12907 72981 12916
rect 72747 12704 72789 12713
rect 72747 12664 72748 12704
rect 72788 12664 72789 12704
rect 72747 12655 72789 12664
rect 72652 12536 72692 12545
rect 73036 12536 73076 14503
rect 73131 14048 73173 14057
rect 73131 14008 73132 14048
rect 73172 14008 73173 14048
rect 73131 13999 73173 14008
rect 73132 13914 73172 13999
rect 73227 13460 73269 13469
rect 73227 13420 73228 13460
rect 73268 13420 73269 13460
rect 73227 13411 73269 13420
rect 72692 12496 72980 12536
rect 72652 12487 72692 12496
rect 72556 12244 72788 12284
rect 72460 11621 72500 11656
rect 72555 11696 72597 11705
rect 72555 11656 72556 11696
rect 72596 11656 72597 11696
rect 72555 11647 72597 11656
rect 72459 11612 72501 11621
rect 72459 11572 72460 11612
rect 72500 11572 72501 11612
rect 72459 11563 72501 11572
rect 72556 11562 72596 11647
rect 72363 11528 72405 11537
rect 72363 11484 72364 11528
rect 72404 11484 72405 11528
rect 72363 11479 72405 11484
rect 72267 11444 72309 11453
rect 72267 11404 72268 11444
rect 72308 11404 72309 11444
rect 72267 11395 72309 11404
rect 72364 11393 72404 11479
rect 72748 11369 72788 12244
rect 72843 11864 72885 11873
rect 72843 11824 72844 11864
rect 72884 11824 72885 11864
rect 72843 11815 72885 11824
rect 72844 11730 72884 11815
rect 72940 11696 72980 12496
rect 73036 12487 73076 12496
rect 73131 11864 73173 11873
rect 73131 11824 73132 11864
rect 73172 11824 73173 11864
rect 73131 11815 73173 11824
rect 73036 11696 73076 11705
rect 72940 11656 73036 11696
rect 73036 11647 73076 11656
rect 73132 11696 73172 11815
rect 73132 11647 73172 11656
rect 73228 11696 73268 13411
rect 73323 12452 73365 12461
rect 73323 12412 73324 12452
rect 73364 12412 73365 12452
rect 73323 12403 73365 12412
rect 73324 11789 73364 12403
rect 73516 11864 73556 14596
rect 73611 14552 73653 14561
rect 73708 14552 73748 15427
rect 73611 14512 73612 14552
rect 73652 14512 73748 14552
rect 73611 14503 73653 14512
rect 73612 14418 73652 14503
rect 73804 14225 73844 16276
rect 73899 16267 73941 16276
rect 74091 16232 74133 16241
rect 74091 16192 74092 16232
rect 74132 16192 74133 16232
rect 74091 16183 74133 16192
rect 74092 16098 74132 16183
rect 74187 16064 74229 16073
rect 74187 16024 74188 16064
rect 74228 16024 74229 16064
rect 74187 16015 74229 16024
rect 74188 15930 74228 16015
rect 74284 15728 74324 17032
rect 74379 15980 74421 15989
rect 74379 15940 74380 15980
rect 74420 15940 74421 15980
rect 74379 15931 74421 15940
rect 73900 15688 74324 15728
rect 73803 14216 73845 14225
rect 73803 14176 73804 14216
rect 73844 14176 73845 14216
rect 73803 14167 73845 14176
rect 73803 14048 73845 14057
rect 73803 14008 73804 14048
rect 73844 14008 73845 14048
rect 73803 13999 73845 14008
rect 73804 13217 73844 13999
rect 73803 13208 73845 13217
rect 73803 13168 73804 13208
rect 73844 13168 73845 13208
rect 73803 13159 73845 13168
rect 73900 13208 73940 15688
rect 74092 15560 74132 15569
rect 74092 14057 74132 15520
rect 74187 14720 74229 14729
rect 74187 14680 74188 14720
rect 74228 14680 74229 14720
rect 74187 14671 74229 14680
rect 74091 14048 74133 14057
rect 74091 14008 74092 14048
rect 74132 14008 74133 14048
rect 74091 13999 74133 14008
rect 74188 13628 74228 14671
rect 74283 14216 74325 14225
rect 74283 14176 74284 14216
rect 74324 14176 74325 14216
rect 74283 14167 74325 14176
rect 74284 14082 74324 14167
rect 74188 13588 74324 13628
rect 73995 13460 74037 13469
rect 73995 13420 73996 13460
rect 74036 13420 74037 13460
rect 73995 13411 74037 13420
rect 73996 13326 74036 13411
rect 74187 13376 74229 13385
rect 74187 13336 74188 13376
rect 74228 13336 74229 13376
rect 74187 13327 74229 13336
rect 73707 12704 73749 12713
rect 73707 12664 73708 12704
rect 73748 12664 73749 12704
rect 73707 12655 73749 12664
rect 73420 11824 73556 11864
rect 73323 11780 73365 11789
rect 73323 11740 73324 11780
rect 73364 11740 73365 11780
rect 73323 11731 73365 11740
rect 73228 11647 73268 11656
rect 73324 11696 73364 11731
rect 73324 11616 73364 11656
rect 73420 11528 73460 11824
rect 73507 11696 73556 11705
rect 73507 11656 73508 11696
rect 73507 11647 73556 11656
rect 73611 11696 73653 11705
rect 73611 11656 73612 11696
rect 73652 11656 73653 11696
rect 73611 11647 73653 11656
rect 73708 11696 73748 12655
rect 73804 12536 73844 13159
rect 73900 12713 73940 13168
rect 74188 13208 74228 13327
rect 74188 13159 74228 13168
rect 73899 12704 73941 12713
rect 73899 12664 73900 12704
rect 73940 12664 73941 12704
rect 73899 12655 73941 12664
rect 73900 12536 73940 12545
rect 73804 12496 73900 12536
rect 73900 12487 73940 12496
rect 73708 11647 73748 11656
rect 73803 11696 73845 11705
rect 73803 11656 73804 11696
rect 73844 11656 73845 11696
rect 73803 11647 73845 11656
rect 73508 11569 73548 11647
rect 73612 11562 73652 11647
rect 73804 11562 73844 11647
rect 73324 11488 73460 11528
rect 73324 11444 73364 11488
rect 72940 11404 73364 11444
rect 72747 11360 72789 11369
rect 72747 11320 72748 11360
rect 72788 11320 72789 11360
rect 72747 11311 72789 11320
rect 72364 11192 72404 11201
rect 72172 11152 72364 11192
rect 72364 11143 72404 11152
rect 72652 11152 72884 11192
rect 72364 10772 72404 10781
rect 72404 10732 72596 10772
rect 72364 10723 72404 10732
rect 71691 10184 71733 10193
rect 71596 10144 71692 10184
rect 71732 10144 71733 10184
rect 72076 10177 72116 10186
rect 72268 10184 72308 10193
rect 71691 10135 71733 10144
rect 71212 10060 71636 10100
rect 71019 10051 71061 10060
rect 71020 6665 71060 10051
rect 71499 9512 71541 9521
rect 71499 9472 71500 9512
rect 71540 9472 71541 9512
rect 71499 9463 71541 9472
rect 71500 8000 71540 9463
rect 71596 9344 71636 10060
rect 71692 10050 71732 10135
rect 72268 10100 72308 10144
rect 71980 10060 72308 10100
rect 72460 10184 72500 10193
rect 71980 9521 72020 10060
rect 72364 10016 72404 10025
rect 72076 9976 72364 10016
rect 71979 9512 72021 9521
rect 71979 9472 71980 9512
rect 72020 9472 72021 9512
rect 71979 9463 72021 9472
rect 72076 9428 72116 9976
rect 72364 9967 72404 9976
rect 72267 9596 72309 9605
rect 72267 9556 72268 9596
rect 72308 9556 72309 9596
rect 72267 9547 72309 9556
rect 72076 9379 72116 9388
rect 72268 9428 72308 9547
rect 72364 9512 72404 9523
rect 72364 9437 72404 9472
rect 72268 9379 72308 9388
rect 72363 9428 72405 9437
rect 72363 9388 72364 9428
rect 72404 9388 72405 9428
rect 72363 9379 72405 9388
rect 72172 9344 72212 9353
rect 71596 9304 72020 9344
rect 71691 8924 71733 8933
rect 71691 8884 71692 8924
rect 71732 8884 71733 8924
rect 71691 8875 71733 8884
rect 71692 8672 71732 8875
rect 71787 8756 71829 8765
rect 71787 8716 71788 8756
rect 71828 8716 71829 8756
rect 71787 8707 71829 8716
rect 71692 8623 71732 8632
rect 71691 8336 71733 8345
rect 71691 8296 71692 8336
rect 71732 8296 71733 8336
rect 71691 8287 71733 8296
rect 71404 7960 71500 8000
rect 71404 7757 71444 7960
rect 71500 7951 71540 7960
rect 71692 8000 71732 8287
rect 71692 7951 71732 7960
rect 71788 8000 71828 8707
rect 71980 8336 72020 9304
rect 72076 8672 72116 8681
rect 72172 8672 72212 9304
rect 72460 8767 72500 10144
rect 72556 10184 72596 10732
rect 72556 10135 72596 10144
rect 72652 9638 72692 11152
rect 72748 11024 72788 11033
rect 72748 10184 72788 10984
rect 72844 11024 72884 11152
rect 72844 10975 72884 10984
rect 72940 11024 72980 11404
rect 73131 11276 73173 11285
rect 73131 11236 73132 11276
rect 73172 11236 73173 11276
rect 73131 11227 73173 11236
rect 72940 10975 72980 10984
rect 73036 11024 73076 11033
rect 73036 10529 73076 10984
rect 73035 10520 73077 10529
rect 73035 10480 73036 10520
rect 73076 10480 73077 10520
rect 73035 10471 73077 10480
rect 73132 10361 73172 11227
rect 74092 11192 74132 11201
rect 73708 11152 74092 11192
rect 73515 10940 73557 10949
rect 73515 10900 73516 10940
rect 73556 10900 73557 10940
rect 73515 10891 73557 10900
rect 73516 10806 73556 10891
rect 73324 10772 73364 10781
rect 73228 10732 73324 10772
rect 73131 10352 73173 10361
rect 73131 10312 73132 10352
rect 73172 10312 73173 10352
rect 73131 10303 73173 10312
rect 72844 10184 72884 10193
rect 73228 10184 73268 10732
rect 73324 10723 73364 10732
rect 73323 10352 73365 10361
rect 73323 10312 73324 10352
rect 73364 10312 73365 10352
rect 73323 10303 73365 10312
rect 72748 10144 72844 10184
rect 72844 10135 72884 10144
rect 73132 10144 73228 10184
rect 72651 9598 72652 9605
rect 72939 9680 72981 9689
rect 72939 9640 72940 9680
rect 72980 9640 72981 9680
rect 72939 9631 72981 9640
rect 73036 9684 73076 9693
rect 72692 9598 72693 9605
rect 72651 9596 72693 9598
rect 72651 9556 72652 9596
rect 72692 9556 72693 9596
rect 72651 9547 72693 9556
rect 72843 9512 72885 9521
rect 72843 9472 72844 9512
rect 72884 9472 72885 9512
rect 72843 9463 72885 9472
rect 72940 9512 72980 9631
rect 72940 9463 72980 9472
rect 72844 9378 72884 9463
rect 73036 9437 73076 9644
rect 73035 9428 73077 9437
rect 73035 9388 73036 9428
rect 73076 9388 73077 9428
rect 73035 9379 73077 9388
rect 72555 8924 72597 8933
rect 72555 8884 72556 8924
rect 72596 8884 72597 8924
rect 72555 8875 72597 8884
rect 72940 8924 72980 8933
rect 73036 8924 73076 9379
rect 72980 8884 73076 8924
rect 72940 8875 72980 8884
rect 72116 8632 72212 8672
rect 72268 8727 72500 8767
rect 72076 8623 72116 8632
rect 72268 8345 72308 8727
rect 72460 8672 72500 8681
rect 72364 8513 72404 8598
rect 72363 8504 72405 8513
rect 72363 8464 72364 8504
rect 72404 8464 72405 8504
rect 72363 8455 72405 8464
rect 71884 8296 72020 8336
rect 72267 8336 72309 8345
rect 72267 8296 72268 8336
rect 72308 8296 72404 8336
rect 71884 8084 71924 8296
rect 72267 8287 72309 8296
rect 71980 8199 72020 8208
rect 72020 8159 72308 8168
rect 71980 8128 72308 8159
rect 71884 8044 72020 8084
rect 71788 7951 71828 7960
rect 71403 7748 71445 7757
rect 71403 7708 71404 7748
rect 71444 7708 71445 7748
rect 71403 7699 71445 7708
rect 71500 7748 71540 7757
rect 71787 7748 71829 7757
rect 71540 7708 71636 7748
rect 71500 7699 71540 7708
rect 71404 7253 71444 7699
rect 71403 7244 71445 7253
rect 71403 7204 71404 7244
rect 71444 7204 71445 7244
rect 71403 7195 71445 7204
rect 71308 7160 71348 7169
rect 71019 6656 71061 6665
rect 71019 6616 71020 6656
rect 71060 6616 71061 6656
rect 71019 6607 71061 6616
rect 71308 6497 71348 7120
rect 71307 6488 71349 6497
rect 71307 6448 71308 6488
rect 71348 6448 71349 6488
rect 71404 6488 71444 7195
rect 71500 6488 71540 6497
rect 71404 6448 71500 6488
rect 71307 6439 71349 6448
rect 71500 6439 71540 6448
rect 71596 6404 71636 7708
rect 71787 7708 71788 7748
rect 71828 7708 71829 7748
rect 71787 7699 71829 7708
rect 71596 6355 71636 6364
rect 71788 6404 71828 7699
rect 71883 7160 71925 7169
rect 71883 7120 71884 7160
rect 71924 7120 71925 7160
rect 71883 7111 71925 7120
rect 71884 6488 71924 7111
rect 71884 6439 71924 6448
rect 71788 6355 71828 6364
rect 71691 6320 71733 6329
rect 71691 6280 71692 6320
rect 71732 6280 71733 6320
rect 71691 6271 71733 6280
rect 71692 6186 71732 6271
rect 70828 6028 70964 6068
rect 70828 2708 70868 6028
rect 71499 5648 71541 5657
rect 71499 5608 71500 5648
rect 71540 5608 71541 5648
rect 71499 5599 71541 5608
rect 70923 5144 70965 5153
rect 70923 5104 70924 5144
rect 70964 5104 70965 5144
rect 70923 5095 70965 5104
rect 70924 4976 70964 5095
rect 70924 4927 70964 4936
rect 71019 4976 71061 4985
rect 71019 4936 71020 4976
rect 71060 4936 71061 4976
rect 71019 4927 71061 4936
rect 71020 4304 71060 4927
rect 71307 4724 71349 4733
rect 71307 4684 71308 4724
rect 71348 4684 71349 4724
rect 71307 4675 71349 4684
rect 70924 4264 71060 4304
rect 70924 3464 70964 4264
rect 71211 4220 71253 4229
rect 71211 4180 71212 4220
rect 71252 4180 71253 4220
rect 71211 4171 71253 4180
rect 71019 4136 71061 4145
rect 71019 4096 71020 4136
rect 71060 4096 71061 4136
rect 71019 4087 71061 4096
rect 71212 4136 71252 4171
rect 71020 4002 71060 4087
rect 71212 4085 71252 4096
rect 71308 4136 71348 4675
rect 71403 4220 71445 4229
rect 71403 4180 71404 4220
rect 71444 4180 71445 4220
rect 71403 4171 71445 4180
rect 71308 4087 71348 4096
rect 71115 3968 71157 3977
rect 71115 3928 71116 3968
rect 71156 3928 71157 3968
rect 71115 3919 71157 3928
rect 71116 3834 71156 3919
rect 70924 2885 70964 3424
rect 71404 3053 71444 4171
rect 71500 4145 71540 5599
rect 71787 4976 71829 4985
rect 71787 4936 71788 4976
rect 71828 4936 71829 4976
rect 71787 4927 71829 4936
rect 71788 4842 71828 4927
rect 71691 4304 71733 4313
rect 71691 4264 71692 4304
rect 71732 4264 71733 4304
rect 71691 4255 71733 4264
rect 71596 4220 71636 4229
rect 71499 4136 71541 4145
rect 71499 4096 71500 4136
rect 71540 4096 71541 4136
rect 71499 4087 71541 4096
rect 71500 3716 71540 4087
rect 71596 3977 71636 4180
rect 71692 4170 71732 4255
rect 71788 4220 71828 4229
rect 71595 3968 71637 3977
rect 71595 3928 71596 3968
rect 71636 3928 71637 3968
rect 71595 3919 71637 3928
rect 71788 3893 71828 4180
rect 71884 4136 71924 4145
rect 71884 3977 71924 4096
rect 71883 3968 71925 3977
rect 71883 3928 71884 3968
rect 71924 3928 71925 3968
rect 71883 3919 71925 3928
rect 71787 3884 71829 3893
rect 71787 3844 71788 3884
rect 71828 3844 71829 3884
rect 71787 3835 71829 3844
rect 71500 3676 71828 3716
rect 71595 3212 71637 3221
rect 71595 3172 71596 3212
rect 71636 3172 71637 3212
rect 71595 3163 71637 3172
rect 71403 3044 71445 3053
rect 71403 3004 71404 3044
rect 71444 3004 71445 3044
rect 71403 2995 71445 3004
rect 71404 2900 71444 2995
rect 70923 2876 70965 2885
rect 70923 2836 70924 2876
rect 70964 2836 70965 2876
rect 71404 2860 71540 2900
rect 70923 2827 70965 2836
rect 70828 2668 71252 2708
rect 71212 2120 71252 2668
rect 71307 2624 71349 2633
rect 71307 2584 71308 2624
rect 71348 2584 71349 2624
rect 71307 2575 71349 2584
rect 71500 2624 71540 2860
rect 71500 2575 71540 2584
rect 71596 2624 71636 3163
rect 71788 2633 71828 3676
rect 71884 3641 71924 3919
rect 71980 3800 72020 8044
rect 72076 8000 72116 8009
rect 72076 6404 72116 7960
rect 72171 8000 72213 8009
rect 72171 7960 72172 8000
rect 72212 7960 72213 8000
rect 72171 7951 72213 7960
rect 72172 7866 72212 7951
rect 72171 7244 72213 7253
rect 72171 7204 72172 7244
rect 72212 7204 72213 7244
rect 72171 7195 72213 7204
rect 72172 6488 72212 7195
rect 72268 7169 72308 8128
rect 72267 7160 72309 7169
rect 72267 7120 72268 7160
rect 72308 7120 72309 7160
rect 72267 7111 72309 7120
rect 72268 6488 72308 6497
rect 72172 6448 72268 6488
rect 72364 6488 72404 8296
rect 72460 7757 72500 8632
rect 72556 8672 72596 8875
rect 72651 8840 72693 8849
rect 72651 8800 72652 8840
rect 72692 8800 72693 8840
rect 72651 8791 72693 8800
rect 72556 8623 72596 8632
rect 72652 8672 72692 8791
rect 72843 8756 72885 8765
rect 72843 8716 72844 8756
rect 72884 8716 72885 8756
rect 72843 8707 72885 8716
rect 72652 8623 72692 8632
rect 72844 8672 72884 8707
rect 72844 8621 72884 8632
rect 72651 8504 72693 8513
rect 72651 8464 72652 8504
rect 72692 8464 72693 8504
rect 72651 8455 72693 8464
rect 72652 8084 72692 8455
rect 72652 8035 72692 8044
rect 73036 8000 73076 8009
rect 73132 8000 73172 10144
rect 73228 10135 73268 10144
rect 73228 9428 73268 9437
rect 73324 9428 73364 10303
rect 73419 9680 73461 9689
rect 73419 9640 73420 9680
rect 73460 9640 73461 9680
rect 73419 9631 73461 9640
rect 73420 9546 73460 9631
rect 73611 9512 73653 9521
rect 73611 9472 73612 9512
rect 73652 9472 73653 9512
rect 73611 9463 73653 9472
rect 73708 9512 73748 11152
rect 74092 11143 74132 11152
rect 74284 10949 74324 13588
rect 73900 10940 73940 10949
rect 74283 10940 74325 10949
rect 73940 10900 74036 10940
rect 73900 10891 73940 10900
rect 73803 10436 73845 10445
rect 73803 10396 73804 10436
rect 73844 10396 73845 10436
rect 73803 10387 73845 10396
rect 73268 9388 73364 9428
rect 73228 8261 73268 9388
rect 73612 9378 73652 9463
rect 73419 9260 73461 9269
rect 73419 9220 73420 9260
rect 73460 9220 73461 9260
rect 73419 9211 73461 9220
rect 73420 9126 73460 9211
rect 73515 9008 73557 9017
rect 73515 8968 73516 9008
rect 73556 8968 73557 9008
rect 73515 8959 73557 8968
rect 73516 8849 73556 8959
rect 73515 8840 73557 8849
rect 73515 8800 73516 8840
rect 73556 8800 73557 8840
rect 73515 8791 73557 8800
rect 73227 8252 73269 8261
rect 73227 8212 73228 8252
rect 73268 8212 73269 8252
rect 73227 8203 73269 8212
rect 73708 8177 73748 9472
rect 73804 9512 73844 10387
rect 73804 9463 73844 9472
rect 73900 9512 73940 9521
rect 73900 9269 73940 9472
rect 73899 9260 73941 9269
rect 73899 9220 73900 9260
rect 73940 9220 73941 9260
rect 73899 9211 73941 9220
rect 73803 8756 73845 8765
rect 73803 8716 73804 8756
rect 73844 8716 73845 8756
rect 73803 8707 73845 8716
rect 73707 8168 73749 8177
rect 73707 8128 73708 8168
rect 73748 8128 73749 8168
rect 73707 8119 73749 8128
rect 73076 7960 73172 8000
rect 73707 8000 73749 8009
rect 73707 7960 73708 8000
rect 73748 7960 73749 8000
rect 72459 7748 72501 7757
rect 72459 7708 72460 7748
rect 72500 7708 72501 7748
rect 72459 7699 72501 7708
rect 72460 7614 72500 7699
rect 73036 7337 73076 7960
rect 73707 7951 73749 7960
rect 73035 7328 73077 7337
rect 73035 7288 73036 7328
rect 73076 7288 73077 7328
rect 73035 7279 73077 7288
rect 73611 7328 73653 7337
rect 73611 7288 73612 7328
rect 73652 7288 73653 7328
rect 73611 7279 73653 7288
rect 73515 7244 73557 7253
rect 73515 7204 73516 7244
rect 73556 7204 73557 7244
rect 73515 7195 73557 7204
rect 72652 7160 72692 7169
rect 72460 6992 72500 7001
rect 72652 6992 72692 7120
rect 72747 7160 72789 7169
rect 72747 7120 72748 7160
rect 72788 7120 72789 7160
rect 72747 7111 72789 7120
rect 72748 7026 72788 7111
rect 73516 7110 73556 7195
rect 72500 6952 72692 6992
rect 73324 6992 73364 7001
rect 72460 6943 72500 6952
rect 72460 6488 72500 6497
rect 72364 6448 72460 6488
rect 72268 6439 72308 6448
rect 72076 6364 72212 6404
rect 72075 5984 72117 5993
rect 72075 5944 72076 5984
rect 72116 5944 72117 5984
rect 72075 5935 72117 5944
rect 72076 4229 72116 5935
rect 72172 5741 72212 6364
rect 72268 6236 72308 6245
rect 72308 6196 72404 6236
rect 72268 6187 72308 6196
rect 72171 5732 72213 5741
rect 72171 5692 72172 5732
rect 72212 5692 72213 5732
rect 72171 5683 72213 5692
rect 72364 5732 72404 6196
rect 72460 5993 72500 6448
rect 72556 6488 72596 6952
rect 72748 6656 72788 6665
rect 72788 6616 73268 6656
rect 72748 6607 72788 6616
rect 73228 6572 73268 6616
rect 73228 6523 73268 6532
rect 72556 6439 72596 6448
rect 72844 6488 72884 6497
rect 72459 5984 72501 5993
rect 72459 5944 72460 5984
rect 72500 5944 72501 5984
rect 72459 5935 72501 5944
rect 72364 5683 72404 5692
rect 72460 5816 72500 5825
rect 72844 5816 72884 6448
rect 72939 6488 72981 6497
rect 72939 6448 72940 6488
rect 72980 6448 72981 6488
rect 72939 6439 72981 6448
rect 73036 6488 73076 6497
rect 72940 6354 72980 6439
rect 73036 6329 73076 6448
rect 73035 6320 73077 6329
rect 73035 6280 73036 6320
rect 73076 6280 73077 6320
rect 73035 6271 73077 6280
rect 72940 5816 72980 5825
rect 72075 4220 72117 4229
rect 72075 4180 72076 4220
rect 72116 4180 72117 4220
rect 72075 4171 72117 4180
rect 72172 4136 72212 5683
rect 72267 5648 72309 5657
rect 72267 5608 72268 5648
rect 72308 5608 72309 5648
rect 72267 5599 72309 5608
rect 72268 5514 72308 5599
rect 72460 5069 72500 5776
rect 72556 5776 72940 5816
rect 72556 5732 72596 5776
rect 72940 5767 72980 5776
rect 73227 5816 73269 5825
rect 73227 5776 73228 5816
rect 73268 5776 73269 5816
rect 73227 5767 73269 5776
rect 72556 5683 72596 5692
rect 72651 5648 72693 5657
rect 72651 5608 72652 5648
rect 72692 5608 72693 5648
rect 72651 5599 72693 5608
rect 73228 5648 73268 5767
rect 73228 5599 73268 5608
rect 73324 5648 73364 6952
rect 73612 6488 73652 7279
rect 73708 7160 73748 7951
rect 73804 7832 73844 8707
rect 73900 8672 73940 9211
rect 73996 9017 74036 10900
rect 74283 10900 74284 10940
rect 74324 10900 74325 10940
rect 74283 10891 74325 10900
rect 74092 10184 74132 10193
rect 73995 9008 74037 9017
rect 73995 8968 73996 9008
rect 74036 8968 74037 9008
rect 73995 8959 74037 8968
rect 73996 8767 74036 8959
rect 73996 8718 74036 8727
rect 74092 8681 74132 10144
rect 74188 8840 74228 8849
rect 74091 8672 74133 8681
rect 73900 8632 74036 8672
rect 73899 8504 73941 8513
rect 73899 8464 73900 8504
rect 73940 8464 73941 8504
rect 73899 8455 73941 8464
rect 73900 8000 73940 8455
rect 73900 7951 73940 7960
rect 73804 7792 73940 7832
rect 73708 7111 73748 7120
rect 73804 7160 73844 7169
rect 73804 6917 73844 7120
rect 73900 7160 73940 7792
rect 73996 7253 74036 8632
rect 74091 8632 74092 8672
rect 74132 8632 74133 8672
rect 74091 8623 74133 8632
rect 74188 8420 74228 8800
rect 74092 8380 74228 8420
rect 73995 7244 74037 7253
rect 73995 7204 73996 7244
rect 74036 7204 74037 7244
rect 73995 7195 74037 7204
rect 73900 7111 73940 7120
rect 73996 7160 74036 7195
rect 73803 6908 73845 6917
rect 73803 6868 73804 6908
rect 73844 6868 73845 6908
rect 73803 6859 73845 6868
rect 73612 6439 73652 6448
rect 73804 6329 73844 6859
rect 73803 6320 73845 6329
rect 73803 6280 73804 6320
rect 73844 6280 73845 6320
rect 73803 6271 73845 6280
rect 72652 5514 72692 5599
rect 73324 5489 73364 5608
rect 73419 5648 73461 5657
rect 73419 5608 73420 5648
rect 73460 5608 73461 5648
rect 73419 5599 73461 5608
rect 73323 5480 73365 5489
rect 73323 5440 73324 5480
rect 73364 5440 73365 5480
rect 73323 5431 73365 5440
rect 73420 5476 73460 5599
rect 73228 5144 73268 5153
rect 73420 5144 73460 5436
rect 73996 5405 74036 7120
rect 74092 6917 74132 8380
rect 74380 8336 74420 15931
rect 74476 13469 74516 17032
rect 74571 13964 74613 13973
rect 74571 13924 74572 13964
rect 74612 13924 74613 13964
rect 74571 13915 74613 13924
rect 74475 13460 74517 13469
rect 74475 13420 74476 13460
rect 74516 13420 74517 13460
rect 74475 13411 74517 13420
rect 74572 13208 74612 13915
rect 74476 13168 74572 13208
rect 74476 11957 74516 13168
rect 74572 13159 74612 13168
rect 74668 12980 74708 17107
rect 74764 16241 74804 17200
rect 74854 17200 74855 17240
rect 74895 17200 74896 17240
rect 74854 17191 74896 17200
rect 75145 17072 75185 17472
rect 75255 17165 75295 17472
rect 75254 17156 75296 17165
rect 75254 17116 75255 17156
rect 75295 17116 75296 17156
rect 75254 17107 75296 17116
rect 75545 17072 75585 17472
rect 75655 17165 75695 17472
rect 75654 17156 75696 17165
rect 75654 17116 75655 17156
rect 75695 17116 75696 17156
rect 75654 17107 75696 17116
rect 75945 17072 75985 17472
rect 74860 17032 75185 17072
rect 75340 17032 75585 17072
rect 75916 17032 75985 17072
rect 76055 17072 76095 17472
rect 76345 17300 76385 17472
rect 76300 17260 76385 17300
rect 76055 17032 76148 17072
rect 74763 16232 74805 16241
rect 74763 16192 74764 16232
rect 74804 16192 74805 16232
rect 74763 16183 74805 16192
rect 74572 12940 74708 12980
rect 74475 11948 74517 11957
rect 74475 11908 74476 11948
rect 74516 11908 74517 11948
rect 74475 11899 74517 11908
rect 74572 8933 74612 12940
rect 74667 11024 74709 11033
rect 74667 10984 74668 11024
rect 74708 10984 74709 11024
rect 74667 10975 74709 10984
rect 74668 10890 74708 10975
rect 74764 10445 74804 16183
rect 74860 12797 74900 17032
rect 75340 16400 75380 17032
rect 75052 16360 75380 16400
rect 74956 15560 74996 15571
rect 74956 15485 74996 15520
rect 74955 15476 74997 15485
rect 74955 15436 74956 15476
rect 74996 15436 74997 15476
rect 74955 15427 74997 15436
rect 75052 15308 75092 16360
rect 75627 16316 75669 16325
rect 75627 16276 75628 16316
rect 75668 16276 75669 16316
rect 75627 16267 75669 16276
rect 75340 16232 75380 16243
rect 75340 16157 75380 16192
rect 75628 16182 75668 16267
rect 75339 16148 75381 16157
rect 75339 16108 75340 16148
rect 75380 16108 75381 16148
rect 75339 16099 75381 16108
rect 75436 16064 75476 16073
rect 75820 16064 75860 16073
rect 75436 15786 75476 16024
rect 75628 16024 75820 16064
rect 75532 15786 75572 15795
rect 75436 15746 75532 15786
rect 75340 15560 75380 15569
rect 75340 15317 75380 15520
rect 75532 15392 75572 15746
rect 75628 15653 75668 16024
rect 75820 16015 75860 16024
rect 75627 15644 75669 15653
rect 75627 15604 75628 15644
rect 75668 15604 75669 15644
rect 75627 15595 75669 15604
rect 75628 15560 75668 15595
rect 75628 15510 75668 15520
rect 75723 15560 75765 15569
rect 75723 15520 75724 15560
rect 75764 15520 75765 15560
rect 75723 15511 75765 15520
rect 75724 15426 75764 15511
rect 75532 15352 75668 15392
rect 74956 15268 75092 15308
rect 75339 15308 75381 15317
rect 75339 15268 75340 15308
rect 75380 15268 75381 15308
rect 74859 12788 74901 12797
rect 74859 12748 74860 12788
rect 74900 12748 74901 12788
rect 74859 12739 74901 12748
rect 74956 12536 74996 15268
rect 75339 15259 75381 15268
rect 75112 15140 75480 15149
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75112 15091 75480 15100
rect 75339 14972 75381 14981
rect 75339 14932 75340 14972
rect 75380 14932 75476 14972
rect 75339 14923 75381 14932
rect 75436 14888 75476 14932
rect 75436 14839 75476 14848
rect 75340 14804 75380 14813
rect 75244 14720 75284 14729
rect 75244 14057 75284 14680
rect 75340 14225 75380 14764
rect 75532 14762 75572 14771
rect 75435 14720 75477 14729
rect 75435 14680 75436 14720
rect 75476 14680 75477 14720
rect 75435 14671 75477 14680
rect 75436 14552 75476 14671
rect 75532 14636 75572 14722
rect 75628 14762 75668 15352
rect 75916 14981 75956 17032
rect 76012 16316 76052 16325
rect 76012 15905 76052 16276
rect 76108 15989 76148 17032
rect 76204 16064 76244 16073
rect 76107 15980 76149 15989
rect 76107 15940 76108 15980
rect 76148 15940 76149 15980
rect 76107 15931 76149 15940
rect 76011 15896 76053 15905
rect 76011 15856 76012 15896
rect 76052 15856 76053 15896
rect 76011 15847 76053 15856
rect 76012 15308 76052 15317
rect 75915 14972 75957 14981
rect 75915 14932 75916 14972
rect 75956 14932 75957 14972
rect 75915 14923 75957 14932
rect 75628 14713 75668 14722
rect 75915 14720 75957 14729
rect 75915 14680 75916 14720
rect 75956 14680 75957 14720
rect 75915 14671 75957 14680
rect 76012 14720 76052 15268
rect 76107 14804 76149 14813
rect 76107 14764 76108 14804
rect 76148 14764 76149 14804
rect 76107 14755 76149 14764
rect 75627 14636 75669 14645
rect 75532 14596 75628 14636
rect 75668 14596 75669 14636
rect 75627 14587 75669 14596
rect 75916 14586 75956 14671
rect 76012 14645 76052 14680
rect 76108 14720 76148 14755
rect 76108 14669 76148 14680
rect 76204 14720 76244 16024
rect 76204 14645 76244 14680
rect 76300 16064 76340 17260
rect 76455 17072 76495 17472
rect 76745 17072 76785 17472
rect 76855 17333 76895 17472
rect 77145 17333 77185 17472
rect 76854 17324 76896 17333
rect 76854 17284 76855 17324
rect 76895 17284 76896 17324
rect 76854 17275 76896 17284
rect 77144 17324 77186 17333
rect 77144 17284 77145 17324
rect 77185 17284 77186 17324
rect 77144 17275 77186 17284
rect 77255 17072 77295 17472
rect 77545 17072 77585 17472
rect 77655 17072 77695 17472
rect 77835 17156 77877 17165
rect 77835 17116 77836 17156
rect 77876 17116 77877 17156
rect 77835 17107 77877 17116
rect 76455 17032 76532 17072
rect 76745 17032 76820 17072
rect 77255 17032 77300 17072
rect 77545 17032 77588 17072
rect 76396 16064 76436 16073
rect 76300 16024 76396 16064
rect 76011 14636 76053 14645
rect 76011 14596 76012 14636
rect 76052 14596 76053 14636
rect 76011 14587 76053 14596
rect 76203 14636 76245 14645
rect 76203 14596 76204 14636
rect 76244 14596 76245 14636
rect 76203 14587 76245 14596
rect 76012 14556 76052 14587
rect 75436 14512 75572 14552
rect 75339 14216 75381 14225
rect 75339 14176 75340 14216
rect 75380 14176 75381 14216
rect 75339 14167 75381 14176
rect 75243 14048 75285 14057
rect 75243 14008 75244 14048
rect 75284 14008 75285 14048
rect 75243 13999 75285 14008
rect 75112 13628 75480 13637
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75112 13579 75480 13588
rect 75435 13208 75477 13217
rect 75435 13168 75436 13208
rect 75476 13168 75477 13208
rect 75435 13159 75477 13168
rect 75436 13074 75476 13159
rect 75532 12872 75572 14512
rect 76300 14494 76340 16024
rect 76396 16015 76436 16024
rect 76396 15560 76436 15569
rect 76396 14729 76436 15520
rect 76492 15317 76532 17032
rect 76780 15737 76820 17032
rect 76779 15728 76821 15737
rect 76779 15688 76780 15728
rect 76820 15688 76821 15728
rect 76779 15679 76821 15688
rect 76971 15644 77013 15653
rect 76971 15604 76972 15644
rect 77012 15604 77013 15644
rect 76971 15595 77013 15604
rect 76683 15560 76725 15569
rect 76683 15520 76684 15560
rect 76724 15520 76725 15560
rect 76683 15511 76725 15520
rect 76780 15560 76820 15571
rect 76491 15308 76533 15317
rect 76491 15268 76492 15308
rect 76532 15268 76533 15308
rect 76491 15259 76533 15268
rect 76395 14720 76437 14729
rect 76395 14680 76396 14720
rect 76436 14680 76437 14720
rect 76395 14671 76437 14680
rect 76684 14720 76724 15511
rect 76780 15485 76820 15520
rect 76779 15476 76821 15485
rect 76779 15436 76780 15476
rect 76820 15436 76821 15476
rect 76779 15427 76821 15436
rect 76684 14671 76724 14680
rect 76780 14720 76820 14729
rect 76780 14645 76820 14680
rect 76875 14720 76917 14729
rect 76875 14680 76876 14720
rect 76916 14680 76917 14720
rect 76875 14671 76917 14680
rect 76972 14720 77012 15595
rect 77012 14680 77204 14720
rect 76972 14671 77012 14680
rect 76779 14636 76821 14645
rect 76779 14596 76780 14636
rect 76820 14596 76821 14636
rect 76779 14587 76821 14596
rect 76204 14454 76340 14494
rect 76204 14384 76244 14454
rect 76108 14344 76244 14384
rect 76352 14384 76720 14393
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 75819 14216 75861 14225
rect 75819 14176 75820 14216
rect 75860 14176 75861 14216
rect 75819 14167 75861 14176
rect 75820 14082 75860 14167
rect 75723 14048 75765 14057
rect 75723 14008 75724 14048
rect 75764 14008 75765 14048
rect 75723 13999 75765 14008
rect 75916 14048 75956 14057
rect 75724 13914 75764 13999
rect 75916 13292 75956 14008
rect 76011 14048 76053 14057
rect 76011 14008 76012 14048
rect 76052 14008 76053 14048
rect 76011 13999 76053 14008
rect 76012 13914 76052 13999
rect 76011 13292 76053 13301
rect 75916 13252 76012 13292
rect 76052 13252 76053 13292
rect 76011 13243 76053 13252
rect 75915 13124 75957 13133
rect 75915 13084 75916 13124
rect 75956 13084 75957 13124
rect 75915 13075 75957 13084
rect 75532 12832 75668 12872
rect 75435 12788 75477 12797
rect 75435 12748 75436 12788
rect 75476 12748 75572 12788
rect 75435 12739 75477 12748
rect 75051 12704 75093 12713
rect 75051 12664 75052 12704
rect 75092 12664 75093 12704
rect 75051 12655 75093 12664
rect 75052 12570 75092 12655
rect 74860 12496 74996 12536
rect 74763 10436 74805 10445
rect 74763 10396 74764 10436
rect 74804 10396 74805 10436
rect 74763 10387 74805 10396
rect 74571 8924 74613 8933
rect 74571 8884 74572 8924
rect 74612 8884 74613 8924
rect 74571 8875 74613 8884
rect 74572 8790 74612 8875
rect 74475 8756 74517 8765
rect 74475 8716 74476 8756
rect 74516 8716 74517 8756
rect 74475 8707 74517 8716
rect 74476 8672 74516 8707
rect 74476 8621 74516 8632
rect 74188 8296 74420 8336
rect 74091 6908 74133 6917
rect 74091 6868 74092 6908
rect 74132 6868 74133 6908
rect 74091 6859 74133 6868
rect 74091 5648 74133 5657
rect 74091 5608 74092 5648
rect 74132 5608 74133 5648
rect 74091 5599 74133 5608
rect 73995 5396 74037 5405
rect 73995 5356 73996 5396
rect 74036 5356 74037 5396
rect 73995 5347 74037 5356
rect 73268 5104 73460 5144
rect 73228 5095 73268 5104
rect 72459 5060 72501 5069
rect 72459 5020 72460 5060
rect 72500 5020 72501 5060
rect 72459 5011 72501 5020
rect 73132 4976 73172 4985
rect 73132 4733 73172 4936
rect 73995 4976 74037 4985
rect 73995 4936 73996 4976
rect 74036 4936 74037 4976
rect 73995 4927 74037 4936
rect 72939 4724 72981 4733
rect 72939 4684 72940 4724
rect 72980 4684 72981 4724
rect 72939 4675 72981 4684
rect 73131 4724 73173 4733
rect 73131 4684 73132 4724
rect 73172 4684 73173 4724
rect 73131 4675 73173 4684
rect 72940 4590 72980 4675
rect 72556 4304 72596 4313
rect 72596 4264 72692 4304
rect 72556 4255 72596 4264
rect 72172 4087 72212 4096
rect 72268 4136 72308 4145
rect 72076 3977 72116 4059
rect 72075 3968 72117 3977
rect 72075 3924 72076 3968
rect 72116 3924 72117 3968
rect 72075 3919 72117 3924
rect 72076 3915 72116 3919
rect 72268 3809 72308 4096
rect 72555 4052 72597 4061
rect 72555 4012 72556 4052
rect 72596 4012 72597 4052
rect 72555 4003 72597 4012
rect 72267 3800 72309 3809
rect 71980 3760 72212 3800
rect 71883 3632 71925 3641
rect 71883 3592 71884 3632
rect 71924 3592 71925 3632
rect 71883 3583 71925 3592
rect 72075 3212 72117 3221
rect 72075 3172 72076 3212
rect 72116 3172 72117 3212
rect 72075 3163 72117 3172
rect 72076 3078 72116 3163
rect 72172 2900 72212 3760
rect 72267 3760 72268 3800
rect 72308 3760 72309 3800
rect 72267 3751 72309 3760
rect 72460 3464 72500 3473
rect 72172 2860 72308 2900
rect 72076 2801 72116 2832
rect 71980 2792 72020 2801
rect 71884 2708 71924 2717
rect 71596 2575 71636 2584
rect 71787 2624 71829 2633
rect 71787 2584 71788 2624
rect 71828 2584 71829 2624
rect 71787 2575 71829 2584
rect 71308 2490 71348 2575
rect 71404 2456 71444 2465
rect 71884 2456 71924 2668
rect 71444 2416 71924 2456
rect 71404 2407 71444 2416
rect 71980 2372 72020 2752
rect 72075 2792 72117 2801
rect 72075 2752 72076 2792
rect 72116 2752 72117 2792
rect 72075 2743 72117 2752
rect 71212 2071 71252 2080
rect 71500 2332 72020 2372
rect 72076 2708 72116 2743
rect 71404 2036 71444 2045
rect 71500 2036 71540 2332
rect 71444 1996 71540 2036
rect 71404 1987 71444 1996
rect 71787 1952 71829 1961
rect 71787 1912 71788 1952
rect 71828 1912 71829 1952
rect 71787 1903 71829 1912
rect 71115 1868 71157 1877
rect 71115 1828 71116 1868
rect 71156 1828 71157 1868
rect 71115 1819 71157 1828
rect 70732 1315 70772 1324
rect 71116 1121 71156 1819
rect 71788 1818 71828 1903
rect 71212 1700 71252 1709
rect 71212 1205 71252 1660
rect 71499 1532 71541 1541
rect 71499 1492 71500 1532
rect 71540 1492 71541 1532
rect 71499 1483 71541 1492
rect 71211 1196 71253 1205
rect 71211 1156 71212 1196
rect 71252 1156 71253 1196
rect 71211 1147 71253 1156
rect 69772 1063 69812 1072
rect 70060 1112 70100 1121
rect 70252 1112 70292 1121
rect 70100 1072 70252 1112
rect 70060 1063 70100 1072
rect 70252 1063 70292 1072
rect 71115 1112 71157 1121
rect 71115 1072 71116 1112
rect 71156 1072 71157 1112
rect 71115 1063 71157 1072
rect 71500 1112 71540 1483
rect 72076 1457 72116 2668
rect 72171 2624 72213 2633
rect 72171 2584 72172 2624
rect 72212 2584 72213 2624
rect 72171 2575 72213 2584
rect 72172 2490 72212 2575
rect 71691 1448 71733 1457
rect 71691 1408 71692 1448
rect 71732 1408 71733 1448
rect 71691 1399 71733 1408
rect 72075 1448 72117 1457
rect 72075 1408 72076 1448
rect 72116 1408 72117 1448
rect 72075 1399 72117 1408
rect 71595 1364 71637 1373
rect 71595 1324 71596 1364
rect 71636 1324 71637 1364
rect 71595 1315 71637 1324
rect 71500 1063 71540 1072
rect 71596 1112 71636 1315
rect 71596 1063 71636 1072
rect 71692 1112 71732 1399
rect 72268 1364 72308 2860
rect 72363 2792 72405 2801
rect 72363 2752 72364 2792
rect 72404 2752 72405 2792
rect 72363 2743 72405 2752
rect 72364 2658 72404 2743
rect 72460 1541 72500 3424
rect 72556 3464 72596 4003
rect 72652 3893 72692 4264
rect 73131 4136 73173 4145
rect 73996 4136 74036 4927
rect 73131 4096 73132 4136
rect 73172 4096 73173 4136
rect 73131 4087 73173 4096
rect 73804 4096 73996 4136
rect 72748 4052 72788 4061
rect 72651 3884 72693 3893
rect 72651 3844 72652 3884
rect 72692 3844 72693 3884
rect 72651 3835 72693 3844
rect 72556 3415 72596 3424
rect 72652 3464 72692 3835
rect 72748 3632 72788 4012
rect 72748 3583 72788 3592
rect 73035 3632 73077 3641
rect 73035 3592 73036 3632
rect 73076 3592 73077 3632
rect 73035 3583 73077 3592
rect 73036 3498 73076 3583
rect 72652 3415 72692 3424
rect 72940 3464 72980 3473
rect 72940 3221 72980 3424
rect 73132 3305 73172 4087
rect 73516 3464 73556 3473
rect 73556 3424 73748 3464
rect 73516 3415 73556 3424
rect 73131 3296 73173 3305
rect 73131 3256 73132 3296
rect 73172 3256 73173 3296
rect 73131 3247 73173 3256
rect 73611 3296 73653 3305
rect 73611 3256 73612 3296
rect 73652 3256 73653 3296
rect 73611 3247 73653 3256
rect 72939 3212 72981 3221
rect 72939 3172 72940 3212
rect 72980 3172 72981 3212
rect 72939 3163 72981 3172
rect 73420 3212 73460 3221
rect 73420 2900 73460 3172
rect 73132 2860 73460 2900
rect 73132 2792 73172 2860
rect 72844 2752 73172 2792
rect 72747 2708 72789 2717
rect 72747 2668 72748 2708
rect 72788 2668 72789 2708
rect 72747 2659 72789 2668
rect 72652 2624 72692 2633
rect 72652 2129 72692 2584
rect 72748 2624 72788 2659
rect 72844 2633 72884 2752
rect 72748 2573 72788 2584
rect 72843 2624 72885 2633
rect 72843 2584 72844 2624
rect 72884 2584 72885 2624
rect 72843 2575 72885 2584
rect 73132 2624 73172 2633
rect 72844 2452 72884 2575
rect 72844 2403 72884 2412
rect 72651 2120 72693 2129
rect 72651 2080 72652 2120
rect 72692 2080 72693 2120
rect 72651 2071 72693 2080
rect 72651 1952 72693 1961
rect 72651 1912 72652 1952
rect 72692 1912 72693 1952
rect 72651 1903 72693 1912
rect 72652 1818 72692 1903
rect 72459 1532 72501 1541
rect 72459 1492 72460 1532
rect 72500 1492 72501 1532
rect 72459 1483 72501 1492
rect 72268 1315 72308 1324
rect 73132 1121 73172 2584
rect 71692 1063 71732 1072
rect 72843 1112 72885 1121
rect 72843 1072 72844 1112
rect 72884 1072 72885 1112
rect 72843 1063 72885 1072
rect 73131 1112 73173 1121
rect 73131 1072 73132 1112
rect 73172 1072 73173 1112
rect 73131 1063 73173 1072
rect 73612 1112 73652 3247
rect 73708 2372 73748 3424
rect 73804 2876 73844 4096
rect 73996 4087 74036 4096
rect 73995 3800 74037 3809
rect 73995 3760 73996 3800
rect 74036 3760 74037 3800
rect 73995 3751 74037 3760
rect 73996 3632 74036 3751
rect 73996 3583 74036 3592
rect 74092 3464 74132 5599
rect 74188 5144 74228 8296
rect 74379 8168 74421 8177
rect 74379 8128 74380 8168
rect 74420 8128 74421 8168
rect 74379 8119 74421 8128
rect 74283 5816 74325 5825
rect 74283 5776 74284 5816
rect 74324 5776 74325 5816
rect 74283 5767 74325 5776
rect 74284 5648 74324 5767
rect 74380 5657 74420 8119
rect 74860 7160 74900 12496
rect 75112 12116 75480 12125
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75112 12067 75480 12076
rect 75051 11948 75093 11957
rect 75051 11908 75052 11948
rect 75092 11908 75093 11948
rect 75051 11899 75093 11908
rect 75052 11024 75092 11899
rect 75052 10975 75092 10984
rect 75112 10604 75480 10613
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75112 10555 75480 10564
rect 75243 10436 75285 10445
rect 75243 10396 75244 10436
rect 75284 10396 75285 10436
rect 75243 10387 75285 10396
rect 75244 10302 75284 10387
rect 75339 10016 75381 10025
rect 75339 9976 75340 10016
rect 75380 9976 75381 10016
rect 75339 9967 75381 9976
rect 75340 9596 75380 9967
rect 75340 9547 75380 9556
rect 75112 9092 75480 9101
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75112 9043 75480 9052
rect 75532 8765 75572 12748
rect 75051 8756 75093 8765
rect 75051 8716 75052 8756
rect 75092 8716 75093 8756
rect 75051 8707 75093 8716
rect 75531 8756 75573 8765
rect 75531 8716 75532 8756
rect 75572 8716 75573 8756
rect 75531 8707 75573 8716
rect 75052 8168 75092 8707
rect 75052 8119 75092 8128
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 75628 7328 75668 12832
rect 75916 11024 75956 13075
rect 76012 11789 76052 13243
rect 76011 11780 76053 11789
rect 76011 11740 76012 11780
rect 76052 11740 76053 11780
rect 76011 11731 76053 11740
rect 75916 10975 75956 10984
rect 76108 10856 76148 14344
rect 76352 14335 76720 14344
rect 76780 14216 76820 14587
rect 76876 14586 76916 14671
rect 76492 14176 76820 14216
rect 76203 14048 76245 14057
rect 76203 14008 76204 14048
rect 76244 14008 76245 14048
rect 76203 13999 76245 14008
rect 76492 14048 76532 14176
rect 76204 13469 76244 13999
rect 76492 13973 76532 14008
rect 76587 14048 76629 14057
rect 76587 14008 76588 14048
rect 76628 14008 76629 14048
rect 76587 13999 76629 14008
rect 76684 14048 76724 14057
rect 76491 13964 76533 13973
rect 76491 13924 76492 13964
rect 76532 13924 76533 13964
rect 76491 13915 76533 13924
rect 76588 13914 76628 13999
rect 76300 13796 76340 13805
rect 76203 13460 76245 13469
rect 76203 13420 76204 13460
rect 76244 13420 76245 13460
rect 76203 13411 76245 13420
rect 76300 12980 76340 13756
rect 76587 13460 76629 13469
rect 76587 13420 76588 13460
rect 76628 13420 76629 13460
rect 76684 13460 76724 14008
rect 76780 14048 76820 14057
rect 76972 14048 77012 14057
rect 76820 14008 76972 14048
rect 76780 13999 76820 14008
rect 76972 13999 77012 14008
rect 76780 13460 76820 13469
rect 76684 13420 76780 13460
rect 76587 13411 76629 13420
rect 76588 13326 76628 13411
rect 76204 12965 76340 12980
rect 76203 12956 76340 12965
rect 76203 12916 76204 12956
rect 76244 12940 76340 12956
rect 76244 12916 76245 12940
rect 76203 12907 76245 12916
rect 76352 12872 76720 12881
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76352 12823 76720 12832
rect 76395 12704 76437 12713
rect 76780 12704 76820 13420
rect 76875 13376 76917 13385
rect 76875 13336 76876 13376
rect 76916 13336 76917 13376
rect 76875 13327 76917 13336
rect 77067 13376 77109 13385
rect 77067 13336 77068 13376
rect 77108 13336 77109 13376
rect 77067 13327 77109 13336
rect 76395 12664 76396 12704
rect 76436 12664 76437 12704
rect 76395 12655 76437 12664
rect 76684 12664 76820 12704
rect 76396 12536 76436 12655
rect 76396 12487 76436 12496
rect 76492 12452 76532 12461
rect 76492 11948 76532 12412
rect 76684 12452 76724 12664
rect 76779 12536 76821 12545
rect 76779 12496 76780 12536
rect 76820 12496 76821 12536
rect 76779 12487 76821 12496
rect 76684 12403 76724 12412
rect 76780 12402 76820 12487
rect 76588 12368 76628 12377
rect 76588 12284 76628 12328
rect 76876 12284 76916 13327
rect 77068 13208 77108 13327
rect 77164 13301 77204 14680
rect 77260 14393 77300 17032
rect 77355 15476 77397 15485
rect 77355 15436 77356 15476
rect 77396 15436 77397 15476
rect 77355 15427 77397 15436
rect 77259 14384 77301 14393
rect 77259 14344 77260 14384
rect 77300 14344 77301 14384
rect 77259 14335 77301 14344
rect 77356 14057 77396 15427
rect 77548 14309 77588 17032
rect 77644 17032 77695 17072
rect 77644 15905 77684 17032
rect 77836 16484 77876 17107
rect 77945 17072 77985 17472
rect 78055 17072 78095 17472
rect 78345 17156 78385 17472
rect 77836 16435 77876 16444
rect 77932 17032 77985 17072
rect 78028 17032 78095 17072
rect 78316 17116 78385 17156
rect 77740 16232 77780 16241
rect 77643 15896 77685 15905
rect 77643 15856 77644 15896
rect 77684 15856 77685 15896
rect 77643 15847 77685 15856
rect 77740 15737 77780 16192
rect 77836 16064 77876 16073
rect 77739 15728 77781 15737
rect 77739 15688 77740 15728
rect 77780 15688 77781 15728
rect 77739 15679 77781 15688
rect 77644 15560 77684 15569
rect 77547 14300 77589 14309
rect 77547 14260 77548 14300
rect 77588 14260 77589 14300
rect 77547 14251 77589 14260
rect 77644 14057 77684 15520
rect 77740 14729 77780 15679
rect 77836 14813 77876 16024
rect 77932 15149 77972 17032
rect 77931 15140 77973 15149
rect 77931 15100 77932 15140
rect 77972 15100 77973 15140
rect 77931 15091 77973 15100
rect 77835 14804 77877 14813
rect 77835 14764 77836 14804
rect 77876 14764 77877 14804
rect 77835 14755 77877 14764
rect 77739 14720 77781 14729
rect 77739 14680 77740 14720
rect 77780 14680 77781 14720
rect 77739 14671 77781 14680
rect 77355 14048 77397 14057
rect 77355 14008 77356 14048
rect 77396 14008 77397 14048
rect 77355 13999 77397 14008
rect 77643 14048 77685 14057
rect 77643 14008 77644 14048
rect 77684 14008 77685 14048
rect 77643 13999 77685 14008
rect 77356 13914 77396 13999
rect 77451 13964 77493 13973
rect 77451 13924 77452 13964
rect 77492 13924 77493 13964
rect 77451 13915 77493 13924
rect 77163 13292 77205 13301
rect 77163 13252 77164 13292
rect 77204 13252 77205 13292
rect 77163 13243 77205 13252
rect 77068 13159 77108 13168
rect 77164 13208 77204 13243
rect 77164 13158 77204 13168
rect 77260 12982 77300 12991
rect 77259 12916 77260 12965
rect 77300 12916 77301 12965
rect 77259 12907 77301 12916
rect 77260 12847 77300 12907
rect 77164 12536 77204 12545
rect 76588 12244 76916 12284
rect 76972 12496 77164 12536
rect 76492 11899 76532 11908
rect 76683 11780 76725 11789
rect 76683 11740 76684 11780
rect 76724 11740 76725 11780
rect 76683 11731 76725 11740
rect 76492 11696 76532 11705
rect 76492 11528 76532 11656
rect 76684 11696 76724 11731
rect 76684 11645 76724 11656
rect 76780 11696 76820 11705
rect 76972 11696 77012 12496
rect 77164 12487 77204 12496
rect 77260 12536 77300 12545
rect 77452 12536 77492 13915
rect 77547 13376 77589 13385
rect 77547 13336 77548 13376
rect 77588 13336 77589 13376
rect 77547 13327 77589 13336
rect 77835 13376 77877 13385
rect 77835 13336 77836 13376
rect 77876 13336 77877 13376
rect 77835 13327 77877 13336
rect 77548 13208 77588 13327
rect 77548 13159 77588 13168
rect 77644 13208 77684 13217
rect 77644 12980 77684 13168
rect 77739 13208 77781 13217
rect 77739 13168 77740 13208
rect 77780 13168 77781 13208
rect 77739 13159 77781 13168
rect 77836 13208 77876 13327
rect 77836 13159 77876 13168
rect 77740 13074 77780 13159
rect 77644 12940 77780 12980
rect 77644 12536 77684 12545
rect 76820 11656 76916 11696
rect 76780 11647 76820 11656
rect 76492 11488 76820 11528
rect 76352 11360 76720 11369
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76352 11311 76720 11320
rect 76780 11108 76820 11488
rect 76876 11192 76916 11656
rect 76972 11647 77012 11656
rect 77067 11192 77109 11201
rect 76876 11152 77068 11192
rect 77108 11152 77109 11192
rect 77067 11143 77109 11152
rect 76780 11068 77012 11108
rect 75916 10816 76148 10856
rect 75819 10100 75861 10109
rect 75819 10060 75820 10100
rect 75860 10060 75861 10100
rect 75819 10051 75861 10060
rect 75532 7288 75668 7328
rect 75724 9512 75764 9521
rect 74956 7160 74996 7169
rect 74860 7120 74956 7160
rect 74956 6665 74996 7120
rect 75051 7076 75093 7085
rect 75051 7036 75052 7076
rect 75092 7036 75093 7076
rect 75051 7027 75093 7036
rect 74955 6656 74997 6665
rect 74955 6616 74956 6656
rect 74996 6616 74997 6656
rect 74955 6607 74997 6616
rect 74476 6488 74516 6497
rect 74516 6448 74708 6488
rect 74476 6439 74516 6448
rect 74475 5816 74517 5825
rect 74475 5776 74476 5816
rect 74516 5776 74517 5816
rect 74475 5767 74517 5776
rect 74284 5599 74324 5608
rect 74379 5648 74421 5657
rect 74379 5608 74380 5648
rect 74420 5608 74421 5648
rect 74379 5599 74421 5608
rect 74476 5648 74516 5767
rect 74476 5599 74516 5608
rect 74572 5648 74612 5657
rect 74380 5514 74420 5599
rect 74572 5489 74612 5608
rect 74571 5480 74613 5489
rect 74476 5440 74572 5480
rect 74612 5440 74613 5480
rect 74380 5144 74420 5153
rect 74188 5104 74380 5144
rect 74380 5095 74420 5104
rect 74284 4976 74324 4985
rect 74284 4313 74324 4936
rect 74380 4724 74420 4733
rect 74283 4304 74325 4313
rect 74092 2900 74132 3424
rect 74188 4264 74284 4304
rect 74324 4264 74325 4304
rect 74188 3464 74228 4264
rect 74283 4255 74325 4264
rect 74380 4061 74420 4684
rect 74379 4052 74421 4061
rect 74379 4012 74380 4052
rect 74420 4012 74421 4052
rect 74379 4003 74421 4012
rect 74188 3415 74228 3424
rect 74284 3464 74324 3473
rect 74476 3464 74516 5440
rect 74571 5431 74613 5440
rect 74668 4985 74708 6448
rect 74956 5825 74996 6607
rect 75052 6497 75092 7027
rect 75051 6488 75093 6497
rect 75051 6448 75052 6488
rect 75092 6448 75093 6488
rect 75051 6439 75093 6448
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 74955 5816 74997 5825
rect 74955 5776 74956 5816
rect 74996 5776 74997 5816
rect 74955 5767 74997 5776
rect 74572 4976 74612 4985
rect 74572 4481 74612 4936
rect 74667 4976 74709 4985
rect 74667 4936 74668 4976
rect 74708 4936 74709 4976
rect 74667 4927 74709 4936
rect 74956 4976 74996 4985
rect 74571 4472 74613 4481
rect 74571 4432 74572 4472
rect 74612 4432 74613 4472
rect 74571 4423 74613 4432
rect 74956 4229 74996 4936
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 75532 4313 75572 7288
rect 75724 7253 75764 9472
rect 75723 7244 75765 7253
rect 75723 7204 75724 7244
rect 75764 7204 75765 7244
rect 75723 7195 75765 7204
rect 75627 7160 75669 7169
rect 75627 7120 75628 7160
rect 75668 7120 75669 7160
rect 75627 7111 75669 7120
rect 75628 7026 75668 7111
rect 75820 7085 75860 10051
rect 75819 7076 75861 7085
rect 75819 7036 75820 7076
rect 75860 7036 75861 7076
rect 75819 7027 75861 7036
rect 75627 6656 75669 6665
rect 75627 6616 75628 6656
rect 75668 6616 75669 6656
rect 75627 6607 75669 6616
rect 75628 6522 75668 6607
rect 75819 4976 75861 4985
rect 75819 4936 75820 4976
rect 75860 4936 75861 4976
rect 75819 4927 75861 4936
rect 75820 4842 75860 4927
rect 75916 4640 75956 10816
rect 76683 10352 76725 10361
rect 76683 10312 76684 10352
rect 76724 10312 76725 10352
rect 76683 10303 76725 10312
rect 76588 10184 76628 10193
rect 76492 10025 76532 10110
rect 76491 10016 76533 10025
rect 76491 9976 76492 10016
rect 76532 9976 76533 10016
rect 76588 10016 76628 10144
rect 76684 10184 76724 10303
rect 76972 10193 77012 11068
rect 77068 11058 77108 11143
rect 77163 11024 77205 11033
rect 77163 10984 77164 11024
rect 77204 10984 77205 11024
rect 77163 10975 77205 10984
rect 77164 10352 77204 10975
rect 77164 10303 77204 10312
rect 77260 10856 77300 12496
rect 77356 12494 77396 12503
rect 77452 12487 77492 12496
rect 77548 12496 77644 12536
rect 77356 12377 77396 12454
rect 77355 12368 77397 12377
rect 77355 12328 77356 12368
rect 77396 12328 77397 12368
rect 77355 12319 77397 12328
rect 77355 12200 77397 12209
rect 77355 12160 77356 12200
rect 77396 12160 77397 12200
rect 77355 12151 77397 12160
rect 77356 11696 77396 12151
rect 77451 11780 77493 11789
rect 77451 11740 77452 11780
rect 77492 11740 77493 11780
rect 77451 11731 77493 11740
rect 77356 11647 77396 11656
rect 77067 10268 77109 10277
rect 77067 10228 77068 10268
rect 77108 10228 77109 10268
rect 77067 10219 77109 10228
rect 77260 10268 77300 10816
rect 77355 10772 77397 10781
rect 77355 10732 77356 10772
rect 77396 10732 77397 10772
rect 77355 10723 77397 10732
rect 77260 10219 77300 10228
rect 76684 10135 76724 10144
rect 76780 10184 76820 10193
rect 76971 10184 77013 10193
rect 76820 10144 76916 10184
rect 76780 10135 76820 10144
rect 76588 9976 76820 10016
rect 76491 9967 76533 9976
rect 76352 9848 76720 9857
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76352 9799 76720 9808
rect 76780 9680 76820 9976
rect 76876 9932 76916 10144
rect 76971 10144 76972 10184
rect 77012 10144 77013 10184
rect 76971 10135 77013 10144
rect 76972 10050 77012 10135
rect 77068 10134 77108 10219
rect 77356 10184 77396 10723
rect 77356 10135 77396 10144
rect 77355 10016 77397 10025
rect 77355 9976 77356 10016
rect 77396 9976 77397 10016
rect 77355 9967 77397 9976
rect 77067 9932 77109 9941
rect 76876 9892 77068 9932
rect 77108 9892 77109 9932
rect 77067 9883 77109 9892
rect 76492 9640 77012 9680
rect 76492 9008 76532 9640
rect 76588 9512 76628 9521
rect 76628 9472 76820 9512
rect 76588 9463 76628 9472
rect 76492 8968 76628 9008
rect 76491 8840 76533 8849
rect 76491 8800 76492 8840
rect 76532 8800 76533 8840
rect 76491 8791 76533 8800
rect 76395 8756 76437 8765
rect 76395 8716 76396 8756
rect 76436 8716 76437 8756
rect 76395 8707 76437 8716
rect 76300 8672 76340 8681
rect 76300 8513 76340 8632
rect 76396 8622 76436 8707
rect 76492 8706 76532 8791
rect 76588 8756 76628 8968
rect 76588 8707 76628 8716
rect 76780 8681 76820 9472
rect 76875 8840 76917 8849
rect 76875 8800 76876 8840
rect 76916 8800 76917 8840
rect 76875 8791 76917 8800
rect 76684 8672 76724 8681
rect 76684 8513 76724 8632
rect 76779 8672 76821 8681
rect 76779 8632 76780 8672
rect 76820 8632 76821 8672
rect 76779 8623 76821 8632
rect 76876 8672 76916 8791
rect 76876 8623 76916 8632
rect 76299 8504 76341 8513
rect 76299 8464 76300 8504
rect 76340 8464 76341 8504
rect 76299 8455 76341 8464
rect 76683 8504 76725 8513
rect 76683 8464 76684 8504
rect 76724 8464 76725 8504
rect 76780 8504 76820 8623
rect 76780 8464 76916 8504
rect 76683 8455 76725 8464
rect 76352 8336 76720 8345
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76352 8287 76720 8296
rect 76492 8000 76532 8009
rect 76011 7244 76053 7253
rect 76011 7204 76012 7244
rect 76052 7204 76053 7244
rect 76011 7195 76053 7204
rect 76012 7160 76052 7195
rect 76492 7169 76532 7960
rect 76588 8000 76628 8009
rect 76012 7109 76052 7120
rect 76491 7160 76533 7169
rect 76491 7120 76492 7160
rect 76532 7120 76533 7160
rect 76491 7111 76533 7120
rect 76588 6992 76628 7960
rect 76683 8000 76725 8009
rect 76683 7960 76684 8000
rect 76724 7960 76725 8000
rect 76683 7951 76725 7960
rect 76780 8000 76820 8009
rect 76684 7866 76724 7951
rect 76780 7169 76820 7960
rect 76779 7160 76821 7169
rect 76779 7120 76780 7160
rect 76820 7120 76821 7160
rect 76779 7111 76821 7120
rect 76876 7160 76916 8464
rect 76972 7832 77012 9640
rect 76972 7783 77012 7792
rect 76876 7111 76916 7120
rect 76971 7160 77013 7169
rect 76971 7120 76972 7160
rect 77012 7120 77013 7160
rect 76971 7111 77013 7120
rect 76588 6952 76820 6992
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 76780 6656 76820 6952
rect 76588 6616 76820 6656
rect 76492 6488 76532 6497
rect 76011 5732 76053 5741
rect 76011 5692 76012 5732
rect 76052 5692 76053 5732
rect 76011 5683 76053 5692
rect 75628 4600 75956 4640
rect 75147 4304 75189 4313
rect 75147 4264 75148 4304
rect 75188 4264 75189 4304
rect 75147 4255 75189 4264
rect 75531 4304 75573 4313
rect 75531 4264 75532 4304
rect 75572 4264 75573 4304
rect 75531 4255 75573 4264
rect 74955 4220 74997 4229
rect 74955 4180 74956 4220
rect 74996 4180 74997 4220
rect 74955 4171 74997 4180
rect 75148 4170 75188 4255
rect 74324 3424 74516 3464
rect 73804 2827 73844 2836
rect 73996 2860 74132 2900
rect 73996 2456 74036 2860
rect 74092 2633 74132 2718
rect 74284 2717 74324 3424
rect 74571 3044 74613 3053
rect 74571 3004 74572 3044
rect 74612 3004 74613 3044
rect 74571 2995 74613 3004
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 74283 2708 74325 2717
rect 74283 2668 74284 2708
rect 74324 2668 74325 2708
rect 74283 2659 74325 2668
rect 74091 2624 74133 2633
rect 74091 2584 74092 2624
rect 74132 2584 74133 2624
rect 74091 2575 74133 2584
rect 74091 2456 74133 2465
rect 73996 2416 74092 2456
rect 74132 2416 74133 2456
rect 74091 2407 74133 2416
rect 73708 2332 73844 2372
rect 73804 2120 73844 2332
rect 73804 2045 73844 2080
rect 73995 2120 74037 2129
rect 73995 2080 73996 2120
rect 74036 2080 74037 2120
rect 73995 2071 74037 2080
rect 73803 2036 73845 2045
rect 73803 1996 73804 2036
rect 73844 1996 73845 2036
rect 73803 1987 73845 1996
rect 73804 1956 73844 1987
rect 73996 1986 74036 2071
rect 74092 1952 74132 2407
rect 74092 1903 74132 1912
rect 74188 1952 74228 1963
rect 74188 1877 74228 1912
rect 74284 1952 74324 2659
rect 74379 2624 74421 2633
rect 74379 2584 74380 2624
rect 74420 2584 74421 2624
rect 74379 2575 74421 2584
rect 74380 1961 74420 2575
rect 74475 2036 74517 2045
rect 74475 1996 74476 2036
rect 74516 1996 74517 2036
rect 74475 1987 74517 1996
rect 74284 1903 74324 1912
rect 74379 1952 74421 1961
rect 74379 1912 74380 1952
rect 74420 1912 74421 1952
rect 74379 1903 74421 1912
rect 74476 1952 74516 1987
rect 74187 1868 74229 1877
rect 74187 1828 74188 1868
rect 74228 1828 74229 1868
rect 74187 1819 74229 1828
rect 74380 1112 74420 1903
rect 74476 1901 74516 1912
rect 74572 1952 74612 2995
rect 75051 2876 75093 2885
rect 75051 2836 75052 2876
rect 75092 2836 75093 2876
rect 75051 2827 75093 2836
rect 74955 2792 74997 2801
rect 74955 2752 74956 2792
rect 74996 2752 74997 2792
rect 74955 2743 74997 2752
rect 74956 2624 74996 2743
rect 75052 2742 75092 2827
rect 75628 2801 75668 4600
rect 75819 4472 75861 4481
rect 75819 4432 75820 4472
rect 75860 4432 75861 4472
rect 75819 4423 75861 4432
rect 75723 4220 75765 4229
rect 75723 4180 75724 4220
rect 75764 4180 75765 4220
rect 75723 4171 75765 4180
rect 75724 2900 75764 4171
rect 75820 4136 75860 4423
rect 75820 4087 75860 4096
rect 75916 4136 75956 4145
rect 75916 3977 75956 4096
rect 76012 4136 76052 5683
rect 76492 5489 76532 6448
rect 76588 6404 76628 6616
rect 76780 6413 76820 6498
rect 76876 6488 76916 6497
rect 76972 6488 77012 7111
rect 77068 7085 77108 9883
rect 77259 9260 77301 9269
rect 77259 9220 77260 9260
rect 77300 9220 77301 9260
rect 77259 9211 77301 9220
rect 77260 8672 77300 9211
rect 77164 8632 77260 8672
rect 77164 7328 77204 8632
rect 77260 8623 77300 8632
rect 77356 8504 77396 9967
rect 77452 9848 77492 11731
rect 77548 11024 77588 12496
rect 77644 12487 77684 12496
rect 77740 12536 77780 12940
rect 77740 12461 77780 12496
rect 77835 12536 77877 12545
rect 77835 12496 77836 12536
rect 77876 12496 77877 12536
rect 77835 12487 77877 12496
rect 77932 12536 77972 12545
rect 77739 12452 77781 12461
rect 77739 12412 77740 12452
rect 77780 12412 77781 12452
rect 77739 12403 77781 12412
rect 77740 12401 77780 12403
rect 77836 12402 77876 12487
rect 77643 11696 77685 11705
rect 77932 11696 77972 12496
rect 77643 11656 77644 11696
rect 77684 11656 77972 11696
rect 77643 11647 77685 11656
rect 77548 10975 77588 10984
rect 77644 11024 77684 11647
rect 77644 10975 77684 10984
rect 77740 11196 77780 11205
rect 77740 10781 77780 11156
rect 77931 11192 77973 11201
rect 77931 11152 77932 11192
rect 77972 11152 77973 11192
rect 77931 11143 77973 11152
rect 77932 11024 77972 11143
rect 78028 11024 78068 17032
rect 78123 14048 78165 14057
rect 78220 14048 78260 14057
rect 78123 14008 78124 14048
rect 78164 14008 78220 14048
rect 78123 13999 78165 14008
rect 78220 13999 78260 14008
rect 78124 13133 78164 13999
rect 78316 13637 78356 17116
rect 78455 17072 78495 17472
rect 78745 17156 78785 17472
rect 78855 17240 78895 17472
rect 78855 17200 79028 17240
rect 78412 17032 78495 17072
rect 78700 17116 78785 17156
rect 78315 13628 78357 13637
rect 78315 13588 78316 13628
rect 78356 13588 78357 13628
rect 78315 13579 78357 13588
rect 78220 13460 78260 13469
rect 78315 13460 78357 13469
rect 78260 13420 78316 13460
rect 78356 13420 78357 13460
rect 78220 13411 78260 13420
rect 78315 13411 78357 13420
rect 78219 13292 78261 13301
rect 78219 13252 78220 13292
rect 78260 13252 78261 13292
rect 78219 13243 78261 13252
rect 78123 13124 78165 13133
rect 78123 13084 78124 13124
rect 78164 13084 78165 13124
rect 78123 13075 78165 13084
rect 78124 12452 78164 13075
rect 78220 12629 78260 13243
rect 78315 13208 78357 13217
rect 78315 13168 78316 13208
rect 78356 13168 78357 13208
rect 78315 13159 78357 13168
rect 78316 13074 78356 13159
rect 78219 12620 78261 12629
rect 78219 12580 78220 12620
rect 78260 12580 78261 12620
rect 78219 12571 78261 12580
rect 78220 12547 78260 12571
rect 78220 12498 78260 12507
rect 78124 12412 78260 12452
rect 78123 12284 78165 12293
rect 78123 12244 78124 12284
rect 78164 12244 78165 12284
rect 78123 12235 78165 12244
rect 78124 12150 78164 12235
rect 78220 11696 78260 12412
rect 78412 12293 78452 17032
rect 78603 16316 78645 16325
rect 78603 16276 78604 16316
rect 78644 16276 78645 16316
rect 78603 16267 78645 16276
rect 78507 16232 78549 16241
rect 78507 16192 78508 16232
rect 78548 16192 78549 16232
rect 78507 16183 78549 16192
rect 78508 16098 78548 16183
rect 78604 16182 78644 16267
rect 78700 14225 78740 17116
rect 78795 15728 78837 15737
rect 78795 15688 78796 15728
rect 78836 15688 78837 15728
rect 78795 15679 78837 15688
rect 78796 15594 78836 15679
rect 78795 15140 78837 15149
rect 78795 15100 78796 15140
rect 78836 15100 78837 15140
rect 78795 15091 78837 15100
rect 78699 14216 78741 14225
rect 78699 14176 78700 14216
rect 78740 14176 78741 14216
rect 78699 14167 78741 14176
rect 78507 14132 78549 14141
rect 78507 14092 78508 14132
rect 78548 14092 78549 14132
rect 78507 14083 78549 14092
rect 78508 13469 78548 14083
rect 78507 13460 78549 13469
rect 78507 13420 78508 13460
rect 78548 13420 78549 13460
rect 78507 13411 78549 13420
rect 78700 13217 78740 14167
rect 78699 13208 78741 13217
rect 78699 13168 78700 13208
rect 78740 13168 78741 13208
rect 78699 13159 78741 13168
rect 78796 12980 78836 15091
rect 78891 14300 78933 14309
rect 78891 14260 78892 14300
rect 78932 14260 78933 14300
rect 78891 14251 78933 14260
rect 78508 12940 78836 12980
rect 78411 12284 78453 12293
rect 78411 12244 78412 12284
rect 78452 12244 78453 12284
rect 78411 12235 78453 12244
rect 78220 11647 78260 11656
rect 78028 10984 78164 11024
rect 77932 10975 77972 10984
rect 77739 10772 77781 10781
rect 77739 10732 77740 10772
rect 77780 10732 77781 10772
rect 77739 10723 77781 10732
rect 78027 10772 78069 10781
rect 78027 10732 78028 10772
rect 78068 10732 78069 10772
rect 78027 10723 78069 10732
rect 78028 10638 78068 10723
rect 77740 10396 78068 10436
rect 77644 10184 77684 10193
rect 77548 10025 77588 10110
rect 77547 10016 77589 10025
rect 77547 9976 77548 10016
rect 77588 9976 77589 10016
rect 77547 9967 77589 9976
rect 77644 9941 77684 10144
rect 77740 10184 77780 10396
rect 77931 10268 77973 10277
rect 77931 10228 77932 10268
rect 77972 10228 77973 10268
rect 77931 10219 77973 10228
rect 77643 9932 77685 9941
rect 77643 9892 77644 9932
rect 77684 9892 77685 9932
rect 77643 9883 77685 9892
rect 77452 9808 77588 9848
rect 77260 8464 77396 8504
rect 77451 8504 77493 8513
rect 77451 8464 77452 8504
rect 77492 8464 77493 8504
rect 77260 8000 77300 8464
rect 77451 8455 77493 8464
rect 77355 8252 77397 8261
rect 77355 8212 77356 8252
rect 77396 8212 77397 8252
rect 77355 8203 77397 8212
rect 77452 8226 77492 8455
rect 77260 7951 77300 7960
rect 77356 8000 77396 8203
rect 77452 8177 77492 8186
rect 77356 7951 77396 7960
rect 77164 7288 77492 7328
rect 77067 7076 77109 7085
rect 77067 7036 77068 7076
rect 77108 7036 77109 7076
rect 77067 7027 77109 7036
rect 76916 6448 77012 6488
rect 77068 6488 77108 6497
rect 76876 6439 76916 6448
rect 76588 5900 76628 6364
rect 76779 6404 76821 6413
rect 76779 6364 76780 6404
rect 76820 6364 76821 6404
rect 76779 6355 76821 6364
rect 76684 6320 76724 6329
rect 76684 6236 76724 6280
rect 77068 6236 77108 6448
rect 76684 6196 77108 6236
rect 77164 5900 77204 5909
rect 76588 5860 77164 5900
rect 77164 5851 77204 5860
rect 76875 5732 76917 5741
rect 76875 5692 76876 5732
rect 76916 5692 76917 5732
rect 76875 5683 76917 5692
rect 76876 5598 76916 5683
rect 76971 5648 77013 5657
rect 76971 5608 76972 5648
rect 77012 5608 77013 5648
rect 76971 5599 77013 5608
rect 76491 5480 76533 5489
rect 76491 5440 76492 5480
rect 76532 5440 76533 5480
rect 76491 5431 76533 5440
rect 76779 5396 76821 5405
rect 76779 5356 76780 5396
rect 76820 5356 76821 5396
rect 76779 5347 76821 5356
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 76107 4304 76149 4313
rect 76107 4264 76108 4304
rect 76148 4264 76149 4304
rect 76107 4255 76149 4264
rect 76300 4304 76340 4313
rect 76012 4087 76052 4096
rect 76108 4136 76148 4255
rect 75915 3968 75957 3977
rect 75915 3928 75916 3968
rect 75956 3928 75957 3968
rect 75915 3919 75957 3928
rect 75724 2860 75860 2900
rect 75627 2792 75669 2801
rect 75627 2752 75628 2792
rect 75668 2752 75669 2792
rect 75627 2743 75669 2752
rect 74956 2575 74996 2584
rect 75052 2456 75092 2465
rect 74956 2416 75052 2456
rect 74764 1961 74804 2046
rect 74572 1903 74612 1912
rect 74763 1952 74805 1961
rect 74763 1912 74764 1952
rect 74804 1912 74805 1952
rect 74763 1903 74805 1912
rect 74763 1784 74805 1793
rect 74763 1744 74764 1784
rect 74804 1744 74805 1784
rect 74763 1735 74805 1744
rect 74764 1650 74804 1735
rect 74956 1373 74996 2416
rect 75052 2407 75092 2416
rect 75628 1961 75668 2743
rect 75723 2624 75765 2633
rect 75723 2584 75724 2624
rect 75764 2584 75765 2624
rect 75723 2575 75765 2584
rect 75435 1952 75477 1961
rect 75435 1912 75436 1952
rect 75476 1912 75477 1952
rect 75435 1903 75477 1912
rect 75627 1952 75669 1961
rect 75627 1912 75628 1952
rect 75668 1912 75669 1952
rect 75627 1903 75669 1912
rect 75436 1818 75476 1903
rect 75532 1868 75572 1879
rect 75532 1793 75572 1828
rect 75724 1868 75764 2575
rect 75820 2129 75860 2860
rect 76108 2624 76148 4096
rect 76300 3977 76340 4264
rect 76587 4136 76629 4145
rect 76587 4096 76588 4136
rect 76628 4096 76629 4136
rect 76587 4087 76629 4096
rect 76684 4136 76724 4145
rect 76780 4136 76820 5347
rect 76972 5144 77012 5599
rect 77260 5228 77300 7288
rect 77355 7160 77397 7169
rect 77355 7120 77356 7160
rect 77396 7120 77397 7160
rect 77355 7111 77397 7120
rect 76972 4901 77012 5104
rect 77164 5188 77300 5228
rect 77356 5228 77396 7111
rect 77452 6488 77492 7288
rect 77452 6439 77492 6448
rect 77548 5909 77588 9808
rect 77740 9680 77780 10144
rect 77740 9631 77780 9640
rect 77836 10184 77876 10193
rect 77836 8588 77876 10144
rect 77932 9680 77972 10219
rect 78028 10184 78068 10396
rect 78124 10361 78164 10984
rect 78123 10352 78165 10361
rect 78123 10312 78124 10352
rect 78164 10312 78165 10352
rect 78123 10303 78165 10312
rect 78124 10218 78164 10303
rect 78028 10100 78068 10144
rect 78508 10100 78548 12940
rect 78603 10940 78645 10949
rect 78603 10900 78604 10940
rect 78644 10900 78645 10940
rect 78603 10891 78645 10900
rect 78028 10060 78548 10100
rect 78028 9680 78068 9689
rect 77932 9640 78028 9680
rect 78028 9631 78068 9640
rect 78124 9640 78356 9680
rect 77740 8548 77876 8588
rect 77932 9512 77972 9521
rect 77644 7916 77684 7927
rect 77644 7841 77684 7876
rect 77643 7832 77685 7841
rect 77643 7792 77644 7832
rect 77684 7792 77685 7832
rect 77643 7783 77685 7792
rect 77740 6992 77780 8548
rect 77835 8420 77877 8429
rect 77835 8380 77836 8420
rect 77876 8380 77877 8420
rect 77835 8371 77877 8380
rect 77836 8168 77876 8371
rect 77836 8119 77876 8128
rect 77932 7841 77972 9472
rect 78124 9512 78164 9640
rect 78124 9463 78164 9472
rect 78220 9512 78260 9521
rect 78220 8765 78260 9472
rect 78316 9008 78356 9640
rect 78604 9428 78644 10891
rect 78604 9379 78644 9388
rect 78411 9260 78453 9269
rect 78411 9220 78412 9260
rect 78452 9220 78453 9260
rect 78411 9211 78453 9220
rect 78412 9126 78452 9211
rect 78316 8968 78452 9008
rect 78315 8840 78357 8849
rect 78315 8800 78316 8840
rect 78356 8800 78357 8840
rect 78315 8791 78357 8800
rect 78219 8756 78261 8765
rect 78219 8716 78220 8756
rect 78260 8716 78261 8756
rect 78219 8707 78261 8716
rect 78123 8672 78165 8681
rect 78123 8632 78124 8672
rect 78164 8632 78165 8672
rect 78123 8623 78165 8632
rect 78124 8538 78164 8623
rect 78027 8504 78069 8513
rect 78027 8464 78028 8504
rect 78068 8464 78069 8504
rect 78027 8455 78069 8464
rect 78028 8168 78068 8455
rect 78028 8119 78068 8128
rect 78124 8000 78164 8009
rect 78220 8000 78260 8707
rect 78164 7960 78260 8000
rect 78124 7951 78164 7960
rect 77931 7832 77973 7841
rect 77931 7792 77932 7832
rect 77972 7792 77973 7832
rect 77931 7783 77973 7792
rect 77836 7748 77876 7757
rect 77836 7169 77876 7708
rect 77835 7160 77877 7169
rect 77835 7120 77836 7160
rect 77876 7120 77877 7160
rect 77835 7111 77877 7120
rect 78219 7160 78261 7169
rect 78219 7120 78220 7160
rect 78260 7120 78261 7160
rect 78219 7111 78261 7120
rect 78123 7076 78165 7085
rect 78123 7036 78124 7076
rect 78164 7036 78165 7076
rect 78123 7027 78165 7036
rect 78027 6992 78069 7001
rect 77740 6952 77876 6992
rect 77739 6404 77781 6413
rect 77739 6364 77740 6404
rect 77780 6364 77781 6404
rect 77739 6355 77781 6364
rect 77547 5900 77589 5909
rect 77547 5860 77548 5900
rect 77588 5860 77589 5900
rect 77547 5851 77589 5860
rect 77547 5732 77589 5741
rect 77547 5692 77548 5732
rect 77588 5692 77589 5732
rect 77547 5683 77589 5692
rect 77451 5648 77493 5657
rect 77451 5608 77452 5648
rect 77492 5608 77493 5648
rect 77451 5599 77493 5608
rect 77548 5648 77588 5683
rect 77452 5514 77492 5599
rect 77548 5405 77588 5608
rect 77643 5480 77685 5489
rect 77643 5436 77644 5480
rect 77684 5436 77685 5480
rect 77643 5431 77685 5436
rect 77547 5396 77589 5405
rect 77547 5356 77548 5396
rect 77588 5356 77589 5396
rect 77547 5347 77589 5356
rect 77644 5345 77684 5431
rect 77356 5188 77684 5228
rect 77164 5060 77204 5188
rect 77082 5020 77204 5060
rect 76971 4892 77013 4901
rect 77082 4892 77122 5020
rect 76971 4852 76972 4892
rect 77012 4852 77013 4892
rect 76971 4843 77013 4852
rect 77068 4852 77122 4892
rect 77164 4934 77204 4943
rect 77260 4934 77300 4987
rect 76875 4388 76917 4397
rect 76875 4348 76876 4388
rect 76916 4348 76917 4388
rect 76875 4339 76917 4348
rect 76724 4096 76820 4136
rect 76684 4087 76724 4096
rect 76588 4002 76628 4087
rect 76299 3968 76341 3977
rect 76299 3928 76300 3968
rect 76340 3928 76341 3968
rect 76299 3919 76341 3928
rect 76780 3910 76820 3919
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 76683 3548 76725 3557
rect 76683 3508 76684 3548
rect 76724 3508 76725 3548
rect 76683 3499 76725 3508
rect 76684 3464 76724 3499
rect 76780 3473 76820 3870
rect 76299 3296 76341 3305
rect 76299 3256 76300 3296
rect 76340 3256 76341 3296
rect 76299 3247 76341 3256
rect 76300 2900 76340 3247
rect 76108 2465 76148 2584
rect 76204 2860 76340 2900
rect 76204 2624 76244 2860
rect 76588 2792 76628 2801
rect 76588 2633 76628 2752
rect 76204 2575 76244 2584
rect 76299 2624 76341 2633
rect 76299 2584 76300 2624
rect 76340 2584 76341 2624
rect 76299 2575 76341 2584
rect 76587 2624 76629 2633
rect 76587 2584 76588 2624
rect 76628 2584 76629 2624
rect 76587 2575 76629 2584
rect 76300 2490 76340 2575
rect 76396 2465 76436 2550
rect 76107 2456 76149 2465
rect 76107 2416 76108 2456
rect 76148 2416 76149 2456
rect 76107 2407 76149 2416
rect 76395 2456 76437 2465
rect 76395 2416 76396 2456
rect 76436 2416 76437 2456
rect 76684 2456 76724 3424
rect 76779 3464 76821 3473
rect 76779 3424 76780 3464
rect 76820 3424 76821 3464
rect 76779 3415 76821 3424
rect 76779 3296 76821 3305
rect 76779 3256 76780 3296
rect 76820 3256 76821 3296
rect 76779 3247 76821 3256
rect 76780 3162 76820 3247
rect 76876 2792 76916 4339
rect 77068 4304 77108 4852
rect 77164 4397 77204 4894
rect 77259 4894 77260 4901
rect 77356 4976 77396 4985
rect 77300 4894 77301 4901
rect 77259 4892 77301 4894
rect 77259 4852 77260 4892
rect 77300 4852 77301 4892
rect 77259 4843 77301 4852
rect 77163 4388 77205 4397
rect 77163 4348 77164 4388
rect 77204 4348 77205 4388
rect 77163 4339 77205 4348
rect 77356 4313 77396 4936
rect 77452 4976 77492 4985
rect 77355 4304 77397 4313
rect 77068 4229 77135 4304
rect 77355 4264 77356 4304
rect 77396 4264 77397 4304
rect 77355 4255 77397 4264
rect 77067 4220 77135 4229
rect 77067 4180 77068 4220
rect 77108 4180 77300 4220
rect 77067 4171 77109 4180
rect 77260 4136 77300 4180
rect 77452 4145 77492 4936
rect 77356 4136 77396 4145
rect 77260 4096 77356 4136
rect 77356 4087 77396 4096
rect 77451 4136 77493 4145
rect 77451 4096 77452 4136
rect 77492 4096 77493 4136
rect 77451 4087 77493 4096
rect 76972 4052 77012 4061
rect 77012 4012 77204 4052
rect 76972 4003 77012 4012
rect 77067 3884 77109 3893
rect 77067 3844 77068 3884
rect 77108 3844 77109 3884
rect 77067 3835 77109 3844
rect 76971 3464 77013 3473
rect 76971 3424 76972 3464
rect 77012 3424 77013 3464
rect 76971 3415 77013 3424
rect 76972 3330 77012 3415
rect 77068 3380 77108 3835
rect 77068 3331 77108 3340
rect 77164 3296 77204 4012
rect 77356 3464 77396 3473
rect 77548 3464 77588 5188
rect 77644 4976 77684 5188
rect 77740 5144 77780 6355
rect 77836 5741 77876 6952
rect 77932 6952 78028 6992
rect 78068 6952 78069 6992
rect 77835 5732 77877 5741
rect 77835 5692 77836 5732
rect 77876 5692 77877 5732
rect 77835 5683 77877 5692
rect 77836 5648 77876 5683
rect 77836 5598 77876 5608
rect 77932 5648 77972 6952
rect 78027 6943 78069 6952
rect 78028 6858 78068 6943
rect 78124 6740 78164 7027
rect 78220 7026 78260 7111
rect 78316 7076 78356 8791
rect 78412 7328 78452 8968
rect 78412 7288 78644 7328
rect 78412 7160 78452 7288
rect 78412 7111 78452 7120
rect 78508 7160 78548 7169
rect 78316 7027 78356 7036
rect 77932 5599 77972 5608
rect 78028 6700 78164 6740
rect 78028 5648 78068 6700
rect 78508 6665 78548 7120
rect 78507 6656 78549 6665
rect 78507 6616 78508 6656
rect 78548 6616 78549 6656
rect 78507 6607 78549 6616
rect 78316 6488 78356 6497
rect 78220 6448 78316 6488
rect 78028 5599 78068 5608
rect 78123 5648 78165 5657
rect 78123 5608 78124 5648
rect 78164 5608 78165 5648
rect 78123 5599 78165 5608
rect 78124 5514 78164 5599
rect 77740 5095 77780 5104
rect 77835 5060 77877 5069
rect 77835 5020 77836 5060
rect 77876 5020 77877 5060
rect 77835 5011 77877 5020
rect 77644 4927 77684 4936
rect 77836 4976 77876 5011
rect 78220 4985 78260 6448
rect 78316 6439 78356 6448
rect 78412 5648 78452 5657
rect 78508 5648 78548 6607
rect 78452 5608 78548 5648
rect 78412 5599 78452 5608
rect 78315 5480 78357 5489
rect 78315 5440 78316 5480
rect 78356 5440 78357 5480
rect 78315 5431 78357 5440
rect 78316 5346 78356 5431
rect 78604 5069 78644 7288
rect 78700 7160 78740 7169
rect 78892 7160 78932 14251
rect 78988 14141 79028 17200
rect 79145 17072 79185 17472
rect 79255 17165 79295 17472
rect 79254 17156 79296 17165
rect 79254 17116 79255 17156
rect 79295 17116 79296 17156
rect 79254 17107 79296 17116
rect 79545 17072 79585 17472
rect 79145 17032 79220 17072
rect 79083 15896 79125 15905
rect 79083 15856 79084 15896
rect 79124 15856 79125 15896
rect 79083 15847 79125 15856
rect 78987 14132 79029 14141
rect 78987 14092 78988 14132
rect 79028 14092 79029 14132
rect 78987 14083 79029 14092
rect 79084 12980 79124 15847
rect 79180 15737 79220 17032
rect 79468 17032 79585 17072
rect 79655 17072 79695 17472
rect 79655 17032 79700 17072
rect 79468 16484 79508 17032
rect 79468 16435 79508 16444
rect 79371 16316 79413 16325
rect 79660 16316 79700 17032
rect 79371 16276 79372 16316
rect 79412 16276 79700 16316
rect 79371 16267 79413 16276
rect 79372 16232 79412 16267
rect 79372 16182 79412 16192
rect 79179 15728 79221 15737
rect 79179 15688 79180 15728
rect 79220 15688 79221 15728
rect 79179 15679 79221 15688
rect 79371 14216 79413 14225
rect 79371 14176 79372 14216
rect 79412 14176 79413 14216
rect 79371 14167 79413 14176
rect 79372 14082 79412 14167
rect 78988 12940 79124 12980
rect 78988 8009 79028 12940
rect 79371 12536 79413 12545
rect 79371 12496 79372 12536
rect 79412 12496 79413 12536
rect 79371 12487 79413 12496
rect 79372 11948 79412 12487
rect 79372 11899 79412 11908
rect 79275 8756 79317 8765
rect 79275 8716 79276 8756
rect 79316 8716 79317 8756
rect 79275 8707 79317 8716
rect 79276 8622 79316 8707
rect 78987 8000 79029 8009
rect 78987 7960 78988 8000
rect 79028 7960 79029 8000
rect 78987 7951 79029 7960
rect 78740 7120 78932 7160
rect 78700 7001 78740 7120
rect 78699 6992 78741 7001
rect 78699 6952 78700 6992
rect 78740 6952 78741 6992
rect 78699 6943 78741 6952
rect 78796 6992 78836 7001
rect 78988 6992 79028 7951
rect 78836 6952 79028 6992
rect 78796 6943 78836 6952
rect 79467 6656 79509 6665
rect 79467 6616 79468 6656
rect 79508 6616 79509 6656
rect 79467 6607 79509 6616
rect 79468 6522 79508 6607
rect 78603 5060 78645 5069
rect 78603 5020 78604 5060
rect 78644 5020 78645 5060
rect 78603 5011 78645 5020
rect 77643 4808 77685 4817
rect 77643 4768 77644 4808
rect 77684 4768 77685 4808
rect 77643 4759 77685 4768
rect 77644 3725 77684 4759
rect 77643 3716 77685 3725
rect 77643 3676 77644 3716
rect 77684 3676 77685 3716
rect 77643 3667 77685 3676
rect 77396 3424 77588 3464
rect 77356 3415 77396 3424
rect 77164 3247 77204 3256
rect 77260 3380 77300 3389
rect 77260 2876 77300 3340
rect 77356 2876 77396 2885
rect 77260 2836 77356 2876
rect 77356 2827 77396 2836
rect 76876 2752 77004 2792
rect 76964 2717 77004 2752
rect 76964 2708 77013 2717
rect 76964 2668 76972 2708
rect 77012 2668 77013 2708
rect 76971 2659 77013 2668
rect 77163 2708 77205 2717
rect 77163 2668 77164 2708
rect 77204 2668 77205 2708
rect 77163 2659 77205 2668
rect 76876 2624 76916 2633
rect 76684 2416 76820 2456
rect 76395 2407 76437 2416
rect 75819 2120 75861 2129
rect 75819 2080 75820 2120
rect 75860 2080 75861 2120
rect 75819 2071 75861 2080
rect 75819 1952 75861 1961
rect 75819 1912 75820 1952
rect 75860 1912 75861 1952
rect 75819 1903 75861 1912
rect 76012 1952 76052 1961
rect 75724 1819 75764 1828
rect 75820 1818 75860 1903
rect 75531 1784 75573 1793
rect 75531 1744 75532 1784
rect 75572 1744 75573 1784
rect 75531 1735 75573 1744
rect 75628 1784 75668 1793
rect 75628 1700 75668 1744
rect 76012 1700 76052 1912
rect 75628 1660 76052 1700
rect 76108 1541 76148 2407
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 76395 2120 76437 2129
rect 76780 2120 76820 2416
rect 76395 2080 76396 2120
rect 76436 2080 76437 2120
rect 76395 2071 76437 2080
rect 76588 2080 76820 2120
rect 76396 1952 76436 2071
rect 76396 1903 76436 1912
rect 76491 1616 76533 1625
rect 76491 1576 76492 1616
rect 76532 1576 76533 1616
rect 76491 1567 76533 1576
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 75627 1532 75669 1541
rect 75627 1492 75628 1532
rect 75668 1492 75669 1532
rect 75627 1483 75669 1492
rect 76107 1532 76149 1541
rect 76107 1492 76108 1532
rect 76148 1492 76149 1532
rect 76107 1483 76149 1492
rect 74955 1364 74997 1373
rect 74955 1324 74956 1364
rect 74996 1324 74997 1364
rect 74955 1315 74997 1324
rect 75628 1364 75668 1483
rect 75628 1315 75668 1324
rect 74476 1112 74516 1121
rect 74380 1072 74476 1112
rect 73612 1063 73652 1072
rect 74476 1063 74516 1072
rect 76492 1112 76532 1567
rect 76588 1205 76628 2080
rect 76683 1532 76725 1541
rect 76683 1492 76684 1532
rect 76724 1492 76725 1532
rect 76683 1483 76725 1492
rect 76587 1196 76629 1205
rect 76587 1156 76588 1196
rect 76628 1156 76629 1196
rect 76587 1147 76629 1156
rect 76492 1063 76532 1072
rect 76588 1112 76628 1147
rect 71116 978 71156 1063
rect 71787 1028 71829 1037
rect 71787 988 71788 1028
rect 71828 988 71829 1028
rect 71787 979 71829 988
rect 71788 894 71828 979
rect 72844 978 72884 1063
rect 76588 1062 76628 1072
rect 76684 1112 76724 1483
rect 76684 1063 76724 1072
rect 76780 1112 76820 1121
rect 76876 1112 76916 2584
rect 76972 2624 77012 2659
rect 76972 2573 77012 2584
rect 77067 2540 77109 2549
rect 77067 2500 77068 2540
rect 77108 2500 77109 2540
rect 77067 2491 77109 2500
rect 76971 2456 77013 2465
rect 76971 2416 76972 2456
rect 77012 2416 77013 2456
rect 76971 2407 77013 2416
rect 76820 1072 76916 1112
rect 76972 1112 77012 2407
rect 77068 2398 77108 2491
rect 77068 1961 77108 2358
rect 77067 1952 77109 1961
rect 77067 1912 77068 1952
rect 77108 1912 77109 1952
rect 77067 1903 77109 1912
rect 77164 1625 77204 2659
rect 77356 2624 77396 2633
rect 77452 2624 77492 3424
rect 77644 3380 77684 3667
rect 77836 3632 77876 4936
rect 77932 4976 77972 4985
rect 78219 4976 78261 4985
rect 77972 4936 78164 4976
rect 77932 4927 77972 4936
rect 78124 4229 78164 4936
rect 78219 4936 78220 4976
rect 78260 4936 78261 4976
rect 78219 4927 78261 4936
rect 78123 4220 78165 4229
rect 78123 4180 78124 4220
rect 78164 4180 78165 4220
rect 78123 4171 78165 4180
rect 77836 3583 77876 3592
rect 78027 3464 78069 3473
rect 78027 3424 78028 3464
rect 78068 3424 78069 3464
rect 78027 3415 78069 3424
rect 78124 3464 78164 4171
rect 78124 3415 78164 3424
rect 78220 4136 78260 4927
rect 79371 4220 79413 4229
rect 79371 4180 79372 4220
rect 79412 4180 79413 4220
rect 79371 4171 79413 4180
rect 77644 3331 77684 3340
rect 78028 3330 78068 3415
rect 77836 3212 77876 3221
rect 77836 2900 77876 3172
rect 77396 2584 77492 2624
rect 77548 2860 77876 2900
rect 77548 2624 77588 2860
rect 77356 2045 77396 2584
rect 77548 2575 77588 2584
rect 77643 2624 77685 2633
rect 77643 2584 77644 2624
rect 77684 2584 77685 2624
rect 77643 2575 77685 2584
rect 77931 2624 77973 2633
rect 77931 2584 77932 2624
rect 77972 2584 77973 2624
rect 77931 2575 77973 2584
rect 77644 2490 77684 2575
rect 77835 2540 77877 2549
rect 77835 2500 77836 2540
rect 77876 2500 77877 2540
rect 77835 2491 77877 2500
rect 77836 2406 77876 2491
rect 77932 2490 77972 2575
rect 77451 2120 77493 2129
rect 77451 2080 77452 2120
rect 77492 2080 77493 2120
rect 77451 2071 77493 2080
rect 77355 2036 77397 2045
rect 77355 1996 77356 2036
rect 77396 1996 77397 2036
rect 77355 1987 77397 1996
rect 77259 1952 77301 1961
rect 77259 1912 77260 1952
rect 77300 1912 77301 1952
rect 77259 1903 77301 1912
rect 77260 1818 77300 1903
rect 77163 1616 77205 1625
rect 77163 1576 77164 1616
rect 77204 1576 77205 1616
rect 77163 1567 77205 1576
rect 76780 1063 76820 1072
rect 76972 1063 77012 1072
rect 77356 1112 77396 1121
rect 77452 1112 77492 2071
rect 78220 1961 78260 4096
rect 79372 4086 79412 4171
rect 78411 2624 78453 2633
rect 78411 2584 78412 2624
rect 78452 2584 78453 2624
rect 78411 2575 78453 2584
rect 78412 2120 78452 2575
rect 78412 2071 78452 2080
rect 78219 1952 78261 1961
rect 78219 1912 78220 1952
rect 78260 1912 78261 1952
rect 78219 1903 78261 1912
rect 77396 1072 77492 1112
rect 78220 1112 78260 1903
rect 79371 1196 79413 1205
rect 79371 1156 79372 1196
rect 79412 1156 79413 1196
rect 79371 1147 79413 1156
rect 77356 1063 77396 1072
rect 78220 1063 78260 1072
rect 79372 1062 79412 1147
rect 73227 1028 73269 1037
rect 73227 988 73228 1028
rect 73268 988 73269 1028
rect 73227 979 73269 988
rect 73228 894 73268 979
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 69580 38368 69620 38408
rect 652 37528 692 37568
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 844 26524 884 26564
rect 652 25768 692 25808
rect 652 24928 692 24968
rect 844 24508 884 24548
rect 652 24088 692 24128
rect 652 23248 692 23288
rect 940 23248 980 23288
rect 844 23080 884 23120
rect 556 22408 596 22448
rect 652 21568 692 21608
rect 1036 21484 1076 21524
rect 56524 37360 56564 37400
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56236 36772 56276 36812
rect 36652 36688 36692 36728
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 29740 29884 29780 29924
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 7180 25516 7220 25556
rect 2380 25180 2420 25220
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 1804 24760 1844 24800
rect 2380 24760 2420 24800
rect 2188 24508 2228 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 1996 23836 2036 23876
rect 2188 23836 2228 23876
rect 1516 23080 1556 23120
rect 1612 22996 1652 23036
rect 1708 20896 1748 20936
rect 652 20728 692 20768
rect 1900 20728 1940 20768
rect 1516 20560 1556 20600
rect 652 19888 692 19928
rect 1228 19468 1268 19508
rect 748 19300 788 19340
rect 1708 20056 1748 20096
rect 652 19048 692 19088
rect 1324 18964 1364 19004
rect 1228 18712 1268 18752
rect 652 18208 692 18248
rect 556 17536 596 17576
rect 460 16024 500 16064
rect 460 7708 500 7748
rect 652 17368 692 17408
rect 652 15688 692 15728
rect 652 14848 692 14888
rect 652 14008 692 14048
rect 652 13168 692 13208
rect 652 12328 692 12368
rect 652 11488 692 11528
rect 652 10732 692 10772
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 652 8128 692 8168
rect 652 7288 692 7328
rect 1612 18712 1652 18752
rect 1804 19972 1844 20012
rect 844 15352 884 15392
rect 1324 17788 1364 17828
rect 1132 17536 1172 17576
rect 1132 17284 1172 17324
rect 1708 17956 1748 17996
rect 1036 16528 1076 16568
rect 844 13252 884 13292
rect 844 13000 884 13040
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 13708 23836 13748 23876
rect 3628 22996 3668 23036
rect 7084 22996 7124 23036
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 3340 21484 3380 21524
rect 2764 21316 2804 21356
rect 3532 21316 3572 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 3532 20980 3572 21020
rect 3340 20896 3380 20936
rect 2860 20812 2900 20852
rect 3244 20812 3284 20852
rect 2764 20644 2804 20684
rect 2764 19468 2804 19508
rect 2188 19300 2228 19340
rect 2092 18628 2132 18668
rect 1996 17284 2036 17324
rect 844 11740 884 11780
rect 844 11488 884 11528
rect 844 10312 884 10352
rect 844 9388 884 9428
rect 1708 16276 1748 16316
rect 1516 15352 1556 15392
rect 1516 13252 1556 13292
rect 1516 13000 1556 13040
rect 1516 11740 1556 11780
rect 1420 11572 1460 11612
rect 1708 15436 1748 15476
rect 1708 13924 1748 13964
rect 1708 13252 1748 13292
rect 1708 12412 1748 12452
rect 1708 11740 1748 11780
rect 940 7708 980 7748
rect 652 6448 692 6488
rect 844 5692 884 5732
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 1516 10312 1556 10352
rect 1708 10228 1748 10268
rect 2668 16948 2708 16988
rect 1612 5692 1652 5732
rect 844 4180 884 4220
rect 1420 4180 1460 4220
rect 652 3928 692 3968
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3916 21568 3956 21608
rect 4588 21568 4628 21608
rect 4012 21484 4052 21524
rect 4492 21484 4532 21524
rect 3820 21148 3860 21188
rect 3916 20980 3956 21020
rect 4108 21316 4148 21356
rect 4012 20896 4052 20936
rect 3724 20476 3764 20516
rect 4012 20476 4052 20516
rect 4012 20140 4052 20180
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 3628 19636 3668 19676
rect 3724 19552 3764 19592
rect 2956 19300 2996 19340
rect 3340 19468 3380 19508
rect 4204 20980 4244 21020
rect 4396 20644 4436 20684
rect 5068 21484 5108 21524
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 4204 20224 4244 20264
rect 4684 20224 4724 20264
rect 4492 20140 4532 20180
rect 4300 20056 4340 20096
rect 4684 19888 4724 19928
rect 4492 19552 4532 19592
rect 3628 19216 3668 19256
rect 5932 21400 5972 21440
rect 5356 21232 5396 21272
rect 5260 20728 5300 20768
rect 5356 20644 5396 20684
rect 7372 21568 7412 21608
rect 7660 21568 7700 21608
rect 6796 20896 6836 20936
rect 7660 20896 7700 20936
rect 6412 20812 6452 20852
rect 6316 20728 6356 20768
rect 5932 20560 5972 20600
rect 5260 20056 5300 20096
rect 5068 19804 5108 19844
rect 5356 19552 5396 19592
rect 4300 19132 4340 19172
rect 3532 18628 3572 18668
rect 3436 18544 3476 18584
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3916 18460 3956 18500
rect 3724 18376 3764 18416
rect 3628 18292 3668 18332
rect 3532 17872 3572 17912
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 2860 15436 2900 15476
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4108 18544 4148 18584
rect 4012 18376 4052 18416
rect 4492 19216 4532 19256
rect 4684 19216 4724 19256
rect 4396 19048 4436 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 4684 18544 4724 18584
rect 4588 18460 4628 18500
rect 4972 19216 5012 19256
rect 4780 18376 4820 18416
rect 5068 18544 5108 18584
rect 6220 20056 6260 20096
rect 6412 20308 6452 20348
rect 6892 20812 6932 20852
rect 7372 20812 7412 20852
rect 6700 20056 6740 20096
rect 6700 19636 6740 19676
rect 5068 17872 5108 17912
rect 4204 17788 4244 17828
rect 4108 17620 4148 17660
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 5164 17704 5204 17744
rect 5068 17284 5108 17324
rect 4012 16948 4052 16988
rect 4012 16192 4052 16232
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3628 10228 3668 10268
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 6508 19048 6548 19088
rect 6892 20056 6932 20096
rect 6796 19552 6836 19592
rect 6892 19468 6932 19508
rect 6796 19216 6836 19256
rect 6220 18460 6260 18500
rect 6124 17620 6164 17660
rect 6028 17368 6068 17408
rect 6412 18376 6452 18416
rect 6220 17284 6260 17324
rect 7084 19468 7124 19508
rect 7468 20728 7508 20768
rect 7564 20140 7604 20180
rect 7276 19300 7316 19340
rect 7468 19048 7508 19088
rect 7564 18964 7604 19004
rect 7468 18712 7508 18752
rect 7948 21568 7988 21608
rect 9004 21568 9044 21608
rect 10540 21568 10580 21608
rect 8140 21400 8180 21440
rect 8140 21232 8180 21272
rect 10156 21064 10196 21104
rect 10252 20896 10292 20936
rect 10156 20812 10196 20852
rect 8428 20728 8468 20768
rect 9292 20140 9332 20180
rect 9772 20140 9812 20180
rect 7948 20056 7988 20096
rect 8140 19804 8180 19844
rect 8524 20056 8564 20096
rect 8428 19804 8468 19844
rect 9964 19804 10004 19844
rect 8620 19636 8660 19676
rect 9868 19636 9908 19676
rect 9388 19468 9428 19508
rect 9772 19468 9812 19508
rect 8332 19216 8372 19256
rect 8044 18964 8084 19004
rect 7084 18628 7124 18668
rect 7564 18628 7604 18668
rect 6988 18376 7028 18416
rect 6796 18208 6836 18248
rect 7372 18544 7412 18584
rect 7660 18544 7700 18584
rect 8332 18460 8372 18500
rect 9004 18460 9044 18500
rect 8140 18376 8180 18416
rect 7852 18292 7892 18332
rect 6604 17620 6644 17660
rect 5260 17032 5300 17072
rect 6796 17284 6836 17324
rect 6316 17200 6356 17240
rect 6124 16948 6164 16988
rect 6316 16192 6356 16232
rect 6508 17032 6548 17072
rect 6700 17032 6740 17072
rect 7084 17284 7124 17324
rect 6988 17200 7028 17240
rect 7084 17032 7124 17072
rect 6988 16276 7028 16316
rect 6124 11740 6164 11780
rect 8140 17788 8180 17828
rect 7564 17536 7604 17576
rect 8332 17704 8372 17744
rect 7468 17368 7508 17408
rect 8140 17368 8180 17408
rect 10060 19216 10100 19256
rect 10252 20140 10292 20180
rect 10444 20224 10484 20264
rect 10636 21064 10676 21104
rect 11020 20812 11060 20852
rect 10636 20056 10676 20096
rect 10924 20560 10964 20600
rect 10828 19804 10868 19844
rect 10252 19384 10292 19424
rect 12460 21568 12500 21608
rect 11596 21400 11636 21440
rect 12940 21232 12980 21272
rect 13612 21232 13652 21272
rect 11692 20896 11732 20936
rect 12076 20140 12116 20180
rect 11116 19552 11156 19592
rect 10444 19216 10484 19256
rect 9868 19048 9908 19088
rect 10252 19084 10292 19088
rect 10252 19048 10292 19084
rect 9772 18712 9812 18752
rect 10732 18628 10772 18668
rect 9964 17704 10004 17744
rect 10732 18376 10772 18416
rect 9868 17620 9908 17660
rect 10060 17116 10100 17156
rect 10348 18292 10388 18332
rect 10636 18292 10676 18332
rect 10252 18040 10292 18080
rect 10156 16948 10196 16988
rect 10060 16864 10100 16904
rect 9484 16276 9524 16316
rect 9388 13924 9428 13964
rect 10348 17536 10388 17576
rect 10348 17116 10388 17156
rect 10444 16864 10484 16904
rect 10924 18544 10964 18584
rect 10828 18040 10868 18080
rect 10732 17704 10772 17744
rect 10924 17704 10964 17744
rect 10828 17620 10868 17660
rect 11116 18712 11156 18752
rect 11212 17956 11252 17996
rect 11980 19216 12020 19256
rect 11788 18544 11828 18584
rect 11308 17704 11348 17744
rect 11500 17620 11540 17660
rect 11020 17536 11060 17576
rect 11020 17032 11060 17072
rect 11500 16948 11540 16988
rect 10540 16276 10580 16316
rect 11020 16276 11060 16316
rect 10348 16024 10388 16064
rect 13612 20980 13652 21020
rect 12940 19468 12980 19508
rect 12364 19384 12404 19424
rect 28780 23752 28820 23792
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 14284 21400 14324 21440
rect 13708 20896 13748 20936
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 13516 19552 13556 19592
rect 13420 19384 13460 19424
rect 12556 19216 12596 19256
rect 12460 18796 12500 18836
rect 12748 19216 12788 19256
rect 12460 18628 12500 18668
rect 13132 19216 13172 19256
rect 13036 18796 13076 18836
rect 12940 18628 12980 18668
rect 12748 18376 12788 18416
rect 13036 18208 13076 18248
rect 12172 17956 12212 17996
rect 13132 17956 13172 17996
rect 13036 17704 13076 17744
rect 13132 17536 13172 17576
rect 13612 18628 13652 18668
rect 31660 27868 31700 27908
rect 31468 27532 31508 27572
rect 31084 22492 31124 22532
rect 30124 22240 30164 22280
rect 29740 21484 29780 21524
rect 30892 21652 30932 21692
rect 30508 21484 30548 21524
rect 30124 21400 30164 21440
rect 29932 21316 29972 21356
rect 27628 20728 27668 20768
rect 28780 20728 28820 20768
rect 16108 20476 16148 20516
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 16972 20056 17012 20096
rect 26956 20056 26996 20096
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 28492 20140 28532 20180
rect 27916 20056 27956 20096
rect 16108 19300 16148 19340
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 15340 18712 15380 18752
rect 13900 18544 13940 18584
rect 14956 18544 14996 18584
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 15244 18376 15284 18416
rect 15436 18292 15476 18332
rect 16972 18544 17012 18584
rect 27628 18544 27668 18584
rect 18124 18376 18164 18416
rect 16108 18208 16148 18248
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 18124 18040 18164 18080
rect 13708 17872 13748 17912
rect 14956 17872 14996 17912
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 12940 17032 12980 17072
rect 13324 17032 13364 17072
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 28300 17200 28340 17240
rect 28780 17200 28820 17240
rect 29164 17200 29204 17240
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 27628 15520 27668 15560
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 11980 13252 12020 13292
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 10252 12412 10292 12452
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 30412 21316 30452 21356
rect 30316 20644 30356 20684
rect 29644 20392 29684 20432
rect 30508 20896 30548 20936
rect 30508 20560 30548 20600
rect 30700 20056 30740 20096
rect 30892 20392 30932 20432
rect 31276 21568 31316 21608
rect 31468 22240 31508 22280
rect 31468 21652 31508 21692
rect 33196 27700 33236 27740
rect 32044 23332 32084 23372
rect 32236 22324 32276 22364
rect 36460 25264 36500 25304
rect 34924 24592 34964 24632
rect 36364 24592 36404 24632
rect 33772 23080 33812 23120
rect 35212 24508 35252 24548
rect 36460 24508 36500 24548
rect 36364 24172 36404 24212
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55468 36184 55508 36224
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 55084 35260 55124 35300
rect 56716 36772 56756 36812
rect 56524 36688 56564 36728
rect 56428 36100 56468 36140
rect 56044 35932 56084 35972
rect 55948 35260 55988 35300
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 51724 34504 51764 34544
rect 52108 34504 52148 34544
rect 50764 34336 50804 34376
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 50476 33664 50516 33704
rect 49324 33412 49364 33452
rect 50476 33412 50516 33452
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 49804 32656 49844 32696
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 46636 30220 46676 30260
rect 47980 30220 48020 30260
rect 48172 30220 48212 30260
rect 40588 29968 40628 30008
rect 40396 29884 40436 29924
rect 40588 29632 40628 29672
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 39916 29296 39956 29336
rect 40684 29296 40724 29336
rect 39724 29044 39764 29084
rect 40108 28876 40148 28916
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 40492 28876 40532 28916
rect 41068 28876 41108 28916
rect 40300 28372 40340 28412
rect 40780 28288 40820 28328
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 39628 27616 39668 27656
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 40204 27112 40244 27152
rect 38380 26944 38420 26984
rect 36940 25936 36980 25976
rect 37708 25264 37748 25304
rect 37804 25096 37844 25136
rect 38668 26776 38708 26816
rect 40396 27028 40436 27068
rect 40108 26944 40148 26984
rect 40492 26944 40532 26984
rect 39436 26776 39476 26816
rect 39724 26776 39764 26816
rect 40012 26860 40052 26900
rect 40876 27616 40916 27656
rect 40780 27196 40820 27236
rect 40588 26860 40628 26900
rect 40780 26860 40820 26900
rect 40204 26776 40244 26816
rect 40108 26608 40148 26648
rect 38668 25936 38708 25976
rect 38188 25096 38228 25136
rect 36652 24424 36692 24464
rect 37228 24256 37268 24296
rect 37036 24088 37076 24128
rect 35596 23668 35636 23708
rect 36364 23668 36404 23708
rect 35308 23164 35348 23204
rect 31756 21652 31796 21692
rect 31852 21568 31892 21608
rect 31756 21484 31796 21524
rect 31660 20728 31700 20768
rect 31372 20644 31412 20684
rect 30988 20224 31028 20264
rect 31180 20224 31220 20264
rect 30796 19888 30836 19928
rect 31372 20140 31412 20180
rect 29836 19132 29876 19172
rect 30892 19048 30932 19088
rect 31468 20056 31508 20096
rect 31852 20560 31892 20600
rect 31756 20224 31796 20264
rect 33196 21988 33236 22028
rect 32428 20728 32468 20768
rect 32236 20560 32276 20600
rect 32140 20140 32180 20180
rect 32812 20728 32852 20768
rect 33004 20728 33044 20768
rect 33484 21988 33524 22028
rect 33292 20728 33332 20768
rect 32812 20560 32852 20600
rect 33484 20728 33524 20768
rect 33388 20392 33428 20432
rect 32524 20224 32564 20264
rect 33964 22324 34004 22364
rect 35884 23332 35924 23372
rect 35788 23164 35828 23204
rect 35692 23080 35732 23120
rect 35500 22156 35540 22196
rect 33964 20812 34004 20852
rect 33676 20560 33716 20600
rect 33196 19888 33236 19928
rect 32428 19300 32468 19340
rect 31564 19132 31604 19172
rect 32236 19132 32276 19172
rect 32236 18544 32276 18584
rect 32428 18208 32468 18248
rect 31948 17956 31988 17996
rect 32140 17956 32180 17996
rect 31756 17788 31796 17828
rect 30220 17704 30260 17744
rect 31180 16780 31220 16820
rect 31660 16360 31700 16400
rect 32236 17872 32276 17912
rect 32140 17704 32180 17744
rect 32620 19216 32660 19256
rect 32812 18628 32852 18668
rect 35308 21568 35348 21608
rect 35500 21568 35540 21608
rect 35404 20896 35444 20936
rect 35212 20728 35252 20768
rect 35980 23248 36020 23288
rect 35980 22408 36020 22448
rect 36748 23584 36788 23624
rect 36748 23416 36788 23456
rect 37036 23416 37076 23456
rect 36940 23248 36980 23288
rect 38092 24592 38132 24632
rect 37900 24088 37940 24128
rect 38092 24004 38132 24044
rect 37612 23920 37652 23960
rect 37996 23920 38036 23960
rect 37324 23584 37364 23624
rect 37228 23164 37268 23204
rect 37036 23080 37076 23120
rect 36748 22492 36788 22532
rect 36268 22240 36308 22280
rect 37228 22324 37268 22364
rect 35692 21988 35732 22028
rect 36748 21988 36788 22028
rect 35788 21316 35828 21356
rect 36556 21316 36596 21356
rect 37132 22240 37172 22280
rect 37036 22072 37076 22112
rect 36940 21652 36980 21692
rect 37228 21652 37268 21692
rect 37036 21568 37076 21608
rect 37132 21316 37172 21356
rect 36268 20728 36308 20768
rect 36172 20560 36212 20600
rect 36748 20560 36788 20600
rect 37036 20728 37076 20768
rect 38092 23836 38132 23876
rect 38284 23836 38324 23876
rect 38476 24676 38516 24716
rect 38572 24592 38612 24632
rect 38476 24088 38516 24128
rect 38476 23668 38516 23708
rect 37804 23332 37844 23372
rect 37516 23248 37556 23288
rect 37420 22324 37460 22364
rect 37708 23164 37748 23204
rect 39628 26104 39668 26144
rect 39532 25936 39572 25976
rect 39436 25852 39476 25892
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 39628 25852 39668 25892
rect 40396 26776 40436 26816
rect 40300 26692 40340 26732
rect 40876 26776 40916 26816
rect 40492 26692 40532 26732
rect 40780 26692 40820 26732
rect 40588 26608 40628 26648
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 40396 26188 40436 26228
rect 39820 25264 39860 25304
rect 40108 25768 40148 25808
rect 39340 25096 39380 25136
rect 39628 25096 39668 25136
rect 38956 24676 38996 24716
rect 38860 24256 38900 24296
rect 38668 24172 38708 24212
rect 38668 24004 38708 24044
rect 39724 24592 39764 24632
rect 39916 24760 39956 24800
rect 39628 24256 39668 24296
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 38860 23920 38900 23960
rect 38764 23584 38804 23624
rect 37420 22072 37460 22112
rect 37612 21988 37652 22028
rect 37420 21652 37460 21692
rect 37708 21568 37748 21608
rect 39244 23836 39284 23876
rect 38956 23668 38996 23708
rect 39436 23584 39476 23624
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 39436 21988 39476 22028
rect 37900 21400 37940 21440
rect 38284 21400 38324 21440
rect 37420 20812 37460 20852
rect 34636 20140 34676 20180
rect 33964 19972 34004 20012
rect 33484 19552 33524 19592
rect 33580 19468 33620 19508
rect 33388 19300 33428 19340
rect 33196 19216 33236 19256
rect 34540 19804 34580 19844
rect 34252 19468 34292 19508
rect 33772 19384 33812 19424
rect 33100 18880 33140 18920
rect 33196 18712 33236 18752
rect 33388 18964 33428 19004
rect 33580 18880 33620 18920
rect 32716 18460 32756 18500
rect 33292 18544 33332 18584
rect 33196 18292 33236 18332
rect 33100 18040 33140 18080
rect 33388 17956 33428 17996
rect 32524 17872 32564 17912
rect 33772 19216 33812 19256
rect 33676 18712 33716 18752
rect 33676 18040 33716 18080
rect 32908 17872 32948 17912
rect 32236 17536 32276 17576
rect 32236 17284 32276 17324
rect 32044 17116 32084 17156
rect 32236 16360 32276 16400
rect 32044 16192 32084 16232
rect 32812 17704 32852 17744
rect 33292 17788 33332 17828
rect 33100 17704 33140 17744
rect 32524 17284 32564 17324
rect 32812 17284 32852 17324
rect 32716 17116 32756 17156
rect 33004 17284 33044 17324
rect 33580 17704 33620 17744
rect 34060 19216 34100 19256
rect 33964 19132 34004 19172
rect 33964 18712 34004 18752
rect 33292 17032 33332 17072
rect 33004 16948 33044 16988
rect 33196 16948 33236 16988
rect 32620 16360 32660 16400
rect 33100 16360 33140 16400
rect 32908 15520 32948 15560
rect 33868 17536 33908 17576
rect 33868 17368 33908 17408
rect 36556 20056 36596 20096
rect 35788 19888 35828 19928
rect 34636 19216 34676 19256
rect 34828 19216 34868 19256
rect 35692 19216 35732 19256
rect 35692 18880 35732 18920
rect 34540 18712 34580 18752
rect 34252 18544 34292 18584
rect 34636 18544 34676 18584
rect 34444 18460 34484 18500
rect 34348 18292 34388 18332
rect 34348 18124 34388 18164
rect 33676 16360 33716 16400
rect 33388 16192 33428 16232
rect 34540 18208 34580 18248
rect 34444 17788 34484 17828
rect 34444 17368 34484 17408
rect 34348 15772 34388 15812
rect 34732 18292 34772 18332
rect 34636 17704 34676 17744
rect 35308 16948 35348 16988
rect 37036 20056 37076 20096
rect 36652 19468 36692 19508
rect 36556 19384 36596 19424
rect 36268 19216 36308 19256
rect 35980 18544 36020 18584
rect 36460 18460 36500 18500
rect 35980 17872 36020 17912
rect 37132 19888 37172 19928
rect 37132 18712 37172 18752
rect 37324 19216 37364 19256
rect 37516 19804 37556 19844
rect 37612 19468 37652 19508
rect 37612 19216 37652 19256
rect 37420 18964 37460 19004
rect 36556 17536 36596 17576
rect 36172 17284 36212 17324
rect 36460 17284 36500 17324
rect 35980 16612 36020 16652
rect 35788 16276 35828 16316
rect 35116 15688 35156 15728
rect 34444 15436 34484 15476
rect 37708 18712 37748 18752
rect 36364 16360 36404 16400
rect 36268 16192 36308 16232
rect 35692 16024 35732 16064
rect 35692 15520 35732 15560
rect 35980 15692 36020 15728
rect 35980 15688 36020 15692
rect 36172 15688 36212 15728
rect 35884 15604 35924 15644
rect 36364 15604 36404 15644
rect 37324 17032 37364 17072
rect 36940 16948 36980 16988
rect 37516 17704 37556 17744
rect 37612 17284 37652 17324
rect 37804 17032 37844 17072
rect 37420 16360 37460 16400
rect 36844 16192 36884 16232
rect 37612 16108 37652 16148
rect 36748 16024 36788 16064
rect 37036 15604 37076 15644
rect 32044 15184 32084 15224
rect 33292 15184 33332 15224
rect 34828 15184 34868 15224
rect 34444 14680 34484 14720
rect 34924 14680 34964 14720
rect 36556 15520 36596 15560
rect 36748 15436 36788 15476
rect 38092 19384 38132 19424
rect 38092 19216 38132 19256
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 39820 23248 39860 23288
rect 40972 26356 41012 26396
rect 40876 26272 40916 26312
rect 40780 25852 40820 25892
rect 42508 28708 42548 28748
rect 41644 28372 41684 28412
rect 41548 27196 41588 27236
rect 41452 26776 41492 26816
rect 41068 26188 41108 26228
rect 40972 25936 41012 25976
rect 40780 25180 40820 25220
rect 40588 25096 40628 25136
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 41068 25096 41108 25136
rect 40876 24844 40916 24884
rect 41068 24676 41108 24716
rect 41356 25348 41396 25388
rect 41260 24592 41300 24632
rect 41260 24004 41300 24044
rect 40876 23920 40916 23960
rect 41068 23920 41108 23960
rect 40972 23836 41012 23876
rect 40108 23668 40148 23708
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 40780 23332 40820 23372
rect 40012 23080 40052 23120
rect 40012 22408 40052 22448
rect 39820 21904 39860 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 40300 21652 40340 21692
rect 41068 23584 41108 23624
rect 40972 22996 41012 23036
rect 40876 22240 40916 22280
rect 40780 21568 40820 21608
rect 40108 21400 40148 21440
rect 40588 20728 40628 20768
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 38668 19552 38708 19592
rect 38860 19468 38900 19508
rect 39244 19384 39284 19424
rect 39532 19384 39572 19424
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 40204 20224 40244 20264
rect 40684 20224 40724 20264
rect 40588 20140 40628 20180
rect 40492 20056 40532 20096
rect 40108 19972 40148 20012
rect 40780 20140 40820 20180
rect 40972 21568 41012 21608
rect 40972 20728 41012 20768
rect 40780 19972 40820 20012
rect 41164 23248 41204 23288
rect 41452 24088 41492 24128
rect 41452 23752 41492 23792
rect 41356 23584 41396 23624
rect 41260 22576 41300 22616
rect 41260 21400 41300 21440
rect 41164 21316 41204 21356
rect 39916 19636 39956 19676
rect 42316 28372 42356 28412
rect 42796 29128 42836 29168
rect 42892 28792 42932 28832
rect 42700 28624 42740 28664
rect 43180 28708 43220 28748
rect 43276 28624 43316 28664
rect 42796 28540 42836 28580
rect 43084 28540 43124 28580
rect 41836 26860 41876 26900
rect 41644 26776 41684 26816
rect 41740 25516 41780 25556
rect 41932 26020 41972 26060
rect 42508 28036 42548 28076
rect 42220 27952 42260 27992
rect 42124 27616 42164 27656
rect 42604 27616 42644 27656
rect 43180 28456 43220 28496
rect 43084 28372 43124 28412
rect 42988 28036 43028 28076
rect 43276 28288 43316 28328
rect 43180 27952 43220 27992
rect 42508 26776 42548 26816
rect 43084 26776 43124 26816
rect 44140 29128 44180 29168
rect 45388 29128 45428 29168
rect 44044 28288 44084 28328
rect 43372 27784 43412 27824
rect 43660 27616 43700 27656
rect 46444 29044 46484 29084
rect 45388 28960 45428 29000
rect 44332 28624 44372 28664
rect 43756 27448 43796 27488
rect 43372 27280 43412 27320
rect 43372 26944 43412 26984
rect 42796 26440 42836 26480
rect 42412 26272 42452 26312
rect 42988 26272 43028 26312
rect 42796 26020 42836 26060
rect 42124 25936 42164 25976
rect 42316 25516 42356 25556
rect 42508 25516 42548 25556
rect 42124 25348 42164 25388
rect 42796 25768 42836 25808
rect 42604 25348 42644 25388
rect 42796 25264 42836 25304
rect 42028 25180 42068 25220
rect 42700 25180 42740 25220
rect 43468 26272 43508 26312
rect 43660 26272 43700 26312
rect 44140 27616 44180 27656
rect 44236 27532 44276 27572
rect 45196 28540 45236 28580
rect 44908 28204 44948 28244
rect 44332 27448 44372 27488
rect 46156 28288 46196 28328
rect 45196 27616 45236 27656
rect 44428 27364 44468 27404
rect 44908 27364 44948 27404
rect 44716 26356 44756 26396
rect 43084 26020 43124 26060
rect 42316 24592 42356 24632
rect 41836 24172 41876 24212
rect 41644 24088 41684 24128
rect 41740 24004 41780 24044
rect 42796 24676 42836 24716
rect 43276 25432 43316 25472
rect 43084 25264 43124 25304
rect 43660 26104 43700 26144
rect 44044 26104 44084 26144
rect 43564 26020 43604 26060
rect 43756 26020 43796 26060
rect 43660 25936 43700 25976
rect 43564 25600 43604 25640
rect 43468 25432 43508 25472
rect 43084 23920 43124 23960
rect 42700 23836 42740 23876
rect 41644 23332 41684 23372
rect 42412 23248 42452 23288
rect 41644 23080 41684 23120
rect 41548 22576 41588 22616
rect 41548 22408 41588 22448
rect 42796 23752 42836 23792
rect 42700 23500 42740 23540
rect 42508 22996 42548 23036
rect 42412 22912 42452 22952
rect 41452 22240 41492 22280
rect 41836 22240 41876 22280
rect 42508 22828 42548 22868
rect 42508 22240 42548 22280
rect 42412 22156 42452 22196
rect 42316 22072 42356 22112
rect 42988 23752 43028 23792
rect 42892 23584 42932 23624
rect 43276 23752 43316 23792
rect 42796 23248 42836 23288
rect 43084 23332 43124 23372
rect 42988 23248 43028 23288
rect 42604 22072 42644 22112
rect 42796 22996 42836 23036
rect 42988 23080 43028 23120
rect 44428 26104 44468 26144
rect 44332 25936 44372 25976
rect 44524 26020 44564 26060
rect 44812 26104 44852 26144
rect 45772 26356 45812 26396
rect 45196 26272 45236 26312
rect 45388 26272 45428 26312
rect 45196 26104 45236 26144
rect 45196 25936 45236 25976
rect 44908 25852 44948 25892
rect 44908 25600 44948 25640
rect 44620 25180 44660 25220
rect 45004 25264 45044 25304
rect 44140 25096 44180 25136
rect 44908 25096 44948 25136
rect 43468 23836 43508 23876
rect 43564 23752 43604 23792
rect 43180 23080 43220 23120
rect 45196 24928 45236 24968
rect 44908 24592 44948 24632
rect 45100 24592 45140 24632
rect 44332 24340 44372 24380
rect 44908 24340 44948 24380
rect 44140 23920 44180 23960
rect 44140 23752 44180 23792
rect 43852 23584 43892 23624
rect 44044 23584 44084 23624
rect 44428 23836 44468 23876
rect 44236 23500 44276 23540
rect 45004 23584 45044 23624
rect 45196 24508 45236 24548
rect 42892 22912 42932 22952
rect 43084 22912 43124 22952
rect 43372 22912 43412 22952
rect 42892 22408 42932 22448
rect 42124 21736 42164 21776
rect 42604 21736 42644 21776
rect 41740 21652 41780 21692
rect 43180 22828 43220 22868
rect 43468 22492 43508 22532
rect 42892 21736 42932 21776
rect 43372 22240 43412 22280
rect 45388 25852 45428 25892
rect 45868 26104 45908 26144
rect 45964 25936 46004 25976
rect 45484 25600 45524 25640
rect 45676 25600 45716 25640
rect 45676 25264 45716 25304
rect 45580 25180 45620 25220
rect 45484 25096 45524 25136
rect 45388 25012 45428 25052
rect 43198 22072 43238 22112
rect 43852 22072 43892 22112
rect 45292 22240 45332 22280
rect 43852 21904 43892 21944
rect 45004 21904 45044 21944
rect 42220 21568 42260 21608
rect 42412 21568 42452 21608
rect 42796 21568 42836 21608
rect 42316 21400 42356 21440
rect 41740 20392 41780 20432
rect 43084 21568 43124 21608
rect 43660 21568 43700 21608
rect 44236 21736 44276 21776
rect 43852 20812 43892 20852
rect 42220 20224 42260 20264
rect 42412 20228 42452 20264
rect 42412 20224 42452 20228
rect 42700 20224 42740 20264
rect 41356 20140 41396 20180
rect 42796 20140 42836 20180
rect 40300 19552 40340 19592
rect 40396 19468 40436 19508
rect 40972 19468 41012 19508
rect 38284 19132 38324 19172
rect 39436 19216 39476 19256
rect 38764 19132 38804 19172
rect 39052 19132 39092 19172
rect 38380 18964 38420 19004
rect 38188 18880 38228 18920
rect 38188 18208 38228 18248
rect 38188 17704 38228 17744
rect 38284 17536 38324 17576
rect 38380 17284 38420 17324
rect 37996 16948 38036 16988
rect 37900 16612 37940 16652
rect 37900 16276 37940 16316
rect 38092 16108 38132 16148
rect 38572 17032 38612 17072
rect 38476 16612 38516 16652
rect 38092 15772 38132 15812
rect 37996 15604 38036 15644
rect 37900 15520 37940 15560
rect 37036 14596 37076 14636
rect 37324 14764 37364 14804
rect 37708 14764 37748 14804
rect 37420 14680 37460 14720
rect 34828 14008 34868 14048
rect 37036 14008 37076 14048
rect 38380 15604 38420 15644
rect 38668 15772 38708 15812
rect 39532 19132 39572 19172
rect 39340 18292 39380 18332
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 39628 18544 39668 18584
rect 40108 19300 40148 19340
rect 39820 19048 39860 19088
rect 40108 18712 40148 18752
rect 39052 17032 39092 17072
rect 39148 16948 39188 16988
rect 38956 16780 38996 16820
rect 38764 15436 38804 15476
rect 38668 14848 38708 14888
rect 38284 14680 38324 14720
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 39340 15520 39380 15560
rect 40108 17452 40148 17492
rect 40300 19216 40340 19256
rect 40780 19300 40820 19340
rect 40684 19216 40724 19256
rect 40492 19084 40532 19088
rect 40492 19048 40532 19084
rect 40780 18964 40820 19004
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 40684 18712 40724 18752
rect 40396 18376 40436 18416
rect 40300 17788 40340 17828
rect 40684 17788 40724 17828
rect 40492 17704 40532 17744
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 39724 17200 39764 17240
rect 40396 17032 40436 17072
rect 39724 16780 39764 16820
rect 41164 19384 41204 19424
rect 41068 18964 41108 19004
rect 40972 18796 41012 18836
rect 40876 18460 40916 18500
rect 41452 19384 41492 19424
rect 41260 18964 41300 19004
rect 41356 18796 41396 18836
rect 41740 19972 41780 20012
rect 42316 19888 42356 19928
rect 41740 19216 41780 19256
rect 42796 19888 42836 19928
rect 42700 19384 42740 19424
rect 42124 19132 42164 19172
rect 42604 19132 42644 19172
rect 41548 18880 41588 18920
rect 42316 18796 42356 18836
rect 41164 18376 41204 18416
rect 40684 16780 40724 16820
rect 40492 16528 40532 16568
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 39628 15604 39668 15644
rect 40876 16780 40916 16820
rect 41068 16192 41108 16232
rect 41164 16024 41204 16064
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 38956 14596 38996 14636
rect 39340 14344 39380 14384
rect 39916 15520 39956 15560
rect 40396 15520 40436 15560
rect 40780 15520 40820 15560
rect 41548 18376 41588 18416
rect 41452 16612 41492 16652
rect 39916 14848 39956 14888
rect 39724 14176 39764 14216
rect 39916 14092 39956 14132
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 39244 13252 39284 13292
rect 38764 13168 38804 13208
rect 39532 13168 39572 13208
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 40780 14260 40820 14300
rect 40396 14180 40436 14216
rect 40396 14176 40436 14180
rect 40300 14092 40340 14132
rect 40684 14092 40724 14132
rect 40204 14008 40244 14048
rect 40588 14008 40628 14048
rect 41068 14176 41108 14216
rect 41356 14344 41396 14384
rect 40876 13924 40916 13964
rect 41260 14008 41300 14048
rect 40108 13252 40148 13292
rect 41356 13168 41396 13208
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 42028 18628 42068 18668
rect 41740 17704 41780 17744
rect 42220 17788 42260 17828
rect 42028 17200 42068 17240
rect 42988 20728 43028 20768
rect 43660 20140 43700 20180
rect 44140 20140 44180 20180
rect 44044 20056 44084 20096
rect 43948 19552 43988 19592
rect 43372 19468 43412 19508
rect 42892 19216 42932 19256
rect 43084 18628 43124 18668
rect 42412 18460 42452 18500
rect 42796 18502 42836 18542
rect 43276 18376 43316 18416
rect 42988 18292 43028 18332
rect 43179 18124 43219 18164
rect 42412 17956 42452 17996
rect 42988 17956 43028 17996
rect 43564 18796 43604 18836
rect 44044 19216 44084 19256
rect 44620 20896 44660 20936
rect 44524 20812 44564 20852
rect 44332 19384 44372 19424
rect 43948 18712 43988 18752
rect 44140 18712 44180 18752
rect 43468 18460 43508 18500
rect 44524 18292 44564 18332
rect 45868 23080 45908 23120
rect 47404 29800 47444 29840
rect 46636 29044 46676 29084
rect 46636 28288 46676 28328
rect 46924 29128 46964 29168
rect 47404 29296 47444 29336
rect 48172 29212 48212 29252
rect 47404 29044 47444 29084
rect 47308 28960 47348 29000
rect 47884 29128 47924 29168
rect 48076 29128 48116 29168
rect 47980 29044 48020 29084
rect 47788 27784 47828 27824
rect 50860 33832 50900 33872
rect 51340 33832 51380 33872
rect 50572 32572 50612 32612
rect 50188 31564 50228 31604
rect 50476 31480 50516 31520
rect 48748 29800 48788 29840
rect 49516 29800 49556 29840
rect 48652 29212 48692 29252
rect 48940 29128 48980 29168
rect 48844 29044 48884 29084
rect 48364 27952 48404 27992
rect 47404 27616 47444 27656
rect 47308 27280 47348 27320
rect 47212 26860 47252 26900
rect 46444 25684 46484 25724
rect 46060 24340 46100 24380
rect 46252 23752 46292 23792
rect 46060 23164 46100 23204
rect 46636 25936 46676 25976
rect 47692 27196 47732 27236
rect 48076 27196 48116 27236
rect 47692 26860 47732 26900
rect 47116 25852 47156 25892
rect 46924 25768 46964 25808
rect 47308 25684 47348 25724
rect 47596 25684 47636 25724
rect 47212 25600 47252 25640
rect 46924 25432 46964 25472
rect 46636 24424 46676 24464
rect 46540 22996 46580 23036
rect 46060 22324 46100 22364
rect 45004 20056 45044 20096
rect 45100 19132 45140 19172
rect 45004 19048 45044 19088
rect 44908 18712 44948 18752
rect 43468 17872 43508 17912
rect 44044 17872 44084 17912
rect 43084 17704 43124 17744
rect 43468 17704 43508 17744
rect 44236 17788 44276 17828
rect 42508 17536 42548 17576
rect 42412 17032 42452 17072
rect 42316 16612 42356 16652
rect 43180 17536 43220 17576
rect 43372 17572 43412 17576
rect 43372 17536 43412 17572
rect 43756 17536 43796 17576
rect 44140 17704 44180 17744
rect 44620 18040 44660 18080
rect 44812 17788 44852 17828
rect 44620 17536 44660 17576
rect 44620 17368 44660 17408
rect 43660 17032 43700 17072
rect 44140 17032 44180 17072
rect 42892 16864 42932 16904
rect 43564 16864 43604 16904
rect 44140 16864 44180 16904
rect 43468 16696 43508 16736
rect 44428 17032 44468 17072
rect 44332 16612 44372 16652
rect 42412 16192 42452 16232
rect 42796 16108 42836 16148
rect 42220 14680 42260 14720
rect 42988 15520 43028 15560
rect 43468 15520 43508 15560
rect 43084 15352 43124 15392
rect 42892 15268 42932 15308
rect 43180 15268 43220 15308
rect 42316 14260 42356 14300
rect 42220 14176 42260 14216
rect 42028 14092 42068 14132
rect 42700 14680 42740 14720
rect 43084 14680 43124 14720
rect 43276 14680 43316 14720
rect 42604 14344 42644 14384
rect 41548 12580 41588 12620
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 41260 11572 41300 11612
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 41740 13252 41780 13292
rect 41836 13168 41876 13208
rect 42892 14092 42932 14132
rect 42796 13924 42836 13964
rect 42796 13756 42836 13796
rect 42412 11572 42452 11612
rect 41452 11236 41492 11276
rect 42700 11320 42740 11360
rect 42604 10984 42644 11024
rect 43852 14344 43892 14384
rect 44428 14260 44468 14300
rect 43276 13924 43316 13964
rect 43660 13924 43700 13964
rect 43084 13756 43124 13796
rect 43276 12496 43316 12536
rect 43276 12160 43316 12200
rect 43468 12160 43508 12200
rect 43564 12076 43604 12116
rect 44716 16948 44756 16988
rect 44812 14428 44852 14468
rect 45100 18712 45140 18752
rect 45868 22072 45908 22112
rect 45964 21736 46004 21776
rect 46540 22324 46580 22364
rect 46156 21736 46196 21776
rect 46540 22156 46580 22196
rect 46828 23080 46868 23120
rect 47404 25432 47444 25472
rect 47788 25432 47828 25472
rect 47116 23836 47156 23876
rect 47116 23164 47156 23204
rect 47308 23752 47348 23792
rect 48076 26776 48116 26816
rect 48556 27616 48596 27656
rect 48364 27364 48404 27404
rect 48556 27280 48596 27320
rect 48172 25936 48212 25976
rect 48460 26776 48500 26816
rect 48364 26692 48404 26732
rect 48268 25516 48308 25556
rect 47980 25180 48020 25220
rect 47500 24592 47540 24632
rect 47692 24592 47732 24632
rect 47596 24508 47636 24548
rect 47500 23752 47540 23792
rect 48172 25264 48212 25304
rect 48268 25180 48308 25220
rect 48460 25264 48500 25304
rect 48268 24508 48308 24548
rect 48844 27700 48884 27740
rect 48748 27616 48788 27656
rect 48844 27448 48884 27488
rect 48652 26356 48692 26396
rect 49900 29800 49940 29840
rect 50380 31312 50420 31352
rect 52204 34420 52244 34460
rect 53068 34420 53108 34460
rect 52300 34336 52340 34376
rect 52108 33664 52148 33704
rect 51916 33496 51956 33536
rect 51532 33412 51572 33452
rect 52012 33412 52052 33452
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 50956 33076 50996 33116
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 52300 33412 52340 33452
rect 51340 32908 51380 32948
rect 51244 32824 51284 32864
rect 50860 32656 50900 32696
rect 52204 33076 52244 33116
rect 51532 32908 51572 32948
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 52972 33832 53012 33872
rect 56140 34588 56180 34628
rect 56620 36268 56660 36308
rect 57004 37360 57044 37400
rect 56908 36940 56948 36980
rect 56716 35848 56756 35888
rect 56620 35764 56660 35804
rect 57580 37360 57620 37400
rect 57292 37276 57332 37316
rect 57484 37192 57524 37232
rect 57964 37192 58004 37232
rect 57580 36940 57620 36980
rect 57484 36688 57524 36728
rect 57292 36268 57332 36308
rect 57100 36184 57140 36224
rect 57100 35848 57140 35888
rect 56620 35596 56660 35636
rect 56812 35596 56852 35636
rect 55948 34504 55988 34544
rect 54124 34336 54164 34376
rect 55180 34336 55220 34376
rect 55468 34336 55508 34376
rect 56044 34336 56084 34376
rect 53452 33664 53492 33704
rect 53836 33664 53876 33704
rect 56140 34252 56180 34292
rect 54316 34084 54356 34124
rect 56044 34084 56084 34124
rect 54316 33832 54356 33872
rect 55084 33832 55124 33872
rect 54124 33412 54164 33452
rect 53068 33076 53108 33116
rect 53836 33076 53876 33116
rect 52972 32992 53012 33032
rect 53644 32908 53684 32948
rect 54028 32908 54068 32948
rect 52012 32572 52052 32612
rect 50956 31480 50996 31520
rect 50764 31228 50804 31268
rect 50956 31228 50996 31268
rect 50188 30640 50228 30680
rect 50380 30304 50420 30344
rect 50668 30640 50708 30680
rect 50476 29632 50516 29672
rect 49708 28960 49748 29000
rect 49516 28876 49556 28916
rect 49132 27364 49172 27404
rect 49228 27112 49268 27152
rect 49420 27112 49460 27152
rect 49036 26692 49076 26732
rect 49132 26608 49172 26648
rect 49036 26104 49076 26144
rect 49036 25852 49076 25892
rect 48940 25768 48980 25808
rect 48940 24592 48980 24632
rect 48844 24424 48884 24464
rect 48556 24088 48596 24128
rect 48364 23416 48404 23456
rect 47212 22240 47252 22280
rect 47020 21820 47060 21860
rect 46924 21736 46964 21776
rect 46924 21568 46964 21608
rect 47404 22156 47444 22196
rect 47212 21652 47252 21692
rect 46444 21484 46484 21524
rect 47500 21484 47540 21524
rect 47404 21316 47444 21356
rect 48748 23752 48788 23792
rect 48652 23416 48692 23456
rect 48844 23416 48884 23456
rect 48940 23080 48980 23120
rect 48844 22240 48884 22280
rect 48460 21820 48500 21860
rect 47692 21316 47732 21356
rect 46060 20812 46100 20852
rect 45772 20056 45812 20096
rect 45580 19384 45620 19424
rect 46540 19468 46580 19508
rect 45484 19300 45524 19340
rect 45868 19216 45908 19256
rect 45772 18964 45812 19004
rect 45292 18880 45332 18920
rect 45196 18460 45236 18500
rect 45388 18460 45428 18500
rect 45100 18292 45140 18332
rect 45100 17704 45140 17744
rect 45004 16948 45044 16988
rect 45484 17032 45524 17072
rect 45388 16696 45428 16736
rect 46348 18880 46388 18920
rect 47212 20728 47252 20768
rect 47788 20728 47828 20768
rect 46828 19636 46868 19676
rect 47884 20140 47924 20180
rect 47500 19552 47540 19592
rect 47212 19468 47252 19508
rect 46732 19384 46772 19424
rect 47116 19384 47156 19424
rect 46732 19216 46772 19256
rect 46636 19132 46676 19172
rect 47020 19132 47060 19172
rect 46924 18880 46964 18920
rect 46156 18292 46196 18332
rect 46540 18712 46580 18752
rect 46444 17704 46484 17744
rect 46348 17452 46388 17492
rect 47020 18544 47060 18584
rect 46732 17704 46772 17744
rect 46252 17032 46292 17072
rect 45004 16360 45044 16400
rect 45580 16024 45620 16064
rect 45964 16780 46004 16820
rect 45964 16528 46004 16568
rect 46060 16276 46100 16316
rect 45868 16060 45908 16064
rect 45868 16024 45908 16060
rect 45868 15856 45908 15896
rect 46252 16192 46292 16232
rect 45004 15268 45044 15308
rect 45676 14764 45716 14804
rect 45388 14596 45428 14636
rect 45580 14680 45620 14720
rect 45484 14428 45524 14468
rect 45868 14596 45908 14636
rect 45772 14344 45812 14384
rect 45196 14176 45236 14216
rect 45100 14092 45140 14132
rect 44620 13084 44660 13124
rect 44044 12664 44084 12704
rect 44620 12664 44660 12704
rect 43948 12580 43988 12620
rect 44428 12580 44468 12620
rect 43756 12496 43796 12536
rect 44044 12328 44084 12368
rect 43852 12244 43892 12284
rect 43660 11740 43700 11780
rect 43276 11320 43316 11360
rect 43852 11488 43892 11528
rect 42796 11068 42836 11108
rect 43276 11068 43316 11108
rect 42988 10984 43028 11024
rect 43372 10900 43412 10940
rect 43372 10732 43412 10772
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 42604 10312 42644 10352
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 43276 10312 43316 10352
rect 43660 11068 43700 11108
rect 43756 10984 43796 11024
rect 44428 12328 44468 12368
rect 45004 13168 45044 13208
rect 44908 13084 44948 13124
rect 44812 13000 44852 13040
rect 44716 12244 44756 12284
rect 44620 12076 44660 12116
rect 44428 11488 44468 11528
rect 44332 11236 44372 11276
rect 44428 11068 44468 11108
rect 44140 10732 44180 10772
rect 43468 10228 43508 10268
rect 43084 10144 43124 10184
rect 43564 10144 43604 10184
rect 44044 10144 44084 10184
rect 44236 10144 44276 10184
rect 43852 10060 43892 10100
rect 42988 9976 43028 10016
rect 29452 9388 29492 9428
rect 31756 9388 31796 9428
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 44620 9304 44660 9344
rect 44812 10144 44852 10184
rect 45292 13168 45332 13208
rect 45580 14008 45620 14048
rect 45868 13168 45908 13208
rect 45484 13000 45524 13040
rect 45868 13000 45908 13040
rect 45388 12748 45428 12788
rect 45100 10312 45140 10352
rect 46924 17368 46964 17408
rect 46636 16276 46676 16316
rect 46828 16948 46868 16988
rect 47980 19972 48020 20012
rect 47500 19132 47540 19172
rect 47308 18544 47348 18584
rect 47212 18292 47252 18332
rect 47116 17368 47156 17408
rect 47020 16864 47060 16904
rect 46924 16528 46964 16568
rect 47116 16780 47156 16820
rect 46924 16192 46964 16232
rect 46732 15856 46772 15896
rect 46636 15604 46676 15644
rect 46348 15436 46388 15476
rect 47596 19048 47636 19088
rect 47500 17704 47540 17744
rect 47404 17452 47444 17492
rect 47308 17032 47348 17072
rect 47404 16948 47444 16988
rect 47212 16612 47252 16652
rect 47308 16276 47348 16316
rect 47596 16192 47636 16232
rect 48268 19300 48308 19340
rect 48748 20056 48788 20096
rect 48556 19300 48596 19340
rect 48076 19242 48116 19256
rect 48076 19216 48116 19242
rect 48844 19048 48884 19088
rect 48652 18796 48692 18836
rect 48556 18544 48596 18584
rect 48556 18040 48596 18080
rect 47980 17620 48020 17660
rect 48748 18040 48788 18080
rect 48748 17872 48788 17912
rect 48652 17704 48692 17744
rect 48556 17536 48596 17576
rect 47404 16024 47444 16064
rect 47500 15520 47540 15560
rect 47788 15520 47828 15560
rect 48268 15520 48308 15560
rect 46828 15436 46868 15476
rect 46924 15352 46964 15392
rect 47308 15436 47348 15476
rect 48076 15436 48116 15476
rect 47884 15352 47924 15392
rect 46636 14764 46676 14804
rect 46828 14764 46868 14804
rect 46252 14260 46292 14300
rect 46060 14176 46100 14216
rect 46348 14176 46388 14216
rect 46156 12832 46196 12872
rect 45964 12748 46004 12788
rect 45964 12580 46004 12620
rect 46060 12496 46100 12536
rect 46732 14092 46772 14132
rect 46540 14008 46580 14048
rect 46924 14344 46964 14384
rect 47020 14176 47060 14216
rect 47212 14260 47252 14300
rect 47116 14008 47156 14048
rect 46732 13336 46772 13376
rect 46828 13168 46868 13208
rect 47020 13336 47060 13376
rect 46540 13084 46580 13124
rect 46444 13000 46484 13040
rect 45772 11824 45812 11864
rect 45676 10984 45716 11024
rect 45868 11488 45908 11528
rect 47980 14008 48020 14048
rect 48268 14344 48308 14384
rect 49132 25516 49172 25556
rect 49228 25264 49268 25304
rect 49132 25180 49172 25220
rect 49804 26524 49844 26564
rect 50380 28624 50420 28664
rect 49996 28288 50036 28328
rect 50284 27280 50324 27320
rect 49996 26104 50036 26144
rect 49900 25516 49940 25556
rect 49804 25432 49844 25472
rect 49228 24760 49268 24800
rect 49420 24760 49460 24800
rect 49228 24256 49268 24296
rect 49132 23080 49172 23120
rect 49324 24088 49364 24128
rect 49324 23920 49364 23960
rect 50092 25264 50132 25304
rect 51340 31564 51380 31604
rect 51436 31312 51476 31352
rect 51436 30976 51476 31016
rect 50956 30220 50996 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 50956 29632 50996 29672
rect 51628 29884 51668 29924
rect 51532 29800 51572 29840
rect 51916 31564 51956 31604
rect 51820 31323 51860 31352
rect 51820 31312 51860 31323
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 52780 32152 52820 32192
rect 53356 32824 53396 32864
rect 53164 32740 53204 32780
rect 53068 31732 53108 31772
rect 52396 31564 52436 31604
rect 52492 31480 52532 31520
rect 52588 31396 52628 31436
rect 52012 31144 52052 31184
rect 51820 31060 51860 31100
rect 51148 29464 51188 29504
rect 52012 30976 52052 31016
rect 50956 29128 50996 29168
rect 50764 29044 50804 29084
rect 51436 29128 51476 29168
rect 51244 28960 51284 29000
rect 51532 29044 51572 29084
rect 50764 28792 50804 28832
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 50860 28624 50900 28664
rect 50860 27028 50900 27068
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 50956 26692 50996 26732
rect 50764 26188 50804 26228
rect 50572 25852 50612 25892
rect 50380 25768 50420 25808
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 50572 25348 50612 25388
rect 51628 28792 51668 28832
rect 52684 31312 52724 31352
rect 52300 31228 52340 31268
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 51916 28624 51956 28664
rect 51820 28288 51860 28328
rect 51724 27112 51764 27152
rect 51724 26608 51764 26648
rect 49804 24508 49844 24548
rect 50284 24760 50324 24800
rect 50668 25264 50708 25304
rect 50476 24760 50516 24800
rect 50476 24424 50516 24464
rect 50764 25096 50804 25136
rect 50668 24088 50708 24128
rect 50572 24004 50612 24044
rect 49420 23500 49460 23540
rect 49900 23332 49940 23372
rect 49324 22408 49364 22448
rect 50476 23752 50516 23792
rect 50380 23500 50420 23540
rect 49804 22576 49844 22616
rect 49612 22240 49652 22280
rect 49708 22072 49748 22112
rect 49132 20140 49172 20180
rect 49516 21316 49556 21356
rect 50092 22408 50132 22448
rect 51148 25096 51188 25136
rect 50956 24508 50996 24548
rect 50956 24088 50996 24128
rect 50860 23332 50900 23372
rect 50668 22996 50708 23036
rect 52204 28960 52244 29000
rect 52012 27784 52052 27824
rect 53068 29884 53108 29924
rect 53548 32824 53588 32864
rect 53452 32740 53492 32780
rect 53644 32656 53684 32696
rect 53452 32488 53492 32528
rect 53356 32404 53396 32444
rect 53356 32152 53396 32192
rect 53644 31480 53684 31520
rect 54604 33328 54644 33368
rect 54412 33076 54452 33116
rect 54412 32824 54452 32864
rect 54796 33412 54836 33452
rect 54700 33160 54740 33200
rect 54700 32824 54740 32864
rect 54028 32572 54068 32612
rect 54604 32404 54644 32444
rect 54508 31732 54548 31772
rect 54796 31816 54836 31856
rect 53932 31396 53972 31436
rect 53836 31228 53876 31268
rect 53836 30556 53876 30596
rect 54124 31312 54164 31352
rect 54028 30304 54068 30344
rect 53356 30220 53396 30260
rect 53932 30220 53972 30260
rect 53164 29800 53204 29840
rect 54220 30136 54260 30176
rect 54316 29800 54356 29840
rect 53260 29044 53300 29084
rect 54316 28876 54356 28916
rect 52780 28456 52820 28496
rect 52492 28372 52532 28412
rect 52396 28288 52436 28328
rect 53068 28456 53108 28496
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 52012 27616 52052 27656
rect 52108 27448 52148 27488
rect 52780 27784 52820 27824
rect 52684 27616 52724 27656
rect 51916 27364 51956 27404
rect 52588 27448 52628 27488
rect 52300 27196 52340 27236
rect 52108 27112 52148 27152
rect 52780 27280 52820 27320
rect 52780 27112 52820 27152
rect 53260 27868 53300 27908
rect 52876 27028 52916 27068
rect 52780 26944 52820 26984
rect 52684 26776 52724 26816
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 52300 25684 52340 25724
rect 52300 25516 52340 25556
rect 51532 25096 51572 25136
rect 51244 24508 51284 24548
rect 51148 24424 51188 24464
rect 51148 24172 51188 24212
rect 50956 22828 50996 22868
rect 50476 22240 50516 22280
rect 50284 21568 50324 21608
rect 50956 22072 50996 22112
rect 50764 21904 50804 21944
rect 50668 21652 50708 21692
rect 50572 21568 50612 21608
rect 50188 21484 50228 21524
rect 51244 24088 51284 24128
rect 51340 24004 51380 24044
rect 51244 23920 51284 23960
rect 51628 24004 51668 24044
rect 51916 25264 51956 25304
rect 51820 24760 51860 24800
rect 52108 25180 52148 25220
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 52300 24760 52340 24800
rect 52108 24508 52148 24548
rect 52300 24508 52340 24548
rect 52012 24172 52052 24212
rect 52204 24424 52244 24464
rect 51916 23500 51956 23540
rect 51724 23164 51764 23204
rect 51532 23080 51572 23120
rect 51244 22996 51284 23036
rect 51340 22828 51380 22868
rect 51532 22828 51572 22868
rect 51244 21568 51284 21608
rect 51148 21484 51188 21524
rect 49612 20140 49652 20180
rect 49420 20056 49460 20096
rect 49612 19300 49652 19340
rect 48940 17788 48980 17828
rect 48940 17536 48980 17576
rect 48748 14680 48788 14720
rect 48652 14260 48692 14300
rect 48364 14092 48404 14132
rect 47788 13252 47828 13292
rect 47692 13168 47732 13208
rect 48460 14008 48500 14048
rect 48076 12832 48116 12872
rect 48076 12664 48116 12704
rect 47212 12496 47252 12536
rect 48268 12748 48308 12788
rect 48172 12580 48212 12620
rect 48652 12496 48692 12536
rect 46924 11824 46964 11864
rect 46252 11572 46292 11612
rect 47116 11236 47156 11276
rect 46252 11068 46292 11108
rect 46348 10984 46388 11024
rect 45772 10312 45812 10352
rect 45388 10228 45428 10268
rect 45004 10144 45044 10184
rect 44908 9892 44948 9932
rect 44428 8800 44468 8840
rect 45964 10228 46004 10268
rect 45772 9808 45812 9848
rect 45484 9388 45524 9428
rect 45292 9304 45332 9344
rect 44908 8800 44948 8840
rect 45100 8716 45140 8756
rect 45292 8632 45332 8672
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 45772 9388 45812 9428
rect 45676 8548 45716 8588
rect 45580 8464 45620 8504
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 45676 7372 45716 7412
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 48940 16024 48980 16064
rect 49420 19048 49460 19088
rect 49612 18712 49652 18752
rect 49132 18544 49172 18584
rect 49420 18460 49460 18500
rect 49324 18376 49364 18416
rect 49132 18292 49172 18332
rect 49708 18292 49748 18332
rect 49324 18124 49364 18164
rect 49132 17788 49172 17828
rect 49900 20140 49940 20180
rect 49996 19636 50036 19676
rect 50092 18810 50132 18836
rect 50092 18796 50132 18810
rect 49900 18544 49940 18584
rect 50572 20812 50612 20852
rect 50380 19888 50420 19928
rect 50764 19636 50804 19676
rect 50668 19216 50708 19256
rect 50380 18880 50420 18920
rect 50380 18712 50420 18752
rect 50572 18376 50612 18416
rect 50476 18292 50516 18332
rect 49900 18124 49940 18164
rect 50188 18124 50228 18164
rect 49420 17872 49460 17912
rect 49708 17872 49748 17912
rect 49324 15688 49364 15728
rect 49036 15604 49076 15644
rect 49132 15520 49172 15560
rect 49132 14176 49172 14216
rect 48940 13924 48980 13964
rect 49036 13756 49076 13796
rect 49612 17704 49652 17744
rect 49516 17536 49556 17576
rect 49804 17368 49844 17408
rect 49708 16864 49748 16904
rect 49996 17788 50036 17828
rect 50188 17704 50228 17744
rect 52012 23332 52052 23372
rect 52108 23080 52148 23120
rect 52492 23836 52532 23876
rect 52492 23332 52532 23372
rect 52396 23164 52436 23204
rect 52588 22996 52628 23036
rect 52588 22828 52628 22868
rect 52684 22744 52724 22784
rect 52396 22492 52436 22532
rect 51916 21736 51956 21776
rect 52396 21652 52436 21692
rect 51628 21316 51668 21356
rect 52204 21568 52244 21608
rect 51916 21316 51956 21356
rect 51820 21232 51860 21272
rect 51532 20896 51572 20936
rect 52492 21568 52532 21608
rect 52588 21400 52628 21440
rect 52492 21064 52532 21104
rect 52300 20980 52340 21020
rect 52492 20896 52532 20936
rect 52204 20728 52244 20768
rect 52588 20728 52628 20768
rect 52108 20476 52148 20516
rect 52300 20560 52340 20600
rect 51436 20140 51476 20180
rect 52204 20140 52244 20180
rect 51148 19888 51188 19928
rect 51916 19972 51956 20012
rect 51532 19636 51572 19676
rect 51340 18796 51380 18836
rect 50956 18712 50996 18752
rect 51148 18628 51188 18668
rect 50956 18544 50996 18584
rect 50860 18460 50900 18500
rect 50764 17872 50804 17912
rect 50092 17368 50132 17408
rect 50092 16948 50132 16988
rect 49612 16192 49652 16232
rect 49996 16192 50036 16232
rect 50572 17536 50612 17576
rect 50284 16780 50324 16820
rect 50764 17704 50804 17744
rect 51052 18376 51092 18416
rect 51244 18124 51284 18164
rect 51436 18460 51476 18500
rect 51052 17788 51092 17828
rect 50380 16696 50420 16736
rect 50380 16528 50420 16568
rect 49804 15604 49844 15644
rect 49420 14932 49460 14972
rect 49324 14680 49364 14720
rect 49516 14260 49556 14300
rect 49324 14092 49364 14132
rect 49516 14092 49556 14132
rect 49420 13504 49460 13544
rect 49132 13168 49172 13208
rect 48940 12244 48980 12284
rect 48844 10900 48884 10940
rect 48268 10816 48308 10856
rect 49900 15436 49940 15476
rect 49996 14680 50036 14720
rect 49708 14260 49748 14300
rect 50092 14260 50132 14300
rect 49804 14008 49844 14048
rect 49804 13336 49844 13376
rect 49804 12748 49844 12788
rect 49516 12664 49556 12704
rect 50188 13840 50228 13880
rect 49900 12664 49940 12704
rect 49708 12580 49748 12620
rect 49996 12496 50036 12536
rect 49900 12412 49940 12452
rect 49324 11068 49364 11108
rect 47788 10396 47828 10436
rect 48940 10396 48980 10436
rect 47116 10144 47156 10184
rect 46444 10060 46484 10100
rect 46636 10060 46676 10100
rect 47020 10060 47060 10100
rect 46252 9976 46292 10016
rect 46060 9808 46100 9848
rect 45964 8716 46004 8756
rect 46252 9556 46292 9596
rect 46156 9472 46196 9512
rect 46060 8632 46100 8672
rect 46636 9892 46676 9932
rect 46540 9472 46580 9512
rect 46828 9556 46868 9596
rect 47020 9556 47060 9596
rect 46732 9472 46772 9512
rect 48364 9892 48404 9932
rect 48268 9724 48308 9764
rect 47212 9472 47252 9512
rect 47788 9472 47828 9512
rect 47596 8800 47636 8840
rect 46444 8632 46484 8672
rect 46348 8548 46388 8588
rect 47788 8716 47828 8756
rect 48460 9808 48500 9848
rect 48364 8968 48404 9008
rect 46924 7708 46964 7748
rect 47596 7708 47636 7748
rect 46828 7372 46868 7412
rect 47884 7624 47924 7664
rect 48076 7540 48116 7580
rect 48364 8548 48404 8588
rect 48268 7960 48308 8000
rect 47884 7120 47924 7160
rect 48748 9556 48788 9596
rect 50668 16780 50708 16820
rect 50572 16696 50612 16736
rect 50764 16696 50804 16736
rect 50860 16612 50900 16652
rect 50668 16528 50708 16568
rect 50572 16024 50612 16064
rect 50476 15604 50516 15644
rect 50380 13756 50420 13796
rect 50284 13336 50324 13376
rect 50380 13168 50420 13208
rect 50284 13000 50324 13040
rect 50188 11236 50228 11276
rect 51340 16696 51380 16736
rect 51244 16612 51284 16652
rect 51052 16108 51092 16148
rect 50956 16024 50996 16064
rect 50860 15604 50900 15644
rect 51148 16024 51188 16064
rect 51628 19216 51668 19256
rect 52012 18964 52052 19004
rect 51820 18628 51860 18668
rect 51724 18460 51764 18500
rect 51820 18376 51860 18416
rect 51628 16780 51668 16820
rect 51628 16192 51668 16232
rect 51436 15856 51476 15896
rect 51052 15436 51092 15476
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 51532 14848 51572 14888
rect 51340 14680 51380 14720
rect 50860 14428 50900 14468
rect 51916 18292 51956 18332
rect 52684 18628 52724 18668
rect 53452 28288 53492 28328
rect 53548 27280 53588 27320
rect 53548 26944 53588 26984
rect 53356 26608 53396 26648
rect 53548 26608 53588 26648
rect 53932 26776 53972 26816
rect 53356 26440 53396 26480
rect 53644 26440 53684 26480
rect 53260 26356 53300 26396
rect 53164 26104 53204 26144
rect 53836 26356 53876 26396
rect 54028 26608 54068 26648
rect 54124 26440 54164 26480
rect 53068 25852 53108 25892
rect 53068 25180 53108 25220
rect 53932 25936 53972 25976
rect 54124 26104 54164 26144
rect 54412 28288 54452 28328
rect 54412 27364 54452 27404
rect 54028 25852 54068 25892
rect 54220 25432 54260 25472
rect 53740 25264 53780 25304
rect 54988 32824 55028 32864
rect 55468 33836 55508 33872
rect 55468 33832 55508 33836
rect 55276 33412 55316 33452
rect 55468 33580 55508 33620
rect 55372 33244 55412 33284
rect 55372 32992 55412 33032
rect 55180 32824 55220 32864
rect 55756 33664 55796 33704
rect 55660 33328 55700 33368
rect 55084 32656 55124 32696
rect 54604 30136 54644 30176
rect 54892 30640 54932 30680
rect 54700 30052 54740 30092
rect 55276 31312 55316 31352
rect 55372 30808 55412 30848
rect 55852 32992 55892 33032
rect 56044 32824 56084 32864
rect 55852 32740 55892 32780
rect 56140 31732 56180 31772
rect 56428 33664 56468 33704
rect 56428 32740 56468 32780
rect 56044 30808 56084 30848
rect 55660 30640 55700 30680
rect 54892 29800 54932 29840
rect 54892 29464 54932 29504
rect 55276 29464 55316 29504
rect 54796 28708 54836 28748
rect 55180 29044 55220 29084
rect 55084 28708 55124 28748
rect 54892 28288 54932 28328
rect 55276 28288 55316 28328
rect 55180 27952 55220 27992
rect 54988 27196 55028 27236
rect 54604 26776 54644 26816
rect 54796 26356 54836 26396
rect 55084 26608 55124 26648
rect 54796 26188 54836 26228
rect 54988 26188 55028 26228
rect 55468 30052 55508 30092
rect 57388 35596 57428 35636
rect 57676 35848 57716 35888
rect 57292 34588 57332 34628
rect 57196 34504 57236 34544
rect 56812 34252 56852 34292
rect 56236 30556 56276 30596
rect 56140 30052 56180 30092
rect 56908 33664 56948 33704
rect 57292 34168 57332 34208
rect 57196 34000 57236 34040
rect 57484 34000 57524 34040
rect 57772 35764 57812 35804
rect 59404 37360 59444 37400
rect 58828 37108 58868 37148
rect 58636 36688 58676 36728
rect 59500 37276 59540 37316
rect 59692 37192 59732 37232
rect 59692 36856 59732 36896
rect 60076 37108 60116 37148
rect 59884 36604 59924 36644
rect 59020 36016 59060 36056
rect 58444 35848 58484 35888
rect 57868 35680 57908 35720
rect 58252 35680 58292 35720
rect 58060 34336 58100 34376
rect 58732 35344 58772 35384
rect 59596 36436 59636 36476
rect 59404 36016 59444 36056
rect 59404 35348 59444 35384
rect 59404 35344 59444 35348
rect 60364 36688 60404 36728
rect 60268 35764 60308 35804
rect 60172 35344 60212 35384
rect 60268 35260 60308 35300
rect 58636 34336 58676 34376
rect 59116 34420 59156 34460
rect 59308 34420 59348 34460
rect 59884 35176 59924 35216
rect 60940 37360 60980 37400
rect 61228 36856 61268 36896
rect 60652 36604 60692 36644
rect 60940 36604 60980 36644
rect 60940 36436 60980 36476
rect 60844 35848 60884 35888
rect 59692 34168 59732 34208
rect 59980 34168 60020 34208
rect 59404 33916 59444 33956
rect 59596 33748 59636 33788
rect 58348 33580 58388 33620
rect 59020 33580 59060 33620
rect 59500 33664 59540 33704
rect 59404 33496 59444 33536
rect 57868 32824 57908 32864
rect 57676 32740 57716 32780
rect 57100 32488 57140 32528
rect 57100 31732 57140 31772
rect 56812 31312 56852 31352
rect 57292 32068 57332 32108
rect 57676 32152 57716 32192
rect 57484 32068 57524 32108
rect 57868 31984 57908 32024
rect 57772 31900 57812 31940
rect 57484 31312 57524 31352
rect 57676 31312 57716 31352
rect 56524 30304 56564 30344
rect 56140 29548 56180 29588
rect 55660 29296 55700 29336
rect 56140 29296 56180 29336
rect 56044 28708 56084 28748
rect 57484 31144 57524 31184
rect 58828 32824 58868 32864
rect 58156 32488 58196 32528
rect 58060 31312 58100 31352
rect 58540 32152 58580 32192
rect 58444 31648 58484 31688
rect 58348 31396 58388 31436
rect 58252 31312 58292 31352
rect 57004 30304 57044 30344
rect 57772 30640 57812 30680
rect 57580 30052 57620 30092
rect 56812 29464 56852 29504
rect 57388 29464 57428 29504
rect 56812 29296 56852 29336
rect 55756 28036 55796 28076
rect 55564 27196 55604 27236
rect 55564 26440 55604 26480
rect 55372 26356 55412 26396
rect 55084 26104 55124 26144
rect 54796 25936 54836 25976
rect 54508 25600 54548 25640
rect 54604 25432 54644 25472
rect 54316 25264 54356 25304
rect 53836 24508 53876 24548
rect 53068 24004 53108 24044
rect 53164 23752 53204 23792
rect 54508 25264 54548 25304
rect 54796 25264 54836 25304
rect 55084 24760 55124 24800
rect 55084 24592 55124 24632
rect 55276 24592 55316 24632
rect 54796 24424 54836 24464
rect 54316 24088 54356 24128
rect 54220 24004 54260 24044
rect 55084 24088 55124 24128
rect 54988 24004 55028 24044
rect 54028 23752 54068 23792
rect 54220 23752 54260 23792
rect 54796 23752 54836 23792
rect 55948 27532 55988 27572
rect 55852 26104 55892 26144
rect 57484 29300 57524 29336
rect 57484 29296 57524 29300
rect 56236 27364 56276 27404
rect 57964 29548 58004 29588
rect 57868 28288 57908 28328
rect 57676 27700 57716 27740
rect 56044 26776 56084 26816
rect 57004 26776 57044 26816
rect 56524 26356 56564 26396
rect 55948 25936 55988 25976
rect 55660 23920 55700 23960
rect 55564 23668 55604 23708
rect 54124 23500 54164 23540
rect 54028 23332 54068 23372
rect 56236 26020 56276 26060
rect 56140 25936 56180 25976
rect 57004 26020 57044 26060
rect 56524 25936 56564 25976
rect 56428 25516 56468 25556
rect 56620 25600 56660 25640
rect 56716 25432 56756 25472
rect 56716 24928 56756 24968
rect 56428 24172 56468 24212
rect 56524 24088 56564 24128
rect 55660 23080 55700 23120
rect 53068 22996 53108 23036
rect 53260 22912 53300 22952
rect 53545 22744 53585 22784
rect 53945 22996 53985 23036
rect 55255 22996 55295 23036
rect 55948 22996 55988 23036
rect 54455 22912 54495 22952
rect 54745 22912 54785 22952
rect 55145 22912 55185 22952
rect 54345 22828 54385 22868
rect 54855 22744 54895 22784
rect 56140 23668 56180 23708
rect 57676 26188 57716 26228
rect 57676 25936 57716 25976
rect 57388 25852 57428 25892
rect 57292 25600 57332 25640
rect 56908 24928 56948 24968
rect 57484 25516 57524 25556
rect 58636 32068 58676 32108
rect 58924 31900 58964 31940
rect 59308 32068 59348 32108
rect 59212 31312 59252 31352
rect 59116 31144 59156 31184
rect 59116 30640 59156 30680
rect 58252 30304 58292 30344
rect 59212 30304 59252 30344
rect 59404 30052 59444 30092
rect 59596 30052 59636 30092
rect 58156 29296 58196 29336
rect 58924 29464 58964 29504
rect 58252 29128 58292 29168
rect 58828 29128 58868 29168
rect 59884 34084 59924 34124
rect 59884 33664 59924 33704
rect 60172 32656 60212 32696
rect 60172 32152 60212 32192
rect 59788 31732 59828 31772
rect 59980 31732 60020 31772
rect 60460 34000 60500 34040
rect 60652 33916 60692 33956
rect 60460 32320 60500 32360
rect 60364 31900 60404 31940
rect 60460 31816 60500 31856
rect 60556 31648 60596 31688
rect 60556 30640 60596 30680
rect 60268 30304 60308 30344
rect 60172 29968 60212 30008
rect 59692 29464 59732 29504
rect 59788 29380 59828 29420
rect 60076 29380 60116 29420
rect 58924 28456 58964 28496
rect 58060 27700 58100 27740
rect 58156 27364 58196 27404
rect 57964 25936 58004 25976
rect 57868 25852 57908 25892
rect 57772 25600 57812 25640
rect 57772 25432 57812 25472
rect 56812 23920 56852 23960
rect 56908 23752 56948 23792
rect 56524 23668 56564 23708
rect 57292 23752 57332 23792
rect 57484 24676 57524 24716
rect 57196 23500 57236 23540
rect 56332 23332 56372 23372
rect 57100 23248 57140 23288
rect 58060 24844 58100 24884
rect 57868 24592 57908 24632
rect 57868 24172 57908 24212
rect 57772 23920 57812 23960
rect 57868 23752 57908 23792
rect 58828 27868 58868 27908
rect 58540 27616 58580 27656
rect 58444 26860 58484 26900
rect 58732 27280 58772 27320
rect 58636 26440 58676 26480
rect 58348 26104 58388 26144
rect 58252 24424 58292 24464
rect 58252 23836 58292 23876
rect 58252 23248 58292 23288
rect 55756 22912 55796 22952
rect 55655 22828 55695 22868
rect 55545 22744 55585 22784
rect 55756 22744 55796 22784
rect 56140 22744 56180 22784
rect 56455 22996 56495 23036
rect 56745 22912 56785 22952
rect 56855 22744 56895 22784
rect 58444 25432 58484 25472
rect 58540 25096 58580 25136
rect 58828 26104 58868 26144
rect 59692 29128 59732 29168
rect 59116 28708 59156 28748
rect 59404 28708 59444 28748
rect 59020 28288 59060 28328
rect 59020 27700 59060 27740
rect 59308 27952 59348 27992
rect 59116 27028 59156 27068
rect 59020 26860 59060 26900
rect 59212 26524 59252 26564
rect 61036 35932 61076 35972
rect 61228 36688 61268 36728
rect 61132 35848 61172 35888
rect 61324 36436 61364 36476
rect 63820 38116 63860 38156
rect 64684 38116 64724 38156
rect 62284 38032 62324 38072
rect 61708 36268 61748 36308
rect 61420 36016 61460 36056
rect 61804 35932 61844 35972
rect 61324 35848 61364 35888
rect 61036 35680 61076 35720
rect 61228 35512 61268 35552
rect 60940 35092 60980 35132
rect 61036 35008 61076 35048
rect 61516 35764 61556 35804
rect 61420 35428 61460 35468
rect 61420 35092 61460 35132
rect 61420 34924 61460 34964
rect 61420 34672 61460 34712
rect 61324 34168 61364 34208
rect 61132 33832 61172 33872
rect 61324 33748 61364 33788
rect 60844 33496 60884 33536
rect 61612 35428 61652 35468
rect 61612 35092 61652 35132
rect 62188 37360 62228 37400
rect 62188 36184 62228 36224
rect 61900 35176 61940 35216
rect 61804 34672 61844 34712
rect 61804 34504 61844 34544
rect 61516 33748 61556 33788
rect 62092 34168 62132 34208
rect 61996 33832 62036 33872
rect 61612 33496 61652 33536
rect 61324 33160 61364 33200
rect 60940 32152 60980 32192
rect 60748 31816 60788 31856
rect 61132 32068 61172 32108
rect 61036 31984 61076 32024
rect 61036 31816 61076 31856
rect 61132 31480 61172 31520
rect 61516 32152 61556 32192
rect 61516 31984 61556 32024
rect 61324 31648 61364 31688
rect 61516 31480 61556 31520
rect 61228 31396 61268 31436
rect 61420 31396 61460 31436
rect 60940 30388 60980 30428
rect 60748 29884 60788 29924
rect 60748 29632 60788 29672
rect 60460 28876 60500 28916
rect 60076 28792 60116 28832
rect 60076 28372 60116 28412
rect 59788 28288 59828 28328
rect 60172 28288 60212 28328
rect 59980 28120 60020 28160
rect 59020 26272 59060 26312
rect 58732 25348 58772 25388
rect 58924 25348 58964 25388
rect 59116 26188 59156 26228
rect 59500 26188 59540 26228
rect 59692 26188 59732 26228
rect 59308 25768 59348 25808
rect 59212 25684 59252 25724
rect 59596 25936 59636 25976
rect 60076 26692 60116 26732
rect 59980 26188 60020 26228
rect 60268 26776 60308 26816
rect 60172 26524 60212 26564
rect 60556 28288 60596 28328
rect 60652 28204 60692 28244
rect 60940 28456 60980 28496
rect 61132 30556 61172 30596
rect 61708 33412 61748 33452
rect 61996 33412 62036 33452
rect 61804 33328 61844 33368
rect 61804 32656 61844 32696
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 62764 37360 62804 37400
rect 62476 35092 62516 35132
rect 62380 34924 62420 34964
rect 62284 34504 62324 34544
rect 62572 34420 62612 34460
rect 62668 34336 62708 34376
rect 62860 35932 62900 35972
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 63724 36184 63764 36224
rect 64396 37444 64436 37484
rect 64492 37360 64532 37400
rect 64780 37192 64820 37232
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 64300 36688 64340 36728
rect 64780 36688 64820 36728
rect 64684 36100 64724 36140
rect 64300 36016 64340 36056
rect 63820 35848 63860 35888
rect 64012 35848 64052 35888
rect 62956 35428 62996 35468
rect 62860 35176 62900 35216
rect 63532 34924 63572 34964
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 63628 34420 63668 34460
rect 62092 31564 62132 31604
rect 61708 31480 61748 31520
rect 61612 31312 61652 31352
rect 61804 31396 61844 31436
rect 61612 30556 61652 30596
rect 61420 30388 61460 30428
rect 61228 30220 61268 30260
rect 61132 29548 61172 29588
rect 60844 28288 60884 28328
rect 61036 28288 61076 28328
rect 60844 27784 60884 27824
rect 60556 26944 60596 26984
rect 60460 26524 60500 26564
rect 60268 26104 60308 26144
rect 61036 27616 61076 27656
rect 60844 27448 60884 27488
rect 60748 27112 60788 27152
rect 60748 26944 60788 26984
rect 60652 26272 60692 26312
rect 59980 25936 60020 25976
rect 59884 25852 59924 25892
rect 59596 25768 59636 25808
rect 59020 24172 59060 24212
rect 59212 25264 59252 25304
rect 59116 23752 59156 23792
rect 59020 23080 59060 23120
rect 59500 25264 59540 25304
rect 59596 25132 59636 25136
rect 59596 25096 59636 25132
rect 59404 24844 59444 24884
rect 59788 24844 59828 24884
rect 59692 24340 59732 24380
rect 59596 23836 59636 23876
rect 59404 23752 59444 23792
rect 59596 23584 59636 23624
rect 59500 23416 59540 23456
rect 60556 25852 60596 25892
rect 60268 25684 60308 25724
rect 59980 25516 60020 25556
rect 60172 25348 60212 25388
rect 60076 25264 60116 25304
rect 59884 24760 59924 24800
rect 59884 24592 59924 24632
rect 59884 23836 59924 23876
rect 59980 23752 60020 23792
rect 60172 24928 60212 24968
rect 59979 23080 60019 23120
rect 57545 22828 57585 22868
rect 57945 22828 57985 22868
rect 57655 22744 57695 22784
rect 58345 22912 58385 22952
rect 59145 22744 59185 22784
rect 59945 22912 59985 22952
rect 60364 25516 60404 25556
rect 60844 26860 60884 26900
rect 60748 25768 60788 25808
rect 60748 25516 60788 25556
rect 60556 25264 60596 25304
rect 60844 25264 60884 25304
rect 60268 24844 60308 24884
rect 60748 24760 60788 24800
rect 60556 24676 60596 24716
rect 60364 23752 60404 23792
rect 60268 23584 60308 23624
rect 60364 23416 60404 23456
rect 60268 22912 60308 22952
rect 61708 29632 61748 29672
rect 61516 29548 61556 29588
rect 62764 32740 62804 32780
rect 62860 32656 62900 32696
rect 63532 34336 63572 34376
rect 63244 33832 63284 33872
rect 63628 33916 63668 33956
rect 63724 33832 63764 33872
rect 63244 33412 63284 33452
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 64012 34924 64052 34964
rect 64012 34504 64052 34544
rect 64588 35848 64628 35888
rect 64876 36184 64916 36224
rect 65452 38032 65492 38072
rect 68332 38200 68372 38240
rect 67756 38116 67796 38156
rect 66508 38032 66548 38072
rect 66892 38032 66932 38072
rect 65836 37948 65876 37988
rect 65260 37444 65300 37484
rect 65164 37360 65204 37400
rect 65548 37360 65588 37400
rect 65932 37360 65972 37400
rect 65452 37192 65492 37232
rect 65164 36184 65204 36224
rect 65068 36100 65108 36140
rect 64876 35848 64916 35888
rect 64972 35680 65012 35720
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 64204 34420 64244 34460
rect 64780 34420 64820 34460
rect 64684 34336 64724 34376
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 64492 33832 64532 33872
rect 64300 33748 64340 33788
rect 63916 33496 63956 33536
rect 63148 33076 63188 33116
rect 63052 32692 63092 32696
rect 63052 32656 63092 32692
rect 62764 32152 62804 32192
rect 63340 32152 63380 32192
rect 63052 32068 63092 32108
rect 63532 32068 63572 32108
rect 63436 31900 63476 31940
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 63244 31396 63284 31436
rect 62572 30640 62612 30680
rect 63532 31312 63572 31352
rect 63436 30472 63476 30512
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 62476 30052 62516 30092
rect 63532 30052 63572 30092
rect 61900 29968 61940 30008
rect 61804 29296 61844 29336
rect 61324 28624 61364 28664
rect 61324 28372 61364 28412
rect 62284 29128 62324 29168
rect 62476 29044 62516 29084
rect 61804 28624 61844 28664
rect 61612 28372 61652 28412
rect 62092 28876 62132 28916
rect 62092 28624 62132 28664
rect 61996 28288 62036 28328
rect 62284 28456 62324 28496
rect 62188 28372 62228 28412
rect 61900 28204 61940 28244
rect 61708 28120 61748 28160
rect 61228 27784 61268 27824
rect 62860 28372 62900 28412
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 63052 28540 63092 28580
rect 62956 28288 62996 28328
rect 62764 28120 62804 28160
rect 61516 27784 61556 27824
rect 61900 27784 61940 27824
rect 61324 27448 61364 27488
rect 61228 27112 61268 27152
rect 61900 27616 61940 27656
rect 62572 27196 62612 27236
rect 62380 26944 62420 26984
rect 61612 26860 61652 26900
rect 62092 26860 62132 26900
rect 61804 26776 61844 26816
rect 61420 26692 61460 26732
rect 61420 26370 61460 26396
rect 61420 26356 61460 26370
rect 61900 26356 61940 26396
rect 61324 26104 61364 26144
rect 61324 25264 61364 25304
rect 61324 24676 61364 24716
rect 61324 24508 61364 24548
rect 61228 24424 61268 24464
rect 61132 24340 61172 24380
rect 61228 23836 61268 23876
rect 61132 23752 61172 23792
rect 61132 23164 61172 23204
rect 61996 25852 62036 25892
rect 62284 26608 62324 26648
rect 62092 25600 62132 25640
rect 61996 25096 62036 25136
rect 62188 24760 62228 24800
rect 61804 24424 61844 24464
rect 61804 24088 61844 24128
rect 61804 23584 61844 23624
rect 62188 24340 62228 24380
rect 62092 24088 62132 24128
rect 61996 23836 62036 23876
rect 62476 24256 62516 24296
rect 62764 26020 62804 26060
rect 62764 25768 62804 25808
rect 62668 25180 62708 25220
rect 64012 33328 64052 33368
rect 63724 32152 63764 32192
rect 63724 31900 63764 31940
rect 64684 33664 64724 33704
rect 65260 36016 65300 36056
rect 66220 36016 66260 36056
rect 65644 35932 65684 35972
rect 65164 34336 65204 34376
rect 65452 35848 65492 35888
rect 65548 35596 65588 35636
rect 65836 35848 65876 35888
rect 65740 35680 65780 35720
rect 65740 35008 65780 35048
rect 65356 34252 65396 34292
rect 65068 33748 65108 33788
rect 64300 33580 64340 33620
rect 64588 33580 64628 33620
rect 64780 33496 64820 33536
rect 64588 33328 64628 33368
rect 64876 33160 64916 33200
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 64012 31816 64052 31856
rect 63916 31312 63956 31352
rect 63724 30388 63764 30428
rect 64012 30220 64052 30260
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 63244 25936 63284 25976
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 63052 25432 63092 25472
rect 62860 24760 62900 24800
rect 62668 24256 62708 24296
rect 61900 23416 61940 23456
rect 61612 23332 61652 23372
rect 60855 22996 60895 23036
rect 60748 22828 60788 22868
rect 62380 23584 62420 23624
rect 61545 22744 61585 22784
rect 62668 23836 62708 23876
rect 62572 23752 62612 23792
rect 62668 23248 62708 23288
rect 62860 24340 62900 24380
rect 62860 24088 62900 24128
rect 62860 23836 62900 23876
rect 62860 23584 62900 23624
rect 63052 24256 63092 24296
rect 62956 23332 62996 23372
rect 61945 22744 61985 22784
rect 63148 24004 63188 24044
rect 63244 23668 63284 23708
rect 63340 23500 63380 23540
rect 63628 27616 63668 27656
rect 64204 32152 64244 32192
rect 64588 32152 64628 32192
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 65356 33580 65396 33620
rect 64876 30136 64916 30176
rect 64396 30052 64436 30092
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 64492 29296 64532 29336
rect 66412 35764 66452 35804
rect 65836 32908 65876 32948
rect 66220 32908 66260 32948
rect 65644 32824 65684 32864
rect 67468 37948 67508 37988
rect 67372 37444 67412 37484
rect 66700 37360 66740 37400
rect 67084 36772 67124 36812
rect 66796 36016 66836 36056
rect 66604 35848 66644 35888
rect 66508 32404 66548 32444
rect 66988 34420 67028 34460
rect 66796 34252 66836 34292
rect 66700 33664 66740 33704
rect 67180 36520 67220 36560
rect 67372 36856 67412 36896
rect 67564 37276 67604 37316
rect 67276 35764 67316 35804
rect 67180 34504 67220 34544
rect 68428 37444 68468 37484
rect 67756 37192 67796 37232
rect 68140 36856 68180 36896
rect 67660 36016 67700 36056
rect 67852 36688 67892 36728
rect 68236 36772 68276 36812
rect 68332 36520 68372 36560
rect 67852 35848 67892 35888
rect 67756 35596 67796 35636
rect 67372 34420 67412 34460
rect 67084 33664 67124 33704
rect 67564 34336 67604 34376
rect 67468 34252 67508 34292
rect 67756 34000 67796 34040
rect 67948 34336 67988 34376
rect 68236 35680 68276 35720
rect 68236 35008 68276 35048
rect 67468 33748 67508 33788
rect 67852 33748 67892 33788
rect 66892 33580 66932 33620
rect 66796 33496 66836 33536
rect 66700 32824 66740 32864
rect 66796 32656 66836 32696
rect 65836 32236 65876 32276
rect 66604 32236 66644 32276
rect 65644 32152 65684 32192
rect 66124 32152 66164 32192
rect 66412 32152 66452 32192
rect 65452 31984 65492 32024
rect 65356 31732 65396 31772
rect 65068 29968 65108 30008
rect 65068 29800 65108 29840
rect 64972 29548 65012 29588
rect 64780 29212 64820 29252
rect 64876 29128 64916 29168
rect 64300 28708 64340 28748
rect 64204 28288 64244 28328
rect 64396 28288 64436 28328
rect 64684 28792 64724 28832
rect 66124 31732 66164 31772
rect 65740 31312 65780 31352
rect 66604 31984 66644 32024
rect 66796 31984 66836 32024
rect 66892 31816 66932 31856
rect 65836 31144 65876 31184
rect 65740 30304 65780 30344
rect 65452 30220 65492 30260
rect 65356 29968 65396 30008
rect 65260 29884 65300 29924
rect 65548 29884 65588 29924
rect 65452 29800 65492 29840
rect 65644 29632 65684 29672
rect 65548 29548 65588 29588
rect 65356 29212 65396 29252
rect 65260 29044 65300 29084
rect 65260 28792 65300 28832
rect 65164 28708 65204 28748
rect 65452 29128 65492 29168
rect 65548 29044 65588 29084
rect 66412 30724 66452 30764
rect 66316 30136 66356 30176
rect 65932 29884 65972 29924
rect 66316 29884 66356 29924
rect 66220 29800 66260 29840
rect 66700 30640 66740 30680
rect 66604 29800 66644 29840
rect 66412 29668 66452 29672
rect 66412 29632 66452 29668
rect 65836 29296 65876 29336
rect 65932 28960 65972 29000
rect 65836 28876 65876 28916
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 64204 27616 64244 27656
rect 63916 26944 63956 26984
rect 64108 26944 64148 26984
rect 63724 26776 63764 26816
rect 63628 26020 63668 26060
rect 63916 26692 63956 26732
rect 64108 26272 64148 26312
rect 65260 28204 65300 28244
rect 65068 27616 65108 27656
rect 64396 26860 64436 26900
rect 64876 27364 64916 27404
rect 64972 26776 65012 26816
rect 64588 26608 64628 26648
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 64684 26272 64724 26312
rect 63724 25432 63764 25472
rect 64108 25348 64148 25388
rect 63628 25264 63668 25304
rect 63532 24592 63572 24632
rect 64108 25096 64148 25136
rect 64588 25180 64628 25220
rect 64972 26524 65012 26564
rect 64876 25936 64916 25976
rect 64780 25096 64820 25136
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 64684 24760 64724 24800
rect 64108 24676 64148 24716
rect 64492 24676 64532 24716
rect 63628 24172 63668 24212
rect 63532 23920 63572 23960
rect 63436 23248 63476 23288
rect 64012 24004 64052 24044
rect 64300 24424 64340 24464
rect 64300 23836 64340 23876
rect 64396 23752 64436 23792
rect 64588 24592 64628 24632
rect 63916 23668 63956 23708
rect 64300 23584 64340 23624
rect 64012 23416 64052 23456
rect 64492 23248 64532 23288
rect 63945 22912 63985 22952
rect 64780 23752 64820 23792
rect 64876 23332 64916 23372
rect 65164 26944 65204 26984
rect 65356 28120 65396 28160
rect 65836 28372 65876 28412
rect 67372 33496 67412 33536
rect 67276 32152 67316 32192
rect 67180 31984 67220 32024
rect 67276 31312 67316 31352
rect 67468 33160 67508 33200
rect 67756 33664 67796 33704
rect 68140 34252 68180 34292
rect 68140 34000 68180 34040
rect 67564 32824 67604 32864
rect 68140 32824 68180 32864
rect 67660 32656 67700 32696
rect 68140 32656 68180 32696
rect 67660 32236 67700 32276
rect 67564 31816 67604 31856
rect 67468 31732 67508 31772
rect 67084 31144 67124 31184
rect 67084 30724 67124 30764
rect 66988 30640 67028 30680
rect 66892 29884 66932 29924
rect 66796 29464 66836 29504
rect 67468 31144 67508 31184
rect 67372 30640 67412 30680
rect 67084 30052 67124 30092
rect 67180 29632 67220 29672
rect 67372 29464 67412 29504
rect 66412 28960 66452 29000
rect 66316 28624 66356 28664
rect 66124 28120 66164 28160
rect 65260 26524 65300 26564
rect 65260 26020 65300 26060
rect 65452 25936 65492 25976
rect 65932 27616 65972 27656
rect 65836 27364 65876 27404
rect 65740 27028 65780 27068
rect 65644 26104 65684 26144
rect 65548 25768 65588 25808
rect 65932 26104 65972 26144
rect 66124 26104 66164 26144
rect 65548 25264 65588 25304
rect 65548 24844 65588 24884
rect 65164 24256 65204 24296
rect 65452 23920 65492 23960
rect 65255 22996 65295 23036
rect 65356 22996 65396 23036
rect 65836 25432 65876 25472
rect 66796 29044 66836 29084
rect 66508 28792 66548 28832
rect 67468 28792 67508 28832
rect 67180 28708 67220 28748
rect 66892 28540 66932 28580
rect 66508 27952 66548 27992
rect 66316 27868 66356 27908
rect 66604 27364 66644 27404
rect 66508 26020 66548 26060
rect 65740 25180 65780 25220
rect 66124 25264 66164 25304
rect 65932 24508 65972 24548
rect 66028 23920 66068 23960
rect 65932 23836 65972 23876
rect 65740 23752 65780 23792
rect 66412 24508 66452 24548
rect 66604 25516 66644 25556
rect 66700 25348 66740 25388
rect 66796 25264 66836 25304
rect 66988 28372 67028 28412
rect 67180 25432 67220 25472
rect 67276 25348 67316 25388
rect 67180 25264 67220 25304
rect 66988 24928 67028 24968
rect 66604 24424 66644 24464
rect 67084 24508 67124 24548
rect 66988 24424 67028 24464
rect 65740 23416 65780 23456
rect 66028 23164 66068 23204
rect 67468 25264 67508 25304
rect 67564 25180 67604 25220
rect 67372 25096 67412 25136
rect 68332 34672 68372 34712
rect 67756 31900 67796 31940
rect 67756 27280 67796 27320
rect 67372 24928 67412 24968
rect 67276 24424 67316 24464
rect 67276 24256 67316 24296
rect 67180 24004 67220 24044
rect 67660 24592 67700 24632
rect 67564 24088 67604 24128
rect 67468 23248 67508 23288
rect 65945 22912 65985 22952
rect 66745 22912 66785 22952
rect 66455 22828 66495 22868
rect 66345 22744 66385 22784
rect 66855 22828 66895 22868
rect 68524 35848 68564 35888
rect 68620 35764 68660 35804
rect 69580 38032 69620 38072
rect 69388 37528 69428 37568
rect 68908 37360 68948 37400
rect 69004 37192 69044 37232
rect 69772 37276 69812 37316
rect 69868 36856 69908 36896
rect 68812 36688 68852 36728
rect 68812 35680 68852 35720
rect 68428 34588 68468 34628
rect 68428 33244 68468 33284
rect 67948 31312 67988 31352
rect 68140 31816 68180 31856
rect 68236 31564 68276 31604
rect 68236 31144 68276 31184
rect 68236 30640 68276 30680
rect 68428 31732 68468 31772
rect 69004 36688 69044 36728
rect 69004 36016 69044 36056
rect 68620 34336 68660 34376
rect 68908 34504 68948 34544
rect 68812 34336 68852 34376
rect 68812 34084 68852 34124
rect 68716 33244 68756 33284
rect 69292 36688 69332 36728
rect 69100 35764 69140 35804
rect 69100 34924 69140 34964
rect 69100 34588 69140 34628
rect 69580 35848 69620 35888
rect 70060 37528 70100 37568
rect 69772 35428 69812 35468
rect 69676 34336 69716 34376
rect 69580 33580 69620 33620
rect 68524 31144 68564 31184
rect 67948 28708 67988 28748
rect 68044 26608 68084 26648
rect 68428 28876 68468 28916
rect 68332 27952 68372 27992
rect 68428 27532 68468 27572
rect 68620 31060 68660 31100
rect 68524 27196 68564 27236
rect 68812 28708 68852 28748
rect 69100 31228 69140 31268
rect 69004 31060 69044 31100
rect 69004 30640 69044 30680
rect 69292 30388 69332 30428
rect 69100 29464 69140 29504
rect 69196 29380 69236 29420
rect 69100 29128 69140 29168
rect 68908 28120 68948 28160
rect 69100 28036 69140 28076
rect 69196 27616 69236 27656
rect 69100 27280 69140 27320
rect 69292 26272 69332 26312
rect 69196 26188 69236 26228
rect 69004 26104 69044 26144
rect 69580 28708 69620 28748
rect 69580 27616 69620 27656
rect 69484 26188 69524 26228
rect 68812 25516 68852 25556
rect 69388 26104 69428 26144
rect 69868 34168 69908 34208
rect 69772 32740 69812 32780
rect 69772 31816 69812 31856
rect 69772 27280 69812 27320
rect 69772 26608 69812 26648
rect 69676 26524 69716 26564
rect 69676 26272 69716 26312
rect 69580 26020 69620 26060
rect 69772 26104 69812 26144
rect 70348 37192 70388 37232
rect 70636 37444 70676 37484
rect 70732 37360 70772 37400
rect 70444 37108 70484 37148
rect 70252 36688 70292 36728
rect 70732 36688 70772 36728
rect 71020 37276 71060 37316
rect 71020 36772 71060 36812
rect 71596 37360 71636 37400
rect 72364 37360 72404 37400
rect 71500 36688 71540 36728
rect 73036 37192 73076 37232
rect 72748 36940 72788 36980
rect 70828 36604 70868 36644
rect 71116 36604 71156 36644
rect 71596 36604 71636 36644
rect 70252 36016 70292 36056
rect 71404 36520 71444 36560
rect 71308 35848 71348 35888
rect 72172 36688 72212 36728
rect 72460 36352 72500 36392
rect 72748 36688 72788 36728
rect 71596 35932 71636 35972
rect 72268 35932 72308 35972
rect 70156 34336 70196 34376
rect 70156 32824 70196 32864
rect 71020 35176 71060 35216
rect 70924 34924 70964 34964
rect 72076 35848 72116 35888
rect 71692 35344 71732 35384
rect 71500 35008 71540 35048
rect 71308 34504 71348 34544
rect 71404 34336 71444 34376
rect 71308 33832 71348 33872
rect 72076 35176 72116 35216
rect 71884 35008 71924 35048
rect 72172 35092 72212 35132
rect 71788 34336 71828 34376
rect 72076 34336 72116 34376
rect 71884 34252 71924 34292
rect 72172 34084 72212 34124
rect 72076 33832 72116 33872
rect 70828 32824 70868 32864
rect 71020 32824 71060 32864
rect 71500 32152 71540 32192
rect 71980 33664 72020 33704
rect 71884 33244 71924 33284
rect 72652 36016 72692 36056
rect 72460 34840 72500 34880
rect 72364 34252 72404 34292
rect 71692 32740 71732 32780
rect 71884 32572 71924 32612
rect 73036 36688 73076 36728
rect 73420 37360 73460 37400
rect 73516 37108 73556 37148
rect 73804 37276 73844 37316
rect 73708 36856 73748 36896
rect 73228 36688 73268 36728
rect 73132 36604 73172 36644
rect 73612 36604 73652 36644
rect 72940 36520 72980 36560
rect 73516 36520 73556 36560
rect 72940 36352 72980 36392
rect 72844 35932 72884 35972
rect 72844 35260 72884 35300
rect 74092 37276 74132 37316
rect 73996 37108 74036 37148
rect 74284 37276 74324 37316
rect 74188 36856 74228 36896
rect 75916 38368 75956 38408
rect 74476 37360 74516 37400
rect 74668 37444 74708 37484
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 75052 37612 75092 37652
rect 75628 37612 75668 37652
rect 76204 37612 76244 37652
rect 75340 37444 75380 37484
rect 74764 37192 74804 37232
rect 73516 35764 73556 35804
rect 73324 35260 73364 35300
rect 72748 34504 72788 34544
rect 72652 34336 72692 34376
rect 72460 33832 72500 33872
rect 72556 33664 72596 33704
rect 73132 35176 73172 35216
rect 72652 33412 72692 33452
rect 73036 33412 73076 33452
rect 73804 36016 73844 36056
rect 73900 35932 73940 35972
rect 74188 36604 74228 36644
rect 74284 36436 74324 36476
rect 74380 36016 74420 36056
rect 74572 36856 74612 36896
rect 74764 36520 74804 36560
rect 74860 35932 74900 35972
rect 74668 35848 74708 35888
rect 74284 35764 74324 35804
rect 74092 35680 74132 35720
rect 73708 35344 73748 35384
rect 73996 35344 74036 35384
rect 73612 34504 73652 34544
rect 73612 34336 73652 34376
rect 74092 34336 74132 34376
rect 73996 33328 74036 33368
rect 73036 33244 73076 33284
rect 72364 32740 72404 32780
rect 72364 32598 72404 32612
rect 72364 32572 72404 32598
rect 72652 32572 72692 32612
rect 72556 32488 72596 32528
rect 72076 32152 72116 32192
rect 71788 32068 71828 32108
rect 71308 31564 71348 31604
rect 70156 31312 70196 31352
rect 69964 30640 70004 30680
rect 70156 30640 70196 30680
rect 69964 30304 70004 30344
rect 70156 28456 70196 28496
rect 70060 28120 70100 28160
rect 69964 27196 70004 27236
rect 70060 26776 70100 26816
rect 69964 26440 70004 26480
rect 69964 26188 70004 26228
rect 69868 25936 69908 25976
rect 69676 25684 69716 25724
rect 70156 26356 70196 26396
rect 71404 31480 71444 31520
rect 70540 30640 70580 30680
rect 71308 30640 71348 30680
rect 71308 30472 71348 30512
rect 71116 30220 71156 30260
rect 70924 30052 70964 30092
rect 70444 29212 70484 29252
rect 70444 28876 70484 28916
rect 70540 28540 70580 28580
rect 71404 30388 71444 30428
rect 71596 31564 71636 31604
rect 71692 30640 71732 30680
rect 71596 30472 71636 30512
rect 72844 32992 72884 33032
rect 72268 31564 72308 31604
rect 72556 31396 72596 31436
rect 72268 31144 72308 31184
rect 71788 30388 71828 30428
rect 72076 30640 72116 30680
rect 71980 30556 72020 30596
rect 71692 30304 71732 30344
rect 71500 30052 71540 30092
rect 71116 29296 71156 29336
rect 71020 29044 71060 29084
rect 70828 28876 70868 28916
rect 71116 28708 71156 28748
rect 70636 28456 70676 28496
rect 70743 28456 70772 28496
rect 70772 28456 70783 28496
rect 71020 28372 71060 28412
rect 71596 29548 71636 29588
rect 71308 29300 71348 29336
rect 71308 29296 71348 29300
rect 71404 29128 71444 29168
rect 71308 29044 71348 29084
rect 71404 28876 71444 28916
rect 71500 28456 71540 28496
rect 70444 28120 70484 28160
rect 70348 27616 70388 27656
rect 69484 25516 69524 25556
rect 68524 25264 68564 25304
rect 68428 25012 68468 25052
rect 68716 24844 68756 24884
rect 68428 24424 68468 24464
rect 68140 24256 68180 24296
rect 67948 24172 67988 24212
rect 67852 23500 67892 23540
rect 67660 23164 67700 23204
rect 68044 23584 68084 23624
rect 68716 24172 68756 24212
rect 68345 22996 68385 23036
rect 68812 24004 68852 24044
rect 68908 23836 68948 23876
rect 68812 23752 68852 23792
rect 69388 25180 69428 25220
rect 69868 25348 69908 25388
rect 69676 25180 69716 25220
rect 70060 25348 70100 25388
rect 70060 25180 70100 25220
rect 69484 24256 69524 24296
rect 69676 24256 69716 24296
rect 69388 23836 69428 23876
rect 69100 23584 69140 23624
rect 69292 23584 69332 23624
rect 69292 23164 69332 23204
rect 70252 25684 70292 25724
rect 71116 27784 71156 27824
rect 71212 27532 71252 27572
rect 70924 26860 70964 26900
rect 71116 26860 71156 26900
rect 70444 26524 70484 26564
rect 70540 26188 70580 26228
rect 70636 26020 70676 26060
rect 70444 25768 70484 25808
rect 70060 23836 70100 23876
rect 70156 23668 70196 23708
rect 69964 23500 70004 23540
rect 70060 23248 70100 23288
rect 70828 26608 70868 26648
rect 70828 26188 70868 26228
rect 70732 25768 70772 25808
rect 71116 26104 71156 26144
rect 71788 30220 71828 30260
rect 72460 31312 72500 31352
rect 72460 31144 72500 31184
rect 72460 30556 72500 30596
rect 72364 30388 72404 30428
rect 72268 30220 72308 30260
rect 72076 29968 72116 30008
rect 72268 29968 72308 30008
rect 72172 29800 72212 29840
rect 71788 29044 71828 29084
rect 71884 28372 71924 28412
rect 72076 28372 72116 28412
rect 71788 28288 71828 28328
rect 72268 29128 72308 29168
rect 72268 28792 72308 28832
rect 72172 28288 72212 28328
rect 71980 28120 72020 28160
rect 71500 27788 71540 27824
rect 71500 27784 71540 27788
rect 71404 27532 71444 27572
rect 71500 27448 71540 27488
rect 71692 27364 71732 27404
rect 72268 27952 72308 27992
rect 71788 27280 71828 27320
rect 71596 27112 71636 27152
rect 71692 26944 71732 26984
rect 72076 26860 72116 26900
rect 71500 26272 71540 26312
rect 72844 31648 72884 31688
rect 73036 31396 73076 31436
rect 72940 31144 72980 31184
rect 74092 32824 74132 32864
rect 73996 31648 74036 31688
rect 73708 31396 73748 31436
rect 72844 30640 72884 30680
rect 72652 30220 72692 30260
rect 73612 31312 73652 31352
rect 73516 31228 73556 31268
rect 73420 30976 73460 31016
rect 73228 30220 73268 30260
rect 73228 30052 73268 30092
rect 72748 29968 72788 30008
rect 72556 29128 72596 29168
rect 72748 28456 72788 28496
rect 73132 29800 73172 29840
rect 73804 31228 73844 31268
rect 73516 30472 73556 30512
rect 73900 30976 73940 31016
rect 74188 31648 74228 31688
rect 73708 30556 73748 30596
rect 73996 30556 74036 30596
rect 73612 30052 73652 30092
rect 73420 29885 73460 29924
rect 73420 29884 73460 29885
rect 73324 29800 73364 29840
rect 73036 28792 73076 28832
rect 72844 28372 72884 28412
rect 72940 28288 72980 28328
rect 72652 27364 72692 27404
rect 72364 26776 72404 26816
rect 71596 26020 71636 26060
rect 72076 26020 72116 26060
rect 71980 25936 72020 25976
rect 71212 25264 71252 25304
rect 71116 25180 71156 25220
rect 71980 25264 72020 25304
rect 71116 24424 71156 24464
rect 70540 22744 70580 22784
rect 70855 22744 70895 22784
rect 71212 24088 71252 24128
rect 71500 23836 71540 23876
rect 71404 23752 71444 23792
rect 71692 24088 71732 24128
rect 71596 23668 71636 23708
rect 71308 23500 71348 23540
rect 71545 22828 71585 22868
rect 71980 25012 72020 25052
rect 72172 25264 72212 25304
rect 72268 25180 72308 25220
rect 71884 24340 71924 24380
rect 72076 24004 72116 24044
rect 71980 23920 72020 23960
rect 72268 24760 72308 24800
rect 74092 30472 74132 30512
rect 73804 30220 73844 30260
rect 73996 29800 74036 29840
rect 73228 28288 73268 28328
rect 73708 28204 73748 28244
rect 73612 28120 73652 28160
rect 73228 27616 73268 27656
rect 73132 27196 73172 27236
rect 72940 27112 72980 27152
rect 72844 26104 72884 26144
rect 73132 26776 73172 26816
rect 72748 26020 72788 26060
rect 72460 25348 72500 25388
rect 72844 25264 72884 25304
rect 72172 23836 72212 23876
rect 73324 26104 73364 26144
rect 73708 26104 73748 26144
rect 73420 25936 73460 25976
rect 73228 25180 73268 25220
rect 73132 25096 73172 25136
rect 73612 25096 73652 25136
rect 72940 24760 72980 24800
rect 72940 24592 72980 24632
rect 72844 24508 72884 24548
rect 72652 23920 72692 23960
rect 72460 23668 72500 23708
rect 72076 23500 72116 23540
rect 72364 23584 72404 23624
rect 72460 23416 72500 23456
rect 72364 23332 72404 23372
rect 71655 22744 71695 22784
rect 71788 22744 71828 22784
rect 72748 23752 72788 23792
rect 73612 24508 73652 24548
rect 73228 23668 73268 23708
rect 73132 23584 73172 23624
rect 72844 23500 72884 23540
rect 73516 23584 73556 23624
rect 73324 23164 73364 23204
rect 73612 23164 73652 23204
rect 73420 22744 73460 22784
rect 73996 28120 74036 28160
rect 73900 25936 73940 25976
rect 73804 23500 73844 23540
rect 74092 24508 74132 24548
rect 74476 35680 74516 35720
rect 74860 35596 74900 35636
rect 76108 37192 76148 37232
rect 76588 37276 76628 37316
rect 75340 37108 75380 37148
rect 75436 36436 75476 36476
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 75916 36688 75956 36728
rect 76492 37192 76532 37232
rect 76204 37108 76244 37148
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 75820 36604 75860 36644
rect 75628 35596 75668 35636
rect 75052 35344 75092 35384
rect 75724 35344 75764 35384
rect 77068 36856 77108 36896
rect 76204 36604 76244 36644
rect 76684 36688 76724 36728
rect 77068 36520 77108 36560
rect 76492 36184 76532 36224
rect 76396 36100 76436 36140
rect 76108 36016 76148 36056
rect 76492 35932 76532 35972
rect 76780 35848 76820 35888
rect 76396 35764 76436 35804
rect 76300 35680 76340 35720
rect 77068 35764 77108 35804
rect 76876 35680 76916 35720
rect 76204 35596 76244 35636
rect 75820 34924 75860 34964
rect 74572 34336 74612 34376
rect 74572 33664 74612 33704
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 76108 34336 76148 34376
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 76300 35344 76340 35384
rect 77260 36604 77300 36644
rect 76876 35176 76916 35216
rect 77068 35176 77108 35216
rect 77260 35176 77300 35216
rect 79180 37276 79220 37316
rect 77548 36184 77588 36224
rect 77452 36100 77492 36140
rect 76780 34924 76820 34964
rect 76300 34840 76340 34880
rect 76876 34840 76916 34880
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 76204 33916 76244 33956
rect 76876 33916 76916 33956
rect 74956 33832 74996 33872
rect 76300 33832 76340 33872
rect 76588 33832 76628 33872
rect 76780 33832 76820 33872
rect 74860 33412 74900 33452
rect 76396 33664 76436 33704
rect 76684 33664 76724 33704
rect 75724 33412 75764 33452
rect 76300 33412 76340 33452
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 74380 31480 74420 31520
rect 74476 31312 74516 31352
rect 74380 31144 74420 31184
rect 74380 27952 74420 27992
rect 74572 28204 74612 28244
rect 74476 27448 74516 27488
rect 74476 26776 74516 26816
rect 74380 26104 74420 26144
rect 74572 26188 74612 26228
rect 74572 26020 74612 26060
rect 74476 24592 74516 24632
rect 74188 23668 74228 23708
rect 74188 23500 74228 23540
rect 74092 22996 74132 23036
rect 73655 22744 73695 22784
rect 73804 22744 73844 22784
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 74956 31312 74996 31352
rect 75436 30640 75476 30680
rect 75052 30472 75092 30512
rect 75532 30388 75572 30428
rect 74956 30220 74996 30260
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 74764 29800 74804 29840
rect 75436 29548 75476 29588
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 74764 27952 74804 27992
rect 74860 27112 74900 27152
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 74956 26692 74996 26732
rect 74860 26608 74900 26648
rect 74764 26020 74804 26060
rect 75244 26440 75284 26480
rect 75436 25936 75476 25976
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 75052 25180 75092 25220
rect 74668 24508 74708 24548
rect 77068 34000 77108 34040
rect 77164 33832 77204 33872
rect 77452 34840 77492 34880
rect 77740 35848 77780 35888
rect 78028 35848 78068 35888
rect 77644 35344 77684 35384
rect 77356 33916 77396 33956
rect 77548 34336 77588 34376
rect 77452 33832 77492 33872
rect 77452 33664 77492 33704
rect 77356 33496 77396 33536
rect 79468 35848 79508 35888
rect 79084 35764 79124 35804
rect 78412 35092 78452 35132
rect 78316 34504 78356 34544
rect 77836 34336 77876 34376
rect 77932 34084 77972 34124
rect 78316 34252 78356 34292
rect 78220 34084 78260 34124
rect 78028 34000 78068 34040
rect 77644 33664 77684 33704
rect 77644 33496 77684 33536
rect 76780 32824 76820 32864
rect 76972 32824 77012 32864
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 76780 32418 76820 32444
rect 76780 32404 76820 32418
rect 76492 32320 76532 32360
rect 75916 32152 75956 32192
rect 76300 31480 76340 31520
rect 76108 31396 76148 31436
rect 76012 31312 76052 31352
rect 76684 32236 76724 32276
rect 76972 32152 77012 32192
rect 76588 31648 76628 31688
rect 76588 31480 76628 31520
rect 77356 32824 77396 32864
rect 77644 32824 77684 32864
rect 77260 31564 77300 31604
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 76300 30640 76340 30680
rect 76012 30472 76052 30512
rect 75724 30388 75764 30428
rect 75628 29968 75668 30008
rect 75820 29968 75860 30008
rect 76876 29968 76916 30008
rect 75916 29296 75956 29336
rect 75820 29212 75860 29252
rect 76780 29884 76820 29924
rect 76684 29800 76724 29840
rect 76204 29716 76244 29756
rect 76876 29716 76916 29756
rect 77260 31060 77300 31100
rect 77548 31648 77588 31688
rect 78220 33664 78260 33704
rect 78220 32824 78260 32864
rect 78124 32404 78164 32444
rect 77932 32236 77972 32276
rect 77836 31564 77876 31604
rect 77644 31312 77684 31352
rect 78124 31900 78164 31940
rect 78028 31396 78068 31436
rect 77740 31228 77780 31268
rect 77452 31060 77492 31100
rect 77260 30556 77300 30596
rect 77452 30556 77492 30596
rect 77260 30220 77300 30260
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 76588 29296 76628 29336
rect 76492 29212 76532 29252
rect 76108 29128 76148 29168
rect 77068 29296 77108 29336
rect 76972 29212 77012 29252
rect 75724 28288 75764 28328
rect 75724 27616 75764 27656
rect 75724 27364 75764 27404
rect 77068 29160 77108 29168
rect 77068 29128 77108 29160
rect 77356 29800 77396 29840
rect 78124 31228 78164 31268
rect 78028 30220 78068 30260
rect 77836 29884 77876 29924
rect 77740 29716 77780 29756
rect 77644 29128 77684 29168
rect 78028 29128 78068 29168
rect 77164 28876 77204 28916
rect 78508 34336 78548 34376
rect 78796 33664 78836 33704
rect 79372 31900 79412 31940
rect 78412 31312 78452 31352
rect 78220 30640 78260 30680
rect 78700 29128 78740 29168
rect 79468 29128 79508 29168
rect 77932 28876 77972 28916
rect 76876 28288 76916 28328
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 76012 27700 76052 27740
rect 76876 27700 76916 27740
rect 76204 27616 76244 27656
rect 76588 27616 76628 27656
rect 75916 27532 75956 27572
rect 76108 27532 76148 27572
rect 76492 27532 76532 27572
rect 76396 27448 76436 27488
rect 76300 27364 76340 27404
rect 75820 26776 75860 26816
rect 75820 26188 75860 26228
rect 75628 25936 75668 25976
rect 76012 26104 76052 26144
rect 75916 25936 75956 25976
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 76588 26272 76628 26312
rect 77260 27532 77300 27572
rect 77452 28036 77492 28076
rect 77548 27616 77588 27656
rect 77740 28288 77780 28328
rect 77836 27616 77876 27656
rect 77356 26776 77396 26816
rect 77836 27364 77876 27404
rect 77740 27028 77780 27068
rect 77932 27028 77972 27068
rect 77836 26608 77876 26648
rect 76204 25936 76244 25976
rect 75916 25264 75956 25304
rect 76684 26104 76724 26144
rect 76300 25264 76340 25304
rect 76492 25264 76532 25304
rect 77260 26104 77300 26144
rect 76876 25936 76916 25976
rect 77740 26440 77780 26480
rect 77644 26272 77684 26312
rect 77356 25264 77396 25304
rect 76972 25180 77012 25220
rect 76876 25096 76916 25136
rect 75532 24928 75572 24968
rect 75532 24760 75572 24800
rect 75244 24676 75284 24716
rect 75436 24676 75476 24716
rect 75148 24508 75188 24548
rect 75628 24592 75668 24632
rect 75436 24424 75476 24464
rect 75244 24340 75284 24380
rect 75052 24256 75092 24296
rect 75532 24340 75572 24380
rect 75148 23752 75188 23792
rect 75436 23668 75476 23708
rect 74860 23584 74900 23624
rect 74572 23500 74612 23540
rect 74345 22996 74385 23036
rect 74055 22744 74095 22784
rect 74188 22744 74228 22784
rect 75148 23500 75188 23540
rect 74745 22744 74785 22784
rect 75255 22996 75295 23036
rect 75820 24928 75860 24968
rect 75916 24508 75956 24548
rect 75820 24088 75860 24128
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 76204 24844 76244 24884
rect 76108 24508 76148 24548
rect 76684 24760 76724 24800
rect 76396 24676 76436 24716
rect 76012 24088 76052 24128
rect 76108 23584 76148 23624
rect 76780 24004 76820 24044
rect 76684 23920 76724 23960
rect 76972 25012 77012 25052
rect 77068 24760 77108 24800
rect 77068 24592 77108 24632
rect 76492 23584 76532 23624
rect 76876 23584 76916 23624
rect 76396 23500 76436 23540
rect 76300 23332 76340 23372
rect 76300 23164 76340 23204
rect 75820 22744 75860 22784
rect 76055 22744 76095 22784
rect 77548 25264 77588 25304
rect 77452 24004 77492 24044
rect 77260 23920 77300 23960
rect 77068 23584 77108 23624
rect 77260 23584 77300 23624
rect 77164 23332 77204 23372
rect 78124 27028 78164 27068
rect 78604 27364 78644 27404
rect 78316 27280 78356 27320
rect 78508 26776 78548 26816
rect 78220 26608 78260 26648
rect 78028 26440 78068 26480
rect 77932 26272 77972 26312
rect 78220 25264 78260 25304
rect 78124 25096 78164 25136
rect 76855 22744 76895 22784
rect 77145 22744 77185 22784
rect 77545 22996 77585 23036
rect 79468 27364 79508 27404
rect 78220 22912 78260 22952
rect 77945 22744 77985 22784
rect 78055 22744 78095 22784
rect 79276 25264 79316 25304
rect 78892 25096 78932 25136
rect 78796 23584 78836 23624
rect 78700 23164 78740 23204
rect 78988 23920 79028 23960
rect 78988 23752 79028 23792
rect 79084 23584 79124 23624
rect 79084 23332 79124 23372
rect 79564 23584 79604 23624
rect 78892 22912 78932 22952
rect 78604 22744 78644 22784
rect 79655 22996 79695 23036
rect 53068 21568 53108 21608
rect 53068 18628 53108 18668
rect 53068 17368 53108 17408
rect 52876 17200 52916 17240
rect 52780 17032 52820 17072
rect 52588 16948 52628 16988
rect 52300 16864 52340 16904
rect 52012 16780 52052 16820
rect 52684 16696 52724 16736
rect 52588 16528 52628 16568
rect 52780 16528 52820 16568
rect 52204 16192 52244 16232
rect 52300 16024 52340 16064
rect 51916 15772 51956 15812
rect 52588 16108 52628 16148
rect 52588 15688 52628 15728
rect 51820 15100 51860 15140
rect 52588 15436 52628 15476
rect 54745 17284 54785 17324
rect 54455 17200 54495 17240
rect 53548 16948 53588 16988
rect 53452 16864 53492 16904
rect 54028 16780 54068 16820
rect 53932 16528 53972 16568
rect 53356 16192 53396 16232
rect 53356 15856 53396 15896
rect 53356 15604 53396 15644
rect 51724 14932 51764 14972
rect 52492 14932 52532 14972
rect 51628 14764 51668 14804
rect 51916 14848 51956 14888
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 51436 13420 51476 13460
rect 51724 13924 51764 13964
rect 50956 13168 50996 13208
rect 51244 13000 51284 13040
rect 50572 12496 50612 12536
rect 50380 11068 50420 11108
rect 49036 9472 49076 9512
rect 48748 8716 48788 8756
rect 49996 10060 50036 10100
rect 49420 9724 49460 9764
rect 49516 9388 49556 9428
rect 49132 8884 49172 8924
rect 48940 8632 48980 8672
rect 49324 8716 49364 8756
rect 48844 8548 48884 8588
rect 48652 8464 48692 8504
rect 49420 8548 49460 8588
rect 49036 8464 49076 8504
rect 48460 7960 48500 8000
rect 49708 9556 49748 9596
rect 49900 8800 49940 8840
rect 49708 8716 49748 8756
rect 50284 10900 50324 10940
rect 51052 12496 51092 12536
rect 51148 12412 51188 12452
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 51628 13168 51668 13208
rect 53548 16192 53588 16232
rect 53452 15184 53492 15224
rect 53452 14932 53492 14972
rect 52012 14596 52052 14636
rect 51916 13840 51956 13880
rect 51820 13420 51860 13460
rect 52108 14512 52148 14552
rect 52780 14548 52820 14552
rect 52780 14512 52820 14548
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 53164 14680 53204 14720
rect 53260 14596 53300 14636
rect 53068 14428 53108 14468
rect 52108 14260 52148 14300
rect 52876 14260 52916 14300
rect 53260 14260 53300 14300
rect 53260 14092 53300 14132
rect 52780 14008 52820 14048
rect 52204 13840 52244 13880
rect 51724 13084 51764 13124
rect 51724 12916 51764 12956
rect 51628 12412 51668 12452
rect 50956 11656 50996 11696
rect 51724 11908 51764 11948
rect 51916 13084 51956 13124
rect 51820 11656 51860 11696
rect 51052 11488 51092 11528
rect 51532 11572 51572 11612
rect 53452 14680 53492 14720
rect 53644 14680 53684 14720
rect 53548 14428 53588 14468
rect 53356 13840 53396 13880
rect 53836 14764 53876 14804
rect 53740 14008 53780 14048
rect 54028 14680 54068 14720
rect 54220 14680 54260 14720
rect 53932 14344 53972 14384
rect 54892 16864 54932 16904
rect 55084 16696 55124 16736
rect 55180 16612 55220 16652
rect 54892 16192 54932 16232
rect 54796 15772 54836 15812
rect 54604 15268 54644 15308
rect 54700 15184 54740 15224
rect 54604 14848 54644 14888
rect 54508 14512 54548 14552
rect 54412 14344 54452 14384
rect 54316 14260 54356 14300
rect 54508 13840 54548 13880
rect 55276 16192 55316 16232
rect 55660 16276 55700 16316
rect 56745 17284 56785 17324
rect 57145 17284 57185 17324
rect 57255 17284 57295 17324
rect 56455 17200 56495 17240
rect 56855 17200 56895 17240
rect 57545 17200 57585 17240
rect 57655 17200 57695 17240
rect 58055 17200 58095 17240
rect 57945 17116 57985 17156
rect 58745 17284 58785 17324
rect 58855 17284 58895 17324
rect 58455 17200 58495 17240
rect 59255 17284 59295 17324
rect 59545 17284 59585 17324
rect 59655 17284 59695 17324
rect 59692 17116 59732 17156
rect 56044 16444 56084 16484
rect 56332 16444 56372 16484
rect 55948 16108 55988 16148
rect 55564 15940 55604 15980
rect 55948 15940 55988 15980
rect 55756 15520 55796 15560
rect 55468 15436 55508 15476
rect 55852 15436 55892 15476
rect 55084 14848 55124 14888
rect 55468 14680 55508 14720
rect 54700 14428 54740 14468
rect 54796 14260 54836 14300
rect 54700 13420 54740 13460
rect 53836 13168 53876 13208
rect 54316 13168 54356 13208
rect 53644 13084 53684 13124
rect 52204 12916 52244 12956
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 52780 12748 52820 12788
rect 52588 12664 52628 12704
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 53740 11908 53780 11948
rect 55372 14008 55412 14048
rect 55756 13756 55796 13796
rect 55180 13420 55220 13460
rect 55564 13420 55604 13460
rect 55276 13168 55316 13208
rect 55468 13084 55508 13124
rect 55084 13000 55124 13040
rect 54796 11824 54836 11864
rect 53356 11740 53396 11780
rect 54124 11236 54164 11276
rect 51628 11152 51668 11192
rect 52780 11152 52820 11192
rect 50860 10816 50900 10856
rect 51340 10732 51380 10772
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 51244 10396 51284 10436
rect 50476 10144 50516 10184
rect 50284 9556 50324 9596
rect 50188 8716 50228 8756
rect 50956 10228 50996 10268
rect 51724 10900 51764 10940
rect 51724 10732 51764 10772
rect 51148 10144 51188 10184
rect 51436 10144 51476 10184
rect 51340 10060 51380 10100
rect 51532 10060 51572 10100
rect 51148 9472 51188 9512
rect 50764 9052 50804 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 50764 8884 50804 8924
rect 51244 8884 51284 8924
rect 50668 8800 50708 8840
rect 49612 8128 49652 8168
rect 50092 8128 50132 8168
rect 50284 8128 50324 8168
rect 50380 7372 50420 7412
rect 50860 8632 50900 8672
rect 51628 8884 51668 8924
rect 51628 8716 51668 8756
rect 52108 10984 52148 11024
rect 52012 10900 52052 10940
rect 52396 10900 52436 10940
rect 52876 10984 52916 11024
rect 52012 10648 52052 10688
rect 52012 10228 52052 10268
rect 51916 10060 51956 10100
rect 52204 10144 52244 10184
rect 52108 9640 52148 9680
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 52012 9472 52052 9512
rect 52108 8800 52148 8840
rect 52300 8800 52340 8840
rect 51724 8406 51764 8420
rect 51724 8380 51764 8406
rect 52876 10480 52916 10520
rect 54124 10480 54164 10520
rect 53452 10312 53492 10352
rect 52972 10060 53012 10100
rect 52876 8716 52916 8756
rect 52588 8632 52628 8672
rect 50668 7960 50708 8000
rect 50572 7372 50612 7412
rect 50188 6700 50228 6740
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 52588 8128 52628 8168
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 50956 6952 50996 6992
rect 51820 7120 51860 7160
rect 51724 6532 51764 6572
rect 50380 6364 50420 6404
rect 55756 13168 55796 13208
rect 56140 15856 56180 15896
rect 56044 15604 56084 15644
rect 56044 14680 56084 14720
rect 56044 14344 56084 14384
rect 57292 16780 57332 16820
rect 56620 16696 56660 16736
rect 57004 16444 57044 16484
rect 59596 17032 59636 17072
rect 58348 16528 58388 16568
rect 58732 16276 58772 16316
rect 56620 15772 56660 15812
rect 57004 16192 57044 16232
rect 56908 15940 56948 15980
rect 56428 15688 56468 15728
rect 56716 15688 56756 15728
rect 57100 15520 57140 15560
rect 56908 15100 56948 15140
rect 56716 14764 56756 14804
rect 56908 14680 56948 14720
rect 56620 14008 56660 14048
rect 56524 13756 56564 13796
rect 56332 13672 56372 13712
rect 55852 13084 55892 13124
rect 55756 13000 55796 13040
rect 55660 12916 55700 12956
rect 55564 12664 55604 12704
rect 56428 13168 56468 13208
rect 56524 13084 56564 13124
rect 56332 13000 56372 13040
rect 55276 11824 55316 11864
rect 55468 11740 55508 11780
rect 55180 11152 55220 11192
rect 55180 10984 55220 11024
rect 54796 10900 54836 10940
rect 55084 10900 55124 10940
rect 54796 10732 54836 10772
rect 54988 10312 55028 10352
rect 55084 10228 55124 10268
rect 54700 10060 54740 10100
rect 53836 9640 53876 9680
rect 53356 9304 53396 9344
rect 53068 7876 53108 7916
rect 52876 7372 52916 7412
rect 52108 6952 52148 6992
rect 52588 6952 52628 6992
rect 51916 6280 51956 6320
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 52684 6616 52724 6656
rect 55180 10060 55220 10100
rect 54796 9976 54836 10016
rect 54508 8632 54548 8672
rect 56044 12580 56084 12620
rect 56236 12668 56276 12704
rect 56236 12664 56276 12668
rect 56140 12496 56180 12536
rect 56140 11992 56180 12032
rect 56044 11908 56084 11948
rect 55948 11656 55988 11696
rect 56428 12580 56468 12620
rect 56620 12580 56660 12620
rect 56716 12496 56756 12536
rect 56812 12412 56852 12452
rect 56236 11908 56276 11948
rect 56524 11908 56564 11948
rect 56620 11824 56660 11864
rect 56428 11740 56468 11780
rect 56332 11656 56372 11696
rect 56044 11488 56084 11528
rect 55564 11320 55604 11360
rect 55948 11320 55988 11360
rect 55468 10144 55508 10184
rect 55756 10984 55796 11024
rect 56140 11320 56180 11360
rect 55948 10816 55988 10856
rect 55948 10648 55988 10688
rect 55852 10228 55892 10268
rect 55372 10060 55412 10100
rect 54892 8632 54932 8672
rect 53836 8128 53876 8168
rect 54124 8128 54164 8168
rect 53548 7876 53588 7916
rect 54316 7960 54356 8000
rect 54700 8132 54740 8168
rect 54700 8128 54740 8132
rect 54796 8044 54836 8084
rect 54412 7876 54452 7916
rect 54220 7708 54260 7748
rect 53452 7456 53492 7496
rect 53356 7288 53396 7328
rect 52588 6448 52628 6488
rect 52876 6616 52916 6656
rect 52972 6364 53012 6404
rect 45772 4936 45812 4976
rect 51724 4768 51764 4808
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 52300 6280 52340 6320
rect 52684 5692 52724 5732
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 52876 5692 52916 5732
rect 52204 4852 52244 4892
rect 53644 7456 53684 7496
rect 53164 6616 53204 6656
rect 53548 6532 53588 6572
rect 53452 6448 53492 6488
rect 53740 7372 53780 7412
rect 54604 7456 54644 7496
rect 54892 7960 54932 8000
rect 54988 7876 55028 7916
rect 54796 7372 54836 7412
rect 54220 6616 54260 6656
rect 53164 6280 53204 6320
rect 53548 6280 53588 6320
rect 52876 4852 52916 4892
rect 52396 4768 52436 4808
rect 52588 4768 52628 4808
rect 54220 5776 54260 5816
rect 53356 4852 53396 4892
rect 53164 4768 53204 4808
rect 55756 8632 55796 8672
rect 55660 8380 55700 8420
rect 55564 7792 55604 7832
rect 55180 7708 55220 7748
rect 55468 7708 55508 7748
rect 55276 7036 55316 7076
rect 54988 6616 55028 6656
rect 55084 6532 55124 6572
rect 55564 6532 55604 6572
rect 55372 6448 55412 6488
rect 55852 7960 55892 8000
rect 56044 9976 56084 10016
rect 56236 10984 56276 11024
rect 56236 10396 56276 10436
rect 56236 10228 56276 10268
rect 56524 10312 56564 10352
rect 56332 10144 56372 10184
rect 56140 9388 56180 9428
rect 56044 8632 56084 8672
rect 56332 9220 56372 9260
rect 56332 8632 56372 8672
rect 56140 8044 56180 8084
rect 56044 7960 56084 8000
rect 58156 16192 58196 16232
rect 57196 13420 57236 13460
rect 57772 15940 57812 15980
rect 57964 15772 58004 15812
rect 57868 15436 57908 15476
rect 58348 15772 58388 15812
rect 58540 15772 58580 15812
rect 58444 15604 58484 15644
rect 58348 15520 58388 15560
rect 58444 15100 58484 15140
rect 57580 14764 57620 14804
rect 57388 14092 57428 14132
rect 57388 13924 57428 13964
rect 57964 14008 58004 14048
rect 57676 13840 57716 13880
rect 57580 13252 57620 13292
rect 57292 13168 57332 13208
rect 57196 12580 57236 12620
rect 58060 13924 58100 13964
rect 58636 15520 58676 15560
rect 58924 15772 58964 15812
rect 58828 15436 58868 15476
rect 58636 15184 58676 15224
rect 59500 16276 59540 16316
rect 59596 16192 59636 16232
rect 59116 15856 59156 15896
rect 59404 15772 59444 15812
rect 59116 15688 59156 15728
rect 59020 15352 59060 15392
rect 58636 14680 58676 14720
rect 58924 14512 58964 14552
rect 59116 14512 59156 14552
rect 58252 13840 58292 13880
rect 58060 13672 58100 13712
rect 57964 13168 58004 13208
rect 57100 12496 57140 12536
rect 57100 11824 57140 11864
rect 57484 10984 57524 11024
rect 57772 10984 57812 11024
rect 56908 10732 56948 10772
rect 56908 10312 56948 10352
rect 57100 9472 57140 9512
rect 57484 9220 57524 9260
rect 57868 9052 57908 9092
rect 56908 8632 56948 8672
rect 56812 7456 56852 7496
rect 55756 6532 55796 6572
rect 55948 6532 55988 6572
rect 55660 6448 55700 6488
rect 56044 6280 56084 6320
rect 54796 5104 54836 5144
rect 54124 4768 54164 4808
rect 54220 4684 54260 4724
rect 53068 4264 53108 4304
rect 53836 4180 53876 4220
rect 55564 5608 55604 5648
rect 57100 7120 57140 7160
rect 56716 7036 56756 7076
rect 56332 6868 56372 6908
rect 56620 6868 56660 6908
rect 55756 5104 55796 5144
rect 55852 4936 55892 4976
rect 54700 4852 54740 4892
rect 55180 4852 55220 4892
rect 54508 4684 54548 4724
rect 56236 5608 56276 5648
rect 58060 12496 58100 12536
rect 58060 12076 58100 12116
rect 58252 11152 58292 11192
rect 58444 11152 58484 11192
rect 58252 10144 58292 10184
rect 58156 9976 58196 10016
rect 58444 10228 58484 10268
rect 57964 7960 58004 8000
rect 57868 7036 57908 7076
rect 57964 6868 58004 6908
rect 57580 6532 57620 6572
rect 56812 6448 56852 6488
rect 56908 6364 56948 6404
rect 56524 5776 56564 5816
rect 56236 4936 56276 4976
rect 56044 4768 56084 4808
rect 55084 4264 55124 4304
rect 54604 4180 54644 4220
rect 54412 4096 54452 4136
rect 52108 3928 52148 3968
rect 54220 3928 54260 3968
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 5164 3592 5204 3632
rect 7372 3592 7412 3632
rect 56332 4096 56372 4136
rect 57484 5608 57524 5648
rect 57004 4936 57044 4976
rect 58252 8632 58292 8672
rect 58828 14344 58868 14384
rect 58732 13840 58772 13880
rect 58828 13672 58868 13712
rect 60055 17116 60095 17156
rect 60455 17200 60495 17240
rect 60855 17200 60895 17240
rect 61036 17116 61076 17156
rect 59692 14764 59732 14804
rect 60076 16948 60116 16988
rect 59788 14176 59828 14216
rect 59212 14008 59252 14048
rect 59212 13840 59252 13880
rect 59116 13420 59156 13460
rect 58924 13168 58964 13208
rect 59116 13084 59156 13124
rect 58636 11992 58676 12032
rect 58636 10900 58676 10940
rect 59116 11656 59156 11696
rect 59788 13756 59828 13796
rect 59692 13420 59732 13460
rect 60076 15772 60116 15812
rect 59980 13924 60020 13964
rect 59980 13504 60020 13544
rect 59596 13168 59636 13208
rect 59500 12664 59540 12704
rect 59308 12496 59348 12536
rect 58732 10144 58772 10184
rect 58636 10060 58676 10100
rect 58732 9472 58772 9512
rect 58540 9052 58580 9092
rect 58636 8800 58676 8840
rect 59692 11152 59732 11192
rect 59596 10564 59636 10604
rect 59788 10648 59828 10688
rect 59500 10144 59540 10184
rect 59116 10060 59156 10100
rect 59308 10060 59348 10100
rect 58924 9976 58964 10016
rect 59020 9892 59060 9932
rect 59404 10012 59444 10016
rect 59404 9976 59444 10012
rect 59596 9976 59636 10016
rect 60172 15352 60212 15392
rect 60172 14764 60212 14804
rect 60748 16612 60788 16652
rect 60748 16360 60788 16400
rect 60364 16276 60404 16316
rect 60460 16192 60500 16232
rect 61255 17284 61295 17324
rect 62055 17284 62095 17324
rect 62455 17200 62495 17240
rect 61132 16360 61172 16400
rect 60556 16108 60596 16148
rect 61036 16108 61076 16148
rect 60940 15856 60980 15896
rect 61420 16024 61460 16064
rect 61420 15856 61460 15896
rect 60940 15520 60980 15560
rect 60460 15016 60500 15056
rect 60364 14764 60404 14804
rect 60268 14260 60308 14300
rect 60652 14848 60692 14888
rect 60556 13924 60596 13964
rect 60460 13756 60500 13796
rect 60172 13588 60212 13628
rect 60172 13420 60212 13460
rect 60364 13420 60404 13460
rect 60268 13336 60308 13376
rect 60076 12664 60116 12704
rect 60844 14596 60884 14636
rect 60748 13840 60788 13880
rect 60364 12916 60404 12956
rect 60652 12916 60692 12956
rect 59980 10564 60020 10604
rect 60172 10984 60212 11024
rect 60172 10228 60212 10268
rect 60268 9976 60308 10016
rect 59116 9052 59156 9092
rect 59116 8800 59156 8840
rect 59020 8548 59060 8588
rect 58348 8128 58388 8168
rect 58444 7960 58484 8000
rect 60172 9388 60212 9428
rect 59308 9052 59348 9092
rect 59404 8132 59444 8168
rect 59404 8128 59444 8132
rect 60652 12496 60692 12536
rect 60652 10816 60692 10856
rect 60556 10564 60596 10604
rect 60460 10228 60500 10268
rect 60460 10060 60500 10100
rect 59692 8128 59732 8168
rect 59500 8044 59540 8084
rect 59308 7960 59348 8000
rect 59596 7960 59636 8000
rect 61132 15520 61172 15560
rect 61228 15436 61268 15476
rect 61612 15016 61652 15056
rect 61036 14848 61076 14888
rect 61324 14848 61364 14888
rect 61420 14680 61460 14720
rect 61324 14176 61364 14216
rect 61036 14092 61076 14132
rect 61228 14008 61268 14048
rect 61228 13000 61268 13040
rect 61036 11824 61076 11864
rect 60940 11068 60980 11108
rect 61324 12748 61364 12788
rect 61132 11236 61172 11276
rect 60844 9304 60884 9344
rect 60748 8884 60788 8924
rect 60556 7960 60596 8000
rect 59884 7120 59924 7160
rect 58828 6952 58868 6992
rect 60844 8044 60884 8084
rect 60652 7036 60692 7076
rect 60076 6952 60116 6992
rect 58348 6448 58388 6488
rect 58348 5776 58388 5816
rect 59404 5692 59444 5732
rect 57964 5524 58004 5564
rect 57772 4768 57812 4808
rect 56524 4180 56564 4220
rect 55084 3424 55124 3464
rect 844 3340 884 3380
rect 2476 3340 2516 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 56044 2752 56084 2792
rect 56716 4096 56756 4136
rect 56428 3928 56468 3968
rect 57388 4180 57428 4220
rect 57100 4096 57140 4136
rect 57292 4096 57332 4136
rect 56524 2752 56564 2792
rect 57676 4096 57716 4136
rect 62956 17116 62996 17156
rect 62764 16864 62804 16904
rect 62572 16528 62612 16568
rect 62284 16108 62324 16148
rect 61996 16024 62036 16064
rect 61900 15688 61940 15728
rect 61900 15436 61940 15476
rect 61900 15268 61940 15308
rect 61804 14848 61844 14888
rect 62284 15436 62324 15476
rect 62476 15268 62516 15308
rect 62092 14680 62132 14720
rect 61996 14512 62036 14552
rect 61708 14176 61748 14216
rect 62092 14092 62132 14132
rect 62860 14932 62900 14972
rect 62380 14512 62420 14552
rect 62284 14008 62324 14048
rect 63820 17200 63860 17240
rect 63244 16444 63284 16484
rect 63628 16780 63668 16820
rect 64455 17284 64495 17324
rect 64345 17200 64385 17240
rect 63916 16696 63956 16736
rect 63916 16444 63956 16484
rect 63436 16108 63476 16148
rect 63148 15940 63188 15980
rect 63532 16024 63572 16064
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 63244 14932 63284 14972
rect 63244 14428 63284 14468
rect 62380 13924 62420 13964
rect 61516 13840 61556 13880
rect 61804 13756 61844 13796
rect 62380 13756 62420 13796
rect 61516 13420 61556 13460
rect 61612 13252 61652 13292
rect 61708 13168 61748 13208
rect 62668 13840 62708 13880
rect 62572 13756 62612 13796
rect 62668 13672 62708 13712
rect 61996 13420 62036 13460
rect 62188 13336 62228 13376
rect 62092 13252 62132 13292
rect 61516 13000 61556 13040
rect 61900 12580 61940 12620
rect 61708 11908 61748 11948
rect 61708 11740 61748 11780
rect 61420 11656 61460 11696
rect 61324 11152 61364 11192
rect 61804 11572 61844 11612
rect 62092 13000 62132 13040
rect 62668 13000 62708 13040
rect 62380 12832 62420 12872
rect 62092 12580 62132 12620
rect 63532 14428 63572 14468
rect 63436 14092 63476 14132
rect 63436 13924 63476 13964
rect 63244 13840 63284 13880
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 62956 13168 62996 13208
rect 63820 16108 63860 16148
rect 64108 15688 64148 15728
rect 63724 14260 63764 14300
rect 64108 14008 64148 14048
rect 63820 13924 63860 13964
rect 63820 13336 63860 13376
rect 63820 13168 63860 13208
rect 63628 13084 63668 13124
rect 63532 12916 63572 12956
rect 62956 12832 62996 12872
rect 63724 12748 63764 12788
rect 61996 11740 62036 11780
rect 63628 12496 63668 12536
rect 62380 11824 62420 11864
rect 62188 11740 62228 11780
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 63148 11656 63188 11696
rect 62284 11572 62324 11612
rect 62092 11152 62132 11192
rect 61900 11068 61940 11108
rect 61900 10816 61940 10856
rect 62092 10900 62132 10940
rect 61996 10732 62036 10772
rect 61132 10396 61172 10436
rect 61900 10144 61940 10184
rect 61132 9388 61172 9428
rect 61420 9388 61460 9428
rect 61324 7960 61364 8000
rect 61036 7120 61076 7160
rect 60748 6532 60788 6572
rect 59884 5944 59924 5984
rect 60076 5860 60116 5900
rect 59884 5524 59924 5564
rect 58252 5440 58292 5480
rect 59788 5440 59828 5480
rect 58060 4936 58100 4976
rect 57964 4180 58004 4220
rect 57292 3424 57332 3464
rect 59788 4936 59828 4976
rect 60940 6448 60980 6488
rect 60556 5020 60596 5060
rect 60460 4936 60500 4976
rect 60748 5020 60788 5060
rect 61132 6448 61172 6488
rect 62764 11156 62804 11192
rect 62764 11152 62804 11156
rect 63340 11572 63380 11612
rect 62476 11068 62516 11108
rect 62284 10732 62324 10772
rect 62188 8884 62228 8924
rect 62092 8212 62132 8252
rect 61804 8044 61844 8084
rect 61612 7036 61652 7076
rect 62188 8044 62228 8084
rect 62284 7708 62324 7748
rect 61708 6700 61748 6740
rect 61132 5860 61172 5900
rect 61036 5440 61076 5480
rect 62092 6700 62132 6740
rect 62188 6532 62228 6572
rect 61900 6448 61940 6488
rect 61324 5440 61364 5480
rect 60172 4012 60212 4052
rect 60076 3928 60116 3968
rect 60364 4096 60404 4136
rect 61036 4348 61076 4388
rect 60748 4264 60788 4304
rect 60652 4012 60692 4052
rect 58636 3424 58676 3464
rect 60172 3508 60212 3548
rect 60076 3424 60116 3464
rect 57484 2836 57524 2876
rect 57868 2836 57908 2876
rect 57100 2752 57140 2792
rect 56716 2584 56756 2624
rect 58540 2752 58580 2792
rect 58732 2584 58772 2624
rect 58924 2584 58964 2624
rect 56332 2500 56372 2540
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 60556 3424 60596 3464
rect 61036 3928 61076 3968
rect 60844 3676 60884 3716
rect 60844 3508 60884 3548
rect 61420 5020 61460 5060
rect 61420 4600 61460 4640
rect 61420 4348 61460 4388
rect 61612 5860 61652 5900
rect 61900 5776 61940 5816
rect 61804 4852 61844 4892
rect 61516 3676 61556 3716
rect 61804 4600 61844 4640
rect 62380 7120 62420 7160
rect 62380 6448 62420 6488
rect 62572 10984 62612 11024
rect 62764 10312 62804 10352
rect 62764 10060 62804 10100
rect 63532 11152 63572 11192
rect 63436 10984 63476 11024
rect 63724 11572 63764 11612
rect 65145 17116 65185 17156
rect 65655 17284 65695 17324
rect 65545 17200 65585 17240
rect 66055 17284 66095 17324
rect 66855 17200 66895 17240
rect 66455 17116 66495 17156
rect 66745 17116 66785 17156
rect 64876 16192 64916 16232
rect 64972 15940 65012 15980
rect 64876 14596 64916 14636
rect 64780 14512 64820 14552
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 65068 15772 65108 15812
rect 66316 17032 66356 17072
rect 67255 17284 67295 17324
rect 67372 17200 67412 17240
rect 67180 17032 67220 17072
rect 65740 16528 65780 16568
rect 65644 16360 65684 16400
rect 65452 16108 65492 16148
rect 65356 15520 65396 15560
rect 65068 15268 65108 15308
rect 65164 15184 65204 15224
rect 65644 15856 65684 15896
rect 65548 15436 65588 15476
rect 65164 14932 65204 14972
rect 65068 14596 65108 14636
rect 65068 14344 65108 14384
rect 64876 13504 64916 13544
rect 64780 12916 64820 12956
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 64204 12412 64244 12452
rect 64780 12412 64820 12452
rect 64396 11824 64436 11864
rect 64876 11656 64916 11696
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 64780 11152 64820 11192
rect 64012 10984 64052 11024
rect 63532 10816 63572 10856
rect 63052 10732 63092 10772
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 62860 9976 62900 10016
rect 62668 8716 62708 8756
rect 62572 7960 62612 8000
rect 61036 2920 61076 2960
rect 60652 2836 60692 2876
rect 60556 2668 60596 2708
rect 60748 2584 60788 2624
rect 60940 2584 60980 2624
rect 61228 2752 61268 2792
rect 61516 2668 61556 2708
rect 61708 2752 61748 2792
rect 61420 2584 61460 2624
rect 61612 2584 61652 2624
rect 61324 2416 61364 2456
rect 58348 1996 58388 2036
rect 59116 1996 59156 2036
rect 60268 1996 60308 2036
rect 59596 1912 59636 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 58732 1492 58772 1532
rect 60268 1492 60308 1532
rect 59884 1072 59924 1112
rect 61132 1912 61172 1952
rect 62476 4264 62516 4304
rect 62284 4096 62324 4136
rect 64972 10564 65012 10604
rect 64684 10396 64724 10436
rect 65740 15520 65780 15560
rect 65452 14512 65492 14552
rect 65644 14512 65684 14552
rect 65260 13168 65300 13208
rect 65164 12496 65204 12536
rect 64684 10228 64724 10268
rect 64012 10144 64052 10184
rect 64876 10144 64916 10184
rect 63148 10060 63188 10100
rect 64204 9976 64244 10016
rect 64396 9976 64436 10016
rect 63532 9640 63572 9680
rect 64012 9640 64052 9680
rect 63340 9304 63380 9344
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 62956 8716 62996 8756
rect 62860 8632 62900 8672
rect 63724 9472 63764 9512
rect 63820 9304 63860 9344
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 64396 9640 64436 9680
rect 64396 9052 64436 9092
rect 63820 8884 63860 8924
rect 64300 8884 64340 8924
rect 63628 8800 63668 8840
rect 63148 8716 63188 8756
rect 63532 8716 63572 8756
rect 63244 8464 63284 8504
rect 63148 8380 63188 8420
rect 63052 8044 63092 8084
rect 63148 7708 63188 7748
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 63532 7120 63572 7160
rect 62764 7036 62804 7076
rect 62668 6952 62708 6992
rect 63532 6700 63572 6740
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 62764 5860 62804 5900
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 63916 8548 63956 8588
rect 65068 9640 65108 9680
rect 64972 9472 65012 9512
rect 64780 9052 64820 9092
rect 64492 8716 64532 8756
rect 64972 8632 65012 8672
rect 64492 8548 64532 8588
rect 64012 8464 64052 8504
rect 64300 8464 64340 8504
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 65068 8548 65108 8588
rect 64588 7288 64628 7328
rect 64780 7120 64820 7160
rect 64012 7036 64052 7076
rect 64396 7036 64436 7076
rect 63724 6616 63764 6656
rect 63052 4264 63092 4304
rect 64204 6952 64244 6992
rect 64588 6952 64628 6992
rect 64108 6616 64148 6656
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 65068 7036 65108 7076
rect 65356 13084 65396 13124
rect 65836 14008 65876 14048
rect 66220 16864 66260 16904
rect 66220 16696 66260 16736
rect 66604 16696 66644 16736
rect 66124 16528 66164 16568
rect 66316 16192 66356 16232
rect 66700 16612 66740 16652
rect 67564 16864 67604 16904
rect 67372 16360 67412 16400
rect 67564 16360 67604 16400
rect 66700 15940 66740 15980
rect 66124 15856 66164 15896
rect 67084 15940 67124 15980
rect 67564 16024 67604 16064
rect 67276 15856 67316 15896
rect 67468 15604 67508 15644
rect 67180 15520 67220 15560
rect 68044 16780 68084 16820
rect 68332 16360 68372 16400
rect 67948 16276 67988 16316
rect 67756 16192 67796 16232
rect 67660 15352 67700 15392
rect 67372 15268 67412 15308
rect 66316 14344 66356 14384
rect 66028 14176 66068 14216
rect 65932 13672 65972 13712
rect 65548 12916 65588 12956
rect 65740 13084 65780 13124
rect 65932 13000 65972 13040
rect 66220 13336 66260 13376
rect 65644 12496 65684 12536
rect 65548 11824 65588 11864
rect 65740 11656 65780 11696
rect 65932 11656 65972 11696
rect 66220 12580 66260 12620
rect 66124 11992 66164 12032
rect 66124 11572 66164 11612
rect 66220 11488 66260 11528
rect 65932 10984 65972 11024
rect 65260 9472 65300 9512
rect 65260 8716 65300 8756
rect 65356 8296 65396 8336
rect 65260 6868 65300 6908
rect 64876 6616 64916 6656
rect 64876 6448 64916 6488
rect 64588 5860 64628 5900
rect 64684 5776 64724 5816
rect 64780 5692 64820 5732
rect 65356 5860 65396 5900
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 65260 5608 65300 5648
rect 66220 11152 66260 11192
rect 66124 10648 66164 10688
rect 65932 9472 65972 9512
rect 65932 8884 65972 8924
rect 66028 8464 66068 8504
rect 65932 8128 65972 8168
rect 66028 7960 66068 8000
rect 66988 14176 67028 14216
rect 66700 13504 66740 13544
rect 66508 13252 66548 13292
rect 66796 13336 66836 13376
rect 67468 14680 67508 14720
rect 67564 14596 67604 14636
rect 67372 13504 67412 13544
rect 67180 13420 67220 13460
rect 67084 13168 67124 13208
rect 66412 13084 66452 13124
rect 66796 13084 66836 13124
rect 66988 13084 67028 13124
rect 66604 12916 66644 12956
rect 66604 12412 66644 12452
rect 67276 13336 67316 13376
rect 67468 13420 67508 13460
rect 67564 13336 67604 13376
rect 67180 12580 67220 12620
rect 67084 11656 67124 11696
rect 67660 13168 67700 13208
rect 67563 13084 67603 13124
rect 68140 16024 68180 16064
rect 68044 15520 68084 15560
rect 68140 15352 68180 15392
rect 67948 14680 67988 14720
rect 68236 14596 68276 14636
rect 68716 16696 68756 16736
rect 68620 16108 68660 16148
rect 68620 15856 68660 15896
rect 68428 15688 68468 15728
rect 68428 15520 68468 15560
rect 68524 15436 68564 15476
rect 68428 14512 68468 14552
rect 68236 13756 68276 13796
rect 68140 13588 68180 13628
rect 68044 13252 68084 13292
rect 68140 13168 68180 13208
rect 68332 13252 68372 13292
rect 68236 13000 68276 13040
rect 67756 12664 67796 12704
rect 67948 12580 67988 12620
rect 67468 11740 67508 11780
rect 66892 11488 66932 11528
rect 66988 11236 67028 11276
rect 66796 10816 66836 10856
rect 66412 10480 66452 10520
rect 66604 10228 66644 10268
rect 66412 10144 66452 10184
rect 66508 10060 66548 10100
rect 66316 8800 66356 8840
rect 66220 8296 66260 8336
rect 66508 8716 66548 8756
rect 66412 8212 66452 8252
rect 66412 7960 66452 8000
rect 66316 7876 66356 7916
rect 65740 7372 65780 7412
rect 65740 7036 65780 7076
rect 65740 6112 65780 6152
rect 65740 5944 65780 5984
rect 65644 5860 65684 5900
rect 65548 5692 65588 5732
rect 65644 5608 65684 5648
rect 65452 5524 65492 5564
rect 62572 3928 62612 3968
rect 62092 3676 62132 3716
rect 61996 3340 62036 3380
rect 63244 3256 63284 3296
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 62092 2920 62132 2960
rect 62764 2920 62804 2960
rect 61036 1072 61076 1112
rect 61900 1912 61940 1952
rect 61324 1828 61364 1868
rect 62668 2836 62708 2876
rect 62476 2752 62516 2792
rect 62284 2584 62324 2624
rect 62572 2668 62612 2708
rect 62188 2452 62228 2456
rect 62188 2416 62228 2452
rect 63628 3928 63668 3968
rect 63340 2668 63380 2708
rect 62860 2584 62900 2624
rect 62956 2416 62996 2456
rect 62764 1996 62804 2036
rect 62764 1660 62804 1700
rect 64588 5104 64628 5144
rect 64972 5104 65012 5144
rect 64876 4936 64916 4976
rect 64972 4852 65012 4892
rect 64492 4264 64532 4304
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 65548 4936 65588 4976
rect 65452 4852 65492 4892
rect 65164 3928 65204 3968
rect 64588 3424 64628 3464
rect 65740 5104 65780 5144
rect 65740 4936 65780 4976
rect 65836 4852 65876 4892
rect 66124 7372 66164 7412
rect 66124 5776 66164 5816
rect 66700 8128 66740 8168
rect 68044 12412 68084 12452
rect 67564 11404 67604 11444
rect 67468 11236 67508 11276
rect 67852 11250 67892 11276
rect 67852 11236 67892 11250
rect 68044 11656 68084 11696
rect 67372 9472 67412 9512
rect 68428 13168 68468 13208
rect 68620 14680 68660 14720
rect 68620 13840 68660 13880
rect 68524 13084 68564 13124
rect 68812 16444 68852 16484
rect 70455 17284 70495 17324
rect 70345 17200 70385 17240
rect 69945 17116 69985 17156
rect 70055 17116 70095 17156
rect 69100 14932 69140 14972
rect 68812 13756 68852 13796
rect 68812 13588 68852 13628
rect 68428 12496 68468 12536
rect 68332 11656 68372 11696
rect 67660 9304 67700 9344
rect 66796 7960 66836 8000
rect 66892 6700 66932 6740
rect 66604 6448 66644 6488
rect 66316 5608 66356 5648
rect 66796 4936 66836 4976
rect 66604 4264 66644 4304
rect 66124 4180 66164 4220
rect 65644 3928 65684 3968
rect 65548 3592 65588 3632
rect 64492 3256 64532 3296
rect 65644 3508 65684 3548
rect 64492 2668 64532 2708
rect 64396 2584 64436 2624
rect 64972 2668 65012 2708
rect 64876 2584 64916 2624
rect 64012 2416 64052 2456
rect 64588 2416 64628 2456
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 63244 2080 63284 2120
rect 64780 2080 64820 2120
rect 65164 2668 65204 2708
rect 65932 3424 65972 3464
rect 66220 3508 66260 3548
rect 66412 3424 66452 3464
rect 67468 8632 67508 8672
rect 68332 10396 68372 10436
rect 68236 10312 68276 10352
rect 68620 12664 68660 12704
rect 69100 14680 69140 14720
rect 69004 13924 69044 13964
rect 69004 13252 69044 13292
rect 68908 13084 68948 13124
rect 69292 16444 69332 16484
rect 69292 16024 69332 16064
rect 69292 14764 69332 14804
rect 69676 16192 69716 16232
rect 69580 16108 69620 16148
rect 69676 15268 69716 15308
rect 69964 16948 70004 16988
rect 70732 16780 70772 16820
rect 71548 17284 71588 17324
rect 71255 17116 71295 17156
rect 72055 17116 72095 17156
rect 70828 16612 70868 16652
rect 69868 16192 69908 16232
rect 69964 15856 70004 15896
rect 69868 15688 69908 15728
rect 69484 14932 69524 14972
rect 69484 14512 69524 14552
rect 69580 13756 69620 13796
rect 69196 12748 69236 12788
rect 68908 12496 68948 12536
rect 68812 12412 68852 12452
rect 68908 10900 68948 10940
rect 68524 10312 68564 10352
rect 68428 10060 68468 10100
rect 68236 9976 68276 10016
rect 67756 8884 67796 8924
rect 67756 5104 67796 5144
rect 67660 3592 67700 3632
rect 67948 8548 67988 8588
rect 68044 8296 68084 8336
rect 68044 7876 68084 7916
rect 68524 9976 68564 10016
rect 68620 9556 68660 9596
rect 69388 12832 69428 12872
rect 69292 10480 69332 10520
rect 68908 10312 68948 10352
rect 69292 10312 69332 10352
rect 68812 9556 68852 9596
rect 68140 7624 68180 7664
rect 68428 7960 68468 8000
rect 68332 7708 68372 7748
rect 68524 7876 68564 7916
rect 68812 8968 68852 9008
rect 69100 10228 69140 10268
rect 69004 8968 69044 9008
rect 68908 8632 68948 8672
rect 69196 10144 69236 10184
rect 69484 12580 69524 12620
rect 69484 11572 69524 11612
rect 70060 15520 70100 15560
rect 70924 16276 70964 16316
rect 71596 16360 71636 16400
rect 71788 16360 71828 16400
rect 71116 16192 71156 16232
rect 70348 15856 70388 15896
rect 70252 15772 70292 15812
rect 69772 14680 69812 14720
rect 69772 14092 69812 14132
rect 69868 13924 69908 13964
rect 70156 14848 70196 14888
rect 70156 14008 70196 14048
rect 69964 13840 70004 13880
rect 70156 13756 70196 13796
rect 69964 13252 70004 13292
rect 69868 13168 69908 13208
rect 70060 12412 70100 12452
rect 69964 10984 70004 11024
rect 69676 10564 69716 10604
rect 70060 10480 70100 10520
rect 70060 10228 70100 10268
rect 69484 9472 69524 9512
rect 69868 8800 69908 8840
rect 69676 8716 69716 8756
rect 69004 8296 69044 8336
rect 68908 8212 68948 8252
rect 70348 15688 70388 15728
rect 70444 15268 70484 15308
rect 70348 14680 70388 14720
rect 70444 14596 70484 14636
rect 70348 14344 70388 14384
rect 70828 15184 70868 15224
rect 70732 14764 70772 14804
rect 70636 14344 70676 14384
rect 70540 14008 70580 14048
rect 70540 13840 70580 13880
rect 70348 13252 70388 13292
rect 70252 11572 70292 11612
rect 70444 11320 70484 11360
rect 70348 10396 70388 10436
rect 71308 15688 71348 15728
rect 70924 14932 70964 14972
rect 71116 14932 71156 14972
rect 71212 14848 71252 14888
rect 71116 14680 71156 14720
rect 71404 14596 71444 14636
rect 70924 14512 70964 14552
rect 70924 14092 70964 14132
rect 71212 13924 71252 13964
rect 70828 13840 70868 13880
rect 70924 13756 70964 13796
rect 70636 13588 70676 13628
rect 70636 13336 70676 13376
rect 70732 13168 70772 13208
rect 70636 12580 70676 12620
rect 70252 10144 70292 10184
rect 70444 9556 70484 9596
rect 70540 9472 70580 9512
rect 70444 8884 70484 8924
rect 70156 8128 70196 8168
rect 69100 7792 69140 7832
rect 68620 7624 68660 7664
rect 68716 7540 68756 7580
rect 69292 7708 69332 7748
rect 67948 6448 67988 6488
rect 68140 6280 68180 6320
rect 68428 6448 68468 6488
rect 68140 5692 68180 5732
rect 68428 5608 68468 5648
rect 68332 5524 68372 5564
rect 68812 6364 68852 6404
rect 69580 6616 69620 6656
rect 69100 6280 69140 6320
rect 68908 5776 68948 5816
rect 69388 5776 69428 5816
rect 68716 5692 68756 5732
rect 68332 4936 68372 4976
rect 68428 4432 68468 4472
rect 68620 4432 68660 4472
rect 68332 4096 68372 4136
rect 66028 2668 66068 2708
rect 66220 2668 66260 2708
rect 66796 2668 66836 2708
rect 63628 1912 63668 1952
rect 65356 1912 65396 1952
rect 63244 1660 63284 1700
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 66220 2080 66260 2120
rect 66220 1912 66260 1952
rect 66892 2584 66932 2624
rect 67564 2584 67604 2624
rect 66700 2416 66740 2456
rect 66796 1996 66836 2036
rect 67660 1996 67700 2036
rect 68140 2416 68180 2456
rect 69292 5608 69332 5648
rect 68812 5524 68852 5564
rect 69004 5524 69044 5564
rect 69196 4936 69236 4976
rect 68908 4264 68948 4304
rect 68716 4012 68756 4052
rect 68428 2584 68468 2624
rect 68812 3592 68852 3632
rect 69196 4096 69236 4136
rect 69004 3676 69044 3716
rect 69196 3340 69236 3380
rect 69676 6448 69716 6488
rect 70828 8632 70868 8672
rect 70828 6616 70868 6656
rect 70540 6448 70580 6488
rect 70732 6448 70772 6488
rect 70156 6364 70196 6404
rect 70444 6364 70484 6404
rect 70060 6280 70100 6320
rect 69772 5692 69812 5732
rect 69676 5524 69716 5564
rect 69676 4264 69716 4304
rect 68812 2416 68852 2456
rect 68620 2178 68660 2204
rect 68620 2164 68660 2178
rect 67756 1912 67796 1952
rect 68044 1912 68084 1952
rect 66220 1660 66260 1700
rect 66604 1660 66644 1700
rect 67372 1660 67412 1700
rect 67180 1156 67220 1196
rect 66796 1072 66836 1112
rect 67948 1744 67988 1784
rect 67756 1072 67796 1112
rect 69100 2164 69140 2204
rect 69196 1996 69236 2036
rect 68620 1744 68660 1784
rect 68524 1660 68564 1700
rect 69484 2584 69524 2624
rect 70348 5608 70388 5648
rect 70156 5104 70196 5144
rect 70540 5020 70580 5060
rect 70060 2836 70100 2876
rect 70156 1996 70196 2036
rect 70060 1912 70100 1952
rect 69772 1660 69812 1700
rect 69580 1492 69620 1532
rect 68428 1072 68468 1112
rect 69484 1072 69524 1112
rect 69676 1156 69716 1196
rect 71020 13588 71060 13628
rect 71116 13504 71156 13544
rect 71404 14008 71444 14048
rect 71116 13168 71156 13208
rect 71308 13336 71348 13376
rect 72076 16192 72116 16232
rect 71980 16024 72020 16064
rect 71884 15184 71924 15224
rect 71596 14008 71636 14048
rect 72268 15772 72308 15812
rect 72172 15688 72212 15728
rect 72460 16612 72500 16652
rect 72460 16444 72500 16484
rect 72556 16276 72596 16316
rect 72556 15940 72596 15980
rect 72364 15604 72404 15644
rect 72076 14848 72116 14888
rect 72268 15520 72308 15560
rect 72460 14596 72500 14636
rect 72172 14512 72212 14552
rect 71692 13924 71732 13964
rect 72268 14344 72308 14384
rect 72268 13924 72308 13964
rect 72172 13336 72212 13376
rect 71404 13084 71444 13124
rect 71596 13168 71636 13208
rect 71980 13168 72020 13208
rect 71788 13084 71828 13124
rect 71020 10060 71060 10100
rect 72076 12916 72116 12956
rect 71980 11824 72020 11864
rect 71884 10984 71924 11024
rect 72076 11488 72116 11528
rect 72556 14344 72596 14384
rect 72460 12916 72500 12956
rect 73132 16612 73172 16652
rect 72844 16528 72884 16568
rect 73132 16360 73172 16400
rect 72844 16276 72884 16316
rect 72748 15688 72788 15728
rect 72940 16108 72980 16148
rect 73420 16444 73460 16484
rect 73516 16360 73556 16400
rect 73420 16276 73460 16316
rect 73420 16024 73460 16064
rect 73612 16024 73652 16064
rect 73228 15940 73268 15980
rect 73132 15688 73172 15728
rect 72844 15436 72884 15476
rect 73439 14932 73479 14972
rect 72748 14848 72788 14888
rect 72652 14176 72692 14216
rect 72652 13168 72692 13208
rect 74188 17200 74228 17240
rect 73996 16444 74036 16484
rect 74668 17116 74708 17156
rect 73900 16276 73940 16316
rect 73708 15772 73748 15812
rect 73708 15436 73748 15476
rect 73439 14680 73479 14720
rect 73036 14512 73076 14552
rect 72844 14176 72884 14216
rect 72940 12916 72980 12956
rect 72748 12664 72788 12704
rect 73132 14008 73172 14048
rect 73228 13420 73268 13460
rect 72556 11656 72596 11696
rect 72460 11572 72500 11612
rect 72364 11524 72404 11528
rect 72364 11488 72404 11524
rect 72268 11404 72308 11444
rect 72844 11824 72884 11864
rect 73132 11824 73172 11864
rect 73324 12412 73364 12452
rect 73612 14512 73652 14552
rect 74092 16192 74132 16232
rect 74188 16024 74228 16064
rect 74380 15940 74420 15980
rect 73804 14176 73844 14216
rect 73804 14008 73844 14048
rect 73804 13168 73844 13208
rect 74188 14680 74228 14720
rect 74092 14008 74132 14048
rect 74284 14176 74324 14216
rect 73996 13420 74036 13460
rect 74188 13336 74228 13376
rect 73708 12664 73748 12704
rect 73324 11740 73364 11780
rect 73508 11656 73516 11696
rect 73516 11656 73548 11696
rect 73612 11656 73652 11696
rect 73900 12664 73940 12704
rect 73804 11656 73844 11696
rect 72748 11320 72788 11360
rect 71692 10144 71732 10184
rect 71500 9472 71540 9512
rect 71980 9472 72020 9512
rect 72268 9556 72308 9596
rect 72364 9388 72404 9428
rect 71692 8884 71732 8924
rect 71788 8716 71828 8756
rect 71692 8296 71732 8336
rect 73132 11236 73172 11276
rect 73036 10480 73076 10520
rect 73516 10900 73556 10940
rect 73132 10312 73172 10352
rect 73324 10312 73364 10352
rect 72940 9640 72980 9680
rect 72652 9556 72692 9596
rect 72844 9472 72884 9512
rect 73036 9388 73076 9428
rect 72556 8884 72596 8924
rect 72364 8464 72404 8504
rect 72268 8296 72308 8336
rect 71404 7708 71444 7748
rect 71404 7204 71444 7244
rect 71020 6616 71060 6656
rect 71308 6448 71348 6488
rect 71788 7708 71828 7748
rect 71884 7120 71924 7160
rect 71692 6280 71732 6320
rect 71500 5608 71540 5648
rect 70924 5104 70964 5144
rect 71020 4936 71060 4976
rect 71308 4684 71348 4724
rect 71212 4180 71252 4220
rect 71020 4096 71060 4136
rect 71404 4180 71444 4220
rect 71116 3928 71156 3968
rect 71788 4936 71828 4976
rect 71692 4264 71732 4304
rect 71500 4096 71540 4136
rect 71596 3928 71636 3968
rect 71884 3928 71924 3968
rect 71788 3844 71828 3884
rect 71596 3172 71636 3212
rect 71404 3004 71444 3044
rect 70924 2836 70964 2876
rect 71308 2584 71348 2624
rect 72172 7960 72212 8000
rect 72172 7204 72212 7244
rect 72268 7120 72308 7160
rect 72652 8800 72692 8840
rect 72844 8716 72884 8756
rect 72652 8464 72692 8504
rect 73420 9640 73460 9680
rect 73612 9472 73652 9512
rect 73804 10396 73844 10436
rect 73420 9220 73460 9260
rect 73516 8968 73556 9008
rect 73516 8800 73556 8840
rect 73228 8212 73268 8252
rect 73900 9220 73940 9260
rect 73804 8716 73844 8756
rect 73708 8128 73748 8168
rect 73708 7960 73748 8000
rect 72460 7708 72500 7748
rect 73036 7288 73076 7328
rect 73612 7288 73652 7328
rect 73516 7204 73556 7244
rect 72748 7120 72788 7160
rect 72076 5944 72116 5984
rect 72172 5692 72212 5732
rect 72460 5944 72500 5984
rect 72940 6448 72980 6488
rect 73036 6280 73076 6320
rect 72076 4180 72116 4220
rect 72268 5608 72308 5648
rect 73228 5776 73268 5816
rect 72652 5608 72692 5648
rect 74284 10900 74324 10940
rect 73996 8968 74036 9008
rect 73900 8464 73940 8504
rect 74092 8632 74132 8672
rect 73996 7204 74036 7244
rect 73804 6868 73844 6908
rect 73804 6280 73844 6320
rect 73420 5608 73460 5648
rect 73324 5440 73364 5480
rect 74572 13924 74612 13964
rect 74476 13420 74516 13460
rect 74855 17200 74895 17240
rect 75255 17116 75295 17156
rect 75655 17116 75695 17156
rect 74764 16192 74804 16232
rect 74476 11908 74516 11948
rect 74668 10984 74708 11024
rect 74956 15436 74996 15476
rect 75628 16276 75668 16316
rect 75340 16108 75380 16148
rect 75628 15604 75668 15644
rect 75724 15520 75764 15560
rect 75340 15268 75380 15308
rect 74860 12748 74900 12788
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 75340 14932 75380 14972
rect 75436 14680 75476 14720
rect 76108 15940 76148 15980
rect 76012 15856 76052 15896
rect 75916 14932 75956 14972
rect 75916 14680 75956 14720
rect 76108 14764 76148 14804
rect 75628 14596 75668 14636
rect 76855 17284 76895 17324
rect 77145 17284 77185 17324
rect 77836 17116 77876 17156
rect 76012 14596 76052 14636
rect 76204 14596 76244 14636
rect 75340 14176 75380 14216
rect 75244 14008 75284 14048
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 75436 13168 75476 13208
rect 76780 15688 76820 15728
rect 76972 15604 77012 15644
rect 76684 15520 76724 15560
rect 76492 15268 76532 15308
rect 76396 14680 76436 14720
rect 76780 15436 76820 15476
rect 76876 14680 76916 14720
rect 76780 14596 76820 14636
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 75820 14176 75860 14216
rect 75724 14008 75764 14048
rect 76012 14008 76052 14048
rect 76012 13252 76052 13292
rect 75916 13084 75956 13124
rect 75436 12748 75476 12788
rect 75052 12664 75092 12704
rect 74764 10396 74804 10436
rect 74572 8884 74612 8924
rect 74476 8716 74516 8756
rect 74092 6868 74132 6908
rect 74092 5608 74132 5648
rect 73996 5356 74036 5396
rect 72460 5020 72500 5060
rect 73996 4936 74036 4976
rect 72940 4684 72980 4724
rect 73132 4684 73172 4724
rect 72076 3964 72116 3968
rect 72076 3928 72116 3964
rect 72556 4012 72596 4052
rect 71884 3592 71924 3632
rect 72076 3172 72116 3212
rect 72268 3760 72308 3800
rect 71788 2584 71828 2624
rect 72076 2752 72116 2792
rect 71788 1912 71828 1952
rect 71116 1828 71156 1868
rect 71500 1492 71540 1532
rect 71212 1156 71252 1196
rect 71116 1072 71156 1112
rect 72172 2584 72212 2624
rect 71692 1408 71732 1448
rect 72076 1408 72116 1448
rect 71596 1324 71636 1364
rect 72364 2752 72404 2792
rect 73132 4096 73172 4136
rect 72652 3844 72692 3884
rect 73036 3592 73076 3632
rect 73132 3256 73172 3296
rect 73612 3256 73652 3296
rect 72940 3172 72980 3212
rect 72748 2668 72788 2708
rect 72844 2584 72884 2624
rect 72652 2080 72692 2120
rect 72652 1912 72692 1952
rect 72460 1492 72500 1532
rect 72844 1072 72884 1112
rect 73132 1072 73172 1112
rect 73996 3760 74036 3800
rect 74380 8128 74420 8168
rect 74284 5776 74324 5816
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 75052 11908 75092 11948
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 75244 10396 75284 10436
rect 75340 9976 75380 10016
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 75052 8716 75092 8756
rect 75532 8716 75572 8756
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 76012 11740 76052 11780
rect 76204 14008 76244 14048
rect 76588 14008 76628 14048
rect 76492 13924 76532 13964
rect 76204 13420 76244 13460
rect 76588 13420 76628 13460
rect 76204 12916 76244 12956
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 76876 13336 76916 13376
rect 77068 13336 77108 13376
rect 76396 12664 76436 12704
rect 76780 12496 76820 12536
rect 77356 15436 77396 15476
rect 77260 14344 77300 14384
rect 77644 15856 77684 15896
rect 77740 15688 77780 15728
rect 77548 14260 77588 14300
rect 77932 15100 77972 15140
rect 77836 14764 77876 14804
rect 77740 14680 77780 14720
rect 77356 14008 77396 14048
rect 77644 14008 77684 14048
rect 77452 13924 77492 13964
rect 77164 13252 77204 13292
rect 77260 12942 77300 12956
rect 77260 12916 77300 12942
rect 76684 11740 76724 11780
rect 77548 13336 77588 13376
rect 77836 13336 77876 13376
rect 77740 13168 77780 13208
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 77068 11152 77108 11192
rect 75820 10060 75860 10100
rect 75052 7036 75092 7076
rect 74956 6616 74996 6656
rect 74476 5776 74516 5816
rect 74380 5608 74420 5648
rect 74572 5440 74612 5480
rect 74284 4264 74324 4304
rect 74380 4012 74420 4052
rect 75052 6448 75092 6488
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 74956 5776 74996 5816
rect 74668 4936 74708 4976
rect 74572 4432 74612 4472
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 75724 7204 75764 7244
rect 75628 7120 75668 7160
rect 75820 7036 75860 7076
rect 75628 6616 75668 6656
rect 75820 4936 75860 4976
rect 76684 10312 76724 10352
rect 76492 9976 76532 10016
rect 77164 10984 77204 11024
rect 77356 12328 77396 12368
rect 77356 12160 77396 12200
rect 77452 11740 77492 11780
rect 77068 10228 77108 10268
rect 77356 10732 77396 10772
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 76972 10144 77012 10184
rect 77356 9976 77396 10016
rect 77068 9892 77108 9932
rect 76492 8800 76532 8840
rect 76396 8716 76436 8756
rect 76876 8800 76916 8840
rect 76780 8632 76820 8672
rect 76300 8464 76340 8504
rect 76684 8464 76724 8504
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 76012 7204 76052 7244
rect 76492 7120 76532 7160
rect 76684 7960 76724 8000
rect 76780 7120 76820 7160
rect 76972 7120 77012 7160
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 76012 5692 76052 5732
rect 75148 4264 75188 4304
rect 75532 4264 75572 4304
rect 74956 4180 74996 4220
rect 74572 3004 74612 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 74284 2668 74324 2708
rect 74092 2584 74132 2624
rect 74092 2416 74132 2456
rect 73996 2080 74036 2120
rect 73804 1996 73844 2036
rect 74380 2584 74420 2624
rect 74476 1996 74516 2036
rect 74380 1912 74420 1952
rect 74188 1828 74228 1868
rect 75052 2836 75092 2876
rect 74956 2752 74996 2792
rect 75820 4432 75860 4472
rect 75724 4180 75764 4220
rect 77260 9220 77300 9260
rect 77836 12496 77876 12536
rect 77740 12412 77780 12452
rect 77644 11656 77684 11696
rect 77932 11152 77972 11192
rect 78124 14008 78164 14048
rect 78316 13588 78356 13628
rect 78316 13420 78356 13460
rect 78220 13252 78260 13292
rect 78124 13084 78164 13124
rect 78316 13168 78356 13208
rect 78220 12580 78260 12620
rect 78124 12244 78164 12284
rect 78604 16276 78644 16316
rect 78508 16192 78548 16232
rect 78796 15688 78836 15728
rect 78796 15100 78836 15140
rect 78700 14176 78740 14216
rect 78508 14092 78548 14132
rect 78508 13420 78548 13460
rect 78700 13168 78740 13208
rect 78892 14260 78932 14300
rect 78412 12244 78452 12284
rect 77740 10732 77780 10772
rect 78028 10732 78068 10772
rect 77548 9976 77588 10016
rect 77932 10228 77972 10268
rect 77644 9892 77684 9932
rect 77452 8464 77492 8504
rect 77356 8212 77396 8252
rect 77068 7036 77108 7076
rect 76780 6364 76820 6404
rect 76876 5692 76916 5732
rect 76972 5608 77012 5648
rect 76492 5440 76532 5480
rect 76780 5356 76820 5396
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 76108 4264 76148 4304
rect 75916 3928 75956 3968
rect 75628 2752 75668 2792
rect 74764 1912 74804 1952
rect 74764 1744 74804 1784
rect 75724 2584 75764 2624
rect 75436 1912 75476 1952
rect 75628 1912 75668 1952
rect 76588 4096 76628 4136
rect 77356 7120 77396 7160
rect 78124 10312 78164 10352
rect 78604 10900 78644 10940
rect 77644 7792 77684 7832
rect 77836 8380 77876 8420
rect 78412 9220 78452 9260
rect 78316 8800 78356 8840
rect 78220 8716 78260 8756
rect 78124 8632 78164 8672
rect 78028 8464 78068 8504
rect 77932 7792 77972 7832
rect 77836 7120 77876 7160
rect 78220 7120 78260 7160
rect 78124 7036 78164 7076
rect 77740 6364 77780 6404
rect 77548 5860 77588 5900
rect 77548 5692 77588 5732
rect 77452 5608 77492 5648
rect 77644 5476 77684 5480
rect 77644 5440 77684 5476
rect 77548 5356 77588 5396
rect 76972 4852 77012 4892
rect 76876 4348 76916 4388
rect 76300 3928 76340 3968
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 76684 3508 76724 3548
rect 76300 3256 76340 3296
rect 76300 2584 76340 2624
rect 76588 2584 76628 2624
rect 76108 2416 76148 2456
rect 76396 2416 76436 2456
rect 76780 3424 76820 3464
rect 76780 3256 76820 3296
rect 77260 4852 77300 4892
rect 77164 4348 77204 4388
rect 77356 4264 77396 4304
rect 77068 4180 77108 4220
rect 77452 4096 77492 4136
rect 77068 3844 77108 3884
rect 76972 3424 77012 3464
rect 78028 6952 78068 6992
rect 77836 5692 77876 5732
rect 78508 6616 78548 6656
rect 78124 5608 78164 5648
rect 77836 5020 77876 5060
rect 78316 5440 78356 5480
rect 79255 17116 79295 17156
rect 79084 15856 79124 15896
rect 78988 14092 79028 14132
rect 79372 16276 79412 16316
rect 79180 15688 79220 15728
rect 79372 14176 79412 14216
rect 79372 12496 79412 12536
rect 79276 8716 79316 8756
rect 78988 7960 79028 8000
rect 78700 6952 78740 6992
rect 79468 6616 79508 6656
rect 78604 5020 78644 5060
rect 77644 4768 77684 4808
rect 77644 3676 77684 3716
rect 76972 2668 77012 2708
rect 77164 2668 77204 2708
rect 75820 2080 75860 2120
rect 75820 1912 75860 1952
rect 75532 1744 75572 1784
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 76396 2080 76436 2120
rect 76492 1576 76532 1616
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 75628 1492 75668 1532
rect 76108 1492 76148 1532
rect 74956 1324 74996 1364
rect 76684 1492 76724 1532
rect 76588 1156 76628 1196
rect 71788 988 71828 1028
rect 77068 2500 77108 2540
rect 76972 2416 77012 2456
rect 77068 1912 77108 1952
rect 78220 4936 78260 4976
rect 78124 4180 78164 4220
rect 78028 3424 78068 3464
rect 79372 4180 79412 4220
rect 77644 2584 77684 2624
rect 77932 2584 77972 2624
rect 77836 2500 77876 2540
rect 77452 2080 77492 2120
rect 77356 1996 77396 2036
rect 77260 1912 77300 1952
rect 77164 1576 77204 1616
rect 78412 2584 78452 2624
rect 78220 1912 78260 1952
rect 79372 1156 79412 1196
rect 73228 988 73268 1028
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 16343 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 16729 38576
rect 28343 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 28729 38576
rect 40343 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 40729 38576
rect 52343 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 52729 38576
rect 64343 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 64729 38576
rect 76343 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 76729 38576
rect 69571 38368 69580 38408
rect 69620 38368 75916 38408
rect 75956 38368 75965 38408
rect 50275 38240 50333 38241
rect 50275 38200 50284 38240
rect 50324 38200 68332 38240
rect 68372 38200 68381 38240
rect 50275 38199 50333 38200
rect 63811 38116 63820 38156
rect 63860 38116 64684 38156
rect 64724 38116 67756 38156
rect 67796 38116 67805 38156
rect 62275 38032 62284 38072
rect 62324 38032 65452 38072
rect 65492 38032 65501 38072
rect 66499 38032 66508 38072
rect 66548 38032 66892 38072
rect 66932 38032 69580 38072
rect 69620 38032 69629 38072
rect 65827 37948 65836 37988
rect 65876 37948 67468 37988
rect 67508 37948 67517 37988
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 15103 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 15489 37820
rect 27103 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 27489 37820
rect 39103 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 39489 37820
rect 51103 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 51489 37820
rect 63103 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 63489 37820
rect 75103 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 75489 37820
rect 75043 37612 75052 37652
rect 75092 37612 75628 37652
rect 75668 37612 76204 37652
rect 76244 37612 76253 37652
rect 0 37568 80 37588
rect 0 37528 652 37568
rect 692 37528 701 37568
rect 69379 37528 69388 37568
rect 69428 37528 70060 37568
rect 70100 37528 70109 37568
rect 0 37508 80 37528
rect 64387 37444 64396 37484
rect 64436 37444 65260 37484
rect 65300 37444 65309 37484
rect 67363 37444 67372 37484
rect 67412 37444 68428 37484
rect 68468 37444 70636 37484
rect 70676 37444 70685 37484
rect 74659 37444 74668 37484
rect 74708 37444 75340 37484
rect 75380 37444 75389 37484
rect 56515 37360 56524 37400
rect 56564 37360 57004 37400
rect 57044 37360 57580 37400
rect 57620 37360 57629 37400
rect 59395 37360 59404 37400
rect 59444 37360 60940 37400
rect 60980 37360 62188 37400
rect 62228 37360 62237 37400
rect 62755 37360 62764 37400
rect 62804 37360 64492 37400
rect 64532 37360 65164 37400
rect 65204 37360 65213 37400
rect 65539 37360 65548 37400
rect 65588 37360 65932 37400
rect 65972 37360 66700 37400
rect 66740 37360 68908 37400
rect 68948 37360 70732 37400
rect 70772 37360 70781 37400
rect 71587 37360 71596 37400
rect 71636 37360 72364 37400
rect 72404 37360 72413 37400
rect 73411 37360 73420 37400
rect 73460 37360 74476 37400
rect 74516 37360 74525 37400
rect 57283 37276 57292 37316
rect 57332 37276 59500 37316
rect 59540 37276 59549 37316
rect 67555 37276 67564 37316
rect 67604 37276 69772 37316
rect 69812 37276 71020 37316
rect 71060 37276 71069 37316
rect 73795 37276 73804 37316
rect 73844 37276 74092 37316
rect 74132 37276 74141 37316
rect 74275 37276 74284 37316
rect 74324 37276 76588 37316
rect 76628 37276 79180 37316
rect 79220 37276 79229 37316
rect 57475 37192 57484 37232
rect 57524 37192 57964 37232
rect 58004 37192 59692 37232
rect 59732 37192 59741 37232
rect 64771 37192 64780 37232
rect 64820 37192 65452 37232
rect 65492 37192 65501 37232
rect 67747 37192 67756 37232
rect 67796 37192 69004 37232
rect 69044 37192 69053 37232
rect 70339 37192 70348 37232
rect 70388 37192 73036 37232
rect 73076 37192 73085 37232
rect 74755 37192 74764 37232
rect 74804 37192 74813 37232
rect 76099 37192 76108 37232
rect 76148 37192 76492 37232
rect 76532 37192 76541 37232
rect 66307 37148 66365 37149
rect 74764 37148 74804 37192
rect 76195 37148 76253 37149
rect 58819 37108 58828 37148
rect 58868 37108 60076 37148
rect 60116 37108 66316 37148
rect 66356 37108 70444 37148
rect 70484 37108 70493 37148
rect 73507 37108 73516 37148
rect 73556 37108 73996 37148
rect 74036 37108 74804 37148
rect 75331 37108 75340 37148
rect 75380 37108 76204 37148
rect 76244 37108 76253 37148
rect 66307 37107 66365 37108
rect 76195 37107 76253 37108
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 16343 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 16729 37064
rect 28343 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 28729 37064
rect 40343 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 40729 37064
rect 52343 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 52729 37064
rect 64343 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 64729 37064
rect 76343 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 76729 37064
rect 56899 36940 56908 36980
rect 56948 36940 57580 36980
rect 57620 36940 57629 36980
rect 72739 36940 72748 36980
rect 72788 36940 73460 36980
rect 73420 36896 73460 36940
rect 74179 36896 74237 36897
rect 59683 36856 59692 36896
rect 59732 36856 61228 36896
rect 61268 36856 61277 36896
rect 67363 36856 67372 36896
rect 67412 36856 68140 36896
rect 68180 36856 69868 36896
rect 69908 36856 69917 36896
rect 73420 36856 73708 36896
rect 73748 36856 73757 36896
rect 74094 36856 74188 36896
rect 74228 36856 74237 36896
rect 74563 36856 74572 36896
rect 74612 36856 77068 36896
rect 77108 36856 77117 36896
rect 74179 36855 74237 36856
rect 74572 36812 74612 36856
rect 56227 36772 56236 36812
rect 56276 36772 56716 36812
rect 56756 36772 56765 36812
rect 67075 36772 67084 36812
rect 67124 36772 68236 36812
rect 68276 36772 68285 36812
rect 71011 36772 71020 36812
rect 71060 36772 74612 36812
rect 0 36728 80 36748
rect 0 36688 36652 36728
rect 36692 36688 36701 36728
rect 56515 36688 56524 36728
rect 56564 36688 57484 36728
rect 57524 36688 58636 36728
rect 58676 36688 58685 36728
rect 60355 36688 60364 36728
rect 60404 36688 61228 36728
rect 61268 36688 61277 36728
rect 64291 36688 64300 36728
rect 64340 36688 64780 36728
rect 64820 36688 64829 36728
rect 67843 36688 67852 36728
rect 67892 36688 68812 36728
rect 68852 36688 68861 36728
rect 68995 36688 69004 36728
rect 69044 36688 69292 36728
rect 69332 36688 69341 36728
rect 70243 36688 70252 36728
rect 70292 36688 70732 36728
rect 70772 36688 71500 36728
rect 71540 36688 71549 36728
rect 72163 36688 72172 36728
rect 72212 36688 72748 36728
rect 72788 36688 72797 36728
rect 73027 36688 73036 36728
rect 73076 36688 73228 36728
rect 73268 36688 73277 36728
rect 75907 36688 75916 36728
rect 75956 36688 76684 36728
rect 76724 36688 76733 36728
rect 0 36668 80 36688
rect 59875 36604 59884 36644
rect 59924 36604 60652 36644
rect 60692 36604 60940 36644
rect 60980 36604 60989 36644
rect 70819 36604 70828 36644
rect 70868 36604 71116 36644
rect 71156 36604 71596 36644
rect 71636 36604 71645 36644
rect 73123 36604 73132 36644
rect 73172 36604 73612 36644
rect 73652 36604 74188 36644
rect 74228 36604 74237 36644
rect 75811 36604 75820 36644
rect 75860 36604 76204 36644
rect 76244 36604 77260 36644
rect 77300 36604 77309 36644
rect 74179 36560 74237 36561
rect 67171 36520 67180 36560
rect 67220 36520 68332 36560
rect 68372 36520 68381 36560
rect 71395 36520 71404 36560
rect 71444 36520 72940 36560
rect 72980 36520 72989 36560
rect 73507 36520 73516 36560
rect 73556 36520 74188 36560
rect 74228 36520 74764 36560
rect 74804 36520 77068 36560
rect 77108 36520 77117 36560
rect 74179 36519 74237 36520
rect 75619 36476 75677 36477
rect 59587 36436 59596 36476
rect 59636 36436 60940 36476
rect 60980 36436 61324 36476
rect 61364 36436 61373 36476
rect 74275 36436 74284 36476
rect 74324 36436 75436 36476
rect 75476 36436 75628 36476
rect 75668 36436 75677 36476
rect 75619 36435 75677 36436
rect 72451 36352 72460 36392
rect 72500 36352 72940 36392
rect 72980 36352 72989 36392
rect 56611 36308 56669 36309
rect 61699 36308 61757 36309
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 15103 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 15489 36308
rect 27103 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 27489 36308
rect 39103 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 39489 36308
rect 51103 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 51489 36308
rect 56526 36268 56620 36308
rect 56660 36268 57292 36308
rect 57332 36268 57341 36308
rect 61614 36268 61708 36308
rect 61748 36268 61757 36308
rect 63103 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 63489 36308
rect 75103 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 75489 36308
rect 56611 36267 56669 36268
rect 61699 36267 61757 36268
rect 55459 36184 55468 36224
rect 55508 36184 57100 36224
rect 57140 36184 57149 36224
rect 62179 36184 62188 36224
rect 62228 36184 63724 36224
rect 63764 36184 63773 36224
rect 64867 36184 64876 36224
rect 64916 36184 65164 36224
rect 65204 36184 65213 36224
rect 76483 36184 76492 36224
rect 76532 36184 77548 36224
rect 77588 36184 77597 36224
rect 56419 36100 56428 36140
rect 56468 36100 56477 36140
rect 64675 36100 64684 36140
rect 64724 36100 65068 36140
rect 65108 36100 66260 36140
rect 76387 36100 76396 36140
rect 76436 36100 77452 36140
rect 77492 36100 77501 36140
rect 56428 35972 56468 36100
rect 61219 36056 61277 36057
rect 66220 36056 66260 36100
rect 59011 36016 59020 36056
rect 59060 36016 59404 36056
rect 59444 36016 59453 36056
rect 61219 36016 61228 36056
rect 61268 36016 61420 36056
rect 61460 36016 61469 36056
rect 64291 36016 64300 36056
rect 64340 36016 65260 36056
rect 65300 36016 65309 36056
rect 66211 36016 66220 36056
rect 66260 36016 66796 36056
rect 66836 36016 66845 36056
rect 67651 36016 67660 36056
rect 67700 36016 69004 36056
rect 69044 36016 70252 36056
rect 70292 36016 70301 36056
rect 72643 36016 72652 36056
rect 72692 36016 73804 36056
rect 73844 36016 73853 36056
rect 74371 36016 74380 36056
rect 74420 36016 74429 36056
rect 76099 36016 76108 36056
rect 76148 36016 76820 36056
rect 61219 36015 61277 36016
rect 74380 35972 74420 36016
rect 76675 35972 76733 35973
rect 56035 35932 56044 35972
rect 56084 35932 56468 35972
rect 61027 35932 61036 35972
rect 61076 35932 61804 35972
rect 61844 35932 61853 35972
rect 62851 35932 62860 35972
rect 62900 35932 65644 35972
rect 65684 35932 65693 35972
rect 71587 35932 71596 35972
rect 71636 35932 72268 35972
rect 72308 35932 72844 35972
rect 72884 35932 72893 35972
rect 73891 35932 73900 35972
rect 73940 35932 74860 35972
rect 74900 35932 74909 35972
rect 76483 35932 76492 35972
rect 76532 35932 76684 35972
rect 76724 35932 76733 35972
rect 76675 35931 76733 35932
rect 0 35828 80 35908
rect 73795 35888 73853 35889
rect 76780 35888 76820 36016
rect 56707 35848 56716 35888
rect 56756 35848 57100 35888
rect 57140 35848 57149 35888
rect 57667 35848 57676 35888
rect 57716 35848 58444 35888
rect 58484 35848 58493 35888
rect 60835 35848 60844 35888
rect 60884 35848 61132 35888
rect 61172 35848 61324 35888
rect 61364 35848 61373 35888
rect 63340 35848 63820 35888
rect 63860 35848 63869 35888
rect 64003 35848 64012 35888
rect 64052 35848 64588 35888
rect 64628 35848 64876 35888
rect 64916 35848 64925 35888
rect 65443 35848 65452 35888
rect 65492 35848 65836 35888
rect 65876 35848 66604 35888
rect 66644 35848 66653 35888
rect 67843 35848 67852 35888
rect 67892 35848 68524 35888
rect 68564 35848 68573 35888
rect 69571 35848 69580 35888
rect 69620 35848 71308 35888
rect 71348 35848 72076 35888
rect 72116 35848 72125 35888
rect 73795 35848 73804 35888
rect 73844 35848 74668 35888
rect 74708 35848 74717 35888
rect 76771 35848 76780 35888
rect 76820 35848 76829 35888
rect 77731 35848 77740 35888
rect 77780 35848 78028 35888
rect 78068 35848 79468 35888
rect 79508 35848 79517 35888
rect 61699 35804 61757 35805
rect 63340 35804 63380 35848
rect 73795 35847 73853 35848
rect 56611 35764 56620 35804
rect 56660 35764 57772 35804
rect 57812 35764 57821 35804
rect 60259 35764 60268 35804
rect 60308 35764 61516 35804
rect 61556 35764 61565 35804
rect 61699 35764 61708 35804
rect 61748 35764 63380 35804
rect 66403 35764 66412 35804
rect 66452 35764 67276 35804
rect 67316 35764 67325 35804
rect 68611 35764 68620 35804
rect 68660 35764 68700 35804
rect 69091 35764 69100 35804
rect 69140 35764 73516 35804
rect 73556 35764 74284 35804
rect 74324 35764 74333 35804
rect 76387 35764 76396 35804
rect 76436 35764 77068 35804
rect 77108 35764 79084 35804
rect 79124 35764 79133 35804
rect 61699 35763 61757 35764
rect 61027 35720 61085 35721
rect 68620 35720 68660 35764
rect 57859 35680 57868 35720
rect 57908 35680 58252 35720
rect 58292 35680 58301 35720
rect 60942 35680 61036 35720
rect 61076 35680 61085 35720
rect 64963 35680 64972 35720
rect 65012 35680 65740 35720
rect 65780 35680 65789 35720
rect 68227 35680 68236 35720
rect 68276 35680 68812 35720
rect 68852 35680 68861 35720
rect 74083 35680 74092 35720
rect 74132 35680 74476 35720
rect 74516 35680 76300 35720
rect 76340 35680 76876 35720
rect 76916 35680 76925 35720
rect 61027 35679 61085 35680
rect 56611 35636 56669 35637
rect 56526 35596 56620 35636
rect 56660 35596 56669 35636
rect 56803 35596 56812 35636
rect 56852 35596 57388 35636
rect 57428 35596 57437 35636
rect 65539 35596 65548 35636
rect 65588 35596 67756 35636
rect 67796 35596 67805 35636
rect 74851 35596 74860 35636
rect 74900 35596 75628 35636
rect 75668 35596 76204 35636
rect 76244 35596 76253 35636
rect 56611 35595 56669 35596
rect 61219 35552 61277 35553
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 16343 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 16729 35552
rect 28343 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 28729 35552
rect 40343 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 40729 35552
rect 52343 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 52729 35552
rect 61134 35512 61228 35552
rect 61268 35512 61277 35552
rect 64343 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 64729 35552
rect 76343 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 76729 35552
rect 61219 35511 61277 35512
rect 61411 35428 61420 35468
rect 61460 35428 61612 35468
rect 61652 35428 62956 35468
rect 62996 35428 69772 35468
rect 69812 35428 69821 35468
rect 58723 35344 58732 35384
rect 58772 35344 59404 35384
rect 59444 35344 60172 35384
rect 60212 35344 60221 35384
rect 71683 35344 71692 35384
rect 71732 35344 73708 35384
rect 73748 35344 73757 35384
rect 73987 35344 73996 35384
rect 74036 35344 75052 35384
rect 75092 35344 75724 35384
rect 75764 35344 75773 35384
rect 76291 35344 76300 35384
rect 76340 35344 77644 35384
rect 77684 35344 77693 35384
rect 61027 35300 61085 35301
rect 55075 35260 55084 35300
rect 55124 35260 55948 35300
rect 55988 35260 55997 35300
rect 60259 35260 60268 35300
rect 60308 35260 61036 35300
rect 61076 35260 61085 35300
rect 72835 35260 72844 35300
rect 72884 35260 73324 35300
rect 73364 35260 73373 35300
rect 61027 35259 61085 35260
rect 73795 35216 73853 35217
rect 76867 35216 76925 35217
rect 59875 35176 59884 35216
rect 59924 35176 61900 35216
rect 61940 35176 62860 35216
rect 62900 35176 62909 35216
rect 71011 35176 71020 35216
rect 71060 35176 72076 35216
rect 72116 35176 72125 35216
rect 72172 35176 73132 35216
rect 73172 35176 73804 35216
rect 73844 35176 73853 35216
rect 76782 35176 76876 35216
rect 76916 35176 76925 35216
rect 77059 35176 77068 35216
rect 77108 35176 77260 35216
rect 77300 35176 77309 35216
rect 72172 35132 72212 35176
rect 73795 35175 73853 35176
rect 76867 35175 76925 35176
rect 76771 35132 76829 35133
rect 60931 35092 60940 35132
rect 60980 35092 61420 35132
rect 61460 35092 61469 35132
rect 61603 35092 61612 35132
rect 61652 35092 62476 35132
rect 62516 35092 62525 35132
rect 72163 35092 72172 35132
rect 72212 35092 72221 35132
rect 76771 35092 76780 35132
rect 76820 35092 78412 35132
rect 78452 35092 78461 35132
rect 0 34988 80 35068
rect 61027 35048 61085 35049
rect 60942 35008 61036 35048
rect 61076 35008 61085 35048
rect 61027 35007 61085 35008
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 15103 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 15489 34796
rect 27103 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 27489 34796
rect 39103 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 39489 34796
rect 51103 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 51489 34796
rect 61324 34712 61364 35092
rect 76771 35091 76829 35092
rect 65731 35008 65740 35048
rect 65780 35008 68236 35048
rect 68276 35008 68285 35048
rect 71491 35008 71500 35048
rect 71540 35008 71884 35048
rect 71924 35008 71933 35048
rect 76771 34964 76829 34965
rect 61411 34924 61420 34964
rect 61460 34924 62380 34964
rect 62420 34924 62429 34964
rect 63523 34924 63532 34964
rect 63572 34924 64012 34964
rect 64052 34924 64061 34964
rect 69091 34924 69100 34964
rect 69140 34924 70924 34964
rect 70964 34924 70973 34964
rect 75811 34924 75820 34964
rect 75860 34924 76780 34964
rect 76820 34924 76829 34964
rect 76771 34923 76829 34924
rect 72451 34840 72460 34880
rect 72500 34840 76300 34880
rect 76340 34840 76349 34880
rect 76867 34840 76876 34880
rect 76916 34840 77452 34880
rect 77492 34840 77501 34880
rect 63103 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 63489 34796
rect 75103 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 75489 34796
rect 61324 34672 61420 34712
rect 61460 34672 61469 34712
rect 61795 34672 61804 34712
rect 61844 34672 68332 34712
rect 68372 34672 68381 34712
rect 56131 34588 56140 34628
rect 56180 34588 57292 34628
rect 57332 34588 57341 34628
rect 68419 34588 68428 34628
rect 68468 34588 69100 34628
rect 69140 34588 69149 34628
rect 51715 34504 51724 34544
rect 51764 34504 52108 34544
rect 52148 34504 52157 34544
rect 55939 34504 55948 34544
rect 55988 34504 57196 34544
rect 57236 34504 57245 34544
rect 61795 34504 61804 34544
rect 61844 34504 62284 34544
rect 62324 34504 62333 34544
rect 62572 34504 64012 34544
rect 64052 34504 64061 34544
rect 67171 34504 67180 34544
rect 67220 34504 67604 34544
rect 68899 34504 68908 34544
rect 68948 34504 71308 34544
rect 71348 34504 71357 34544
rect 72739 34504 72748 34544
rect 72788 34504 73612 34544
rect 73652 34504 73661 34544
rect 77548 34504 78316 34544
rect 78356 34504 78365 34544
rect 62572 34460 62612 34504
rect 52195 34420 52204 34460
rect 52244 34420 53068 34460
rect 53108 34420 53117 34460
rect 59107 34420 59116 34460
rect 59156 34420 59308 34460
rect 59348 34420 60116 34460
rect 62563 34420 62572 34460
rect 62612 34420 62621 34460
rect 63619 34420 63628 34460
rect 63668 34420 64204 34460
rect 64244 34420 64780 34460
rect 64820 34420 64829 34460
rect 66979 34420 66988 34460
rect 67028 34420 67372 34460
rect 67412 34420 67421 34460
rect 50755 34336 50764 34376
rect 50804 34336 52300 34376
rect 52340 34336 52349 34376
rect 54115 34336 54124 34376
rect 54164 34336 55180 34376
rect 55220 34336 55229 34376
rect 55459 34336 55468 34376
rect 55508 34336 55517 34376
rect 56035 34336 56044 34376
rect 56084 34336 58060 34376
rect 58100 34336 58109 34376
rect 58627 34336 58636 34376
rect 58676 34336 60020 34376
rect 0 34148 80 34228
rect 55468 34124 55508 34336
rect 56131 34252 56140 34292
rect 56180 34252 56812 34292
rect 56852 34252 56861 34292
rect 59980 34208 60020 34336
rect 60076 34292 60116 34420
rect 67564 34376 67604 34504
rect 77548 34376 77588 34504
rect 62659 34336 62668 34376
rect 62708 34336 63532 34376
rect 63572 34336 63581 34376
rect 64675 34336 64684 34376
rect 64724 34336 65164 34376
rect 65204 34336 65213 34376
rect 67555 34336 67564 34376
rect 67604 34336 67613 34376
rect 67939 34336 67948 34376
rect 67988 34336 68620 34376
rect 68660 34336 68669 34376
rect 68803 34336 68812 34376
rect 68852 34336 69676 34376
rect 69716 34336 70156 34376
rect 70196 34336 70205 34376
rect 71395 34336 71404 34376
rect 71444 34336 71788 34376
rect 71828 34336 71837 34376
rect 72067 34336 72076 34376
rect 72116 34336 72652 34376
rect 72692 34336 72701 34376
rect 73603 34336 73612 34376
rect 73652 34336 74092 34376
rect 74132 34336 74572 34376
rect 74612 34336 76108 34376
rect 76148 34336 77548 34376
rect 77588 34336 77597 34376
rect 77827 34336 77836 34376
rect 77876 34336 78508 34376
rect 78548 34336 78557 34376
rect 64684 34292 64724 34336
rect 77347 34292 77405 34293
rect 60076 34252 64724 34292
rect 65347 34252 65356 34292
rect 65396 34252 66796 34292
rect 66836 34252 66845 34292
rect 67459 34252 67468 34292
rect 67508 34252 68140 34292
rect 68180 34252 68189 34292
rect 71875 34252 71884 34292
rect 71924 34252 72364 34292
rect 72404 34252 72413 34292
rect 77347 34252 77356 34292
rect 77396 34252 78316 34292
rect 78356 34252 78365 34292
rect 66796 34208 66836 34252
rect 77347 34251 77405 34252
rect 57283 34168 57292 34208
rect 57332 34168 59692 34208
rect 59732 34168 59741 34208
rect 59971 34168 59980 34208
rect 60020 34168 60029 34208
rect 61315 34168 61324 34208
rect 61364 34168 62092 34208
rect 62132 34168 62141 34208
rect 66796 34168 69868 34208
rect 69908 34168 69917 34208
rect 61324 34124 61364 34168
rect 77923 34124 77981 34125
rect 54307 34084 54316 34124
rect 54356 34084 56044 34124
rect 56084 34084 56093 34124
rect 59875 34084 59884 34124
rect 59924 34084 61364 34124
rect 68803 34084 68812 34124
rect 68852 34084 72172 34124
rect 72212 34084 72221 34124
rect 77838 34084 77932 34124
rect 77972 34084 78220 34124
rect 78260 34084 78269 34124
rect 77923 34083 77981 34084
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 16343 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 16729 34040
rect 28343 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 28729 34040
rect 40343 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 40729 34040
rect 52343 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 52729 34040
rect 57187 34000 57196 34040
rect 57236 34000 57484 34040
rect 57524 34000 60460 34040
rect 60500 34000 60509 34040
rect 64343 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 64729 34040
rect 67747 34000 67756 34040
rect 67796 34000 68140 34040
rect 68180 34000 68189 34040
rect 76343 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 76729 34040
rect 77059 34000 77068 34040
rect 77108 34000 78028 34040
rect 78068 34000 78077 34040
rect 59395 33916 59404 33956
rect 59444 33916 60652 33956
rect 60692 33916 63628 33956
rect 63668 33916 63677 33956
rect 76195 33916 76204 33956
rect 76244 33916 76628 33956
rect 76867 33916 76876 33956
rect 76916 33916 77356 33956
rect 77396 33916 77405 33956
rect 76588 33872 76628 33916
rect 50851 33832 50860 33872
rect 50900 33832 51340 33872
rect 51380 33832 52972 33872
rect 53012 33832 54316 33872
rect 54356 33832 54365 33872
rect 55075 33832 55084 33872
rect 55124 33832 55468 33872
rect 55508 33832 55517 33872
rect 61123 33832 61132 33872
rect 61172 33832 61996 33872
rect 62036 33832 63244 33872
rect 63284 33832 63293 33872
rect 63715 33832 63724 33872
rect 63764 33832 64492 33872
rect 64532 33832 64541 33872
rect 71299 33832 71308 33872
rect 71348 33832 72076 33872
rect 72116 33832 72460 33872
rect 72500 33832 72509 33872
rect 74947 33832 74956 33872
rect 74996 33832 76300 33872
rect 76340 33832 76349 33872
rect 76579 33832 76588 33872
rect 76628 33832 76637 33872
rect 76771 33832 76780 33872
rect 76820 33832 77164 33872
rect 77204 33832 77452 33872
rect 77492 33832 77501 33872
rect 59587 33748 59596 33788
rect 59636 33748 61324 33788
rect 61364 33748 61516 33788
rect 61556 33748 61565 33788
rect 64291 33748 64300 33788
rect 64340 33748 65068 33788
rect 65108 33748 65117 33788
rect 67459 33748 67468 33788
rect 67508 33748 67852 33788
rect 67892 33748 67901 33788
rect 77155 33704 77213 33705
rect 50467 33664 50476 33704
rect 50516 33664 52108 33704
rect 52148 33664 53452 33704
rect 53492 33664 53836 33704
rect 53876 33664 55756 33704
rect 55796 33664 56428 33704
rect 56468 33664 56908 33704
rect 56948 33664 56957 33704
rect 59491 33664 59500 33704
rect 59540 33664 59884 33704
rect 59924 33664 59933 33704
rect 64675 33664 64684 33704
rect 64724 33664 66700 33704
rect 66740 33664 66749 33704
rect 67075 33664 67084 33704
rect 67124 33664 67756 33704
rect 67796 33664 67805 33704
rect 71971 33664 71980 33704
rect 72020 33664 72556 33704
rect 72596 33664 74572 33704
rect 74612 33664 74621 33704
rect 76387 33664 76396 33704
rect 76436 33664 76684 33704
rect 76724 33664 77164 33704
rect 77204 33664 77213 33704
rect 77443 33664 77452 33704
rect 77492 33664 77644 33704
rect 77684 33664 77693 33704
rect 78211 33664 78220 33704
rect 78260 33664 78796 33704
rect 78836 33664 78845 33704
rect 77155 33663 77213 33664
rect 55459 33580 55468 33620
rect 55508 33580 58348 33620
rect 58388 33580 58397 33620
rect 59011 33580 59020 33620
rect 59060 33580 64300 33620
rect 64340 33580 64349 33620
rect 64579 33580 64588 33620
rect 64628 33580 65356 33620
rect 65396 33580 65405 33620
rect 66883 33580 66892 33620
rect 66932 33580 69580 33620
rect 69620 33580 69629 33620
rect 50476 33496 51916 33536
rect 51956 33496 51965 33536
rect 59395 33496 59404 33536
rect 59444 33496 60844 33536
rect 60884 33496 61612 33536
rect 61652 33496 61661 33536
rect 63907 33496 63916 33536
rect 63956 33496 64780 33536
rect 64820 33496 64829 33536
rect 66787 33496 66796 33536
rect 66836 33496 67372 33536
rect 67412 33496 67421 33536
rect 77347 33496 77356 33536
rect 77396 33496 77644 33536
rect 77684 33496 77693 33536
rect 50476 33452 50516 33496
rect 77347 33452 77405 33453
rect 49315 33412 49324 33452
rect 49364 33412 50476 33452
rect 50516 33412 50525 33452
rect 51523 33412 51532 33452
rect 51572 33412 52012 33452
rect 52052 33412 52061 33452
rect 52291 33412 52300 33452
rect 52340 33412 54124 33452
rect 54164 33412 54173 33452
rect 54787 33412 54796 33452
rect 54836 33412 55276 33452
rect 55316 33412 55325 33452
rect 61699 33412 61708 33452
rect 61748 33412 61996 33452
rect 62036 33412 62045 33452
rect 63235 33412 63244 33452
rect 63284 33412 64916 33452
rect 72643 33412 72652 33452
rect 72692 33412 72701 33452
rect 73027 33412 73036 33452
rect 73076 33412 74860 33452
rect 74900 33412 75724 33452
rect 75764 33412 75773 33452
rect 76291 33412 76300 33452
rect 76340 33412 77356 33452
rect 77396 33412 77405 33452
rect 0 33308 80 33388
rect 61219 33368 61277 33369
rect 54595 33328 54604 33368
rect 54644 33328 55660 33368
rect 55700 33328 55709 33368
rect 61219 33328 61228 33368
rect 61268 33328 61804 33368
rect 61844 33328 61853 33368
rect 64003 33328 64012 33368
rect 64052 33328 64588 33368
rect 64628 33328 64637 33368
rect 61219 33327 61277 33328
rect 55363 33284 55421 33285
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 15103 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 15489 33284
rect 27103 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 27489 33284
rect 39103 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 39489 33284
rect 51103 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 51489 33284
rect 55278 33244 55372 33284
rect 55412 33244 55421 33284
rect 63103 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 63489 33284
rect 55363 33243 55421 33244
rect 64876 33200 64916 33412
rect 72652 33368 72692 33412
rect 77347 33411 77405 33412
rect 72652 33328 73996 33368
rect 74036 33328 74045 33368
rect 68419 33244 68428 33284
rect 68468 33244 68716 33284
rect 68756 33244 71884 33284
rect 71924 33244 73036 33284
rect 73076 33244 73085 33284
rect 75103 33244 75112 33284
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75480 33244 75489 33284
rect 54508 33160 54700 33200
rect 54740 33160 54749 33200
rect 61315 33160 61324 33200
rect 61364 33160 61940 33200
rect 64867 33160 64876 33200
rect 64916 33160 67468 33200
rect 67508 33160 67517 33200
rect 54508 33116 54548 33160
rect 50947 33076 50956 33116
rect 50996 33076 52204 33116
rect 52244 33076 53012 33116
rect 53059 33076 53068 33116
rect 53108 33076 53836 33116
rect 53876 33076 53885 33116
rect 54403 33076 54412 33116
rect 54452 33076 54548 33116
rect 61900 33116 61940 33160
rect 61900 33076 63148 33116
rect 63188 33076 63197 33116
rect 52972 33032 53012 33076
rect 72835 33032 72893 33033
rect 52963 32992 52972 33032
rect 53012 32992 53021 33032
rect 55363 32992 55372 33032
rect 55412 32992 55852 33032
rect 55892 32992 55901 33032
rect 72750 32992 72844 33032
rect 72884 32992 72893 33032
rect 72835 32991 72893 32992
rect 51331 32908 51340 32948
rect 51380 32908 51532 32948
rect 51572 32908 53644 32948
rect 53684 32908 53693 32948
rect 54019 32908 54028 32948
rect 54068 32908 56084 32948
rect 65827 32908 65836 32948
rect 65876 32908 66220 32948
rect 66260 32908 66269 32948
rect 56044 32864 56084 32908
rect 51235 32824 51244 32864
rect 51284 32824 53356 32864
rect 53396 32824 53405 32864
rect 53539 32824 53548 32864
rect 53588 32824 54412 32864
rect 54452 32824 54461 32864
rect 54691 32824 54700 32864
rect 54740 32824 54988 32864
rect 55028 32824 55180 32864
rect 55220 32824 55229 32864
rect 56035 32824 56044 32864
rect 56084 32824 57868 32864
rect 57908 32824 58828 32864
rect 58868 32824 58877 32864
rect 65635 32824 65644 32864
rect 65684 32824 66700 32864
rect 66740 32824 66749 32864
rect 67555 32824 67564 32864
rect 67604 32824 68140 32864
rect 68180 32824 68189 32864
rect 70147 32824 70156 32864
rect 70196 32824 70828 32864
rect 70868 32824 70877 32864
rect 71011 32824 71020 32864
rect 71060 32824 74092 32864
rect 74132 32824 74141 32864
rect 76771 32824 76780 32864
rect 76820 32824 76972 32864
rect 77012 32824 77356 32864
rect 77396 32824 77405 32864
rect 77635 32824 77644 32864
rect 77684 32824 78220 32864
rect 78260 32824 78269 32864
rect 72355 32780 72413 32781
rect 53155 32740 53164 32780
rect 53204 32740 53452 32780
rect 53492 32740 53501 32780
rect 55843 32740 55852 32780
rect 55892 32740 56428 32780
rect 56468 32740 57676 32780
rect 57716 32740 57725 32780
rect 62755 32740 62764 32780
rect 62804 32740 62813 32780
rect 69763 32740 69772 32780
rect 69812 32740 71692 32780
rect 71732 32740 71741 32780
rect 72270 32740 72364 32780
rect 72404 32740 72413 32780
rect 55363 32696 55421 32697
rect 62764 32696 62804 32740
rect 72355 32739 72413 32740
rect 49795 32656 49804 32696
rect 49844 32656 50860 32696
rect 50900 32656 50909 32696
rect 53635 32656 53644 32696
rect 53684 32656 55084 32696
rect 55124 32656 55372 32696
rect 55412 32656 55421 32696
rect 60163 32656 60172 32696
rect 60212 32656 61804 32696
rect 61844 32656 62804 32696
rect 62851 32656 62860 32696
rect 62900 32656 63052 32696
rect 63092 32656 63101 32696
rect 66787 32656 66796 32696
rect 66836 32656 67660 32696
rect 67700 32656 68140 32696
rect 68180 32656 68189 32696
rect 55363 32655 55421 32656
rect 50563 32572 50572 32612
rect 50612 32572 52012 32612
rect 52052 32572 54028 32612
rect 54068 32572 54077 32612
rect 71875 32572 71884 32612
rect 71924 32572 72364 32612
rect 72404 32572 72652 32612
rect 72692 32572 72701 32612
rect 0 32468 80 32548
rect 73603 32528 73661 32529
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 16343 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 16729 32528
rect 28343 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 28729 32528
rect 40343 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 40729 32528
rect 52343 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 52729 32528
rect 53443 32488 53452 32528
rect 53492 32488 57100 32528
rect 57140 32488 58156 32528
rect 58196 32488 58205 32528
rect 64343 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 64729 32528
rect 72547 32488 72556 32528
rect 72596 32488 73612 32528
rect 73652 32488 73661 32528
rect 76343 32488 76352 32528
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76720 32488 76729 32528
rect 73603 32487 73661 32488
rect 53347 32404 53356 32444
rect 53396 32404 54604 32444
rect 54644 32404 66508 32444
rect 66548 32404 66557 32444
rect 76771 32404 76780 32444
rect 76820 32404 78124 32444
rect 78164 32404 78173 32444
rect 76780 32360 76820 32404
rect 60451 32320 60460 32360
rect 60500 32320 66068 32360
rect 76483 32320 76492 32360
rect 76532 32320 76820 32360
rect 64204 32236 65836 32276
rect 65876 32236 65885 32276
rect 63523 32192 63581 32193
rect 64204 32192 64244 32236
rect 52771 32152 52780 32192
rect 52820 32152 53356 32192
rect 53396 32152 53405 32192
rect 57667 32152 57676 32192
rect 57716 32152 58540 32192
rect 58580 32152 58589 32192
rect 60163 32152 60172 32192
rect 60212 32152 60940 32192
rect 60980 32152 60989 32192
rect 61507 32152 61516 32192
rect 61556 32152 62764 32192
rect 62804 32152 62813 32192
rect 63331 32152 63340 32192
rect 63380 32152 63532 32192
rect 63572 32152 63581 32192
rect 63715 32152 63724 32192
rect 63764 32152 64204 32192
rect 64244 32152 64253 32192
rect 64579 32152 64588 32192
rect 64628 32152 65644 32192
rect 65684 32152 65693 32192
rect 61516 32108 61556 32152
rect 63523 32151 63581 32152
rect 66028 32108 66068 32320
rect 77923 32276 77981 32277
rect 66595 32236 66604 32276
rect 66644 32236 67660 32276
rect 67700 32236 67709 32276
rect 76675 32236 76684 32276
rect 76724 32236 77932 32276
rect 77972 32236 77981 32276
rect 77923 32235 77981 32236
rect 66115 32152 66124 32192
rect 66164 32152 66412 32192
rect 66452 32152 67276 32192
rect 67316 32152 67325 32192
rect 71491 32152 71500 32192
rect 71540 32152 72076 32192
rect 72116 32152 72125 32192
rect 75907 32152 75916 32192
rect 75956 32152 76972 32192
rect 77012 32152 77021 32192
rect 72835 32108 72893 32109
rect 57283 32068 57292 32108
rect 57332 32068 57341 32108
rect 57475 32068 57484 32108
rect 57524 32068 58636 32108
rect 58676 32068 58685 32108
rect 59299 32068 59308 32108
rect 59348 32068 61132 32108
rect 61172 32068 61556 32108
rect 63043 32068 63052 32108
rect 63092 32068 63532 32108
rect 63572 32068 63581 32108
rect 66028 32068 67892 32108
rect 71779 32068 71788 32108
rect 71828 32068 72844 32108
rect 72884 32068 72893 32108
rect 57292 32024 57332 32068
rect 57292 31984 57868 32024
rect 57908 31984 57917 32024
rect 61027 31984 61036 32024
rect 61076 31984 61516 32024
rect 61556 31984 61565 32024
rect 65443 31984 65452 32024
rect 65492 31984 66604 32024
rect 66644 31984 66653 32024
rect 66787 31984 66796 32024
rect 66836 31984 67180 32024
rect 67220 31984 67229 32024
rect 67852 31940 67892 32068
rect 72835 32067 72893 32068
rect 57763 31900 57772 31940
rect 57812 31900 58924 31940
rect 58964 31900 60364 31940
rect 60404 31900 60413 31940
rect 63427 31900 63436 31940
rect 63476 31900 63724 31940
rect 63764 31900 63773 31940
rect 63916 31900 67756 31940
rect 67796 31900 67805 31940
rect 67852 31900 69812 31940
rect 78115 31900 78124 31940
rect 78164 31900 79372 31940
rect 79412 31900 79421 31940
rect 56419 31856 56477 31857
rect 63916 31856 63956 31900
rect 69772 31856 69812 31900
rect 54787 31816 54796 31856
rect 54836 31816 56428 31856
rect 56468 31816 56477 31856
rect 60451 31816 60460 31856
rect 60500 31816 60748 31856
rect 60788 31816 61036 31856
rect 61076 31816 61085 31856
rect 61132 31816 63956 31856
rect 64003 31816 64012 31856
rect 64052 31816 66892 31856
rect 66932 31816 67564 31856
rect 67604 31816 68140 31856
rect 68180 31816 68189 31856
rect 69763 31816 69772 31856
rect 69812 31816 69821 31856
rect 56419 31815 56477 31816
rect 53059 31772 53117 31773
rect 61132 31772 61172 31816
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 15103 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 15489 31772
rect 27103 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 27489 31772
rect 39103 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 39489 31772
rect 51103 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 51489 31772
rect 52974 31732 53068 31772
rect 53108 31732 53117 31772
rect 54499 31732 54508 31772
rect 54548 31732 56140 31772
rect 56180 31732 57100 31772
rect 57140 31732 57149 31772
rect 59779 31732 59788 31772
rect 59828 31732 59837 31772
rect 59971 31732 59980 31772
rect 60020 31732 61172 31772
rect 63103 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 63489 31772
rect 65347 31732 65356 31772
rect 65396 31732 66124 31772
rect 66164 31732 66173 31772
rect 67459 31732 67468 31772
rect 67508 31732 68428 31772
rect 68468 31732 68477 31772
rect 75103 31732 75112 31772
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75480 31732 75489 31772
rect 53059 31731 53117 31732
rect 0 31628 80 31708
rect 59788 31688 59828 31732
rect 72835 31688 72893 31689
rect 58435 31648 58444 31688
rect 58484 31648 59828 31688
rect 60547 31648 60556 31688
rect 60596 31648 61324 31688
rect 61364 31648 61373 31688
rect 72750 31648 72844 31688
rect 72884 31648 72893 31688
rect 73987 31648 73996 31688
rect 74036 31648 74188 31688
rect 74228 31648 74237 31688
rect 76579 31648 76588 31688
rect 76628 31648 77548 31688
rect 77588 31648 77597 31688
rect 72835 31647 72893 31648
rect 50179 31564 50188 31604
rect 50228 31564 51340 31604
rect 51380 31564 51389 31604
rect 51907 31564 51916 31604
rect 51956 31564 52396 31604
rect 52436 31564 52445 31604
rect 62083 31564 62092 31604
rect 62132 31564 68236 31604
rect 68276 31564 68285 31604
rect 71299 31564 71308 31604
rect 71348 31564 71596 31604
rect 71636 31564 72268 31604
rect 72308 31564 77260 31604
rect 77300 31564 77836 31604
rect 77876 31564 77885 31604
rect 62659 31520 62717 31521
rect 73315 31520 73373 31521
rect 50467 31480 50476 31520
rect 50516 31480 50956 31520
rect 50996 31480 51005 31520
rect 52483 31480 52492 31520
rect 52532 31480 53644 31520
rect 53684 31480 53693 31520
rect 61123 31480 61132 31520
rect 61172 31480 61516 31520
rect 61556 31480 61565 31520
rect 61699 31480 61708 31520
rect 61748 31480 62668 31520
rect 62708 31480 62717 31520
rect 71395 31480 71404 31520
rect 71444 31480 73324 31520
rect 73364 31480 74380 31520
rect 74420 31480 74429 31520
rect 76291 31480 76300 31520
rect 76340 31480 76588 31520
rect 76628 31480 76637 31520
rect 62659 31479 62717 31480
rect 73315 31479 73373 31480
rect 63523 31436 63581 31437
rect 52579 31396 52588 31436
rect 52628 31396 53932 31436
rect 53972 31396 53981 31436
rect 57484 31396 58348 31436
rect 58388 31396 58397 31436
rect 61219 31396 61228 31436
rect 61268 31396 61420 31436
rect 61460 31396 61804 31436
rect 61844 31396 61853 31436
rect 63235 31396 63244 31436
rect 63284 31396 63532 31436
rect 63572 31396 63581 31436
rect 72547 31396 72556 31436
rect 72596 31396 73036 31436
rect 73076 31396 73085 31436
rect 73699 31396 73708 31436
rect 73748 31396 76052 31436
rect 76099 31396 76108 31436
rect 76148 31396 78028 31436
rect 78068 31396 78077 31436
rect 57484 31352 57524 31396
rect 63523 31395 63581 31396
rect 61123 31352 61181 31353
rect 63907 31352 63965 31353
rect 73603 31352 73661 31353
rect 76012 31352 76052 31396
rect 77251 31352 77309 31353
rect 50371 31312 50380 31352
rect 50420 31312 51436 31352
rect 51476 31312 51485 31352
rect 51811 31312 51820 31352
rect 51860 31312 51869 31352
rect 52675 31312 52684 31352
rect 52724 31312 54124 31352
rect 54164 31312 55276 31352
rect 55316 31312 55325 31352
rect 56803 31312 56812 31352
rect 56852 31312 57484 31352
rect 57524 31312 57533 31352
rect 57667 31312 57676 31352
rect 57716 31312 58060 31352
rect 58100 31312 58109 31352
rect 58243 31312 58252 31352
rect 58292 31312 59212 31352
rect 59252 31312 59261 31352
rect 61123 31312 61132 31352
rect 61172 31312 61612 31352
rect 61652 31312 63532 31352
rect 63572 31312 63581 31352
rect 63822 31312 63916 31352
rect 63956 31312 65740 31352
rect 65780 31312 65789 31352
rect 67267 31312 67276 31352
rect 67316 31312 67325 31352
rect 67939 31312 67948 31352
rect 67988 31312 70156 31352
rect 70196 31312 70205 31352
rect 72451 31312 72460 31352
rect 72500 31312 73460 31352
rect 51820 31268 51860 31312
rect 61123 31311 61181 31312
rect 63907 31311 63965 31312
rect 67276 31268 67316 31312
rect 73420 31268 73460 31312
rect 73603 31312 73612 31352
rect 73652 31312 73746 31352
rect 73804 31312 74476 31352
rect 74516 31312 74956 31352
rect 74996 31312 75005 31352
rect 76003 31312 76012 31352
rect 76052 31312 77260 31352
rect 77300 31312 77644 31352
rect 77684 31312 78412 31352
rect 78452 31312 78461 31352
rect 73603 31311 73661 31312
rect 73804 31268 73844 31312
rect 77251 31311 77309 31312
rect 50755 31228 50764 31268
rect 50804 31228 50956 31268
rect 50996 31228 52300 31268
rect 52340 31228 53836 31268
rect 53876 31228 53885 31268
rect 67276 31228 69100 31268
rect 69140 31228 69149 31268
rect 73420 31228 73516 31268
rect 73556 31228 73565 31268
rect 73795 31228 73804 31268
rect 73844 31228 73853 31268
rect 77731 31228 77740 31268
rect 77780 31228 78124 31268
rect 78164 31228 78173 31268
rect 51820 31144 52012 31184
rect 52052 31144 52061 31184
rect 57475 31144 57484 31184
rect 57524 31144 59116 31184
rect 59156 31144 65836 31184
rect 65876 31144 65885 31184
rect 67075 31144 67084 31184
rect 67124 31144 67468 31184
rect 67508 31144 67517 31184
rect 68227 31144 68236 31184
rect 68276 31144 68524 31184
rect 68564 31144 68573 31184
rect 72259 31144 72268 31184
rect 72308 31144 72460 31184
rect 72500 31144 72509 31184
rect 72931 31144 72940 31184
rect 72980 31144 74380 31184
rect 74420 31144 74429 31184
rect 51820 31100 51860 31144
rect 51811 31060 51820 31100
rect 51860 31060 51869 31100
rect 68611 31060 68620 31100
rect 68660 31060 69004 31100
rect 69044 31060 69053 31100
rect 77251 31060 77260 31100
rect 77300 31060 77452 31100
rect 77492 31060 77501 31100
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 16343 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 16729 31016
rect 28343 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 28729 31016
rect 40343 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 40729 31016
rect 51427 30976 51436 31016
rect 51476 30976 52012 31016
rect 52052 30976 52061 31016
rect 52343 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 52729 31016
rect 64343 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 64729 31016
rect 73411 30976 73420 31016
rect 73460 30976 73900 31016
rect 73940 30976 73949 31016
rect 76343 30976 76352 31016
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76720 30976 76729 31016
rect 0 30788 80 30868
rect 55363 30808 55372 30848
rect 55412 30808 56044 30848
rect 56084 30808 56093 30848
rect 66403 30724 66412 30764
rect 66452 30724 67084 30764
rect 67124 30724 67133 30764
rect 50179 30640 50188 30680
rect 50228 30640 50668 30680
rect 50708 30640 50717 30680
rect 54883 30640 54892 30680
rect 54932 30640 55660 30680
rect 55700 30640 57772 30680
rect 57812 30640 59116 30680
rect 59156 30640 60556 30680
rect 60596 30640 62572 30680
rect 62612 30640 62621 30680
rect 66691 30640 66700 30680
rect 66740 30640 66988 30680
rect 67028 30640 67372 30680
rect 67412 30640 67421 30680
rect 68227 30640 68236 30680
rect 68276 30640 69004 30680
rect 69044 30640 69964 30680
rect 70004 30640 70013 30680
rect 70147 30640 70156 30680
rect 70196 30640 70540 30680
rect 70580 30640 71308 30680
rect 71348 30640 71357 30680
rect 71683 30640 71692 30680
rect 71732 30640 72076 30680
rect 72116 30640 72125 30680
rect 72835 30640 72844 30680
rect 72884 30640 75436 30680
rect 75476 30640 75485 30680
rect 76291 30640 76300 30680
rect 76340 30640 78220 30680
rect 78260 30640 78269 30680
rect 61123 30596 61181 30597
rect 75436 30596 75476 30640
rect 53827 30556 53836 30596
rect 53876 30556 56236 30596
rect 56276 30556 56285 30596
rect 61038 30556 61132 30596
rect 61172 30556 61612 30596
rect 61652 30556 61661 30596
rect 71971 30556 71980 30596
rect 72020 30556 72460 30596
rect 72500 30556 72509 30596
rect 73699 30556 73708 30596
rect 73748 30556 73996 30596
rect 74036 30556 74045 30596
rect 75436 30556 77260 30596
rect 77300 30556 77452 30596
rect 77492 30556 77501 30596
rect 61123 30555 61181 30556
rect 64003 30512 64061 30513
rect 63427 30472 63436 30512
rect 63476 30472 64012 30512
rect 64052 30472 64061 30512
rect 71299 30472 71308 30512
rect 71348 30472 71596 30512
rect 71636 30472 71645 30512
rect 73507 30472 73516 30512
rect 73556 30472 74092 30512
rect 74132 30472 74141 30512
rect 75043 30472 75052 30512
rect 75092 30472 76012 30512
rect 76052 30472 76061 30512
rect 64003 30471 64061 30472
rect 62659 30428 62717 30429
rect 72355 30428 72413 30429
rect 60931 30388 60940 30428
rect 60980 30388 61420 30428
rect 61460 30388 61469 30428
rect 62659 30388 62668 30428
rect 62708 30388 63724 30428
rect 63764 30388 63773 30428
rect 69283 30388 69292 30428
rect 69332 30388 71404 30428
rect 71444 30388 71788 30428
rect 71828 30388 71837 30428
rect 72270 30388 72364 30428
rect 72404 30388 72413 30428
rect 75523 30388 75532 30428
rect 75572 30388 75724 30428
rect 75764 30388 75773 30428
rect 62659 30387 62717 30388
rect 72355 30387 72413 30388
rect 51811 30344 51869 30345
rect 50371 30304 50380 30344
rect 50420 30304 51820 30344
rect 51860 30304 51869 30344
rect 54019 30304 54028 30344
rect 54068 30304 56524 30344
rect 56564 30304 57004 30344
rect 57044 30304 58252 30344
rect 58292 30304 58301 30344
rect 59203 30304 59212 30344
rect 59252 30304 60268 30344
rect 60308 30304 65740 30344
rect 65780 30304 65789 30344
rect 69955 30304 69964 30344
rect 70004 30304 71692 30344
rect 71732 30304 71741 30344
rect 51811 30303 51869 30304
rect 61219 30260 61277 30261
rect 73795 30260 73853 30261
rect 74947 30260 75005 30261
rect 77251 30260 77309 30261
rect 78019 30260 78077 30261
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 15103 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 15489 30260
rect 27103 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 27489 30260
rect 39103 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 39489 30260
rect 46627 30220 46636 30260
rect 46676 30220 47980 30260
rect 48020 30220 48029 30260
rect 48163 30220 48172 30260
rect 48212 30220 50956 30260
rect 50996 30220 51005 30260
rect 51103 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 51489 30260
rect 53347 30220 53356 30260
rect 53396 30220 53932 30260
rect 53972 30220 53981 30260
rect 61134 30220 61228 30260
rect 61268 30220 61277 30260
rect 63103 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 63489 30260
rect 64003 30220 64012 30260
rect 64052 30220 65452 30260
rect 65492 30220 65501 30260
rect 71107 30220 71116 30260
rect 71156 30220 71788 30260
rect 71828 30220 72268 30260
rect 72308 30220 72317 30260
rect 72643 30220 72652 30260
rect 72692 30220 73228 30260
rect 73268 30220 73277 30260
rect 73710 30220 73804 30260
rect 73844 30220 73853 30260
rect 74862 30220 74956 30260
rect 74996 30220 75005 30260
rect 75103 30220 75112 30260
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75480 30220 75489 30260
rect 77166 30220 77260 30260
rect 77300 30220 77309 30260
rect 77934 30220 78028 30260
rect 78068 30220 78077 30260
rect 61219 30219 61277 30220
rect 73795 30219 73853 30220
rect 74947 30219 75005 30220
rect 77251 30219 77309 30220
rect 78019 30219 78077 30220
rect 54211 30136 54220 30176
rect 54260 30136 54604 30176
rect 54644 30136 54653 30176
rect 64867 30136 64876 30176
rect 64916 30136 66316 30176
rect 66356 30136 66365 30176
rect 54691 30052 54700 30092
rect 54740 30052 55468 30092
rect 55508 30052 56140 30092
rect 56180 30052 57580 30092
rect 57620 30052 57629 30092
rect 59395 30052 59404 30092
rect 59444 30052 59596 30092
rect 59636 30052 62476 30092
rect 62516 30052 62525 30092
rect 63523 30052 63532 30092
rect 63572 30052 64396 30092
rect 64436 30052 67084 30092
rect 67124 30052 67133 30092
rect 70915 30052 70924 30092
rect 70964 30052 71500 30092
rect 71540 30052 71549 30092
rect 73219 30052 73228 30092
rect 73268 30052 73612 30092
rect 73652 30052 73661 30092
rect 0 29948 80 30028
rect 40579 29968 40588 30008
rect 40628 29968 60172 30008
rect 60212 29968 60221 30008
rect 61891 29968 61900 30008
rect 61940 29968 61949 30008
rect 65059 29968 65068 30008
rect 65108 29968 65356 30008
rect 65396 29968 65405 30008
rect 72067 29968 72076 30008
rect 72116 29968 72268 30008
rect 72308 29968 72748 30008
rect 72788 29968 72797 30008
rect 75619 29968 75628 30008
rect 75668 29968 75820 30008
rect 75860 29968 76876 30008
rect 76916 29968 76925 30008
rect 53155 29924 53213 29925
rect 61900 29924 61940 29968
rect 29731 29884 29740 29924
rect 29780 29884 40396 29924
rect 40436 29884 40445 29924
rect 51619 29884 51628 29924
rect 51668 29884 53068 29924
rect 53108 29884 53164 29924
rect 53204 29884 53232 29924
rect 60739 29884 60748 29924
rect 60788 29884 61940 29924
rect 65251 29884 65260 29924
rect 65300 29884 65340 29924
rect 65539 29884 65548 29924
rect 65588 29884 65932 29924
rect 65972 29884 65981 29924
rect 66307 29884 66316 29924
rect 66356 29884 66892 29924
rect 66932 29884 66941 29924
rect 73411 29884 73420 29924
rect 73460 29884 76780 29924
rect 76820 29884 77836 29924
rect 77876 29884 77885 29924
rect 53155 29883 53213 29884
rect 65260 29840 65300 29884
rect 47395 29800 47404 29840
rect 47444 29800 48748 29840
rect 48788 29800 49516 29840
rect 49556 29800 49900 29840
rect 49940 29800 49949 29840
rect 51523 29800 51532 29840
rect 51572 29800 53164 29840
rect 53204 29800 53213 29840
rect 54307 29800 54316 29840
rect 54356 29800 54892 29840
rect 54932 29800 54941 29840
rect 65059 29800 65068 29840
rect 65108 29800 65452 29840
rect 65492 29800 65501 29840
rect 66211 29800 66220 29840
rect 66260 29800 66604 29840
rect 66644 29800 66653 29840
rect 72163 29800 72172 29840
rect 72212 29800 73132 29840
rect 73172 29800 73181 29840
rect 73315 29800 73324 29840
rect 73364 29800 73996 29840
rect 74036 29800 74764 29840
rect 74804 29800 74813 29840
rect 76675 29800 76684 29840
rect 76724 29800 77356 29840
rect 77396 29800 77405 29840
rect 39907 29672 39965 29673
rect 51532 29672 51572 29800
rect 76195 29716 76204 29756
rect 76244 29716 76876 29756
rect 76916 29716 77740 29756
rect 77780 29716 77789 29756
rect 39907 29632 39916 29672
rect 39956 29632 40588 29672
rect 40628 29632 40637 29672
rect 50467 29632 50476 29672
rect 50516 29632 50956 29672
rect 50996 29632 51572 29672
rect 60739 29632 60748 29672
rect 60788 29632 61708 29672
rect 61748 29632 61757 29672
rect 65635 29632 65644 29672
rect 65684 29632 66412 29672
rect 66452 29632 67180 29672
rect 67220 29632 67229 29672
rect 39907 29631 39965 29632
rect 56131 29548 56140 29588
rect 56180 29548 57964 29588
rect 58004 29548 58964 29588
rect 61123 29548 61132 29588
rect 61172 29548 61516 29588
rect 61556 29548 64972 29588
rect 65012 29548 65548 29588
rect 65588 29548 65597 29588
rect 71587 29548 71596 29588
rect 71636 29548 75436 29588
rect 75476 29548 75485 29588
rect 58924 29504 58964 29548
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 16343 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 16729 29504
rect 28343 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 28729 29504
rect 40343 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 40729 29504
rect 51139 29464 51148 29504
rect 51188 29464 51197 29504
rect 52343 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 52729 29504
rect 54883 29464 54892 29504
rect 54932 29464 55276 29504
rect 55316 29464 56812 29504
rect 56852 29464 57388 29504
rect 57428 29464 57437 29504
rect 58915 29464 58924 29504
rect 58964 29464 58973 29504
rect 59683 29464 59692 29504
rect 59732 29464 63380 29504
rect 64343 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 64729 29504
rect 66787 29464 66796 29504
rect 66836 29464 67372 29504
rect 67412 29464 69100 29504
rect 69140 29464 69149 29504
rect 76343 29464 76352 29504
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76720 29464 76729 29504
rect 51148 29336 51188 29464
rect 63340 29420 63380 29464
rect 59779 29380 59788 29420
rect 59828 29380 60076 29420
rect 60116 29380 63284 29420
rect 63340 29380 69196 29420
rect 69236 29380 69245 29420
rect 63244 29336 63284 29380
rect 64195 29336 64253 29337
rect 65827 29336 65885 29337
rect 39907 29296 39916 29336
rect 39956 29296 40684 29336
rect 40724 29296 47404 29336
rect 47444 29296 47453 29336
rect 51148 29296 55660 29336
rect 55700 29296 56140 29336
rect 56180 29296 56189 29336
rect 56803 29296 56812 29336
rect 56852 29296 57484 29336
rect 57524 29296 58156 29336
rect 58196 29296 58205 29336
rect 61795 29296 61804 29336
rect 61844 29296 61853 29336
rect 63244 29296 64204 29336
rect 64244 29296 64492 29336
rect 64532 29296 64541 29336
rect 65742 29296 65836 29336
rect 65876 29296 65885 29336
rect 71107 29296 71116 29336
rect 71156 29296 71308 29336
rect 71348 29296 71357 29336
rect 75907 29296 75916 29336
rect 75956 29296 76588 29336
rect 76628 29296 76637 29336
rect 76972 29296 77068 29336
rect 77108 29296 77117 29336
rect 48163 29212 48172 29252
rect 48212 29212 48652 29252
rect 48692 29212 48701 29252
rect 0 29108 80 29188
rect 42787 29128 42796 29168
rect 42836 29128 44140 29168
rect 44180 29128 44189 29168
rect 45379 29128 45388 29168
rect 45428 29128 46924 29168
rect 46964 29128 47884 29168
rect 47924 29128 47933 29168
rect 48067 29128 48076 29168
rect 48116 29128 48940 29168
rect 48980 29128 48989 29168
rect 50947 29128 50956 29168
rect 50996 29128 51436 29168
rect 51476 29128 51485 29168
rect 39907 29084 39965 29085
rect 50371 29084 50429 29085
rect 51532 29084 51572 29296
rect 61804 29168 61844 29296
rect 64195 29295 64253 29296
rect 65827 29295 65885 29296
rect 76972 29252 77012 29296
rect 64771 29212 64780 29252
rect 64820 29212 65356 29252
rect 65396 29212 65405 29252
rect 70435 29212 70444 29252
rect 70484 29212 72596 29252
rect 75811 29212 75820 29252
rect 75860 29212 76492 29252
rect 76532 29212 76541 29252
rect 76963 29212 76972 29252
rect 77012 29212 77021 29252
rect 72556 29168 72596 29212
rect 58243 29128 58252 29168
rect 58292 29128 58828 29168
rect 58868 29128 58877 29168
rect 59683 29128 59692 29168
rect 59732 29128 62284 29168
rect 62324 29128 62333 29168
rect 64867 29128 64876 29168
rect 64916 29128 65452 29168
rect 65492 29128 65501 29168
rect 69091 29128 69100 29168
rect 69140 29128 71156 29168
rect 71395 29128 71404 29168
rect 71444 29128 72268 29168
rect 72308 29128 72317 29168
rect 72547 29128 72556 29168
rect 72596 29128 72605 29168
rect 76099 29128 76108 29168
rect 76148 29128 77068 29168
rect 77108 29128 77117 29168
rect 77635 29128 77644 29168
rect 77684 29128 78028 29168
rect 78068 29128 78700 29168
rect 78740 29128 79468 29168
rect 79508 29128 79517 29168
rect 39715 29044 39724 29084
rect 39764 29044 39916 29084
rect 39956 29044 39965 29084
rect 46435 29044 46444 29084
rect 46484 29044 46636 29084
rect 46676 29044 46685 29084
rect 47395 29044 47404 29084
rect 47444 29044 47980 29084
rect 48020 29044 48029 29084
rect 48835 29044 48844 29084
rect 48884 29044 50380 29084
rect 50420 29044 50764 29084
rect 50804 29044 50813 29084
rect 51523 29044 51532 29084
rect 51572 29044 51581 29084
rect 53251 29044 53260 29084
rect 53300 29044 55180 29084
rect 55220 29044 55229 29084
rect 62467 29044 62476 29084
rect 62516 29044 65260 29084
rect 65300 29044 65309 29084
rect 65539 29044 65548 29084
rect 65588 29044 66796 29084
rect 66836 29044 66845 29084
rect 70444 29044 71020 29084
rect 71060 29044 71069 29084
rect 39907 29043 39965 29044
rect 50371 29043 50429 29044
rect 45379 28960 45388 29000
rect 45428 28960 47308 29000
rect 47348 28960 47357 29000
rect 49699 28960 49708 29000
rect 49748 28960 51244 29000
rect 51284 28960 52204 29000
rect 52244 28960 52253 29000
rect 65923 28960 65932 29000
rect 65972 28960 66412 29000
rect 66452 28960 66461 29000
rect 70444 28916 70484 29044
rect 71116 29000 71156 29128
rect 71299 29044 71308 29084
rect 71348 29044 71788 29084
rect 71828 29044 71837 29084
rect 71116 28960 71444 29000
rect 71404 28916 71444 28960
rect 77923 28916 77981 28917
rect 40099 28876 40108 28916
rect 40148 28876 40492 28916
rect 40532 28876 41068 28916
rect 41108 28876 41117 28916
rect 49507 28876 49516 28916
rect 49556 28876 54316 28916
rect 54356 28876 54365 28916
rect 60451 28876 60460 28916
rect 60500 28876 62092 28916
rect 62132 28876 65836 28916
rect 65876 28876 65885 28916
rect 68419 28876 68428 28916
rect 68468 28876 70444 28916
rect 70484 28876 70493 28916
rect 70819 28876 70828 28916
rect 70868 28876 71156 28916
rect 71395 28876 71404 28916
rect 71444 28876 71453 28916
rect 77155 28876 77164 28916
rect 77204 28876 77932 28916
rect 77972 28876 77981 28916
rect 42883 28832 42941 28833
rect 65260 28832 65300 28876
rect 71011 28832 71069 28833
rect 42798 28792 42892 28832
rect 42932 28792 42941 28832
rect 50755 28792 50764 28832
rect 50804 28792 51628 28832
rect 51668 28792 51677 28832
rect 59404 28792 60076 28832
rect 60116 28792 60125 28832
rect 62956 28792 64684 28832
rect 64724 28792 64733 28832
rect 65251 28792 65260 28832
rect 65300 28792 65340 28832
rect 66499 28792 66508 28832
rect 66548 28792 67468 28832
rect 67508 28792 71020 28832
rect 71060 28792 71069 28832
rect 42883 28791 42941 28792
rect 59404 28748 59444 28792
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 15103 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 15489 28748
rect 27103 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 27489 28748
rect 39103 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 39489 28748
rect 42499 28708 42508 28748
rect 42548 28708 43180 28748
rect 43220 28708 43229 28748
rect 51103 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 51489 28748
rect 54787 28708 54796 28748
rect 54836 28708 55084 28748
rect 55124 28708 56044 28748
rect 56084 28708 59116 28748
rect 59156 28708 59165 28748
rect 59395 28708 59404 28748
rect 59444 28708 59453 28748
rect 42691 28624 42700 28664
rect 42740 28624 43220 28664
rect 43267 28624 43276 28664
rect 43316 28624 44332 28664
rect 44372 28624 44381 28664
rect 50371 28624 50380 28664
rect 50420 28624 50860 28664
rect 50900 28624 51916 28664
rect 51956 28624 51965 28664
rect 61315 28624 61324 28664
rect 61364 28624 61804 28664
rect 61844 28624 62092 28664
rect 62132 28624 62141 28664
rect 43180 28580 43220 28624
rect 43267 28580 43325 28581
rect 62956 28580 62996 28792
rect 71011 28791 71069 28792
rect 71116 28748 71156 28876
rect 77923 28875 77981 28876
rect 72259 28792 72268 28832
rect 72308 28792 73036 28832
rect 73076 28792 73085 28832
rect 63103 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 63489 28748
rect 64291 28708 64300 28748
rect 64340 28708 65164 28748
rect 65204 28708 67180 28748
rect 67220 28708 67948 28748
rect 67988 28708 68812 28748
rect 68852 28708 69580 28748
rect 69620 28708 69629 28748
rect 71107 28708 71116 28748
rect 71156 28708 71165 28748
rect 75103 28708 75112 28748
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75480 28708 75489 28748
rect 66307 28664 66365 28665
rect 66222 28624 66316 28664
rect 66356 28624 66365 28664
rect 66307 28623 66365 28624
rect 65827 28580 65885 28581
rect 73315 28580 73373 28581
rect 42787 28540 42796 28580
rect 42836 28540 43084 28580
rect 43124 28540 43133 28580
rect 43180 28540 43276 28580
rect 43316 28540 43325 28580
rect 45187 28540 45196 28580
rect 45236 28540 53300 28580
rect 62956 28540 63052 28580
rect 63092 28540 63101 28580
rect 65827 28540 65836 28580
rect 65876 28540 66892 28580
rect 66932 28540 66941 28580
rect 70531 28540 70540 28580
rect 70580 28540 73324 28580
rect 73364 28540 73373 28580
rect 43267 28539 43325 28540
rect 52195 28496 52253 28497
rect 53260 28496 53300 28540
rect 65827 28539 65885 28540
rect 73315 28539 73373 28540
rect 70915 28496 70973 28497
rect 41644 28456 43180 28496
rect 43220 28456 43229 28496
rect 52195 28456 52204 28496
rect 52244 28456 52780 28496
rect 52820 28456 53068 28496
rect 53108 28456 53117 28496
rect 53260 28456 58924 28496
rect 58964 28456 58973 28496
rect 60931 28456 60940 28496
rect 60980 28456 62284 28496
rect 62324 28456 62333 28496
rect 70147 28456 70156 28496
rect 70196 28456 70636 28496
rect 70676 28456 70685 28496
rect 70734 28456 70743 28496
rect 70783 28456 70924 28496
rect 70964 28456 70973 28496
rect 71491 28456 71500 28496
rect 71540 28456 72748 28496
rect 72788 28456 72797 28496
rect 41644 28412 41684 28456
rect 52195 28455 52253 28456
rect 70915 28455 70973 28456
rect 40291 28372 40300 28412
rect 40340 28372 41644 28412
rect 41684 28372 41693 28412
rect 42307 28372 42316 28412
rect 42356 28372 43084 28412
rect 43124 28372 43133 28412
rect 52483 28372 52492 28412
rect 52532 28372 52541 28412
rect 60067 28372 60076 28412
rect 60116 28372 61324 28412
rect 61364 28372 61612 28412
rect 61652 28372 61661 28412
rect 62179 28372 62188 28412
rect 62228 28372 62860 28412
rect 62900 28372 64436 28412
rect 65827 28372 65836 28412
rect 65876 28372 66988 28412
rect 67028 28372 67037 28412
rect 71011 28372 71020 28412
rect 71060 28372 71884 28412
rect 71924 28372 71933 28412
rect 72067 28372 72076 28412
rect 72116 28372 72844 28412
rect 72884 28372 72893 28412
rect 0 28268 80 28348
rect 52492 28328 52532 28372
rect 64396 28328 64436 28372
rect 40771 28288 40780 28328
rect 40820 28288 43276 28328
rect 43316 28288 44044 28328
rect 44084 28288 46156 28328
rect 46196 28288 46636 28328
rect 46676 28288 49996 28328
rect 50036 28288 50045 28328
rect 51811 28288 51820 28328
rect 51860 28288 52396 28328
rect 52436 28288 52445 28328
rect 52492 28288 53452 28328
rect 53492 28288 53501 28328
rect 54403 28288 54412 28328
rect 54452 28288 54892 28328
rect 54932 28288 55276 28328
rect 55316 28288 57868 28328
rect 57908 28288 57917 28328
rect 59011 28288 59020 28328
rect 59060 28288 59788 28328
rect 59828 28288 59837 28328
rect 60163 28288 60172 28328
rect 60212 28288 60556 28328
rect 60596 28288 60844 28328
rect 60884 28288 60893 28328
rect 61027 28288 61036 28328
rect 61076 28288 61996 28328
rect 62036 28288 62045 28328
rect 62947 28288 62956 28328
rect 62996 28288 64204 28328
rect 64244 28288 64253 28328
rect 64387 28288 64396 28328
rect 64436 28288 65300 28328
rect 71779 28288 71788 28328
rect 71828 28288 72172 28328
rect 72212 28288 72221 28328
rect 72931 28288 72940 28328
rect 72980 28288 72989 28328
rect 73219 28288 73228 28328
rect 73268 28288 75724 28328
rect 75764 28288 75773 28328
rect 76867 28288 76876 28328
rect 76916 28288 77740 28328
rect 77780 28288 77789 28328
rect 50083 28244 50141 28245
rect 65260 28244 65300 28288
rect 72940 28244 72980 28288
rect 44899 28204 44908 28244
rect 44948 28204 50092 28244
rect 50132 28204 53300 28244
rect 60643 28204 60652 28244
rect 60692 28204 61900 28244
rect 61940 28204 61949 28244
rect 65251 28204 65260 28244
rect 65300 28204 65309 28244
rect 72940 28204 73708 28244
rect 73748 28204 74572 28244
rect 74612 28204 74621 28244
rect 50083 28203 50141 28204
rect 53260 28160 53300 28204
rect 53260 28120 59980 28160
rect 60020 28120 60029 28160
rect 61699 28120 61708 28160
rect 61748 28120 62764 28160
rect 62804 28120 62813 28160
rect 65347 28120 65356 28160
rect 65396 28120 66124 28160
rect 66164 28120 66173 28160
rect 68899 28120 68908 28160
rect 68948 28120 70060 28160
rect 70100 28120 70444 28160
rect 70484 28120 70493 28160
rect 71971 28120 71980 28160
rect 72020 28120 73612 28160
rect 73652 28120 73996 28160
rect 74036 28120 74045 28160
rect 77251 28076 77309 28077
rect 42499 28036 42508 28076
rect 42548 28036 42988 28076
rect 43028 28036 43037 28076
rect 48172 28036 55756 28076
rect 55796 28036 55805 28076
rect 69091 28036 69100 28076
rect 69140 28036 77260 28076
rect 77300 28036 77452 28076
rect 77492 28036 77501 28076
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 16343 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 16729 27992
rect 28343 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 28729 27992
rect 40343 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 40729 27992
rect 42211 27952 42220 27992
rect 42260 27952 43180 27992
rect 43220 27952 43229 27992
rect 48172 27908 48212 28036
rect 77251 28035 77309 28036
rect 48355 27992 48413 27993
rect 53347 27992 53405 27993
rect 48355 27952 48364 27992
rect 48404 27952 48498 27992
rect 52343 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 52729 27992
rect 53260 27952 53356 27992
rect 53396 27952 53405 27992
rect 55171 27952 55180 27992
rect 55220 27952 59308 27992
rect 59348 27952 59357 27992
rect 64343 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 64729 27992
rect 66499 27952 66508 27992
rect 66548 27952 68332 27992
rect 68372 27952 72268 27992
rect 72308 27952 72317 27992
rect 74371 27952 74380 27992
rect 74420 27952 74764 27992
rect 74804 27952 74813 27992
rect 76343 27952 76352 27992
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76720 27952 76729 27992
rect 48355 27951 48413 27952
rect 53260 27908 53300 27952
rect 53347 27951 53405 27952
rect 31651 27868 31660 27908
rect 31700 27868 48212 27908
rect 53251 27868 53260 27908
rect 53300 27868 53309 27908
rect 58819 27868 58828 27908
rect 58868 27868 66316 27908
rect 66356 27868 66365 27908
rect 43363 27824 43421 27825
rect 43278 27784 43372 27824
rect 43412 27784 43421 27824
rect 47779 27784 47788 27824
rect 47828 27784 47837 27824
rect 52003 27784 52012 27824
rect 52052 27784 52780 27824
rect 52820 27784 52829 27824
rect 60835 27784 60844 27824
rect 60884 27784 61228 27824
rect 61268 27784 61277 27824
rect 61507 27784 61516 27824
rect 61556 27784 61900 27824
rect 61940 27784 61949 27824
rect 71107 27784 71116 27824
rect 71156 27784 71500 27824
rect 71540 27784 71549 27824
rect 43363 27783 43421 27784
rect 33187 27700 33196 27740
rect 33236 27700 47348 27740
rect 42883 27656 42941 27657
rect 39619 27616 39628 27656
rect 39668 27616 40876 27656
rect 40916 27616 42124 27656
rect 42164 27616 42173 27656
rect 42595 27616 42604 27656
rect 42644 27616 42892 27656
rect 42932 27616 42941 27656
rect 43651 27616 43660 27656
rect 43700 27616 44140 27656
rect 44180 27616 45196 27656
rect 45236 27616 45245 27656
rect 42883 27615 42941 27616
rect 47308 27572 47348 27700
rect 47788 27656 47828 27784
rect 62851 27740 62909 27741
rect 48835 27700 48844 27740
rect 48884 27700 53300 27740
rect 57667 27700 57676 27740
rect 57716 27700 58060 27740
rect 58100 27700 59020 27740
rect 59060 27700 62860 27740
rect 62900 27700 62909 27740
rect 76003 27700 76012 27740
rect 76052 27700 76876 27740
rect 76916 27700 76925 27740
rect 53260 27656 53300 27700
rect 62851 27699 62909 27700
rect 47395 27616 47404 27656
rect 47444 27616 47828 27656
rect 48547 27616 48556 27656
rect 48596 27616 48748 27656
rect 48788 27616 48797 27656
rect 52003 27616 52012 27656
rect 52052 27616 52684 27656
rect 52724 27616 52733 27656
rect 53260 27616 58540 27656
rect 58580 27616 58589 27656
rect 61027 27616 61036 27656
rect 61076 27616 61900 27656
rect 61940 27616 61949 27656
rect 63619 27616 63628 27656
rect 63668 27616 64204 27656
rect 64244 27616 64253 27656
rect 65059 27616 65068 27656
rect 65108 27616 65932 27656
rect 65972 27616 65981 27656
rect 69187 27616 69196 27656
rect 69236 27616 69580 27656
rect 69620 27616 70348 27656
rect 70388 27616 73228 27656
rect 73268 27616 73277 27656
rect 75715 27616 75724 27656
rect 75764 27616 76204 27656
rect 76244 27616 76253 27656
rect 76579 27616 76588 27656
rect 76628 27616 77548 27656
rect 77588 27616 77836 27656
rect 77876 27616 77885 27656
rect 73315 27572 73373 27573
rect 31459 27532 31468 27572
rect 31508 27532 44236 27572
rect 44276 27532 44285 27572
rect 47308 27532 55948 27572
rect 55988 27532 55997 27572
rect 68419 27532 68428 27572
rect 68468 27532 71212 27572
rect 71252 27532 71404 27572
rect 71444 27532 71453 27572
rect 71500 27532 73324 27572
rect 73364 27532 75916 27572
rect 75956 27532 76108 27572
rect 76148 27532 76157 27572
rect 76483 27532 76492 27572
rect 76532 27532 77260 27572
rect 77300 27532 77309 27572
rect 0 27428 80 27508
rect 71500 27488 71540 27532
rect 73315 27531 73373 27532
rect 43747 27448 43756 27488
rect 43796 27448 44332 27488
rect 44372 27448 48844 27488
rect 48884 27448 48893 27488
rect 52099 27448 52108 27488
rect 52148 27448 52588 27488
rect 52628 27448 52637 27488
rect 60835 27448 60844 27488
rect 60884 27448 61324 27488
rect 61364 27448 61373 27488
rect 71491 27448 71500 27488
rect 71540 27448 71549 27488
rect 74467 27448 74476 27488
rect 74516 27448 76396 27488
rect 76436 27448 76445 27488
rect 44419 27364 44428 27404
rect 44468 27364 44908 27404
rect 44948 27364 44957 27404
rect 48355 27364 48364 27404
rect 48404 27364 49132 27404
rect 49172 27364 49181 27404
rect 51907 27364 51916 27404
rect 51956 27364 54412 27404
rect 54452 27364 54461 27404
rect 56227 27364 56236 27404
rect 56276 27364 58156 27404
rect 58196 27364 64876 27404
rect 64916 27364 64925 27404
rect 65827 27364 65836 27404
rect 65876 27364 66604 27404
rect 66644 27364 66653 27404
rect 71683 27364 71692 27404
rect 71732 27364 72652 27404
rect 72692 27364 72701 27404
rect 75715 27364 75724 27404
rect 75764 27364 76300 27404
rect 76340 27364 76349 27404
rect 77827 27364 77836 27404
rect 77876 27364 78604 27404
rect 78644 27364 79468 27404
rect 79508 27364 79517 27404
rect 48355 27320 48413 27321
rect 68707 27320 68765 27321
rect 69091 27320 69149 27321
rect 43363 27280 43372 27320
rect 43412 27280 47308 27320
rect 47348 27280 47357 27320
rect 48355 27280 48364 27320
rect 48404 27280 48556 27320
rect 48596 27280 48605 27320
rect 50275 27280 50284 27320
rect 50324 27280 52780 27320
rect 52820 27280 53300 27320
rect 53539 27280 53548 27320
rect 53588 27280 58732 27320
rect 58772 27280 58781 27320
rect 67747 27280 67756 27320
rect 67796 27280 68716 27320
rect 68756 27280 68765 27320
rect 69006 27280 69100 27320
rect 69140 27280 69149 27320
rect 48355 27279 48413 27280
rect 42883 27236 42941 27237
rect 52195 27236 52253 27237
rect 53260 27236 53300 27280
rect 68707 27279 68765 27280
rect 69091 27279 69149 27280
rect 69667 27320 69725 27321
rect 71299 27320 71357 27321
rect 69667 27280 69676 27320
rect 69716 27280 69772 27320
rect 69812 27280 69821 27320
rect 71299 27280 71308 27320
rect 71348 27280 71788 27320
rect 71828 27280 71837 27320
rect 73420 27280 78316 27320
rect 78356 27280 78365 27320
rect 69667 27279 69725 27280
rect 71299 27279 71357 27280
rect 68803 27236 68861 27237
rect 73420 27236 73460 27280
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 15103 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 15489 27236
rect 27103 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 27489 27236
rect 39103 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 39489 27236
rect 40771 27196 40780 27236
rect 40820 27196 41548 27236
rect 41588 27196 41597 27236
rect 42883 27196 42892 27236
rect 42932 27196 47692 27236
rect 47732 27196 48076 27236
rect 48116 27196 48125 27236
rect 51103 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 51489 27236
rect 52195 27196 52204 27236
rect 52244 27196 52300 27236
rect 52340 27196 52349 27236
rect 53260 27196 54988 27236
rect 55028 27196 55037 27236
rect 55555 27196 55564 27236
rect 55604 27196 62572 27236
rect 62612 27196 62621 27236
rect 63103 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 63489 27236
rect 68515 27196 68524 27236
rect 68564 27196 68812 27236
rect 68852 27196 68861 27236
rect 69955 27196 69964 27236
rect 70004 27196 73132 27236
rect 73172 27196 73460 27236
rect 75103 27196 75112 27236
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75480 27196 75489 27236
rect 42883 27195 42941 27196
rect 52195 27195 52253 27196
rect 68803 27195 68861 27196
rect 74851 27152 74909 27153
rect 40195 27112 40204 27152
rect 40244 27112 40820 27152
rect 49219 27112 49228 27152
rect 49268 27112 49420 27152
rect 49460 27112 51724 27152
rect 51764 27112 52108 27152
rect 52148 27112 52780 27152
rect 52820 27112 52829 27152
rect 60739 27112 60748 27152
rect 60788 27112 61228 27152
rect 61268 27112 61277 27152
rect 71587 27112 71596 27152
rect 71636 27112 72940 27152
rect 72980 27112 72989 27152
rect 74766 27112 74860 27152
rect 74900 27112 74909 27152
rect 40195 27068 40253 27069
rect 40195 27028 40204 27068
rect 40244 27028 40396 27068
rect 40436 27028 40445 27068
rect 40195 27027 40253 27028
rect 40099 26984 40157 26985
rect 38371 26944 38380 26984
rect 38420 26944 40108 26984
rect 40148 26944 40492 26984
rect 40532 26944 40541 26984
rect 40099 26943 40157 26944
rect 40780 26900 40820 27112
rect 74851 27111 74909 27112
rect 52963 27068 53021 27069
rect 50851 27028 50860 27068
rect 50900 27028 52876 27068
rect 52916 27028 52972 27068
rect 53012 27028 53040 27068
rect 59107 27028 59116 27068
rect 59156 27028 65740 27068
rect 65780 27028 65789 27068
rect 77731 27028 77740 27068
rect 77780 27028 77932 27068
rect 77972 27028 78124 27068
rect 78164 27028 78173 27068
rect 52963 27027 53021 27028
rect 71683 26984 71741 26985
rect 43180 26944 43372 26984
rect 43412 26944 43421 26984
rect 52771 26944 52780 26984
rect 52820 26944 53548 26984
rect 53588 26944 53597 26984
rect 60547 26944 60556 26984
rect 60596 26944 60748 26984
rect 60788 26944 60797 26984
rect 62371 26944 62380 26984
rect 62420 26944 63916 26984
rect 63956 26944 63965 26984
rect 64099 26944 64108 26984
rect 64148 26944 65164 26984
rect 65204 26944 65213 26984
rect 71598 26944 71692 26984
rect 71732 26944 71741 26984
rect 40003 26860 40012 26900
rect 40052 26860 40588 26900
rect 40628 26860 40637 26900
rect 40771 26860 40780 26900
rect 40820 26860 41836 26900
rect 41876 26860 41885 26900
rect 43180 26816 43220 26944
rect 71683 26943 71741 26944
rect 58435 26900 58493 26901
rect 61603 26900 61661 26901
rect 64195 26900 64253 26901
rect 70915 26900 70973 26901
rect 47203 26860 47212 26900
rect 47252 26860 47692 26900
rect 47732 26860 47741 26900
rect 58350 26860 58444 26900
rect 58484 26860 58493 26900
rect 59011 26860 59020 26900
rect 59060 26860 60844 26900
rect 60884 26860 60893 26900
rect 61518 26860 61612 26900
rect 61652 26860 62092 26900
rect 62132 26860 62141 26900
rect 64195 26860 64204 26900
rect 64244 26860 64396 26900
rect 64436 26860 64445 26900
rect 70830 26860 70924 26900
rect 70964 26860 70973 26900
rect 71107 26860 71116 26900
rect 71156 26860 72076 26900
rect 72116 26860 72125 26900
rect 58435 26859 58493 26860
rect 61603 26859 61661 26860
rect 64195 26859 64253 26860
rect 70915 26859 70973 26860
rect 38659 26776 38668 26816
rect 38708 26776 39436 26816
rect 39476 26776 39485 26816
rect 39715 26776 39724 26816
rect 39764 26776 40204 26816
rect 40244 26776 40253 26816
rect 40387 26776 40396 26816
rect 40436 26776 40876 26816
rect 40916 26776 40925 26816
rect 41443 26776 41452 26816
rect 41492 26776 41644 26816
rect 41684 26776 42508 26816
rect 42548 26776 42557 26816
rect 43075 26776 43084 26816
rect 43124 26776 43220 26816
rect 48067 26776 48076 26816
rect 48116 26776 48460 26816
rect 48500 26776 48509 26816
rect 52675 26776 52684 26816
rect 52724 26776 53932 26816
rect 53972 26776 53981 26816
rect 54595 26776 54604 26816
rect 54644 26776 56044 26816
rect 56084 26776 57004 26816
rect 57044 26776 57053 26816
rect 60259 26776 60268 26816
rect 60308 26776 61804 26816
rect 61844 26776 61853 26816
rect 63715 26776 63724 26816
rect 63764 26776 64972 26816
rect 65012 26776 65021 26816
rect 70051 26776 70060 26816
rect 70100 26776 72364 26816
rect 72404 26776 73132 26816
rect 73172 26776 73460 26816
rect 74467 26776 74476 26816
rect 74516 26776 75820 26816
rect 75860 26776 75869 26816
rect 77347 26776 77356 26816
rect 77396 26776 78508 26816
rect 78548 26776 78557 26816
rect 40003 26732 40061 26733
rect 63916 26732 63956 26776
rect 73420 26732 73460 26776
rect 40003 26692 40012 26732
rect 40052 26692 40300 26732
rect 40340 26692 40349 26732
rect 40483 26692 40492 26732
rect 40532 26692 40780 26732
rect 40820 26692 40829 26732
rect 48355 26692 48364 26732
rect 48404 26692 49036 26732
rect 49076 26692 50956 26732
rect 50996 26692 57695 26732
rect 60067 26692 60076 26732
rect 60116 26692 61420 26732
rect 61460 26692 63380 26732
rect 63907 26692 63916 26732
rect 63956 26692 63996 26732
rect 73420 26692 74956 26732
rect 74996 26692 75005 26732
rect 40003 26691 40061 26692
rect 0 26588 80 26668
rect 49123 26648 49181 26649
rect 57655 26648 57695 26692
rect 63340 26648 63380 26692
rect 71683 26648 71741 26649
rect 75820 26648 75860 26776
rect 40099 26608 40108 26648
rect 40148 26608 40588 26648
rect 40628 26608 40637 26648
rect 49038 26608 49132 26648
rect 49172 26608 49181 26648
rect 51715 26608 51724 26648
rect 51764 26608 53356 26648
rect 53396 26608 53548 26648
rect 53588 26608 53597 26648
rect 54019 26608 54028 26648
rect 54068 26608 55084 26648
rect 55124 26608 55133 26648
rect 57655 26608 62284 26648
rect 62324 26608 62333 26648
rect 63340 26608 64588 26648
rect 64628 26608 64637 26648
rect 68035 26608 68044 26648
rect 68084 26608 69772 26648
rect 69812 26608 69821 26648
rect 70819 26608 70828 26648
rect 70868 26608 71692 26648
rect 71732 26608 74860 26648
rect 74900 26608 74909 26648
rect 75820 26608 77836 26648
rect 77876 26608 78220 26648
rect 78260 26608 78269 26648
rect 49123 26607 49181 26608
rect 71683 26607 71741 26608
rect 835 26524 844 26564
rect 884 26524 49804 26564
rect 49844 26524 49853 26564
rect 59203 26524 59212 26564
rect 59252 26524 59292 26564
rect 60163 26524 60172 26564
rect 60212 26524 60460 26564
rect 60500 26524 64916 26564
rect 64963 26524 64972 26564
rect 65012 26524 65260 26564
rect 65300 26524 65309 26564
rect 69667 26524 69676 26564
rect 69716 26524 70444 26564
rect 70484 26524 70493 26564
rect 49891 26480 49949 26481
rect 52963 26480 53021 26481
rect 59212 26480 59252 26524
rect 64876 26480 64916 26524
rect 69763 26480 69821 26481
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 16343 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 16729 26480
rect 28343 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 28729 26480
rect 40343 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 40729 26480
rect 42787 26440 42796 26480
rect 42836 26440 49900 26480
rect 49940 26440 49949 26480
rect 52343 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 52729 26480
rect 52963 26440 52972 26480
rect 53012 26440 53356 26480
rect 53396 26440 53405 26480
rect 53635 26440 53644 26480
rect 53684 26440 54124 26480
rect 54164 26440 55564 26480
rect 55604 26440 55613 26480
rect 58627 26440 58636 26480
rect 58676 26440 63380 26480
rect 64343 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 64729 26480
rect 64876 26440 69772 26480
rect 69812 26440 69964 26480
rect 70004 26440 70013 26480
rect 70156 26440 75244 26480
rect 75284 26440 75293 26480
rect 76343 26440 76352 26480
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76720 26440 76729 26480
rect 77731 26440 77740 26480
rect 77780 26440 78028 26480
rect 78068 26440 78077 26480
rect 49891 26439 49949 26440
rect 52963 26439 53021 26440
rect 43267 26396 43325 26397
rect 63340 26396 63380 26440
rect 69763 26439 69821 26440
rect 70156 26396 70196 26440
rect 40963 26356 40972 26396
rect 41012 26356 43276 26396
rect 43316 26356 44716 26396
rect 44756 26356 45772 26396
rect 45812 26356 48652 26396
rect 48692 26356 48701 26396
rect 53251 26356 53260 26396
rect 53300 26356 53836 26396
rect 53876 26356 53885 26396
rect 54787 26356 54796 26396
rect 54836 26356 55372 26396
rect 55412 26356 56524 26396
rect 56564 26356 56573 26396
rect 61411 26356 61420 26396
rect 61460 26356 61900 26396
rect 61940 26356 61949 26396
rect 63340 26356 70156 26396
rect 70196 26356 70205 26396
rect 43267 26355 43325 26356
rect 69283 26312 69341 26313
rect 40867 26272 40876 26312
rect 40916 26272 42412 26312
rect 42452 26272 42461 26312
rect 42979 26272 42988 26312
rect 43028 26272 43468 26312
rect 43508 26272 43517 26312
rect 43651 26272 43660 26312
rect 43700 26272 45196 26312
rect 45236 26272 45245 26312
rect 45379 26272 45388 26312
rect 45428 26272 59020 26312
rect 59060 26272 59069 26312
rect 60460 26272 60652 26312
rect 60692 26272 64108 26312
rect 64148 26272 64684 26312
rect 64724 26272 64733 26312
rect 69198 26272 69292 26312
rect 69332 26272 69341 26312
rect 69667 26272 69676 26312
rect 69716 26272 71500 26312
rect 71540 26272 71549 26312
rect 76579 26272 76588 26312
rect 76628 26272 77644 26312
rect 77684 26272 77932 26312
rect 77972 26272 77981 26312
rect 42412 26228 42452 26272
rect 60460 26228 60500 26272
rect 69283 26271 69341 26272
rect 40387 26188 40396 26228
rect 40436 26188 41068 26228
rect 41108 26188 41204 26228
rect 42412 26188 48212 26228
rect 50755 26188 50764 26228
rect 50804 26188 54796 26228
rect 54836 26188 54845 26228
rect 54979 26188 54988 26228
rect 55028 26188 57676 26228
rect 57716 26188 57725 26228
rect 59107 26188 59116 26228
rect 59156 26188 59500 26228
rect 59540 26188 59549 26228
rect 59683 26188 59692 26228
rect 59732 26188 59980 26228
rect 60020 26188 60500 26228
rect 69187 26188 69196 26228
rect 69236 26188 69484 26228
rect 69524 26188 69964 26228
rect 70004 26188 70540 26228
rect 70580 26188 70828 26228
rect 70868 26188 70877 26228
rect 74563 26188 74572 26228
rect 74612 26188 75820 26228
rect 75860 26188 75869 26228
rect 41059 26144 41117 26145
rect 39619 26104 39628 26144
rect 39668 26104 41068 26144
rect 41108 26104 41117 26144
rect 41164 26144 41204 26188
rect 41164 26104 43660 26144
rect 43700 26104 44044 26144
rect 44084 26104 44093 26144
rect 44419 26104 44428 26144
rect 44468 26104 44812 26144
rect 44852 26104 44861 26144
rect 45187 26104 45196 26144
rect 45236 26104 45868 26144
rect 45908 26104 45917 26144
rect 41059 26103 41117 26104
rect 48172 26060 48212 26188
rect 77251 26144 77309 26145
rect 49027 26104 49036 26144
rect 49076 26104 49996 26144
rect 50036 26104 50045 26144
rect 53155 26104 53164 26144
rect 53204 26104 54124 26144
rect 54164 26104 54173 26144
rect 55075 26104 55084 26144
rect 55124 26104 55852 26144
rect 55892 26104 55901 26144
rect 55948 26104 58348 26144
rect 58388 26104 58397 26144
rect 58819 26104 58828 26144
rect 58868 26104 60268 26144
rect 60308 26104 60317 26144
rect 61315 26104 61324 26144
rect 61364 26104 61373 26144
rect 65635 26104 65644 26144
rect 65684 26104 65932 26144
rect 65972 26104 65981 26144
rect 66115 26104 66124 26144
rect 66164 26104 69004 26144
rect 69044 26104 69053 26144
rect 69379 26104 69388 26144
rect 69428 26104 69524 26144
rect 69763 26104 69772 26144
rect 69812 26104 71116 26144
rect 71156 26104 71165 26144
rect 72835 26104 72844 26144
rect 72884 26104 73324 26144
rect 73364 26104 73708 26144
rect 73748 26104 74380 26144
rect 74420 26104 74429 26144
rect 76003 26104 76012 26144
rect 76052 26104 76684 26144
rect 76724 26104 76733 26144
rect 77166 26104 77260 26144
rect 77300 26104 77309 26144
rect 55948 26060 55988 26104
rect 41923 26020 41932 26060
rect 41972 26020 42796 26060
rect 42836 26020 42845 26060
rect 43075 26020 43084 26060
rect 43124 26020 43564 26060
rect 43604 26020 43613 26060
rect 43747 26020 43756 26060
rect 43796 26020 44524 26060
rect 44564 26020 44573 26060
rect 48172 26020 55988 26060
rect 56227 26020 56236 26060
rect 56276 26020 57004 26060
rect 57044 26020 57053 26060
rect 36931 25936 36940 25976
rect 36980 25936 38668 25976
rect 38708 25936 38717 25976
rect 39523 25936 39532 25976
rect 39572 25936 40972 25976
rect 41012 25936 41021 25976
rect 42115 25936 42124 25976
rect 42164 25936 43660 25976
rect 43700 25936 43709 25976
rect 44323 25936 44332 25976
rect 44372 25936 45196 25976
rect 45236 25936 45245 25976
rect 45955 25936 45964 25976
rect 46004 25936 46636 25976
rect 46676 25936 48172 25976
rect 48212 25936 48221 25976
rect 53923 25936 53932 25976
rect 53972 25936 54796 25976
rect 54836 25936 54845 25976
rect 55939 25936 55948 25976
rect 55988 25936 56140 25976
rect 56180 25936 56524 25976
rect 56564 25936 56573 25976
rect 57667 25936 57676 25976
rect 57716 25936 57964 25976
rect 58004 25936 58013 25976
rect 59587 25936 59596 25976
rect 59636 25936 59980 25976
rect 60020 25936 60029 25976
rect 43363 25892 43421 25893
rect 53347 25892 53405 25893
rect 61324 25892 61364 26104
rect 62755 26020 62764 26060
rect 62804 26020 63628 26060
rect 63668 26020 65260 26060
rect 65300 26020 66508 26060
rect 66548 26020 66557 26060
rect 63235 25936 63244 25976
rect 63284 25936 64876 25976
rect 64916 25936 65452 25976
rect 65492 25936 65501 25976
rect 69484 25892 69524 26104
rect 77251 26103 77309 26104
rect 69571 26020 69580 26060
rect 69620 26020 70004 26060
rect 70627 26020 70636 26060
rect 70676 26020 71596 26060
rect 71636 26020 71645 26060
rect 72067 26020 72076 26060
rect 72116 26020 72748 26060
rect 72788 26020 72797 26060
rect 74563 26020 74572 26060
rect 74612 26020 74764 26060
rect 74804 26020 74813 26060
rect 69859 25976 69917 25977
rect 69774 25936 69868 25976
rect 69908 25936 69917 25976
rect 69964 25976 70004 26020
rect 69964 25936 70772 25976
rect 71971 25936 71980 25976
rect 72020 25936 73420 25976
rect 73460 25936 73900 25976
rect 73940 25936 73949 25976
rect 75427 25936 75436 25976
rect 75476 25936 75628 25976
rect 75668 25936 75677 25976
rect 75907 25936 75916 25976
rect 75956 25936 76204 25976
rect 76244 25936 76876 25976
rect 76916 25936 76925 25976
rect 69859 25935 69917 25936
rect 39427 25852 39436 25892
rect 39476 25852 39628 25892
rect 39668 25852 39677 25892
rect 40771 25852 40780 25892
rect 40820 25852 43372 25892
rect 43412 25852 43421 25892
rect 43363 25851 43421 25852
rect 43468 25852 44908 25892
rect 44948 25852 44957 25892
rect 45379 25852 45388 25892
rect 45428 25852 47116 25892
rect 47156 25852 47165 25892
rect 49027 25852 49036 25892
rect 49076 25852 50572 25892
rect 50612 25852 50621 25892
rect 53059 25852 53068 25892
rect 53108 25852 53356 25892
rect 53396 25852 53405 25892
rect 54019 25852 54028 25892
rect 54068 25852 57388 25892
rect 57428 25852 57437 25892
rect 57859 25852 57868 25892
rect 57908 25852 59884 25892
rect 59924 25852 59933 25892
rect 60547 25852 60556 25892
rect 60596 25852 61996 25892
rect 62036 25852 62045 25892
rect 69484 25852 70484 25892
rect 0 25808 80 25828
rect 40003 25808 40061 25809
rect 0 25768 652 25808
rect 692 25768 701 25808
rect 40003 25768 40012 25808
rect 40052 25768 40108 25808
rect 40148 25768 40157 25808
rect 42787 25768 42796 25808
rect 42836 25768 43220 25808
rect 0 25748 80 25768
rect 40003 25767 40061 25768
rect 43180 25724 43220 25768
rect 43468 25724 43508 25852
rect 53347 25851 53405 25852
rect 54028 25808 54068 25852
rect 70444 25808 70484 25852
rect 70732 25808 70772 25936
rect 46915 25768 46924 25808
rect 46964 25768 48940 25808
rect 48980 25768 48989 25808
rect 50371 25768 50380 25808
rect 50420 25768 54068 25808
rect 59299 25768 59308 25808
rect 59348 25768 59596 25808
rect 59636 25768 59645 25808
rect 60739 25768 60748 25808
rect 60788 25768 62764 25808
rect 62804 25768 65548 25808
rect 65588 25768 65597 25808
rect 70435 25768 70444 25808
rect 70484 25768 70493 25808
rect 70723 25768 70732 25808
rect 70772 25768 70781 25808
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 15103 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 15489 25724
rect 27103 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 27489 25724
rect 39103 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 39489 25724
rect 43180 25684 43508 25724
rect 43756 25684 46444 25724
rect 46484 25684 47308 25724
rect 47348 25684 47596 25724
rect 47636 25684 47645 25724
rect 51103 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 51489 25724
rect 52291 25684 52300 25724
rect 52340 25684 56660 25724
rect 59203 25684 59212 25724
rect 59252 25684 60268 25724
rect 60308 25684 60317 25724
rect 63103 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 63489 25724
rect 69667 25684 69676 25724
rect 69716 25684 70252 25724
rect 70292 25684 70301 25724
rect 75103 25684 75112 25724
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75480 25684 75489 25724
rect 42883 25640 42941 25641
rect 42883 25600 42892 25640
rect 42932 25600 43564 25640
rect 43604 25600 43613 25640
rect 42883 25599 42941 25600
rect 43756 25556 43796 25684
rect 54499 25640 54557 25641
rect 56620 25640 56660 25684
rect 44899 25600 44908 25640
rect 44948 25600 45484 25640
rect 45524 25600 45533 25640
rect 45667 25600 45676 25640
rect 45716 25600 47212 25640
rect 47252 25600 53300 25640
rect 54414 25600 54508 25640
rect 54548 25600 54557 25640
rect 56611 25600 56620 25640
rect 56660 25600 57292 25640
rect 57332 25600 57772 25640
rect 57812 25600 57821 25640
rect 62083 25600 62092 25640
rect 62132 25600 70100 25640
rect 51523 25556 51581 25557
rect 53260 25556 53300 25600
rect 54499 25599 54557 25600
rect 66595 25556 66653 25557
rect 7171 25516 7180 25556
rect 7220 25516 41740 25556
rect 41780 25516 41789 25556
rect 42307 25516 42316 25556
rect 42356 25516 42508 25556
rect 42548 25516 43796 25556
rect 48259 25516 48268 25556
rect 48308 25516 49132 25556
rect 49172 25516 49181 25556
rect 49891 25516 49900 25556
rect 49940 25516 51532 25556
rect 51572 25516 52300 25556
rect 52340 25516 52349 25556
rect 53260 25516 56276 25556
rect 56419 25516 56428 25556
rect 56468 25516 57484 25556
rect 57524 25516 57533 25556
rect 59971 25516 59980 25556
rect 60020 25516 60364 25556
rect 60404 25516 60748 25556
rect 60788 25516 60797 25556
rect 66510 25516 66604 25556
rect 66644 25516 66653 25556
rect 68803 25516 68812 25556
rect 68852 25516 69484 25556
rect 69524 25516 69533 25556
rect 51523 25515 51581 25516
rect 51907 25472 51965 25473
rect 43267 25432 43276 25472
rect 43316 25432 43468 25472
rect 43508 25432 46924 25472
rect 46964 25432 46973 25472
rect 47395 25432 47404 25472
rect 47444 25432 47788 25472
rect 47828 25432 47837 25472
rect 49795 25432 49804 25472
rect 49844 25432 51916 25472
rect 51956 25432 51965 25472
rect 54211 25432 54220 25472
rect 54260 25432 54604 25472
rect 54644 25432 54653 25472
rect 51907 25431 51965 25432
rect 41347 25348 41356 25388
rect 41396 25348 42124 25388
rect 42164 25348 42604 25388
rect 42644 25348 50572 25388
rect 50612 25348 50621 25388
rect 36451 25264 36460 25304
rect 36500 25264 37708 25304
rect 37748 25264 37757 25304
rect 39811 25264 39820 25304
rect 39860 25264 42796 25304
rect 42836 25264 43084 25304
rect 43124 25264 43133 25304
rect 44995 25264 45004 25304
rect 45044 25264 45676 25304
rect 45716 25264 45725 25304
rect 48163 25264 48172 25304
rect 48212 25264 48460 25304
rect 48500 25264 48509 25304
rect 40291 25220 40349 25221
rect 45571 25220 45629 25221
rect 49132 25220 49172 25348
rect 56236 25304 56276 25516
rect 66595 25515 66653 25516
rect 56707 25432 56716 25472
rect 56756 25432 57772 25472
rect 57812 25432 58444 25472
rect 58484 25432 58493 25472
rect 63043 25432 63052 25472
rect 63092 25432 63724 25472
rect 63764 25432 63773 25472
rect 65827 25432 65836 25472
rect 65876 25432 67180 25472
rect 67220 25432 67229 25472
rect 58723 25388 58781 25389
rect 69763 25388 69821 25389
rect 70060 25388 70100 25600
rect 58638 25348 58732 25388
rect 58772 25348 58781 25388
rect 58915 25348 58924 25388
rect 58964 25348 60172 25388
rect 60212 25348 64052 25388
rect 64099 25348 64108 25388
rect 64148 25348 66700 25388
rect 66740 25348 67276 25388
rect 67316 25348 67325 25388
rect 69763 25348 69772 25388
rect 69812 25348 69868 25388
rect 69908 25348 69917 25388
rect 70051 25348 70060 25388
rect 70100 25348 72460 25388
rect 72500 25348 72509 25388
rect 58723 25347 58781 25348
rect 64012 25304 64052 25348
rect 69763 25347 69821 25348
rect 75043 25304 75101 25305
rect 49219 25264 49228 25304
rect 49268 25264 50092 25304
rect 50132 25264 50141 25304
rect 50659 25264 50668 25304
rect 50708 25264 51916 25304
rect 51956 25264 53740 25304
rect 53780 25264 54316 25304
rect 54356 25264 54365 25304
rect 54499 25264 54508 25304
rect 54548 25264 54796 25304
rect 54836 25264 54845 25304
rect 56236 25264 59212 25304
rect 59252 25264 59261 25304
rect 59491 25264 59500 25304
rect 59540 25264 60076 25304
rect 60116 25264 60556 25304
rect 60596 25264 60605 25304
rect 60835 25264 60844 25304
rect 60884 25264 61324 25304
rect 61364 25264 63628 25304
rect 63668 25264 63677 25304
rect 64012 25264 64244 25304
rect 65539 25264 65548 25304
rect 65588 25264 66124 25304
rect 66164 25264 66796 25304
rect 66836 25264 66845 25304
rect 67171 25264 67180 25304
rect 67220 25264 67229 25304
rect 67459 25264 67468 25304
rect 67508 25264 68524 25304
rect 68564 25264 68573 25304
rect 71203 25264 71212 25304
rect 71252 25264 71980 25304
rect 72020 25264 72029 25304
rect 72163 25264 72172 25304
rect 72212 25264 72844 25304
rect 72884 25264 72893 25304
rect 75043 25264 75052 25304
rect 75092 25264 75916 25304
rect 75956 25264 76300 25304
rect 76340 25264 76349 25304
rect 76483 25264 76492 25304
rect 76532 25264 77356 25304
rect 77396 25264 77405 25304
rect 77539 25264 77548 25304
rect 77588 25264 78220 25304
rect 78260 25264 79276 25304
rect 79316 25264 79325 25304
rect 50563 25220 50621 25221
rect 2371 25180 2380 25220
rect 2420 25180 40300 25220
rect 40340 25180 40349 25220
rect 40771 25180 40780 25220
rect 40820 25180 42028 25220
rect 42068 25180 42700 25220
rect 42740 25180 44084 25220
rect 44611 25180 44620 25220
rect 44660 25180 45580 25220
rect 45620 25180 45629 25220
rect 47971 25180 47980 25220
rect 48020 25180 48268 25220
rect 48308 25180 48317 25220
rect 49123 25180 49132 25220
rect 49172 25180 49181 25220
rect 50563 25180 50572 25220
rect 50612 25180 52108 25220
rect 52148 25180 52157 25220
rect 53059 25180 53068 25220
rect 53108 25180 62668 25220
rect 62708 25180 62717 25220
rect 40291 25179 40349 25180
rect 41059 25136 41117 25137
rect 37795 25096 37804 25136
rect 37844 25096 38188 25136
rect 38228 25096 38237 25136
rect 39331 25096 39340 25136
rect 39380 25096 39628 25136
rect 39668 25096 40588 25136
rect 40628 25096 40637 25136
rect 40974 25096 41068 25136
rect 41108 25096 41117 25136
rect 40588 25052 40628 25096
rect 41059 25095 41117 25096
rect 44044 25052 44084 25180
rect 45571 25179 45629 25180
rect 50563 25179 50621 25180
rect 50572 25136 50612 25179
rect 44131 25096 44140 25136
rect 44180 25096 44908 25136
rect 44948 25096 44957 25136
rect 45475 25096 45484 25136
rect 45524 25096 50612 25136
rect 50755 25136 50813 25137
rect 50755 25096 50764 25136
rect 50804 25096 50898 25136
rect 51139 25096 51148 25136
rect 51188 25096 51532 25136
rect 51572 25096 51581 25136
rect 58531 25096 58540 25136
rect 58580 25096 59596 25136
rect 59636 25096 59645 25136
rect 61987 25096 61996 25136
rect 62036 25096 64108 25136
rect 64148 25096 64157 25136
rect 50755 25095 50813 25096
rect 64204 25052 64244 25264
rect 67180 25220 67220 25264
rect 75043 25263 75101 25264
rect 67555 25220 67613 25221
rect 64579 25180 64588 25220
rect 64628 25180 65740 25220
rect 65780 25180 67220 25220
rect 67470 25180 67564 25220
rect 67604 25180 67613 25220
rect 69379 25180 69388 25220
rect 69428 25180 69676 25220
rect 69716 25180 70060 25220
rect 70100 25180 71116 25220
rect 71156 25180 72268 25220
rect 72308 25180 72317 25220
rect 73219 25180 73228 25220
rect 73268 25180 75052 25220
rect 75092 25180 75101 25220
rect 76963 25180 76972 25220
rect 77012 25180 77021 25220
rect 67555 25179 67613 25180
rect 76771 25136 76829 25137
rect 76972 25136 77012 25180
rect 64771 25096 64780 25136
rect 64820 25096 67372 25136
rect 67412 25096 67421 25136
rect 71980 25096 73132 25136
rect 73172 25096 73612 25136
rect 73652 25096 73661 25136
rect 76771 25096 76780 25136
rect 76820 25096 76876 25136
rect 76916 25096 76925 25136
rect 76972 25096 78124 25136
rect 78164 25096 78892 25136
rect 78932 25096 78941 25136
rect 71980 25052 72020 25096
rect 76771 25095 76829 25096
rect 77251 25052 77309 25053
rect 40588 25012 43220 25052
rect 44044 25012 45388 25052
rect 45428 25012 45437 25052
rect 64204 25012 68428 25052
rect 68468 25012 68756 25052
rect 71971 25012 71980 25052
rect 72020 25012 72029 25052
rect 76963 25012 76972 25052
rect 77012 25012 77260 25052
rect 77300 25012 77309 25052
rect 0 24968 80 24988
rect 43180 24968 43220 25012
rect 52771 24968 52829 24969
rect 56131 24968 56189 24969
rect 57571 24968 57629 24969
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 16343 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 16729 24968
rect 28343 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 28729 24968
rect 40343 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 40729 24968
rect 43180 24928 45196 24968
rect 45236 24928 45245 24968
rect 52343 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 52729 24968
rect 52771 24928 52780 24968
rect 52820 24928 56140 24968
rect 56180 24928 56189 24968
rect 56707 24928 56716 24968
rect 56756 24928 56908 24968
rect 56948 24928 56957 24968
rect 57571 24928 57580 24968
rect 57620 24928 60172 24968
rect 60212 24928 60221 24968
rect 64343 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 64729 24968
rect 66979 24928 66988 24968
rect 67028 24928 67372 24968
rect 67412 24928 67421 24968
rect 0 24908 80 24928
rect 52771 24927 52829 24928
rect 56131 24927 56189 24928
rect 57571 24927 57629 24928
rect 68716 24884 68756 25012
rect 77251 25011 77309 25012
rect 75523 24928 75532 24968
rect 75572 24928 75820 24968
rect 75860 24928 75869 24968
rect 76343 24928 76352 24968
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76720 24928 76729 24968
rect 40867 24844 40876 24884
rect 40916 24844 58060 24884
rect 58100 24844 58109 24884
rect 59395 24844 59404 24884
rect 59444 24844 59788 24884
rect 59828 24844 59837 24884
rect 60259 24844 60268 24884
rect 60308 24844 65548 24884
rect 65588 24844 65597 24884
rect 68707 24844 68716 24884
rect 68756 24844 76204 24884
rect 76244 24844 76253 24884
rect 1795 24760 1804 24800
rect 1844 24760 2380 24800
rect 2420 24760 2429 24800
rect 39907 24760 39916 24800
rect 39956 24760 43220 24800
rect 49219 24760 49228 24800
rect 49268 24760 49420 24800
rect 49460 24760 49469 24800
rect 50275 24760 50284 24800
rect 50324 24760 50476 24800
rect 50516 24760 50525 24800
rect 51811 24760 51820 24800
rect 51860 24760 52300 24800
rect 52340 24760 52349 24800
rect 55075 24760 55084 24800
rect 55124 24760 57620 24800
rect 59875 24760 59884 24800
rect 59924 24760 60748 24800
rect 60788 24760 62188 24800
rect 62228 24760 62237 24800
rect 62851 24760 62860 24800
rect 62900 24760 64684 24800
rect 64724 24760 64733 24800
rect 72259 24760 72268 24800
rect 72308 24760 72940 24800
rect 72980 24760 75532 24800
rect 75572 24760 76684 24800
rect 76724 24760 76733 24800
rect 77059 24760 77068 24800
rect 77108 24760 77117 24800
rect 43180 24716 43220 24760
rect 57580 24716 57620 24760
rect 38467 24676 38476 24716
rect 38516 24676 38956 24716
rect 38996 24676 39005 24716
rect 41059 24676 41068 24716
rect 41108 24676 42796 24716
rect 42836 24676 42845 24716
rect 43180 24676 57484 24716
rect 57524 24676 57533 24716
rect 57580 24676 60556 24716
rect 60596 24676 60605 24716
rect 61315 24676 61324 24716
rect 61364 24676 61373 24716
rect 61324 24632 61364 24676
rect 34915 24592 34924 24632
rect 34964 24592 36364 24632
rect 36404 24592 38092 24632
rect 38132 24592 38572 24632
rect 38612 24592 39724 24632
rect 39764 24592 41260 24632
rect 41300 24592 42316 24632
rect 42356 24592 44908 24632
rect 44948 24592 45100 24632
rect 45140 24592 47500 24632
rect 47540 24592 47692 24632
rect 47732 24592 47741 24632
rect 48931 24592 48940 24632
rect 48980 24592 55084 24632
rect 55124 24592 55133 24632
rect 55267 24592 55276 24632
rect 55316 24592 57868 24632
rect 57908 24592 57917 24632
rect 59875 24592 59884 24632
rect 59924 24592 61364 24632
rect 62188 24632 62228 24760
rect 77068 24716 77108 24760
rect 64099 24676 64108 24716
rect 64148 24676 64492 24716
rect 64532 24676 64541 24716
rect 75235 24676 75244 24716
rect 75284 24676 75436 24716
rect 75476 24676 75485 24716
rect 76387 24676 76396 24716
rect 76436 24676 77108 24716
rect 62188 24592 63532 24632
rect 63572 24592 64588 24632
rect 64628 24592 67660 24632
rect 67700 24592 72940 24632
rect 72980 24592 74476 24632
rect 74516 24592 74525 24632
rect 75619 24592 75628 24632
rect 75668 24592 77068 24632
rect 77108 24592 77117 24632
rect 51907 24548 51965 24549
rect 835 24508 844 24548
rect 884 24508 2188 24548
rect 2228 24508 2237 24548
rect 35203 24508 35212 24548
rect 35252 24508 36460 24548
rect 36500 24508 36509 24548
rect 45187 24508 45196 24548
rect 45236 24508 47596 24548
rect 47636 24508 48268 24548
rect 48308 24508 48317 24548
rect 49795 24508 49804 24548
rect 49844 24508 50956 24548
rect 50996 24508 51244 24548
rect 51284 24508 51293 24548
rect 51907 24508 51916 24548
rect 51956 24508 52108 24548
rect 52148 24508 52157 24548
rect 52291 24508 52300 24548
rect 52340 24508 53836 24548
rect 53876 24508 61324 24548
rect 61364 24508 61373 24548
rect 65923 24508 65932 24548
rect 65972 24508 66412 24548
rect 66452 24508 67084 24548
rect 67124 24508 67133 24548
rect 72835 24508 72844 24548
rect 72884 24508 73612 24548
rect 73652 24508 74092 24548
rect 74132 24508 74141 24548
rect 74659 24508 74668 24548
rect 74708 24508 75092 24548
rect 75139 24508 75148 24548
rect 75188 24508 75916 24548
rect 75956 24508 76108 24548
rect 76148 24508 76157 24548
rect 41347 24464 41405 24465
rect 46636 24464 46676 24508
rect 51907 24507 51965 24508
rect 58243 24464 58301 24465
rect 67555 24464 67613 24465
rect 69283 24464 69341 24465
rect 75052 24464 75092 24508
rect 36643 24424 36652 24464
rect 36692 24424 41356 24464
rect 41396 24424 41405 24464
rect 46627 24424 46636 24464
rect 46676 24424 46685 24464
rect 48835 24424 48844 24464
rect 48884 24424 50476 24464
rect 50516 24424 50525 24464
rect 51139 24424 51148 24464
rect 51188 24424 52204 24464
rect 52244 24424 54796 24464
rect 54836 24424 54845 24464
rect 58158 24424 58252 24464
rect 58292 24424 58301 24464
rect 61219 24424 61228 24464
rect 61268 24424 61804 24464
rect 61844 24424 64300 24464
rect 64340 24424 64349 24464
rect 66595 24424 66604 24464
rect 66644 24424 66988 24464
rect 67028 24424 67037 24464
rect 67267 24424 67276 24464
rect 67316 24424 67564 24464
rect 67604 24424 68428 24464
rect 68468 24424 68477 24464
rect 69283 24424 69292 24464
rect 69332 24424 71116 24464
rect 71156 24424 71165 24464
rect 75052 24424 75436 24464
rect 75476 24424 75485 24464
rect 41347 24423 41405 24424
rect 58243 24423 58301 24424
rect 67555 24423 67613 24424
rect 69283 24423 69341 24424
rect 66595 24380 66653 24381
rect 44323 24340 44332 24380
rect 44372 24340 44908 24380
rect 44948 24340 46060 24380
rect 46100 24340 59692 24380
rect 59732 24340 59741 24380
rect 61123 24340 61132 24380
rect 61172 24340 62188 24380
rect 62228 24340 62860 24380
rect 62900 24340 62909 24380
rect 66595 24340 66604 24380
rect 66644 24340 71884 24380
rect 71924 24340 71933 24380
rect 75235 24340 75244 24380
rect 75284 24340 75532 24380
rect 75572 24340 75581 24380
rect 66595 24339 66653 24340
rect 50371 24296 50429 24297
rect 69859 24296 69917 24297
rect 75043 24296 75101 24297
rect 37219 24256 37228 24296
rect 37268 24256 38860 24296
rect 38900 24256 39628 24296
rect 39668 24256 39677 24296
rect 49219 24256 49228 24296
rect 49268 24256 50380 24296
rect 50420 24256 62476 24296
rect 62516 24256 62525 24296
rect 62659 24256 62668 24296
rect 62708 24256 63052 24296
rect 63092 24256 63101 24296
rect 65155 24256 65164 24296
rect 65204 24256 67276 24296
rect 67316 24256 67325 24296
rect 68131 24256 68140 24296
rect 68180 24256 69484 24296
rect 69524 24256 69533 24296
rect 69667 24256 69676 24296
rect 69716 24256 69868 24296
rect 69908 24256 69917 24296
rect 74958 24256 75052 24296
rect 75092 24256 75101 24296
rect 50371 24255 50429 24256
rect 69859 24255 69917 24256
rect 75043 24255 75101 24256
rect 40195 24212 40253 24213
rect 56227 24212 56285 24213
rect 56419 24212 56477 24213
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 15103 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 15489 24212
rect 27103 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 27489 24212
rect 36355 24172 36364 24212
rect 36404 24172 38668 24212
rect 38708 24172 38717 24212
rect 39103 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 39489 24212
rect 40195 24172 40204 24212
rect 40244 24172 41836 24212
rect 41876 24172 51148 24212
rect 51188 24172 52012 24212
rect 52052 24172 52061 24212
rect 53260 24172 56236 24212
rect 56276 24172 56285 24212
rect 56334 24172 56428 24212
rect 56468 24172 56477 24212
rect 40195 24171 40253 24172
rect 0 24128 80 24148
rect 53260 24128 53300 24172
rect 56227 24171 56285 24172
rect 56419 24171 56477 24172
rect 56611 24212 56669 24213
rect 64003 24212 64061 24213
rect 68707 24212 68765 24213
rect 56611 24172 56620 24212
rect 56660 24172 57620 24212
rect 57859 24172 57868 24212
rect 57908 24172 59020 24212
rect 59060 24172 63628 24212
rect 63668 24172 63677 24212
rect 64003 24172 64012 24212
rect 64052 24172 67948 24212
rect 67988 24172 67997 24212
rect 68622 24172 68716 24212
rect 68756 24172 68765 24212
rect 56611 24171 56669 24172
rect 57580 24128 57620 24172
rect 64003 24171 64061 24172
rect 68707 24171 68765 24172
rect 62659 24128 62717 24129
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 37027 24088 37036 24128
rect 37076 24088 37900 24128
rect 37940 24088 38476 24128
rect 38516 24088 38525 24128
rect 41443 24088 41452 24128
rect 41492 24088 41644 24128
rect 41684 24088 41693 24128
rect 48547 24088 48556 24128
rect 48596 24088 49324 24128
rect 49364 24088 49373 24128
rect 50659 24088 50668 24128
rect 50708 24088 50956 24128
rect 50996 24088 51005 24128
rect 51235 24088 51244 24128
rect 51284 24088 53300 24128
rect 54307 24088 54316 24128
rect 54356 24088 55084 24128
rect 55124 24088 56524 24128
rect 56564 24088 56573 24128
rect 57580 24088 61804 24128
rect 61844 24088 61853 24128
rect 62083 24088 62092 24128
rect 62132 24088 62668 24128
rect 62708 24088 62717 24128
rect 62851 24088 62860 24128
rect 62900 24088 67564 24128
rect 67604 24088 67613 24128
rect 71203 24088 71212 24128
rect 71252 24088 71692 24128
rect 71732 24088 71741 24128
rect 75811 24088 75820 24128
rect 75860 24088 76012 24128
rect 76052 24088 76061 24128
rect 0 24068 80 24088
rect 62659 24087 62717 24088
rect 53059 24044 53117 24045
rect 64003 24044 64061 24045
rect 38083 24004 38092 24044
rect 38132 24004 38668 24044
rect 38708 24004 38717 24044
rect 41251 24004 41260 24044
rect 41300 24004 41740 24044
rect 41780 24004 41789 24044
rect 50563 24004 50572 24044
rect 50612 24004 51340 24044
rect 51380 24004 51628 24044
rect 51668 24004 51677 24044
rect 52974 24004 53068 24044
rect 53108 24004 53117 24044
rect 54211 24004 54220 24044
rect 54260 24004 54988 24044
rect 55028 24004 63148 24044
rect 63188 24004 63197 24044
rect 63918 24004 64012 24044
rect 64052 24004 64061 24044
rect 67171 24004 67180 24044
rect 67220 24004 68812 24044
rect 68852 24004 72076 24044
rect 72116 24004 72125 24044
rect 73420 24004 76780 24044
rect 76820 24004 77452 24044
rect 77492 24004 77501 24044
rect 53059 24003 53117 24004
rect 64003 24003 64061 24004
rect 52771 23960 52829 23961
rect 55651 23960 55709 23961
rect 37603 23920 37612 23960
rect 37652 23920 37996 23960
rect 38036 23920 38045 23960
rect 38851 23920 38860 23960
rect 38900 23920 40876 23960
rect 40916 23920 40925 23960
rect 41059 23920 41068 23960
rect 41108 23920 43084 23960
rect 43124 23920 43133 23960
rect 44131 23920 44140 23960
rect 44180 23920 44220 23960
rect 49315 23920 49324 23960
rect 49364 23920 51244 23960
rect 51284 23920 51293 23960
rect 51724 23920 52780 23960
rect 52820 23920 52829 23960
rect 55566 23920 55660 23960
rect 55700 23920 55709 23960
rect 56803 23920 56812 23960
rect 56852 23920 57772 23960
rect 57812 23920 63532 23960
rect 63572 23920 63581 23960
rect 63628 23920 65452 23960
rect 65492 23920 65501 23960
rect 66019 23920 66028 23960
rect 66068 23920 71980 23960
rect 72020 23920 72652 23960
rect 72692 23920 72701 23960
rect 44140 23876 44180 23920
rect 51724 23876 51764 23920
rect 52771 23919 52829 23920
rect 55651 23919 55709 23920
rect 53155 23876 53213 23877
rect 63628 23876 63668 23920
rect 73420 23876 73460 24004
rect 76675 23920 76684 23960
rect 76724 23920 77260 23960
rect 77300 23920 78988 23960
rect 79028 23920 79037 23960
rect 1987 23836 1996 23876
rect 2036 23836 2188 23876
rect 2228 23836 13708 23876
rect 13748 23836 13757 23876
rect 38083 23836 38092 23876
rect 38132 23836 38284 23876
rect 38324 23836 39244 23876
rect 39284 23836 39293 23876
rect 40963 23836 40972 23876
rect 41012 23836 42700 23876
rect 42740 23836 42749 23876
rect 42796 23836 43468 23876
rect 43508 23836 44428 23876
rect 44468 23836 44477 23876
rect 47107 23836 47116 23876
rect 47156 23836 51764 23876
rect 52483 23836 52492 23876
rect 52532 23836 53164 23876
rect 53204 23836 58252 23876
rect 58292 23836 58301 23876
rect 59587 23836 59596 23876
rect 59636 23836 59884 23876
rect 59924 23836 61228 23876
rect 61268 23836 61277 23876
rect 61987 23836 61996 23876
rect 62036 23836 62668 23876
rect 62708 23836 62717 23876
rect 62851 23836 62860 23876
rect 62900 23836 63668 23876
rect 64291 23836 64300 23876
rect 64340 23836 65932 23876
rect 65972 23836 65981 23876
rect 68899 23836 68908 23876
rect 68948 23836 69388 23876
rect 69428 23836 70060 23876
rect 70100 23836 71500 23876
rect 71540 23836 72172 23876
rect 72212 23836 73460 23876
rect 42796 23792 42836 23836
rect 53155 23835 53213 23836
rect 48739 23792 48797 23793
rect 50755 23792 50813 23793
rect 53827 23792 53885 23793
rect 68803 23792 68861 23793
rect 75139 23792 75197 23793
rect 78979 23792 79037 23793
rect 28771 23752 28780 23792
rect 28820 23752 41452 23792
rect 41492 23752 41501 23792
rect 42787 23752 42796 23792
rect 42836 23752 42845 23792
rect 42979 23752 42988 23792
rect 43028 23752 43276 23792
rect 43316 23752 43325 23792
rect 43555 23752 43564 23792
rect 43604 23752 44140 23792
rect 44180 23752 44189 23792
rect 46243 23752 46252 23792
rect 46292 23752 47308 23792
rect 47348 23752 47357 23792
rect 47491 23752 47500 23792
rect 47540 23752 48748 23792
rect 48788 23752 48797 23792
rect 50467 23752 50476 23792
rect 50516 23752 50764 23792
rect 50804 23752 50813 23792
rect 53155 23752 53164 23792
rect 53204 23752 53836 23792
rect 53876 23752 53885 23792
rect 54019 23752 54028 23792
rect 54068 23752 54220 23792
rect 54260 23752 54269 23792
rect 54787 23752 54796 23792
rect 54836 23752 56908 23792
rect 56948 23752 56957 23792
rect 57283 23752 57292 23792
rect 57332 23752 57868 23792
rect 57908 23752 57917 23792
rect 59107 23752 59116 23792
rect 59156 23752 59404 23792
rect 59444 23752 59453 23792
rect 59971 23752 59980 23792
rect 60020 23752 60364 23792
rect 60404 23752 60413 23792
rect 61123 23752 61132 23792
rect 61172 23752 62572 23792
rect 62612 23752 63380 23792
rect 64387 23752 64396 23792
rect 64436 23752 64780 23792
rect 64820 23752 65740 23792
rect 65780 23752 65789 23792
rect 68718 23752 68812 23792
rect 68852 23752 68861 23792
rect 71395 23752 71404 23792
rect 71444 23752 72748 23792
rect 72788 23752 73460 23792
rect 75054 23752 75148 23792
rect 75188 23752 75197 23792
rect 78894 23752 78988 23792
rect 79028 23752 79037 23792
rect 48739 23751 48797 23752
rect 50755 23751 50813 23752
rect 53827 23751 53885 23752
rect 50371 23708 50429 23709
rect 35587 23668 35596 23708
rect 35636 23668 36364 23708
rect 36404 23668 36413 23708
rect 38467 23668 38476 23708
rect 38516 23668 38956 23708
rect 38996 23668 40108 23708
rect 40148 23668 40157 23708
rect 50371 23668 50380 23708
rect 50420 23668 55564 23708
rect 55604 23668 56140 23708
rect 56180 23668 56189 23708
rect 56515 23668 56524 23708
rect 56564 23668 63244 23708
rect 63284 23668 63293 23708
rect 50371 23667 50429 23668
rect 63340 23624 63380 23752
rect 68803 23751 68861 23752
rect 63907 23708 63965 23709
rect 63822 23668 63916 23708
rect 63956 23668 64436 23708
rect 70147 23668 70156 23708
rect 70196 23668 71596 23708
rect 71636 23668 72460 23708
rect 72500 23668 73228 23708
rect 73268 23668 73277 23708
rect 63907 23667 63965 23668
rect 64396 23624 64436 23668
rect 69091 23624 69149 23625
rect 73420 23624 73460 23752
rect 75139 23751 75197 23752
rect 78979 23751 79037 23752
rect 74179 23668 74188 23708
rect 74228 23668 75436 23708
rect 75476 23668 75485 23708
rect 74851 23624 74909 23625
rect 77347 23624 77405 23625
rect 36739 23584 36748 23624
rect 36788 23584 37324 23624
rect 37364 23584 38764 23624
rect 38804 23584 39436 23624
rect 39476 23584 39485 23624
rect 41059 23584 41068 23624
rect 41108 23584 41356 23624
rect 41396 23584 41405 23624
rect 42883 23584 42892 23624
rect 42932 23584 43852 23624
rect 43892 23584 43901 23624
rect 44035 23584 44044 23624
rect 44084 23584 45004 23624
rect 45044 23584 59540 23624
rect 59587 23584 59596 23624
rect 59636 23584 60268 23624
rect 60308 23584 60317 23624
rect 61795 23584 61804 23624
rect 61844 23584 62380 23624
rect 62420 23584 62860 23624
rect 62900 23584 62909 23624
rect 63340 23584 64300 23624
rect 64340 23584 64349 23624
rect 64396 23584 68044 23624
rect 68084 23584 68093 23624
rect 69006 23584 69100 23624
rect 69140 23584 69149 23624
rect 69283 23584 69292 23624
rect 69332 23584 72364 23624
rect 72404 23584 73132 23624
rect 73172 23584 73181 23624
rect 73420 23584 73516 23624
rect 73556 23584 73565 23624
rect 74766 23584 74860 23624
rect 74900 23584 74909 23624
rect 76099 23584 76108 23624
rect 76148 23584 76492 23624
rect 76532 23584 76541 23624
rect 76867 23584 76876 23624
rect 76916 23584 77068 23624
rect 77108 23584 77117 23624
rect 77251 23584 77260 23624
rect 77300 23584 77356 23624
rect 77396 23584 77405 23624
rect 78787 23584 78796 23624
rect 78836 23584 79084 23624
rect 79124 23584 79564 23624
rect 79604 23584 79613 23624
rect 43363 23540 43421 23541
rect 42691 23500 42700 23540
rect 42740 23500 43372 23540
rect 43412 23500 44236 23540
rect 44276 23500 44285 23540
rect 49411 23500 49420 23540
rect 49460 23500 50380 23540
rect 50420 23500 50429 23540
rect 51907 23500 51916 23540
rect 51956 23500 54124 23540
rect 54164 23500 57196 23540
rect 57236 23500 57245 23540
rect 43363 23499 43421 23500
rect 59500 23456 59540 23584
rect 69091 23583 69149 23584
rect 74851 23583 74909 23584
rect 77347 23583 77405 23584
rect 60739 23540 60797 23541
rect 71299 23540 71357 23541
rect 76195 23540 76253 23541
rect 60739 23500 60748 23540
rect 60788 23500 63340 23540
rect 63380 23500 63389 23540
rect 67843 23500 67852 23540
rect 67892 23500 69964 23540
rect 70004 23500 70013 23540
rect 71214 23500 71308 23540
rect 71348 23500 71357 23540
rect 72067 23500 72076 23540
rect 72116 23500 72844 23540
rect 72884 23500 72893 23540
rect 73795 23500 73804 23540
rect 73844 23500 74188 23540
rect 74228 23500 74237 23540
rect 74563 23500 74572 23540
rect 74612 23500 75148 23540
rect 75188 23500 75197 23540
rect 76195 23500 76204 23540
rect 76244 23500 76396 23540
rect 76436 23500 76445 23540
rect 60739 23499 60797 23500
rect 71299 23499 71357 23500
rect 76195 23499 76253 23500
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 16343 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 16729 23456
rect 28343 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 28729 23456
rect 36739 23416 36748 23456
rect 36788 23416 37036 23456
rect 37076 23416 37085 23456
rect 40343 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 40729 23456
rect 48355 23416 48364 23456
rect 48404 23416 48652 23456
rect 48692 23416 48844 23456
rect 48884 23416 57524 23456
rect 59491 23416 59500 23456
rect 59540 23416 59549 23456
rect 60355 23416 60364 23456
rect 60404 23416 61900 23456
rect 61940 23416 64012 23456
rect 64052 23416 64061 23456
rect 65731 23416 65740 23456
rect 65780 23416 72460 23456
rect 72500 23416 72509 23456
rect 52771 23372 52829 23373
rect 57484 23372 57524 23416
rect 32035 23332 32044 23372
rect 32084 23332 35884 23372
rect 35924 23332 37804 23372
rect 37844 23332 37853 23372
rect 40771 23332 40780 23372
rect 40820 23332 41644 23372
rect 41684 23332 41693 23372
rect 42412 23332 43084 23372
rect 43124 23332 43133 23372
rect 49891 23332 49900 23372
rect 49940 23332 50860 23372
rect 50900 23332 50909 23372
rect 52003 23332 52012 23372
rect 52052 23332 52492 23372
rect 52532 23332 52541 23372
rect 52771 23332 52780 23372
rect 52820 23332 54028 23372
rect 54068 23332 54077 23372
rect 56323 23332 56332 23372
rect 56372 23332 57236 23372
rect 57484 23332 61612 23372
rect 61652 23332 61661 23372
rect 62947 23332 62956 23372
rect 62996 23332 64876 23372
rect 64916 23332 72364 23372
rect 72404 23332 72413 23372
rect 76291 23332 76300 23372
rect 76340 23332 77164 23372
rect 77204 23332 79084 23372
rect 79124 23332 79133 23372
rect 0 23288 80 23308
rect 39811 23288 39869 23289
rect 42412 23288 42452 23332
rect 52771 23331 52829 23332
rect 57196 23288 57236 23332
rect 57859 23288 57917 23289
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 931 23248 940 23288
rect 980 23248 35980 23288
rect 36020 23248 36029 23288
rect 36931 23248 36940 23288
rect 36980 23248 37516 23288
rect 37556 23248 39820 23288
rect 39860 23248 39869 23288
rect 41155 23248 41164 23288
rect 41204 23248 42412 23288
rect 42452 23248 42461 23288
rect 42787 23248 42796 23288
rect 42836 23248 42845 23288
rect 42979 23248 42988 23288
rect 43028 23248 57100 23288
rect 57140 23248 57149 23288
rect 57196 23248 57868 23288
rect 57908 23248 57917 23288
rect 58243 23248 58252 23288
rect 58292 23248 61268 23288
rect 62659 23248 62668 23288
rect 62708 23248 63436 23288
rect 63476 23248 64492 23288
rect 64532 23248 64541 23288
rect 67459 23248 67468 23288
rect 67508 23248 70060 23288
rect 70100 23248 70109 23288
rect 0 23228 80 23248
rect 39811 23247 39869 23248
rect 42796 23204 42836 23248
rect 57859 23247 57917 23248
rect 61228 23204 61268 23248
rect 69667 23204 69725 23205
rect 75619 23204 75677 23205
rect 35299 23164 35308 23204
rect 35348 23164 35788 23204
rect 35828 23164 37228 23204
rect 37268 23164 37277 23204
rect 37699 23164 37708 23204
rect 37748 23164 41780 23204
rect 42796 23164 43412 23204
rect 46051 23164 46060 23204
rect 46100 23164 47116 23204
rect 47156 23164 47165 23204
rect 51715 23164 51724 23204
rect 51764 23164 52396 23204
rect 52436 23164 61132 23204
rect 61172 23164 61181 23204
rect 61228 23164 66028 23204
rect 66068 23164 66077 23204
rect 67651 23164 67660 23204
rect 67700 23164 67709 23204
rect 69283 23164 69292 23204
rect 69332 23164 69676 23204
rect 69716 23164 69725 23204
rect 73315 23164 73324 23204
rect 73364 23164 73612 23204
rect 73652 23164 73661 23204
rect 75619 23164 75628 23204
rect 75668 23164 76300 23204
rect 76340 23164 76349 23204
rect 78691 23164 78700 23204
rect 78740 23164 78836 23204
rect 41740 23120 41780 23164
rect 835 23080 844 23120
rect 884 23080 1516 23120
rect 1556 23080 1565 23120
rect 33763 23080 33772 23120
rect 33812 23080 35692 23120
rect 35732 23080 37036 23120
rect 37076 23080 37085 23120
rect 40003 23080 40012 23120
rect 40052 23080 41644 23120
rect 41684 23080 41693 23120
rect 41740 23080 42988 23120
rect 43028 23080 43037 23120
rect 43084 23080 43180 23120
rect 43220 23080 43248 23120
rect 1603 22996 1612 23036
rect 1652 22996 3628 23036
rect 3668 22996 7084 23036
rect 7124 22996 7133 23036
rect 40963 22996 40972 23036
rect 41012 22996 42508 23036
rect 42548 22996 42796 23036
rect 42836 22996 42845 23036
rect 43084 22952 43124 23080
rect 43372 22952 43412 23164
rect 51523 23120 51581 23121
rect 45859 23080 45868 23120
rect 45908 23080 46828 23120
rect 46868 23080 46877 23120
rect 48931 23080 48940 23120
rect 48980 23080 49132 23120
rect 49172 23080 49181 23120
rect 51438 23080 51532 23120
rect 51572 23080 51581 23120
rect 51523 23079 51581 23080
rect 51811 23120 51869 23121
rect 55171 23120 55229 23121
rect 62659 23120 62717 23121
rect 67660 23120 67700 23164
rect 69667 23163 69725 23164
rect 75619 23163 75677 23164
rect 51811 23080 51820 23120
rect 51860 23080 52108 23120
rect 52148 23080 52157 23120
rect 52684 23080 54895 23120
rect 51811 23079 51869 23080
rect 46531 22996 46540 23036
rect 46580 22996 50668 23036
rect 50708 22996 50717 23036
rect 51235 22996 51244 23036
rect 51284 22996 52588 23036
rect 52628 22996 52637 23036
rect 52684 22952 52724 23080
rect 53443 23036 53501 23037
rect 53059 22996 53068 23036
rect 53108 22996 53396 23036
rect 53356 22952 53396 22996
rect 53443 22996 53452 23036
rect 53492 22996 53945 23036
rect 53985 22996 53994 23036
rect 53443 22995 53501 22996
rect 54691 22952 54749 22953
rect 42403 22912 42412 22952
rect 42452 22912 42892 22952
rect 42932 22912 42941 22952
rect 43075 22912 43084 22952
rect 43124 22912 43133 22952
rect 43363 22912 43372 22952
rect 43412 22912 43421 22952
rect 51532 22912 52724 22952
rect 53164 22912 53260 22952
rect 53300 22912 53309 22952
rect 53356 22912 54455 22952
rect 54495 22912 54504 22952
rect 54650 22912 54700 22952
rect 54740 22912 54745 22952
rect 54785 22912 54794 22952
rect 51532 22868 51572 22912
rect 53164 22868 53204 22912
rect 54691 22911 54749 22912
rect 42499 22828 42508 22868
rect 42548 22828 43180 22868
rect 43220 22828 43229 22868
rect 50947 22828 50956 22868
rect 50996 22828 51340 22868
rect 51380 22828 51389 22868
rect 51523 22828 51532 22868
rect 51572 22828 51581 22868
rect 52579 22828 52588 22868
rect 52628 22828 53204 22868
rect 53251 22868 53309 22869
rect 54855 22868 54895 23080
rect 55171 23080 55180 23120
rect 55220 23080 55260 23120
rect 55651 23080 55660 23120
rect 55700 23080 56180 23120
rect 59011 23080 59020 23120
rect 59060 23080 59979 23120
rect 60019 23080 60028 23120
rect 62659 23080 62668 23120
rect 62708 23080 67700 23120
rect 55171 23079 55229 23080
rect 55180 23036 55220 23079
rect 56140 23036 56180 23080
rect 62659 23079 62717 23080
rect 78796 23060 78836 23164
rect 57091 23036 57149 23037
rect 62851 23036 62909 23037
rect 74947 23036 75005 23037
rect 78019 23036 78077 23037
rect 55180 22996 55255 23036
rect 55295 22996 55304 23036
rect 55939 22996 55948 23036
rect 55988 22996 55997 23036
rect 56140 22996 56455 23036
rect 56495 22996 56504 23036
rect 57091 22996 57100 23036
rect 57140 22996 60855 23036
rect 60895 22996 60904 23036
rect 62851 22996 62860 23036
rect 62900 22996 65255 23036
rect 65295 22996 65304 23036
rect 65347 22996 65356 23036
rect 65396 22996 68345 23036
rect 68385 22996 68394 23036
rect 74083 22996 74092 23036
rect 74132 22996 74345 23036
rect 74385 22996 74394 23036
rect 74947 22996 74956 23036
rect 74996 22996 75255 23036
rect 75295 22996 75304 23036
rect 77536 22996 77545 23036
rect 77585 22996 78028 23036
rect 78068 22996 78077 23036
rect 78700 23036 78836 23060
rect 78700 22996 79655 23036
rect 79695 22996 79704 23036
rect 55171 22952 55229 22953
rect 55747 22952 55805 22953
rect 55136 22912 55145 22952
rect 55220 22912 55280 22952
rect 55662 22912 55756 22952
rect 55796 22912 55805 22952
rect 55948 22952 55988 22996
rect 57091 22995 57149 22996
rect 62851 22995 62909 22996
rect 74947 22995 75005 22996
rect 78019 22995 78077 22996
rect 57955 22952 58013 22953
rect 59011 22952 59069 22953
rect 64771 22952 64829 22953
rect 66307 22952 66365 22953
rect 55948 22912 56745 22952
rect 56785 22912 56794 22952
rect 57955 22912 57964 22952
rect 58004 22912 58345 22952
rect 58385 22912 58394 22952
rect 59011 22912 59020 22952
rect 59060 22912 59945 22952
rect 59985 22912 59994 22952
rect 60259 22912 60268 22952
rect 60308 22912 63945 22952
rect 63985 22912 63994 22952
rect 64771 22912 64780 22952
rect 64820 22912 65945 22952
rect 65985 22912 65994 22952
rect 66307 22912 66316 22952
rect 66356 22912 66745 22952
rect 66785 22912 66794 22952
rect 78211 22912 78220 22952
rect 78260 22912 78892 22952
rect 78932 22912 78941 22952
rect 55171 22911 55229 22912
rect 55747 22911 55805 22912
rect 57955 22911 58013 22912
rect 59011 22911 59069 22912
rect 64771 22911 64829 22912
rect 66307 22911 66365 22912
rect 56227 22868 56285 22869
rect 57763 22868 57821 22869
rect 60739 22868 60797 22869
rect 53251 22828 53260 22868
rect 53300 22828 54345 22868
rect 54385 22828 54394 22868
rect 54855 22828 55655 22868
rect 55695 22828 55704 22868
rect 56227 22828 56236 22868
rect 56276 22828 57545 22868
rect 57585 22828 57594 22868
rect 57763 22828 57772 22868
rect 57812 22828 57945 22868
rect 57985 22828 57994 22868
rect 60654 22828 60748 22868
rect 60788 22828 60797 22868
rect 53251 22827 53309 22828
rect 56227 22827 56285 22828
rect 57763 22827 57821 22828
rect 60739 22827 60797 22828
rect 66211 22868 66269 22869
rect 66595 22868 66653 22869
rect 71011 22868 71069 22869
rect 66211 22828 66220 22868
rect 66260 22828 66455 22868
rect 66495 22828 66504 22868
rect 66595 22828 66604 22868
rect 66644 22828 66855 22868
rect 66895 22828 66904 22868
rect 71011 22828 71020 22868
rect 71060 22828 71545 22868
rect 71585 22828 71594 22868
rect 66211 22827 66269 22828
rect 66595 22827 66653 22828
rect 71011 22827 71069 22828
rect 54883 22784 54941 22785
rect 55555 22784 55613 22785
rect 55843 22784 55901 22785
rect 57667 22784 57725 22785
rect 59107 22784 59165 22785
rect 60451 22784 60509 22785
rect 61891 22784 61949 22785
rect 66499 22784 66557 22785
rect 71875 22784 71933 22785
rect 76867 22784 76925 22785
rect 77155 22784 77213 22785
rect 77923 22784 77981 22785
rect 52675 22744 52684 22784
rect 52724 22744 53545 22784
rect 53585 22744 53594 22784
rect 54846 22744 54855 22784
rect 54932 22744 54990 22784
rect 55536 22744 55545 22784
rect 55604 22744 55680 22784
rect 55747 22744 55756 22784
rect 55796 22744 55852 22784
rect 55892 22744 55901 22784
rect 56131 22744 56140 22784
rect 56180 22744 56855 22784
rect 56895 22744 56904 22784
rect 57581 22744 57655 22784
rect 57716 22744 57725 22784
rect 59050 22744 59116 22784
rect 59185 22744 59194 22784
rect 60451 22744 60460 22784
rect 60500 22744 61545 22784
rect 61585 22744 61594 22784
rect 61850 22744 61900 22784
rect 61940 22744 61945 22784
rect 61985 22744 61994 22784
rect 66336 22744 66345 22784
rect 66385 22744 66508 22784
rect 66548 22744 66557 22784
rect 70531 22744 70540 22784
rect 70580 22744 70855 22784
rect 70895 22744 70904 22784
rect 71646 22744 71655 22784
rect 71695 22744 71788 22784
rect 71828 22744 71884 22784
rect 71924 22744 71933 22784
rect 73411 22744 73420 22784
rect 73460 22744 73655 22784
rect 73695 22744 73704 22784
rect 73795 22744 73804 22784
rect 73844 22744 74055 22784
rect 74095 22744 74104 22784
rect 74179 22744 74188 22784
rect 74228 22744 74745 22784
rect 74785 22744 74794 22784
rect 75811 22744 75820 22784
rect 75860 22744 76055 22784
rect 76095 22744 76104 22784
rect 76781 22744 76855 22784
rect 76916 22744 76925 22784
rect 77069 22744 77145 22784
rect 77204 22744 77213 22784
rect 77850 22744 77932 22784
rect 77985 22744 77994 22784
rect 78046 22744 78055 22784
rect 78095 22744 78604 22784
rect 78644 22744 78653 22784
rect 54883 22743 54941 22744
rect 55555 22743 55613 22744
rect 55843 22743 55901 22744
rect 57667 22743 57725 22744
rect 59107 22743 59165 22744
rect 60451 22743 60509 22744
rect 61891 22743 61949 22744
rect 66499 22743 66557 22744
rect 71875 22743 71933 22744
rect 76867 22743 76925 22744
rect 77155 22743 77213 22744
rect 77923 22743 77981 22744
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 15103 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 15489 22700
rect 27103 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 27489 22700
rect 39103 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 39489 22700
rect 41251 22576 41260 22616
rect 41300 22576 41548 22616
rect 41588 22576 41597 22616
rect 49795 22576 49804 22616
rect 49844 22576 49853 22616
rect 43459 22532 43517 22533
rect 31075 22492 31084 22532
rect 31124 22492 36748 22532
rect 36788 22492 36797 22532
rect 43374 22492 43468 22532
rect 43508 22492 43517 22532
rect 43459 22491 43517 22492
rect 0 22448 80 22468
rect 49804 22448 49844 22576
rect 52387 22532 52445 22533
rect 52302 22492 52396 22532
rect 52436 22492 52445 22532
rect 52387 22491 52445 22492
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 35971 22408 35980 22448
rect 36020 22408 40012 22448
rect 40052 22408 40061 22448
rect 41539 22408 41548 22448
rect 41588 22408 42892 22448
rect 42932 22408 42941 22448
rect 49315 22408 49324 22448
rect 49364 22408 50092 22448
rect 50132 22408 50141 22448
rect 0 22388 80 22408
rect 32227 22324 32236 22364
rect 32276 22324 33964 22364
rect 34004 22324 34013 22364
rect 37219 22324 37228 22364
rect 37268 22324 37420 22364
rect 37460 22324 37469 22364
rect 46051 22324 46060 22364
rect 46100 22324 46540 22364
rect 46580 22324 46589 22364
rect 30115 22240 30124 22280
rect 30164 22240 31468 22280
rect 31508 22240 31517 22280
rect 36259 22240 36268 22280
rect 36308 22240 37132 22280
rect 37172 22240 37181 22280
rect 40867 22240 40876 22280
rect 40916 22240 41452 22280
rect 41492 22240 41501 22280
rect 41827 22240 41836 22280
rect 41876 22240 42508 22280
rect 42548 22240 42557 22280
rect 43363 22240 43372 22280
rect 43412 22240 45292 22280
rect 45332 22240 45341 22280
rect 47203 22240 47212 22280
rect 47252 22240 48844 22280
rect 48884 22240 48893 22280
rect 49603 22240 49612 22280
rect 49652 22240 50476 22280
rect 50516 22240 50525 22280
rect 40099 22196 40157 22197
rect 42403 22196 42461 22197
rect 51619 22196 51677 22197
rect 35491 22156 35500 22196
rect 35540 22156 40108 22196
rect 40148 22156 40157 22196
rect 42318 22156 42412 22196
rect 42452 22156 42461 22196
rect 46531 22156 46540 22196
rect 46580 22156 47404 22196
rect 47444 22156 47453 22196
rect 47500 22156 51628 22196
rect 51668 22156 51677 22196
rect 40099 22155 40157 22156
rect 42403 22155 42461 22156
rect 38851 22112 38909 22113
rect 37027 22072 37036 22112
rect 37076 22072 37420 22112
rect 37460 22072 38860 22112
rect 38900 22072 38909 22112
rect 42307 22072 42316 22112
rect 42356 22072 42604 22112
rect 42644 22072 42653 22112
rect 43189 22072 43198 22112
rect 43238 22072 43852 22112
rect 43892 22072 45868 22112
rect 45908 22072 45917 22112
rect 38851 22071 38909 22072
rect 47500 22028 47540 22156
rect 51619 22155 51677 22156
rect 49699 22072 49708 22112
rect 49748 22072 50956 22112
rect 50996 22072 51005 22112
rect 33187 21988 33196 22028
rect 33236 21988 33484 22028
rect 33524 21988 35692 22028
rect 35732 21988 35741 22028
rect 36739 21988 36748 22028
rect 36788 21988 37612 22028
rect 37652 21988 37661 22028
rect 39427 21988 39436 22028
rect 39476 21988 47540 22028
rect 37612 21944 37652 21988
rect 50764 21944 50804 22072
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 16343 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 16729 21944
rect 28343 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 28729 21944
rect 37612 21904 39820 21944
rect 39860 21904 39869 21944
rect 40343 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 40729 21944
rect 43843 21904 43852 21944
rect 43892 21904 45004 21944
rect 45044 21904 45053 21944
rect 50755 21904 50764 21944
rect 50804 21904 50813 21944
rect 47011 21820 47020 21860
rect 47060 21820 48460 21860
rect 48500 21820 48509 21860
rect 42115 21736 42124 21776
rect 42164 21736 42604 21776
rect 42644 21736 42653 21776
rect 42883 21736 42892 21776
rect 42932 21736 44236 21776
rect 44276 21736 44285 21776
rect 45955 21736 45964 21776
rect 46004 21736 46156 21776
rect 46196 21736 46924 21776
rect 46964 21736 46973 21776
rect 50572 21736 51916 21776
rect 51956 21736 51965 21776
rect 40099 21692 40157 21693
rect 30883 21652 30892 21692
rect 30932 21652 31468 21692
rect 31508 21652 31517 21692
rect 31747 21652 31756 21692
rect 31796 21652 36940 21692
rect 36980 21652 36989 21692
rect 37219 21652 37228 21692
rect 37268 21652 37420 21692
rect 37460 21652 37469 21692
rect 40099 21652 40108 21692
rect 40148 21652 40300 21692
rect 40340 21652 40349 21692
rect 41731 21652 41740 21692
rect 41780 21652 42260 21692
rect 40099 21651 40157 21652
rect 0 21608 80 21628
rect 3907 21608 3965 21609
rect 4579 21608 4637 21609
rect 7363 21608 7421 21609
rect 42220 21608 42260 21652
rect 46924 21652 47212 21692
rect 47252 21652 47261 21692
rect 46924 21608 46964 21652
rect 50572 21608 50612 21736
rect 99920 21692 100000 21726
rect 50659 21652 50668 21692
rect 50708 21652 52396 21692
rect 52436 21652 52445 21692
rect 99888 21652 100000 21692
rect 51244 21608 51284 21652
rect 52195 21608 52253 21609
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 3822 21568 3916 21608
rect 3956 21568 3965 21608
rect 4494 21568 4588 21608
rect 4628 21568 4637 21608
rect 7278 21568 7372 21608
rect 7412 21568 7660 21608
rect 7700 21568 7709 21608
rect 7939 21568 7948 21608
rect 7988 21568 9004 21608
rect 9044 21568 10540 21608
rect 10580 21568 12460 21608
rect 12500 21568 12509 21608
rect 31267 21568 31276 21608
rect 31316 21568 31852 21608
rect 31892 21568 35308 21608
rect 35348 21568 35500 21608
rect 35540 21568 35549 21608
rect 37027 21568 37036 21608
rect 37076 21568 37708 21608
rect 37748 21568 37757 21608
rect 40771 21568 40780 21608
rect 40820 21568 40972 21608
rect 41012 21568 41021 21608
rect 42211 21568 42220 21608
rect 42260 21568 42269 21608
rect 42403 21568 42412 21608
rect 42452 21568 42796 21608
rect 42836 21568 42845 21608
rect 43075 21568 43084 21608
rect 43124 21568 43660 21608
rect 43700 21568 43709 21608
rect 46915 21568 46924 21608
rect 46964 21568 46973 21608
rect 50275 21568 50284 21608
rect 50324 21568 50572 21608
rect 50612 21568 50621 21608
rect 51235 21568 51244 21608
rect 51284 21568 51293 21608
rect 52110 21568 52204 21608
rect 52244 21568 52253 21608
rect 52483 21568 52492 21608
rect 52532 21568 53068 21608
rect 53108 21568 53117 21608
rect 99920 21586 100000 21652
rect 0 21548 80 21568
rect 3907 21567 3965 21568
rect 4579 21567 4637 21568
rect 7363 21567 7421 21568
rect 52195 21567 52253 21568
rect 43459 21524 43517 21525
rect 51811 21524 51869 21525
rect 1027 21484 1036 21524
rect 1076 21484 3340 21524
rect 3380 21484 3389 21524
rect 4003 21484 4012 21524
rect 4052 21484 4492 21524
rect 4532 21484 5068 21524
rect 5108 21484 5117 21524
rect 7180 21484 29740 21524
rect 29780 21484 29789 21524
rect 30499 21484 30508 21524
rect 30548 21484 31756 21524
rect 31796 21484 31805 21524
rect 42316 21484 43468 21524
rect 43508 21484 43517 21524
rect 46435 21484 46444 21524
rect 46484 21484 47500 21524
rect 47540 21484 47549 21524
rect 50179 21484 50188 21524
rect 50228 21484 51148 21524
rect 51188 21484 51820 21524
rect 51860 21484 51869 21524
rect 7180 21440 7220 21484
rect 42316 21440 42356 21484
rect 43459 21483 43517 21484
rect 51811 21483 51869 21484
rect 53059 21440 53117 21441
rect 5923 21400 5932 21440
rect 5972 21400 7220 21440
rect 8131 21400 8140 21440
rect 8180 21400 11596 21440
rect 11636 21400 14284 21440
rect 14324 21400 14333 21440
rect 17260 21400 30124 21440
rect 30164 21400 30173 21440
rect 33100 21400 37900 21440
rect 37940 21400 37949 21440
rect 38275 21400 38284 21440
rect 38324 21400 40108 21440
rect 40148 21400 41260 21440
rect 41300 21400 41309 21440
rect 42307 21400 42316 21440
rect 42356 21400 42365 21440
rect 43180 21400 52588 21440
rect 52628 21400 53068 21440
rect 53108 21400 53117 21440
rect 17260 21356 17300 21400
rect 33100 21356 33140 21400
rect 43180 21356 43220 21400
rect 53059 21399 53117 21400
rect 51619 21356 51677 21357
rect 51907 21356 51965 21357
rect 52963 21356 53021 21357
rect 2755 21316 2764 21356
rect 2804 21316 3532 21356
rect 3572 21316 4108 21356
rect 4148 21316 17300 21356
rect 29923 21316 29932 21356
rect 29972 21316 30412 21356
rect 30452 21316 33140 21356
rect 35779 21316 35788 21356
rect 35828 21316 36556 21356
rect 36596 21316 37132 21356
rect 37172 21316 37181 21356
rect 41155 21316 41164 21356
rect 41204 21316 43220 21356
rect 47395 21316 47404 21356
rect 47444 21316 47692 21356
rect 47732 21316 49516 21356
rect 49556 21316 49565 21356
rect 51534 21316 51628 21356
rect 51668 21316 51677 21356
rect 51822 21316 51916 21356
rect 51956 21316 52972 21356
rect 53012 21316 53021 21356
rect 51619 21315 51677 21316
rect 51907 21315 51965 21316
rect 52963 21315 53021 21316
rect 51715 21272 51773 21273
rect 5347 21232 5356 21272
rect 5396 21232 8140 21272
rect 8180 21232 8189 21272
rect 12931 21232 12940 21272
rect 12980 21232 13612 21272
rect 13652 21232 51724 21272
rect 51764 21232 51820 21272
rect 51860 21232 51869 21272
rect 51715 21231 51773 21232
rect 51619 21188 51677 21189
rect 52675 21188 52733 21189
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 3811 21148 3820 21188
rect 3860 21148 3869 21188
rect 15103 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 15489 21188
rect 27103 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 27489 21188
rect 39103 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 39489 21188
rect 51619 21148 51628 21188
rect 51668 21148 52684 21188
rect 52724 21148 52733 21188
rect 3820 21020 3860 21148
rect 51619 21147 51677 21148
rect 52675 21147 52733 21148
rect 10147 21064 10156 21104
rect 10196 21064 10636 21104
rect 10676 21064 52492 21104
rect 52532 21064 52541 21104
rect 52291 21020 52349 21021
rect 3523 20980 3532 21020
rect 3572 20980 3860 21020
rect 3907 20980 3916 21020
rect 3956 20980 4204 21020
rect 4244 20980 4253 21020
rect 13603 20980 13612 21020
rect 13652 20980 52300 21020
rect 52340 20980 52349 21020
rect 52291 20979 52349 20980
rect 52483 20936 52541 20937
rect 1699 20896 1708 20936
rect 1748 20896 3340 20936
rect 3380 20896 4012 20936
rect 4052 20896 4061 20936
rect 6787 20896 6796 20936
rect 6836 20896 7660 20936
rect 7700 20896 7709 20936
rect 10243 20896 10252 20936
rect 10292 20896 11692 20936
rect 11732 20896 11741 20936
rect 13699 20896 13708 20936
rect 13748 20896 30508 20936
rect 30548 20896 30557 20936
rect 33004 20896 35404 20936
rect 35444 20896 35453 20936
rect 44611 20896 44620 20936
rect 44660 20896 51532 20936
rect 51572 20896 51581 20936
rect 52398 20896 52492 20936
rect 52532 20896 52541 20936
rect 2851 20812 2860 20852
rect 2900 20812 3244 20852
rect 3284 20812 6412 20852
rect 6452 20812 6461 20852
rect 6883 20812 6892 20852
rect 6932 20812 7372 20852
rect 7412 20812 7421 20852
rect 10147 20812 10156 20852
rect 10196 20812 11020 20852
rect 11060 20812 11069 20852
rect 0 20768 80 20788
rect 33004 20768 33044 20896
rect 52483 20895 52541 20896
rect 50563 20852 50621 20853
rect 33955 20812 33964 20852
rect 34004 20812 37420 20852
rect 37460 20812 37469 20852
rect 43843 20812 43852 20852
rect 43892 20812 44524 20852
rect 44564 20812 46060 20852
rect 46100 20812 46109 20852
rect 50478 20812 50572 20852
rect 50612 20812 50621 20852
rect 50563 20811 50621 20812
rect 52099 20768 52157 20769
rect 52771 20768 52829 20769
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 1891 20728 1900 20768
rect 1940 20728 5260 20768
rect 5300 20728 6316 20768
rect 6356 20728 7468 20768
rect 7508 20728 7517 20768
rect 8419 20728 8428 20768
rect 8468 20728 27628 20768
rect 27668 20728 28780 20768
rect 28820 20728 28829 20768
rect 31651 20728 31660 20768
rect 31700 20728 32428 20768
rect 32468 20728 32477 20768
rect 32803 20728 32812 20768
rect 32852 20728 33004 20768
rect 33044 20728 33053 20768
rect 33283 20728 33292 20768
rect 33332 20728 33484 20768
rect 33524 20728 35212 20768
rect 35252 20728 35261 20768
rect 36259 20728 36268 20768
rect 36308 20728 37036 20768
rect 37076 20728 37085 20768
rect 40579 20728 40588 20768
rect 40628 20728 40972 20768
rect 41012 20728 42988 20768
rect 43028 20728 43037 20768
rect 47203 20728 47212 20768
rect 47252 20728 47788 20768
rect 47828 20728 47837 20768
rect 52099 20728 52108 20768
rect 52148 20728 52204 20768
rect 52244 20728 52253 20768
rect 52579 20728 52588 20768
rect 52628 20728 52780 20768
rect 52820 20728 52829 20768
rect 0 20708 80 20728
rect 52099 20727 52157 20728
rect 52771 20727 52829 20728
rect 2755 20644 2764 20684
rect 2804 20644 4396 20684
rect 4436 20644 5356 20684
rect 5396 20644 5405 20684
rect 30307 20644 30316 20684
rect 30356 20644 31372 20684
rect 31412 20644 32948 20684
rect 10915 20600 10973 20601
rect 32908 20600 32948 20644
rect 52291 20600 52349 20601
rect 52579 20600 52637 20601
rect 1507 20560 1516 20600
rect 1556 20560 5932 20600
rect 5972 20560 5981 20600
rect 10830 20560 10924 20600
rect 10964 20560 10973 20600
rect 30499 20560 30508 20600
rect 30548 20560 31852 20600
rect 31892 20560 31901 20600
rect 32227 20560 32236 20600
rect 32276 20560 32812 20600
rect 32852 20560 32861 20600
rect 32908 20560 33676 20600
rect 33716 20560 36172 20600
rect 36212 20560 36748 20600
rect 36788 20560 36797 20600
rect 52206 20560 52300 20600
rect 52340 20560 52588 20600
rect 52628 20560 52637 20600
rect 10915 20559 10973 20560
rect 52291 20559 52349 20560
rect 52579 20559 52637 20560
rect 3715 20476 3724 20516
rect 3764 20476 4012 20516
rect 4052 20476 4061 20516
rect 16099 20476 16108 20516
rect 16148 20476 52108 20516
rect 52148 20476 52157 20516
rect 42787 20432 42845 20433
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 16343 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 16729 20432
rect 28343 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 28729 20432
rect 29635 20392 29644 20432
rect 29684 20392 30892 20432
rect 30932 20392 33388 20432
rect 33428 20392 33437 20432
rect 40343 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 40729 20432
rect 41731 20392 41740 20432
rect 41780 20392 42796 20432
rect 42836 20392 42845 20432
rect 42787 20391 42845 20392
rect 52771 20348 52829 20349
rect 6403 20308 6412 20348
rect 6452 20308 52780 20348
rect 52820 20308 52829 20348
rect 52771 20307 52829 20308
rect 4195 20224 4204 20264
rect 4244 20224 4684 20264
rect 4724 20224 4733 20264
rect 10435 20224 10444 20264
rect 10484 20224 10493 20264
rect 30979 20224 30988 20264
rect 31028 20224 31037 20264
rect 31171 20224 31180 20264
rect 31220 20224 31756 20264
rect 31796 20224 32524 20264
rect 32564 20224 32573 20264
rect 40195 20224 40204 20264
rect 40244 20224 40684 20264
rect 40724 20224 40733 20264
rect 41548 20224 42220 20264
rect 42260 20224 42269 20264
rect 42403 20224 42412 20264
rect 42452 20224 42700 20264
rect 42740 20224 42749 20264
rect 10444 20180 10484 20224
rect 30988 20180 31028 20224
rect 41548 20180 41588 20224
rect 4003 20140 4012 20180
rect 4052 20140 4492 20180
rect 4532 20140 4541 20180
rect 7555 20140 7564 20180
rect 7604 20140 9292 20180
rect 9332 20140 9772 20180
rect 9812 20140 9821 20180
rect 10243 20140 10252 20180
rect 10292 20140 12076 20180
rect 12116 20140 12125 20180
rect 28483 20140 28492 20180
rect 28532 20140 31372 20180
rect 31412 20140 32140 20180
rect 32180 20140 34636 20180
rect 34676 20140 34685 20180
rect 40579 20140 40588 20180
rect 40628 20140 40780 20180
rect 40820 20140 40829 20180
rect 41347 20140 41356 20180
rect 41396 20140 41588 20180
rect 42412 20096 42452 20224
rect 42787 20180 42845 20181
rect 42702 20140 42796 20180
rect 42836 20140 42845 20180
rect 43651 20140 43660 20180
rect 43700 20140 44140 20180
rect 44180 20140 47884 20180
rect 47924 20140 47933 20180
rect 49123 20140 49132 20180
rect 49172 20140 49612 20180
rect 49652 20140 49900 20180
rect 49940 20140 51436 20180
rect 51476 20140 51485 20180
rect 51724 20140 52204 20180
rect 52244 20140 52253 20180
rect 42787 20139 42845 20140
rect 1699 20056 1708 20096
rect 1748 20056 4300 20096
rect 4340 20056 5260 20096
rect 5300 20056 6220 20096
rect 6260 20056 6269 20096
rect 6691 20056 6700 20096
rect 6740 20056 6892 20096
rect 6932 20056 7948 20096
rect 7988 20056 7997 20096
rect 8515 20056 8524 20096
rect 8564 20056 10636 20096
rect 10676 20056 10685 20096
rect 16963 20056 16972 20096
rect 17012 20056 26956 20096
rect 26996 20056 27916 20096
rect 27956 20056 27965 20096
rect 30691 20056 30700 20096
rect 30740 20056 31468 20096
rect 31508 20056 31517 20096
rect 36547 20056 36556 20096
rect 36596 20056 37036 20096
rect 37076 20056 37085 20096
rect 40483 20056 40492 20096
rect 40532 20056 42452 20096
rect 44035 20056 44044 20096
rect 44084 20056 45004 20096
rect 45044 20056 45053 20096
rect 45763 20056 45772 20096
rect 45812 20056 48748 20096
rect 48788 20056 49420 20096
rect 49460 20056 49469 20096
rect 8524 20012 8564 20056
rect 40099 20012 40157 20013
rect 51724 20012 51764 20140
rect 51907 20012 51965 20013
rect 99920 20012 100000 20089
rect 1795 19972 1804 20012
rect 1844 19972 8564 20012
rect 23020 19972 33964 20012
rect 34004 19972 34013 20012
rect 40014 19972 40108 20012
rect 40148 19972 40157 20012
rect 40771 19972 40780 20012
rect 40820 19972 41740 20012
rect 41780 19972 41789 20012
rect 47971 19972 47980 20012
rect 48020 19972 51764 20012
rect 51822 19972 51916 20012
rect 51956 19972 51965 20012
rect 99888 19972 100000 20012
rect 0 19928 80 19948
rect 23020 19928 23060 19972
rect 40099 19971 40157 19972
rect 51907 19971 51965 19972
rect 99920 19949 100000 19972
rect 42403 19928 42461 19929
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 4675 19888 4684 19928
rect 4724 19888 23060 19928
rect 30787 19888 30796 19928
rect 30836 19888 33196 19928
rect 33236 19888 35788 19928
rect 35828 19888 37132 19928
rect 37172 19888 37181 19928
rect 42307 19888 42316 19928
rect 42356 19888 42412 19928
rect 42452 19888 42796 19928
rect 42836 19888 42845 19928
rect 50371 19888 50380 19928
rect 50420 19888 51148 19928
rect 51188 19888 51197 19928
rect 0 19868 80 19888
rect 42403 19887 42461 19888
rect 5059 19804 5068 19844
rect 5108 19804 8140 19844
rect 8180 19804 8428 19844
rect 8468 19804 9964 19844
rect 10004 19804 10828 19844
rect 10868 19804 10877 19844
rect 34531 19804 34540 19844
rect 34580 19804 37516 19844
rect 37556 19804 37565 19844
rect 47011 19676 47069 19677
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 3619 19636 3628 19676
rect 3668 19636 6700 19676
rect 6740 19636 8620 19676
rect 8660 19636 9868 19676
rect 9908 19636 9917 19676
rect 15103 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 15489 19676
rect 27103 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 27489 19676
rect 39103 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 39489 19676
rect 39907 19636 39916 19676
rect 39956 19636 46828 19676
rect 46868 19636 47020 19676
rect 47060 19636 47069 19676
rect 49987 19636 49996 19676
rect 50036 19636 50764 19676
rect 50804 19636 51532 19676
rect 51572 19636 51581 19676
rect 39916 19592 39956 19636
rect 47011 19635 47069 19636
rect 3340 19552 3724 19592
rect 3764 19552 3773 19592
rect 4483 19552 4492 19592
rect 4532 19552 5356 19592
rect 5396 19552 6796 19592
rect 6836 19552 7220 19592
rect 11107 19552 11116 19592
rect 11156 19552 13516 19592
rect 13556 19552 33484 19592
rect 33524 19552 33533 19592
rect 38659 19552 38668 19592
rect 38708 19552 39956 19592
rect 40291 19552 40300 19592
rect 40340 19552 43948 19592
rect 43988 19552 47500 19592
rect 47540 19552 47549 19592
rect 3340 19508 3380 19552
rect 1219 19468 1228 19508
rect 1268 19468 2764 19508
rect 2804 19468 2813 19508
rect 3331 19468 3340 19508
rect 3380 19468 3389 19508
rect 6883 19468 6892 19508
rect 6932 19468 7084 19508
rect 7124 19468 7133 19508
rect 7180 19424 7220 19552
rect 37027 19508 37085 19509
rect 9379 19468 9388 19508
rect 9428 19468 9772 19508
rect 9812 19468 12940 19508
rect 12980 19468 12989 19508
rect 33571 19468 33580 19508
rect 33620 19468 34252 19508
rect 34292 19468 34301 19508
rect 36643 19468 36652 19508
rect 36692 19468 37036 19508
rect 37076 19468 37612 19508
rect 37652 19468 37661 19508
rect 38851 19468 38860 19508
rect 38900 19468 40396 19508
rect 40436 19468 40972 19508
rect 41012 19468 43372 19508
rect 43412 19468 43421 19508
rect 46531 19468 46540 19508
rect 46580 19468 47212 19508
rect 47252 19468 47261 19508
rect 37027 19467 37085 19468
rect 7180 19384 10252 19424
rect 10292 19384 10301 19424
rect 12355 19384 12364 19424
rect 12404 19384 13420 19424
rect 13460 19384 13469 19424
rect 33763 19384 33772 19424
rect 33812 19384 33821 19424
rect 36547 19384 36556 19424
rect 36596 19384 38092 19424
rect 38132 19384 38141 19424
rect 39235 19384 39244 19424
rect 39284 19384 39293 19424
rect 39523 19384 39532 19424
rect 39572 19384 41164 19424
rect 41204 19384 41213 19424
rect 41443 19384 41452 19424
rect 41492 19384 42700 19424
rect 42740 19384 42749 19424
rect 44323 19384 44332 19424
rect 44372 19384 45580 19424
rect 45620 19384 45629 19424
rect 46723 19384 46732 19424
rect 46772 19384 47116 19424
rect 47156 19384 47165 19424
rect 7276 19340 7316 19384
rect 33772 19340 33812 19384
rect 39244 19340 39284 19384
rect 739 19300 748 19340
rect 788 19300 2188 19340
rect 2228 19300 2956 19340
rect 2996 19300 3005 19340
rect 7267 19300 7276 19340
rect 7316 19300 7325 19340
rect 12556 19300 16108 19340
rect 16148 19300 16157 19340
rect 32419 19300 32428 19340
rect 32468 19300 33388 19340
rect 33428 19300 33437 19340
rect 33772 19300 38132 19340
rect 39244 19300 40108 19340
rect 40148 19300 40780 19340
rect 40820 19300 40829 19340
rect 45475 19300 45484 19340
rect 45524 19300 48268 19340
rect 48308 19300 48317 19340
rect 48547 19300 48556 19340
rect 48596 19300 49612 19340
rect 49652 19300 49661 19340
rect 12556 19256 12596 19300
rect 38092 19256 38132 19300
rect 41347 19256 41405 19257
rect 48076 19256 48116 19300
rect 3619 19216 3628 19256
rect 3668 19216 4492 19256
rect 4532 19216 4541 19256
rect 4675 19216 4684 19256
rect 4724 19216 4972 19256
rect 5012 19216 5021 19256
rect 6787 19216 6796 19256
rect 6836 19216 8332 19256
rect 8372 19216 8381 19256
rect 10051 19216 10060 19256
rect 10100 19216 10444 19256
rect 10484 19216 10493 19256
rect 11971 19216 11980 19256
rect 12020 19216 12556 19256
rect 12596 19216 12605 19256
rect 12739 19216 12748 19256
rect 12788 19216 13132 19256
rect 13172 19216 13181 19256
rect 32611 19216 32620 19256
rect 32660 19216 33196 19256
rect 33236 19216 33772 19256
rect 33812 19216 33821 19256
rect 34051 19216 34060 19256
rect 34100 19216 34636 19256
rect 34676 19216 34828 19256
rect 34868 19216 35692 19256
rect 35732 19216 35741 19256
rect 36259 19216 36268 19256
rect 36308 19216 37324 19256
rect 37364 19216 37612 19256
rect 37652 19216 37661 19256
rect 38083 19216 38092 19256
rect 38132 19216 39436 19256
rect 39476 19216 39485 19256
rect 40291 19216 40300 19256
rect 40340 19216 40684 19256
rect 40724 19216 40733 19256
rect 41347 19216 41356 19256
rect 41396 19216 41740 19256
rect 41780 19216 41789 19256
rect 42883 19216 42892 19256
rect 42932 19216 44044 19256
rect 44084 19216 44093 19256
rect 45859 19216 45868 19256
rect 45908 19216 46732 19256
rect 46772 19216 46781 19256
rect 48067 19216 48076 19256
rect 48116 19216 48156 19256
rect 50659 19216 50668 19256
rect 50708 19216 51628 19256
rect 51668 19216 51677 19256
rect 41347 19215 41405 19216
rect 4291 19132 4300 19172
rect 4340 19132 29836 19172
rect 29876 19132 31564 19172
rect 31604 19132 31613 19172
rect 32227 19132 32236 19172
rect 32276 19132 33964 19172
rect 34004 19132 34013 19172
rect 38275 19132 38284 19172
rect 38324 19132 38764 19172
rect 38804 19132 38813 19172
rect 39043 19132 39052 19172
rect 39092 19132 39532 19172
rect 39572 19132 41204 19172
rect 42115 19132 42124 19172
rect 42164 19132 42604 19172
rect 42644 19132 42653 19172
rect 43180 19132 45100 19172
rect 45140 19132 45149 19172
rect 46627 19132 46636 19172
rect 46676 19132 46685 19172
rect 47011 19132 47020 19172
rect 47060 19132 47500 19172
rect 47540 19132 47549 19172
rect 0 19088 80 19108
rect 32236 19088 32276 19132
rect 41164 19088 41204 19132
rect 43180 19088 43220 19132
rect 46636 19088 46676 19132
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 4387 19048 4396 19088
rect 4436 19048 6508 19088
rect 6548 19048 7468 19088
rect 7508 19048 7517 19088
rect 9859 19048 9868 19088
rect 9908 19048 10252 19088
rect 10292 19048 10301 19088
rect 30883 19048 30892 19088
rect 30932 19048 32276 19088
rect 39811 19048 39820 19088
rect 39860 19048 40492 19088
rect 40532 19048 41108 19088
rect 41164 19048 43220 19088
rect 44995 19048 45004 19088
rect 45044 19048 47596 19088
rect 47636 19048 48844 19088
rect 48884 19048 49420 19088
rect 49460 19048 49469 19088
rect 0 19028 80 19048
rect 34339 19004 34397 19005
rect 41068 19004 41108 19048
rect 42979 19004 43037 19005
rect 1315 18964 1324 19004
rect 1364 18964 7564 19004
rect 7604 18964 7613 19004
rect 8035 18964 8044 19004
rect 8084 18964 23060 19004
rect 33379 18964 33388 19004
rect 33428 18964 34348 19004
rect 34388 18964 34397 19004
rect 37411 18964 37420 19004
rect 37460 18964 38380 19004
rect 38420 18964 40780 19004
rect 40820 18964 40829 19004
rect 41059 18964 41068 19004
rect 41108 18964 41117 19004
rect 41251 18964 41260 19004
rect 41300 18964 42988 19004
rect 43028 18964 45772 19004
rect 45812 18964 45821 19004
rect 47020 18964 52012 19004
rect 52052 18964 52061 19004
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 16343 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 16729 18920
rect 23020 18836 23060 18964
rect 34339 18963 34397 18964
rect 42979 18963 43037 18964
rect 28343 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 28729 18920
rect 33091 18880 33100 18920
rect 33140 18880 33580 18920
rect 33620 18880 33629 18920
rect 35683 18880 35692 18920
rect 35732 18880 38188 18920
rect 38228 18880 38237 18920
rect 40343 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 40729 18920
rect 41539 18880 41548 18920
rect 41588 18880 43604 18920
rect 45283 18880 45292 18920
rect 45332 18880 46348 18920
rect 46388 18880 46924 18920
rect 46964 18880 46973 18920
rect 43564 18836 43604 18880
rect 47020 18836 47060 18964
rect 50371 18920 50429 18921
rect 50286 18880 50380 18920
rect 50420 18880 50429 18920
rect 50371 18879 50429 18880
rect 12364 18796 12460 18836
rect 12500 18796 13036 18836
rect 13076 18796 13085 18836
rect 23020 18796 40972 18836
rect 41012 18796 41021 18836
rect 41347 18796 41356 18836
rect 41396 18796 42316 18836
rect 42356 18796 42365 18836
rect 43555 18796 43564 18836
rect 43604 18796 47060 18836
rect 48643 18796 48652 18836
rect 48692 18796 50092 18836
rect 50132 18796 51340 18836
rect 51380 18796 51389 18836
rect 1219 18712 1228 18752
rect 1268 18712 1612 18752
rect 1652 18712 1661 18752
rect 7459 18712 7468 18752
rect 7508 18712 9772 18752
rect 9812 18712 11116 18752
rect 11156 18712 11165 18752
rect 12364 18668 12404 18796
rect 15331 18712 15340 18752
rect 15380 18712 15389 18752
rect 32716 18712 32948 18752
rect 33187 18712 33196 18752
rect 33236 18712 33676 18752
rect 33716 18712 33725 18752
rect 33955 18712 33964 18752
rect 34004 18712 34540 18752
rect 34580 18712 34589 18752
rect 37123 18712 37132 18752
rect 37172 18712 37708 18752
rect 37748 18712 37757 18752
rect 40099 18712 40108 18752
rect 40148 18712 40684 18752
rect 40724 18712 40733 18752
rect 43939 18712 43948 18752
rect 43988 18712 44140 18752
rect 44180 18712 44908 18752
rect 44948 18712 44957 18752
rect 45091 18712 45100 18752
rect 45140 18712 46540 18752
rect 46580 18712 46589 18752
rect 49603 18712 49612 18752
rect 49652 18712 50380 18752
rect 50420 18712 50429 18752
rect 50947 18712 50956 18752
rect 50996 18712 51092 18752
rect 15340 18668 15380 18712
rect 32716 18668 32756 18712
rect 32908 18668 32948 18712
rect 41731 18668 41789 18669
rect 2083 18628 2092 18668
rect 2132 18628 3532 18668
rect 3572 18628 3581 18668
rect 7075 18628 7084 18668
rect 7124 18628 7220 18668
rect 7180 18584 7220 18628
rect 7468 18628 7564 18668
rect 7604 18628 10732 18668
rect 10772 18628 10781 18668
rect 10924 18628 12404 18668
rect 12451 18628 12460 18668
rect 12500 18628 12940 18668
rect 12980 18628 13612 18668
rect 13652 18628 13661 18668
rect 15340 18628 32756 18668
rect 32803 18628 32812 18668
rect 32852 18628 32861 18668
rect 32908 18628 41740 18668
rect 41780 18628 41789 18668
rect 42019 18628 42028 18668
rect 42068 18628 43084 18668
rect 43124 18628 43133 18668
rect 3427 18544 3436 18584
rect 3476 18544 4108 18584
rect 4148 18544 4157 18584
rect 4675 18544 4684 18584
rect 4724 18544 5068 18584
rect 5108 18544 5117 18584
rect 7180 18544 7372 18584
rect 7412 18544 7421 18584
rect 7468 18500 7508 18628
rect 7651 18584 7709 18585
rect 10924 18584 10964 18628
rect 32227 18584 32285 18585
rect 7566 18544 7660 18584
rect 7700 18544 7709 18584
rect 10915 18544 10924 18584
rect 10964 18544 10973 18584
rect 11779 18544 11788 18584
rect 11828 18544 13900 18584
rect 13940 18544 14956 18584
rect 14996 18544 16972 18584
rect 17012 18544 17021 18584
rect 17260 18544 27628 18584
rect 27668 18544 27677 18584
rect 32142 18544 32236 18584
rect 32276 18544 32285 18584
rect 32812 18584 32852 18628
rect 41731 18627 41789 18628
rect 40867 18584 40925 18585
rect 51052 18584 51092 18712
rect 51139 18628 51148 18668
rect 51188 18628 51820 18668
rect 51860 18628 52684 18668
rect 52724 18628 53068 18668
rect 53108 18628 53117 18668
rect 32812 18544 33292 18584
rect 33332 18544 33341 18584
rect 34243 18544 34252 18584
rect 34292 18544 34301 18584
rect 34627 18544 34636 18584
rect 34676 18544 35980 18584
rect 36020 18544 36029 18584
rect 39619 18544 39628 18584
rect 39668 18544 40876 18584
rect 40916 18544 40925 18584
rect 47011 18544 47020 18584
rect 47060 18544 47308 18584
rect 47348 18544 47357 18584
rect 48547 18544 48556 18584
rect 48596 18544 49132 18584
rect 49172 18544 49181 18584
rect 49891 18544 49900 18584
rect 49940 18544 50956 18584
rect 50996 18544 51005 18584
rect 51052 18544 51860 18584
rect 7651 18543 7709 18544
rect 17260 18500 17300 18544
rect 32227 18543 32285 18544
rect 34252 18500 34292 18544
rect 40867 18543 40925 18544
rect 42787 18502 42796 18542
rect 42836 18502 42932 18542
rect 42892 18500 42932 18502
rect 3907 18460 3916 18500
rect 3956 18460 4588 18500
rect 4628 18460 4637 18500
rect 6211 18460 6220 18500
rect 6260 18460 7508 18500
rect 8323 18460 8332 18500
rect 8372 18460 9004 18500
rect 9044 18460 17300 18500
rect 32707 18460 32716 18500
rect 32756 18460 34292 18500
rect 34435 18460 34444 18500
rect 34484 18460 36460 18500
rect 36500 18460 36509 18500
rect 40867 18460 40876 18500
rect 40916 18460 42412 18500
rect 42452 18460 42461 18500
rect 42892 18460 43468 18500
rect 43508 18460 45196 18500
rect 45236 18460 45388 18500
rect 45428 18460 45437 18500
rect 49411 18460 49420 18500
rect 49460 18460 50860 18500
rect 50900 18460 50909 18500
rect 51427 18460 51436 18500
rect 51476 18460 51724 18500
rect 51764 18460 51773 18500
rect 40771 18416 40829 18417
rect 43651 18416 43709 18417
rect 3715 18376 3724 18416
rect 3764 18376 4012 18416
rect 4052 18376 4061 18416
rect 4771 18376 4780 18416
rect 4820 18376 6412 18416
rect 6452 18376 6461 18416
rect 6979 18376 6988 18416
rect 7028 18376 8140 18416
rect 8180 18376 8189 18416
rect 10723 18376 10732 18416
rect 10772 18376 12748 18416
rect 12788 18376 15244 18416
rect 15284 18376 15293 18416
rect 18115 18376 18124 18416
rect 18164 18376 36308 18416
rect 40387 18376 40396 18416
rect 40436 18376 40780 18416
rect 40820 18376 40829 18416
rect 41155 18376 41164 18416
rect 41204 18376 41548 18416
rect 41588 18376 43276 18416
rect 43316 18376 43660 18416
rect 43700 18376 43709 18416
rect 34723 18332 34781 18333
rect 3619 18292 3628 18332
rect 3668 18292 7852 18332
rect 7892 18292 7901 18332
rect 10339 18292 10348 18332
rect 10388 18292 10636 18332
rect 10676 18292 15436 18332
rect 15476 18292 15485 18332
rect 33100 18292 33196 18332
rect 33236 18292 33245 18332
rect 34339 18292 34348 18332
rect 34388 18292 34732 18332
rect 34772 18292 34781 18332
rect 0 18248 80 18268
rect 7555 18248 7613 18249
rect 33100 18248 33140 18292
rect 34723 18291 34781 18292
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 6787 18208 6796 18248
rect 6836 18208 7564 18248
rect 7604 18208 7613 18248
rect 13027 18208 13036 18248
rect 13076 18208 16108 18248
rect 16148 18208 16157 18248
rect 32419 18208 32428 18248
rect 32468 18208 34540 18248
rect 34580 18208 34589 18248
rect 0 18188 80 18208
rect 7555 18207 7613 18208
rect 34339 18164 34397 18165
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 15103 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 15489 18164
rect 27103 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 27489 18164
rect 34254 18124 34348 18164
rect 34388 18124 34397 18164
rect 34339 18123 34397 18124
rect 36268 18080 36308 18376
rect 40771 18375 40829 18376
rect 43651 18375 43709 18376
rect 47491 18416 47549 18417
rect 51820 18416 51860 18544
rect 47491 18376 47500 18416
rect 47540 18376 49324 18416
rect 49364 18376 49373 18416
rect 50563 18376 50572 18416
rect 50612 18376 51052 18416
rect 51092 18376 51101 18416
rect 51811 18376 51820 18416
rect 51860 18376 51869 18416
rect 47491 18375 47549 18376
rect 42979 18332 43037 18333
rect 44611 18332 44669 18333
rect 39331 18292 39340 18332
rect 39380 18292 39389 18332
rect 42894 18292 42988 18332
rect 43028 18292 43037 18332
rect 44515 18292 44524 18332
rect 44564 18292 44620 18332
rect 44660 18292 44669 18332
rect 45091 18292 45100 18332
rect 45140 18292 46156 18332
rect 46196 18292 47212 18332
rect 47252 18292 47261 18332
rect 49123 18292 49132 18332
rect 49172 18292 49708 18332
rect 49748 18292 49757 18332
rect 50467 18292 50476 18332
rect 50516 18292 51916 18332
rect 51956 18292 51965 18332
rect 39340 18248 39380 18292
rect 42979 18291 43037 18292
rect 44611 18291 44669 18292
rect 51907 18248 51965 18249
rect 38179 18208 38188 18248
rect 38228 18208 51916 18248
rect 51956 18208 51965 18248
rect 51907 18207 51965 18208
rect 48931 18164 48989 18165
rect 39103 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 39489 18164
rect 43170 18124 43179 18164
rect 43219 18124 48940 18164
rect 48980 18124 48989 18164
rect 49315 18124 49324 18164
rect 49364 18124 49900 18164
rect 49940 18124 49949 18164
rect 50179 18124 50188 18164
rect 50228 18124 51244 18164
rect 51284 18124 51293 18164
rect 48931 18123 48989 18124
rect 10243 18040 10252 18080
rect 10292 18040 10828 18080
rect 10868 18040 18124 18080
rect 18164 18040 18173 18080
rect 33091 18040 33100 18080
rect 33140 18040 33676 18080
rect 33716 18040 33725 18080
rect 36268 18040 44620 18080
rect 44660 18040 44669 18080
rect 48547 18040 48556 18080
rect 48596 18040 48748 18080
rect 48788 18040 48797 18080
rect 51811 17996 51869 17997
rect 1699 17956 1708 17996
rect 1748 17956 11212 17996
rect 11252 17956 11261 17996
rect 12163 17956 12172 17996
rect 12212 17956 13132 17996
rect 13172 17956 13181 17996
rect 31939 17956 31948 17996
rect 31988 17956 31997 17996
rect 32131 17956 32140 17996
rect 32180 17956 33388 17996
rect 33428 17956 33437 17996
rect 42403 17956 42412 17996
rect 42452 17956 42988 17996
rect 43028 17956 43037 17996
rect 43084 17956 51820 17996
rect 51860 17956 51869 17996
rect 11212 17912 11252 17956
rect 31948 17912 31988 17956
rect 43084 17912 43124 17956
rect 51811 17955 51869 17956
rect 3523 17872 3532 17912
rect 3572 17872 5068 17912
rect 5108 17872 5117 17912
rect 11212 17872 13708 17912
rect 13748 17872 14956 17912
rect 14996 17872 15005 17912
rect 31948 17872 32236 17912
rect 32276 17872 32285 17912
rect 32515 17872 32524 17912
rect 32564 17872 32908 17912
rect 32948 17872 33140 17912
rect 35971 17872 35980 17912
rect 36020 17872 43124 17912
rect 43459 17872 43468 17912
rect 43508 17872 44044 17912
rect 44084 17872 44093 17912
rect 48739 17872 48748 17912
rect 48788 17872 49420 17912
rect 49460 17872 49708 17912
rect 49748 17872 49757 17912
rect 50755 17872 50764 17912
rect 50804 17872 50813 17912
rect 31747 17828 31805 17829
rect 1315 17788 1324 17828
rect 1364 17788 4204 17828
rect 4244 17788 4253 17828
rect 8131 17788 8140 17828
rect 8180 17788 10964 17828
rect 31662 17788 31756 17828
rect 31796 17788 31805 17828
rect 33100 17828 33140 17872
rect 40195 17828 40253 17829
rect 49795 17828 49853 17829
rect 50764 17828 50804 17872
rect 33100 17788 33292 17828
rect 33332 17788 34444 17828
rect 34484 17788 34493 17828
rect 40195 17788 40204 17828
rect 40244 17788 40300 17828
rect 40340 17788 40349 17828
rect 40675 17788 40684 17828
rect 40724 17788 42220 17828
rect 42260 17788 44236 17828
rect 44276 17788 44812 17828
rect 44852 17788 44861 17828
rect 48931 17788 48940 17828
rect 48980 17788 49132 17828
rect 49172 17788 49181 17828
rect 49795 17788 49804 17828
rect 49844 17788 49996 17828
rect 50036 17788 50045 17828
rect 50764 17788 51052 17828
rect 51092 17788 51101 17828
rect 10924 17744 10964 17788
rect 31747 17787 31805 17788
rect 40195 17787 40253 17788
rect 49795 17787 49853 17788
rect 33091 17744 33149 17745
rect 43459 17744 43517 17745
rect 5155 17704 5164 17744
rect 5204 17704 8332 17744
rect 8372 17704 8381 17744
rect 9955 17704 9964 17744
rect 10004 17704 10732 17744
rect 10772 17704 10781 17744
rect 10915 17704 10924 17744
rect 10964 17704 11308 17744
rect 11348 17704 13036 17744
rect 13076 17704 13085 17744
rect 30211 17704 30220 17744
rect 30260 17704 32140 17744
rect 32180 17704 32189 17744
rect 32803 17704 32812 17744
rect 32852 17704 33100 17744
rect 33140 17704 33149 17744
rect 33571 17704 33580 17744
rect 33620 17704 34636 17744
rect 34676 17704 34685 17744
rect 37507 17704 37516 17744
rect 37556 17704 38188 17744
rect 38228 17704 38237 17744
rect 40483 17704 40492 17744
rect 40532 17704 41740 17744
rect 41780 17704 43084 17744
rect 43124 17704 43133 17744
rect 43374 17704 43468 17744
rect 43508 17704 43517 17744
rect 44131 17704 44140 17744
rect 44180 17704 45100 17744
rect 45140 17704 45149 17744
rect 46435 17704 46444 17744
rect 46484 17704 46732 17744
rect 46772 17704 46781 17744
rect 47491 17704 47500 17744
rect 47540 17704 48652 17744
rect 48692 17704 48701 17744
rect 49603 17704 49612 17744
rect 49652 17704 50188 17744
rect 50228 17704 50764 17744
rect 50804 17704 50813 17744
rect 33091 17703 33149 17704
rect 43459 17703 43517 17704
rect 4099 17620 4108 17660
rect 4148 17620 6124 17660
rect 6164 17620 6604 17660
rect 6644 17620 9868 17660
rect 9908 17620 10828 17660
rect 10868 17620 10877 17660
rect 11491 17620 11500 17660
rect 11540 17620 47980 17660
rect 48020 17620 48029 17660
rect 7555 17576 7613 17577
rect 38275 17576 38333 17577
rect 547 17536 556 17576
rect 596 17536 1132 17576
rect 1172 17536 1181 17576
rect 7470 17536 7564 17576
rect 7604 17536 7613 17576
rect 10339 17536 10348 17576
rect 10388 17536 11020 17576
rect 11060 17536 13132 17576
rect 13172 17536 13181 17576
rect 32227 17536 32236 17576
rect 32276 17536 33868 17576
rect 33908 17536 33917 17576
rect 36547 17536 36556 17576
rect 36596 17536 38284 17576
rect 38324 17536 38333 17576
rect 7555 17535 7613 17536
rect 38275 17535 38333 17536
rect 40771 17576 40829 17577
rect 40771 17536 40780 17576
rect 40820 17536 42508 17576
rect 42548 17536 42557 17576
rect 43171 17536 43180 17576
rect 43220 17536 43372 17576
rect 43412 17536 43421 17576
rect 43747 17536 43756 17576
rect 43796 17536 44620 17576
rect 44660 17536 44669 17576
rect 48547 17536 48556 17576
rect 48596 17536 48940 17576
rect 48980 17536 48989 17576
rect 49507 17536 49516 17576
rect 49556 17536 50572 17576
rect 50612 17536 50621 17576
rect 40771 17535 40829 17536
rect 53059 17492 53117 17493
rect 40099 17452 40108 17492
rect 40148 17452 43220 17492
rect 46339 17452 46348 17492
rect 46388 17452 47404 17492
rect 47444 17452 53068 17492
rect 53108 17452 53117 17492
rect 0 17408 80 17428
rect 43180 17408 43220 17452
rect 53059 17451 53117 17452
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 6019 17368 6028 17408
rect 6068 17368 7468 17408
rect 7508 17368 8140 17408
rect 8180 17368 8189 17408
rect 16343 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 16729 17408
rect 28343 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 28729 17408
rect 33859 17368 33868 17408
rect 33908 17368 34444 17408
rect 34484 17368 34493 17408
rect 40343 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 40729 17408
rect 43180 17368 44620 17408
rect 44660 17368 44669 17408
rect 46915 17368 46924 17408
rect 46964 17368 47116 17408
rect 47156 17368 47165 17408
rect 49795 17368 49804 17408
rect 49844 17368 50092 17408
rect 50132 17368 50141 17408
rect 53059 17368 53068 17408
rect 53108 17368 53117 17408
rect 0 17348 80 17368
rect 53068 17324 53108 17368
rect 56131 17324 56189 17325
rect 56899 17324 56957 17325
rect 57283 17324 57341 17325
rect 57571 17324 57629 17325
rect 59011 17324 59069 17325
rect 59395 17324 59453 17325
rect 59683 17324 59741 17325
rect 60835 17324 60893 17325
rect 61891 17324 61949 17325
rect 63907 17324 63965 17325
rect 64771 17324 64829 17325
rect 66019 17324 66077 17325
rect 66211 17324 66269 17325
rect 69091 17324 69149 17325
rect 71011 17324 71069 17325
rect 77155 17324 77213 17325
rect 1123 17284 1132 17324
rect 1172 17284 1996 17324
rect 2036 17284 2045 17324
rect 5059 17284 5068 17324
rect 5108 17284 6220 17324
rect 6260 17284 6269 17324
rect 6787 17284 6796 17324
rect 6836 17284 7084 17324
rect 7124 17284 7133 17324
rect 32227 17284 32236 17324
rect 32276 17284 32524 17324
rect 32564 17284 32573 17324
rect 32803 17284 32812 17324
rect 32852 17284 33004 17324
rect 33044 17284 33053 17324
rect 36163 17284 36172 17324
rect 36212 17284 36460 17324
rect 36500 17284 37612 17324
rect 37652 17284 38380 17324
rect 38420 17284 38429 17324
rect 53068 17284 54745 17324
rect 54785 17284 54794 17324
rect 56131 17284 56140 17324
rect 56180 17284 56745 17324
rect 56785 17284 56794 17324
rect 56899 17284 56908 17324
rect 56948 17284 57145 17324
rect 57185 17284 57194 17324
rect 57246 17284 57255 17324
rect 57332 17284 57390 17324
rect 57571 17284 57580 17324
rect 57620 17284 58745 17324
rect 58785 17284 58794 17324
rect 58846 17284 58855 17324
rect 58895 17284 58964 17324
rect 56131 17283 56189 17284
rect 56899 17283 56957 17284
rect 57283 17283 57341 17284
rect 57571 17283 57629 17284
rect 58924 17241 58964 17284
rect 59011 17284 59020 17324
rect 59060 17284 59255 17324
rect 59295 17284 59304 17324
rect 59395 17284 59404 17324
rect 59444 17284 59545 17324
rect 59585 17284 59594 17324
rect 59646 17284 59655 17324
rect 59732 17284 59790 17324
rect 60835 17284 60844 17324
rect 60884 17284 61255 17324
rect 61295 17284 61304 17324
rect 61891 17284 61900 17324
rect 61940 17284 62055 17324
rect 62095 17284 62104 17324
rect 63907 17284 63916 17324
rect 63956 17284 64455 17324
rect 64495 17284 64504 17324
rect 64771 17284 64780 17324
rect 64820 17284 65655 17324
rect 65695 17284 65704 17324
rect 65960 17284 66028 17324
rect 66095 17284 66104 17324
rect 66211 17284 66220 17324
rect 66260 17284 67255 17324
rect 67295 17284 67304 17324
rect 69091 17284 69100 17324
rect 69140 17284 70455 17324
rect 70495 17284 70504 17324
rect 71011 17284 71020 17324
rect 71060 17284 71548 17324
rect 71588 17284 71597 17324
rect 76780 17284 76855 17324
rect 76895 17284 76904 17324
rect 77136 17284 77145 17324
rect 77204 17284 77280 17324
rect 59011 17283 59069 17284
rect 59395 17283 59453 17284
rect 59683 17283 59741 17284
rect 60835 17283 60893 17284
rect 61891 17283 61949 17284
rect 63907 17283 63965 17284
rect 64771 17283 64829 17284
rect 66019 17283 66077 17284
rect 66211 17283 66269 17284
rect 69091 17283 69149 17284
rect 71011 17283 71069 17284
rect 76780 17241 76820 17284
rect 77155 17283 77213 17284
rect 53251 17240 53309 17241
rect 56419 17240 56477 17241
rect 56707 17240 56765 17241
rect 57379 17240 57437 17241
rect 57667 17240 57725 17241
rect 58051 17240 58109 17241
rect 58435 17240 58493 17241
rect 58915 17240 58973 17241
rect 6307 17200 6316 17240
rect 6356 17200 6988 17240
rect 7028 17200 7037 17240
rect 28291 17200 28300 17240
rect 28340 17200 28780 17240
rect 28820 17200 29164 17240
rect 29204 17200 29213 17240
rect 39715 17200 39724 17240
rect 39764 17200 42028 17240
rect 42068 17200 52876 17240
rect 52916 17200 52925 17240
rect 53251 17200 53260 17240
rect 53300 17200 54455 17240
rect 54495 17200 54504 17240
rect 56360 17200 56428 17240
rect 56495 17200 56504 17240
rect 56707 17200 56716 17240
rect 56756 17200 56855 17240
rect 56895 17200 56904 17240
rect 57379 17200 57388 17240
rect 57428 17200 57545 17240
rect 57585 17200 57594 17240
rect 57646 17200 57655 17240
rect 57716 17200 57790 17240
rect 58046 17200 58055 17240
rect 58100 17200 58190 17240
rect 58360 17200 58444 17240
rect 58495 17200 58504 17240
rect 58915 17200 58924 17240
rect 58964 17200 58973 17240
rect 53251 17199 53309 17200
rect 56419 17199 56477 17200
rect 56707 17199 56765 17200
rect 57379 17199 57437 17200
rect 57667 17199 57725 17200
rect 58051 17199 58109 17200
rect 58435 17199 58493 17200
rect 58915 17199 58973 17200
rect 59203 17240 59261 17241
rect 60643 17240 60701 17241
rect 61987 17240 62045 17241
rect 65251 17240 65309 17241
rect 66499 17240 66557 17241
rect 76771 17240 76829 17241
rect 59203 17200 59212 17240
rect 59252 17200 60455 17240
rect 60495 17200 60504 17240
rect 60643 17200 60652 17240
rect 60692 17200 60855 17240
rect 60895 17200 60904 17240
rect 61987 17200 61996 17240
rect 62036 17200 62455 17240
rect 62495 17200 62504 17240
rect 63811 17200 63820 17240
rect 63860 17200 64345 17240
rect 64385 17200 64394 17240
rect 65251 17200 65260 17240
rect 65300 17200 65545 17240
rect 65585 17200 65594 17240
rect 66499 17200 66508 17240
rect 66548 17200 66855 17240
rect 66895 17200 66904 17240
rect 67363 17200 67372 17240
rect 67412 17200 70345 17240
rect 70385 17200 70394 17240
rect 74179 17200 74188 17240
rect 74228 17200 74855 17240
rect 74895 17200 74904 17240
rect 76771 17200 76780 17240
rect 76820 17200 76829 17240
rect 59203 17199 59261 17200
rect 60643 17199 60701 17200
rect 61987 17199 62045 17200
rect 65251 17199 65309 17200
rect 66499 17199 66557 17200
rect 76771 17199 76829 17200
rect 54691 17156 54749 17157
rect 65155 17156 65213 17157
rect 66307 17156 66365 17157
rect 66691 17156 66749 17157
rect 68419 17156 68477 17157
rect 70147 17156 70205 17157
rect 72547 17156 72605 17157
rect 75811 17156 75869 17157
rect 6508 17116 10060 17156
rect 10100 17116 10348 17156
rect 10388 17116 10397 17156
rect 32035 17116 32044 17156
rect 32084 17116 32716 17156
rect 32756 17116 32765 17156
rect 54691 17116 54700 17156
rect 54740 17116 57945 17156
rect 57985 17116 57994 17156
rect 59683 17116 59692 17156
rect 59732 17116 60055 17156
rect 60095 17116 60104 17156
rect 61027 17116 61036 17156
rect 61076 17116 62956 17156
rect 62996 17116 65012 17156
rect 65136 17116 65145 17156
rect 65204 17116 65280 17156
rect 66307 17116 66316 17156
rect 66356 17116 66455 17156
rect 66495 17116 66504 17156
rect 66650 17116 66700 17156
rect 66740 17116 66745 17156
rect 66785 17116 66794 17156
rect 68419 17116 68428 17156
rect 68468 17116 69945 17156
rect 69985 17116 69994 17156
rect 70046 17116 70055 17156
rect 70095 17116 70156 17156
rect 70196 17116 70205 17156
rect 6508 17072 6548 17116
rect 54691 17115 54749 17116
rect 32227 17072 32285 17073
rect 42403 17072 42461 17073
rect 43651 17072 43709 17073
rect 5251 17032 5260 17072
rect 5300 17032 6508 17072
rect 6548 17032 6557 17072
rect 6691 17032 6700 17072
rect 6740 17032 7084 17072
rect 7124 17032 7133 17072
rect 11011 17032 11020 17072
rect 11060 17032 12940 17072
rect 12980 17032 13324 17072
rect 13364 17032 13373 17072
rect 32227 17032 32236 17072
rect 32276 17032 33292 17072
rect 33332 17032 37324 17072
rect 37364 17032 37373 17072
rect 37795 17032 37804 17072
rect 37844 17032 38132 17072
rect 38563 17032 38572 17072
rect 38612 17032 39052 17072
rect 39092 17032 40396 17072
rect 40436 17032 40445 17072
rect 42318 17032 42412 17072
rect 42452 17032 42461 17072
rect 43566 17032 43660 17072
rect 43700 17032 44140 17072
rect 44180 17032 44189 17072
rect 44419 17032 44428 17072
rect 44468 17032 45484 17072
rect 45524 17032 45533 17072
rect 46243 17032 46252 17072
rect 46292 17032 47308 17072
rect 47348 17032 47357 17072
rect 49900 17032 52780 17072
rect 52820 17032 52829 17072
rect 59587 17032 59596 17072
rect 59636 17032 64916 17072
rect 32227 17031 32285 17032
rect 35299 16988 35357 16989
rect 37987 16988 38045 16989
rect 2659 16948 2668 16988
rect 2708 16948 4012 16988
rect 4052 16948 4061 16988
rect 6115 16948 6124 16988
rect 6164 16948 10156 16988
rect 10196 16948 11500 16988
rect 11540 16948 11549 16988
rect 32995 16948 33004 16988
rect 33044 16948 33196 16988
rect 33236 16948 35308 16988
rect 35348 16948 35357 16988
rect 36931 16948 36940 16988
rect 36980 16948 37996 16988
rect 38036 16948 38045 16988
rect 38092 16988 38132 17032
rect 42403 17031 42461 17032
rect 43651 17031 43709 17032
rect 40771 16988 40829 16989
rect 38092 16948 39148 16988
rect 39188 16948 40780 16988
rect 40820 16948 40829 16988
rect 44707 16948 44716 16988
rect 44756 16948 45004 16988
rect 45044 16948 45053 16988
rect 46819 16948 46828 16988
rect 46868 16948 47404 16988
rect 47444 16948 47453 16988
rect 35299 16947 35357 16948
rect 37987 16947 38045 16948
rect 40771 16947 40829 16948
rect 10051 16864 10060 16904
rect 10100 16864 10444 16904
rect 10484 16864 10493 16904
rect 42883 16864 42892 16904
rect 42932 16864 43220 16904
rect 43555 16864 43564 16904
rect 43604 16864 44140 16904
rect 44180 16864 44189 16904
rect 47011 16864 47020 16904
rect 47060 16864 49708 16904
rect 49748 16864 49757 16904
rect 40675 16820 40733 16821
rect 40867 16820 40925 16821
rect 31171 16780 31180 16820
rect 31220 16780 38956 16820
rect 38996 16780 39724 16820
rect 39764 16780 39773 16820
rect 40590 16780 40684 16820
rect 40724 16780 40733 16820
rect 40782 16780 40876 16820
rect 40916 16780 40925 16820
rect 40675 16779 40733 16780
rect 40867 16779 40925 16780
rect 43180 16736 43220 16864
rect 45955 16780 45964 16820
rect 46004 16780 47116 16820
rect 47156 16780 47165 16820
rect 49900 16736 49940 17032
rect 50371 16988 50429 16989
rect 50083 16948 50092 16988
rect 50132 16948 50380 16988
rect 50420 16948 50429 16988
rect 52579 16948 52588 16988
rect 52628 16948 53548 16988
rect 53588 16948 53597 16988
rect 60067 16948 60076 16988
rect 60116 16948 64724 16988
rect 50371 16947 50429 16948
rect 52291 16864 52300 16904
rect 52340 16864 53452 16904
rect 53492 16864 53501 16904
rect 54883 16864 54892 16904
rect 54932 16864 62764 16904
rect 62804 16864 62813 16904
rect 50275 16780 50284 16820
rect 50324 16780 50668 16820
rect 50708 16780 51628 16820
rect 51668 16780 51677 16820
rect 52003 16780 52012 16820
rect 52052 16780 54028 16820
rect 54068 16780 54077 16820
rect 57283 16780 57292 16820
rect 57332 16780 63628 16820
rect 63668 16780 63677 16820
rect 64684 16736 64724 16948
rect 64876 16820 64916 17032
rect 64972 16988 65012 17116
rect 65155 17115 65213 17116
rect 66307 17115 66365 17116
rect 66691 17115 66749 17116
rect 68419 17115 68477 17116
rect 70147 17115 70205 17116
rect 71212 17116 71255 17156
rect 71295 17116 71304 17156
rect 72046 17116 72055 17156
rect 72095 17116 72556 17156
rect 72596 17116 72605 17156
rect 74659 17116 74668 17156
rect 74708 17116 75255 17156
rect 75295 17116 75304 17156
rect 75646 17116 75655 17156
rect 75695 17116 75820 17156
rect 75860 17116 75869 17156
rect 77827 17116 77836 17156
rect 77876 17116 79255 17156
rect 79295 17116 79304 17156
rect 66787 17072 66845 17073
rect 71212 17072 71252 17116
rect 72547 17115 72605 17116
rect 75811 17115 75869 17116
rect 66307 17032 66316 17072
rect 66356 17032 66796 17072
rect 66836 17032 66845 17072
rect 67171 17032 67180 17072
rect 67220 17032 67229 17072
rect 69964 17032 71252 17072
rect 66787 17031 66845 17032
rect 67180 16988 67220 17032
rect 69964 16988 70004 17032
rect 64972 16948 67220 16988
rect 69955 16948 69964 16988
rect 70004 16948 70013 16988
rect 66211 16864 66220 16904
rect 66260 16864 67564 16904
rect 67604 16864 67613 16904
rect 64876 16780 68044 16820
rect 68084 16780 68093 16820
rect 69196 16780 70732 16820
rect 70772 16780 70781 16820
rect 69196 16736 69236 16780
rect 43180 16696 43468 16736
rect 43508 16696 43517 16736
rect 45379 16696 45388 16736
rect 45428 16696 49940 16736
rect 50371 16696 50380 16736
rect 50420 16696 50572 16736
rect 50612 16696 50621 16736
rect 50755 16696 50764 16736
rect 50804 16696 51340 16736
rect 51380 16696 52684 16736
rect 52724 16696 55084 16736
rect 55124 16696 55133 16736
rect 56611 16696 56620 16736
rect 56660 16696 63916 16736
rect 63956 16696 63965 16736
rect 64684 16696 66220 16736
rect 66260 16696 66269 16736
rect 66595 16696 66604 16736
rect 66644 16696 68716 16736
rect 68756 16696 69236 16736
rect 61027 16652 61085 16653
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 15103 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 15489 16652
rect 27103 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 27489 16652
rect 35971 16612 35980 16652
rect 36020 16612 37900 16652
rect 37940 16612 38476 16652
rect 38516 16612 38525 16652
rect 39103 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 39489 16652
rect 41443 16612 41452 16652
rect 41492 16612 42316 16652
rect 42356 16612 44332 16652
rect 44372 16612 47060 16652
rect 47203 16612 47212 16652
rect 47252 16612 50804 16652
rect 50851 16612 50860 16652
rect 50900 16612 51244 16652
rect 51284 16612 55180 16652
rect 55220 16612 55229 16652
rect 60739 16612 60748 16652
rect 60788 16612 61036 16652
rect 61076 16612 61085 16652
rect 66691 16612 66700 16652
rect 66740 16612 70828 16652
rect 70868 16612 70877 16652
rect 72451 16612 72460 16652
rect 72500 16612 73132 16652
rect 73172 16612 73181 16652
rect 0 16568 80 16588
rect 47020 16568 47060 16612
rect 47491 16568 47549 16569
rect 0 16528 1036 16568
rect 1076 16528 1085 16568
rect 40483 16528 40492 16568
rect 40532 16528 43220 16568
rect 45955 16528 45964 16568
rect 46004 16528 46924 16568
rect 46964 16528 46973 16568
rect 47020 16528 47500 16568
rect 47540 16528 47549 16568
rect 0 16508 80 16528
rect 43180 16484 43220 16528
rect 47491 16527 47549 16528
rect 49795 16568 49853 16569
rect 50764 16568 50804 16612
rect 61027 16611 61085 16612
rect 65731 16568 65789 16569
rect 49795 16528 49804 16568
rect 49844 16528 50380 16568
rect 50420 16528 50668 16568
rect 50708 16528 50717 16568
rect 50764 16528 52588 16568
rect 52628 16528 52637 16568
rect 52771 16528 52780 16568
rect 52820 16528 53932 16568
rect 53972 16528 53981 16568
rect 55756 16528 58348 16568
rect 58388 16528 58397 16568
rect 62563 16528 62572 16568
rect 62612 16528 63380 16568
rect 65646 16528 65740 16568
rect 65780 16528 65789 16568
rect 66115 16528 66124 16568
rect 66164 16528 72844 16568
rect 72884 16528 72893 16568
rect 49795 16527 49853 16528
rect 55756 16484 55796 16528
rect 56323 16484 56381 16485
rect 63340 16484 63380 16528
rect 65731 16527 65789 16528
rect 43180 16444 55796 16484
rect 56035 16444 56044 16484
rect 56084 16444 56093 16484
rect 56238 16444 56332 16484
rect 56372 16444 56381 16484
rect 56995 16444 57004 16484
rect 57044 16444 63244 16484
rect 63284 16444 63293 16484
rect 63340 16444 63916 16484
rect 63956 16444 68812 16484
rect 68852 16444 68861 16484
rect 69283 16444 69292 16484
rect 69332 16444 72460 16484
rect 72500 16444 72509 16484
rect 73411 16444 73420 16484
rect 73460 16444 73996 16484
rect 74036 16444 74045 16484
rect 56044 16400 56084 16444
rect 56323 16443 56381 16444
rect 60739 16400 60797 16401
rect 31651 16360 31660 16400
rect 31700 16360 32236 16400
rect 32276 16360 32285 16400
rect 32611 16360 32620 16400
rect 32660 16360 33100 16400
rect 33140 16360 33676 16400
rect 33716 16360 36364 16400
rect 36404 16360 37420 16400
rect 37460 16360 37469 16400
rect 44995 16360 45004 16400
rect 45044 16360 56084 16400
rect 60654 16360 60748 16400
rect 60788 16360 60797 16400
rect 60739 16359 60797 16360
rect 60931 16400 60989 16401
rect 71779 16400 71837 16401
rect 60931 16360 60940 16400
rect 60980 16360 61132 16400
rect 61172 16360 61181 16400
rect 65635 16360 65644 16400
rect 65684 16360 67372 16400
rect 67412 16360 67421 16400
rect 67555 16360 67564 16400
rect 67604 16360 68332 16400
rect 68372 16360 68381 16400
rect 69676 16360 71596 16400
rect 71636 16360 71645 16400
rect 71779 16360 71788 16400
rect 71828 16360 71922 16400
rect 73123 16360 73132 16400
rect 73172 16360 73516 16400
rect 73556 16360 73565 16400
rect 60931 16359 60989 16360
rect 1699 16276 1708 16316
rect 1748 16276 6988 16316
rect 7028 16276 9484 16316
rect 9524 16276 9533 16316
rect 10531 16276 10540 16316
rect 10580 16276 11020 16316
rect 11060 16276 11069 16316
rect 35779 16276 35788 16316
rect 35828 16276 37900 16316
rect 37940 16276 37949 16316
rect 46051 16276 46060 16316
rect 46100 16276 46636 16316
rect 46676 16276 46685 16316
rect 47299 16276 47308 16316
rect 47348 16276 55660 16316
rect 55700 16276 55709 16316
rect 58723 16276 58732 16316
rect 58772 16276 59500 16316
rect 59540 16276 60364 16316
rect 60404 16276 67948 16316
rect 67988 16276 67997 16316
rect 60451 16232 60509 16233
rect 69676 16232 69716 16360
rect 71779 16359 71837 16360
rect 70915 16316 70973 16317
rect 70830 16276 70924 16316
rect 70964 16276 70973 16316
rect 72547 16276 72556 16316
rect 72596 16276 72844 16316
rect 72884 16276 72893 16316
rect 73411 16276 73420 16316
rect 73460 16276 73900 16316
rect 73940 16276 73949 16316
rect 73996 16276 75628 16316
rect 75668 16276 75677 16316
rect 78595 16276 78604 16316
rect 78644 16276 79372 16316
rect 79412 16276 79421 16316
rect 70915 16275 70973 16276
rect 70819 16232 70877 16233
rect 73996 16232 74036 16276
rect 78499 16232 78557 16233
rect 4003 16192 4012 16232
rect 4052 16192 6316 16232
rect 6356 16192 6365 16232
rect 32035 16192 32044 16232
rect 32084 16192 33388 16232
rect 33428 16192 33437 16232
rect 36259 16192 36268 16232
rect 36308 16192 36844 16232
rect 36884 16192 36893 16232
rect 41059 16192 41068 16232
rect 41108 16192 42412 16232
rect 42452 16192 42461 16232
rect 46243 16192 46252 16232
rect 46292 16192 46924 16232
rect 46964 16192 46973 16232
rect 47587 16192 47596 16232
rect 47636 16192 49612 16232
rect 49652 16192 49661 16232
rect 49987 16192 49996 16232
rect 50036 16192 51628 16232
rect 51668 16192 51677 16232
rect 52195 16192 52204 16232
rect 52244 16192 53356 16232
rect 53396 16192 53405 16232
rect 53539 16192 53548 16232
rect 53588 16192 54892 16232
rect 54932 16192 54941 16232
rect 55267 16192 55276 16232
rect 55316 16192 57004 16232
rect 57044 16192 57053 16232
rect 58147 16192 58156 16232
rect 58196 16192 59596 16232
rect 59636 16192 59645 16232
rect 60366 16192 60460 16232
rect 60500 16192 60509 16232
rect 64867 16192 64876 16232
rect 64916 16192 66316 16232
rect 66356 16192 66365 16232
rect 67747 16192 67756 16232
rect 67796 16192 69676 16232
rect 69716 16192 69725 16232
rect 69859 16192 69868 16232
rect 69908 16192 70828 16232
rect 70868 16192 71116 16232
rect 71156 16192 71165 16232
rect 72067 16192 72076 16232
rect 72116 16192 74036 16232
rect 74083 16192 74092 16232
rect 74132 16192 74764 16232
rect 74804 16192 74813 16232
rect 78414 16192 78508 16232
rect 78548 16192 78557 16232
rect 60451 16191 60509 16192
rect 70819 16191 70877 16192
rect 78499 16191 78557 16192
rect 42787 16148 42845 16149
rect 71011 16148 71069 16149
rect 74851 16148 74909 16149
rect 37603 16108 37612 16148
rect 37652 16108 38092 16148
rect 38132 16108 38141 16148
rect 42702 16108 42796 16148
rect 42836 16108 42845 16148
rect 51043 16108 51052 16148
rect 51092 16108 52436 16148
rect 52579 16108 52588 16148
rect 52628 16108 55948 16148
rect 55988 16108 55997 16148
rect 60547 16108 60556 16148
rect 60596 16108 61036 16148
rect 61076 16108 61085 16148
rect 61132 16108 62284 16148
rect 62324 16108 62333 16148
rect 63427 16108 63436 16148
rect 63476 16108 63820 16148
rect 63860 16108 65452 16148
rect 65492 16108 68620 16148
rect 68660 16108 68669 16148
rect 69571 16108 69580 16148
rect 69620 16108 71020 16148
rect 71060 16108 71069 16148
rect 72931 16108 72940 16148
rect 72980 16108 74860 16148
rect 74900 16108 75340 16148
rect 75380 16108 75389 16148
rect 42787 16107 42845 16108
rect 36739 16064 36797 16065
rect 41155 16064 41213 16065
rect 51139 16064 51197 16065
rect 451 16024 460 16064
rect 500 16024 10348 16064
rect 10388 16024 10397 16064
rect 35683 16024 35692 16064
rect 35732 16024 36748 16064
rect 36788 16024 36797 16064
rect 41070 16024 41164 16064
rect 41204 16024 41213 16064
rect 45571 16024 45580 16064
rect 45620 16024 45868 16064
rect 45908 16024 45917 16064
rect 47395 16024 47404 16064
rect 47444 16024 48940 16064
rect 48980 16024 48989 16064
rect 50563 16024 50572 16064
rect 50612 16024 50956 16064
rect 50996 16024 51005 16064
rect 51054 16024 51148 16064
rect 51188 16024 51197 16064
rect 36739 16023 36797 16024
rect 41155 16023 41213 16024
rect 48940 15980 48980 16024
rect 51139 16023 51197 16024
rect 52195 16064 52253 16065
rect 52396 16064 52436 16108
rect 61132 16064 61172 16108
rect 71011 16107 71069 16108
rect 74851 16107 74909 16108
rect 61411 16064 61469 16065
rect 52195 16024 52204 16064
rect 52244 16024 52300 16064
rect 52340 16024 52349 16064
rect 52396 16024 61172 16064
rect 61326 16024 61420 16064
rect 61460 16024 61469 16064
rect 61987 16024 61996 16064
rect 62036 16024 63532 16064
rect 63572 16024 67564 16064
rect 67604 16024 67613 16064
rect 68131 16024 68140 16064
rect 68180 16024 69292 16064
rect 69332 16024 69341 16064
rect 71971 16024 71980 16064
rect 72020 16024 73420 16064
rect 73460 16024 73469 16064
rect 73603 16024 73612 16064
rect 73652 16024 74188 16064
rect 74228 16024 74237 16064
rect 52195 16023 52253 16024
rect 61411 16023 61469 16024
rect 66595 15980 66653 15981
rect 48940 15940 55564 15980
rect 55604 15940 55613 15980
rect 55939 15940 55948 15980
rect 55988 15940 56908 15980
rect 56948 15940 57772 15980
rect 57812 15940 63148 15980
rect 63188 15940 63197 15980
rect 64963 15940 64972 15980
rect 65012 15940 66260 15980
rect 53155 15896 53213 15897
rect 59107 15896 59165 15897
rect 64972 15896 65012 15940
rect 66220 15896 66260 15940
rect 66595 15940 66604 15980
rect 66644 15940 66700 15980
rect 66740 15940 66749 15980
rect 67075 15940 67084 15980
rect 67124 15940 72556 15980
rect 72596 15940 73228 15980
rect 73268 15940 73277 15980
rect 74371 15940 74380 15980
rect 74420 15940 76108 15980
rect 76148 15940 76157 15980
rect 66595 15939 66653 15940
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 16343 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 16729 15896
rect 28343 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 28729 15896
rect 40343 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 40729 15896
rect 45859 15856 45868 15896
rect 45908 15856 46732 15896
rect 46772 15856 46781 15896
rect 51427 15856 51436 15896
rect 51476 15856 53164 15896
rect 53204 15856 53213 15896
rect 53347 15856 53356 15896
rect 53396 15856 56140 15896
rect 56180 15856 56189 15896
rect 59022 15856 59116 15896
rect 59156 15856 59165 15896
rect 60931 15856 60940 15896
rect 60980 15856 61420 15896
rect 61460 15856 65012 15896
rect 65635 15856 65644 15896
rect 65684 15856 66124 15896
rect 66164 15856 66173 15896
rect 66220 15856 67276 15896
rect 67316 15856 67325 15896
rect 68611 15856 68620 15896
rect 68660 15856 69964 15896
rect 70004 15856 70013 15896
rect 70339 15856 70348 15896
rect 70388 15856 76012 15896
rect 76052 15856 76061 15896
rect 77635 15856 77644 15896
rect 77684 15856 79084 15896
rect 79124 15856 79133 15896
rect 53155 15855 53213 15856
rect 59107 15855 59165 15856
rect 56131 15812 56189 15813
rect 70348 15812 70388 15856
rect 34339 15772 34348 15812
rect 34388 15772 38092 15812
rect 38132 15772 38668 15812
rect 38708 15772 38717 15812
rect 51907 15772 51916 15812
rect 51956 15772 54796 15812
rect 54836 15772 54845 15812
rect 56131 15772 56140 15812
rect 56180 15772 56620 15812
rect 56660 15772 56669 15812
rect 57955 15772 57964 15812
rect 58004 15772 58348 15812
rect 58388 15772 58397 15812
rect 58531 15772 58540 15812
rect 58580 15772 58924 15812
rect 58964 15772 58973 15812
rect 59116 15772 59404 15812
rect 59444 15772 60076 15812
rect 60116 15772 65068 15812
rect 65108 15772 70252 15812
rect 70292 15772 70388 15812
rect 72259 15772 72268 15812
rect 72308 15772 73708 15812
rect 73748 15772 73757 15812
rect 56131 15771 56189 15772
rect 0 15728 80 15748
rect 53251 15728 53309 15729
rect 59116 15728 59156 15772
rect 64099 15728 64157 15729
rect 77059 15728 77117 15729
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 35107 15688 35116 15728
rect 35156 15688 35980 15728
rect 36020 15688 36172 15728
rect 36212 15688 36221 15728
rect 49315 15688 49324 15728
rect 49364 15688 52588 15728
rect 52628 15688 52637 15728
rect 53251 15688 53260 15728
rect 53300 15688 56428 15728
rect 56468 15688 56477 15728
rect 56707 15688 56716 15728
rect 56756 15688 58580 15728
rect 59107 15688 59116 15728
rect 59156 15688 59165 15728
rect 60652 15688 61900 15728
rect 61940 15688 61949 15728
rect 64014 15688 64108 15728
rect 64148 15688 64157 15728
rect 0 15668 80 15688
rect 53251 15687 53309 15688
rect 37027 15644 37085 15645
rect 41155 15644 41213 15645
rect 53155 15644 53213 15645
rect 58540 15644 58580 15688
rect 60547 15644 60605 15645
rect 35875 15604 35884 15644
rect 35924 15604 36364 15644
rect 36404 15604 36413 15644
rect 36942 15604 37036 15644
rect 37076 15604 37085 15644
rect 37987 15604 37996 15644
rect 38036 15604 38380 15644
rect 38420 15604 38429 15644
rect 39619 15604 39628 15644
rect 39668 15604 41164 15644
rect 41204 15604 41213 15644
rect 46627 15604 46636 15644
rect 46676 15604 49036 15644
rect 49076 15604 49085 15644
rect 49795 15604 49804 15644
rect 49844 15604 50476 15644
rect 50516 15604 50860 15644
rect 50900 15604 50909 15644
rect 53155 15604 53164 15644
rect 53204 15604 53356 15644
rect 53396 15604 53405 15644
rect 56035 15604 56044 15644
rect 56084 15604 58444 15644
rect 58484 15604 58493 15644
rect 58540 15604 60556 15644
rect 60596 15604 60605 15644
rect 37027 15603 37085 15604
rect 41155 15603 41213 15604
rect 53155 15603 53213 15604
rect 60547 15603 60605 15604
rect 47491 15560 47549 15561
rect 47779 15560 47837 15561
rect 51139 15560 51197 15561
rect 60652 15560 60692 15688
rect 64099 15687 64157 15688
rect 67468 15688 68428 15728
rect 68468 15688 68477 15728
rect 69859 15688 69868 15728
rect 69908 15688 70348 15728
rect 70388 15688 70397 15728
rect 71299 15688 71308 15728
rect 71348 15688 72172 15728
rect 72212 15688 72748 15728
rect 72788 15688 73132 15728
rect 73172 15688 73181 15728
rect 76771 15688 76780 15728
rect 76820 15688 77068 15728
rect 77108 15688 77117 15728
rect 77731 15688 77740 15728
rect 77780 15688 78796 15728
rect 78836 15688 79180 15728
rect 79220 15688 79229 15728
rect 67468 15644 67508 15688
rect 77059 15687 77117 15688
rect 63340 15604 67468 15644
rect 67508 15604 67517 15644
rect 68428 15604 72364 15644
rect 72404 15604 72413 15644
rect 75619 15604 75628 15644
rect 75668 15604 76972 15644
rect 77012 15604 77021 15644
rect 60931 15560 60989 15561
rect 63340 15560 63380 15604
rect 68428 15560 68468 15604
rect 27619 15520 27628 15560
rect 27668 15520 32908 15560
rect 32948 15520 35692 15560
rect 35732 15520 36556 15560
rect 36596 15520 37900 15560
rect 37940 15520 39340 15560
rect 39380 15520 39916 15560
rect 39956 15520 39965 15560
rect 40387 15520 40396 15560
rect 40436 15520 40780 15560
rect 40820 15520 42988 15560
rect 43028 15520 43468 15560
rect 43508 15520 43517 15560
rect 47406 15520 47500 15560
rect 47540 15520 47549 15560
rect 47694 15520 47788 15560
rect 47828 15520 48268 15560
rect 48308 15520 48317 15560
rect 49123 15520 49132 15560
rect 49172 15520 51148 15560
rect 51188 15520 51197 15560
rect 55747 15520 55756 15560
rect 55796 15520 57100 15560
rect 57140 15520 58348 15560
rect 58388 15520 58397 15560
rect 58627 15520 58636 15560
rect 58676 15520 60692 15560
rect 60846 15520 60940 15560
rect 60980 15520 60989 15560
rect 61123 15520 61132 15560
rect 61172 15520 63380 15560
rect 65347 15520 65356 15560
rect 65396 15520 65740 15560
rect 65780 15520 67180 15560
rect 67220 15520 68044 15560
rect 68084 15520 68093 15560
rect 68419 15520 68428 15560
rect 68468 15520 68477 15560
rect 70051 15520 70060 15560
rect 70100 15520 72268 15560
rect 72308 15520 72317 15560
rect 75715 15520 75724 15560
rect 75764 15520 76684 15560
rect 76724 15520 76733 15560
rect 47491 15519 47549 15520
rect 47779 15519 47837 15520
rect 51139 15519 51197 15520
rect 60931 15519 60989 15520
rect 62275 15476 62333 15477
rect 1699 15436 1708 15476
rect 1748 15436 2860 15476
rect 2900 15436 2909 15476
rect 34435 15436 34444 15476
rect 34484 15436 36748 15476
rect 36788 15436 38764 15476
rect 38804 15436 38813 15476
rect 46339 15436 46348 15476
rect 46388 15436 46828 15476
rect 46868 15436 46877 15476
rect 47299 15436 47308 15476
rect 47348 15436 48076 15476
rect 48116 15436 48125 15476
rect 49891 15436 49900 15476
rect 49940 15436 51052 15476
rect 51092 15436 51101 15476
rect 52579 15436 52588 15476
rect 52628 15436 55468 15476
rect 55508 15436 55852 15476
rect 55892 15436 57868 15476
rect 57908 15436 57917 15476
rect 58819 15436 58828 15476
rect 58868 15436 61228 15476
rect 61268 15436 61900 15476
rect 61940 15436 61949 15476
rect 62190 15436 62284 15476
rect 62324 15436 62333 15476
rect 62275 15435 62333 15436
rect 64963 15476 65021 15477
rect 64963 15436 64972 15476
rect 65012 15436 65548 15476
rect 65588 15436 65597 15476
rect 64963 15435 65021 15436
rect 47875 15392 47933 15393
rect 68428 15392 68468 15520
rect 68515 15436 68524 15476
rect 68564 15436 72844 15476
rect 72884 15436 72893 15476
rect 73699 15436 73708 15476
rect 73748 15436 74956 15476
rect 74996 15436 76780 15476
rect 76820 15436 77356 15476
rect 77396 15436 77405 15476
rect 835 15352 844 15392
rect 884 15352 1516 15392
rect 1556 15352 1565 15392
rect 43075 15352 43084 15392
rect 43124 15352 46924 15392
rect 46964 15352 46973 15392
rect 47790 15352 47884 15392
rect 47924 15352 47933 15392
rect 47875 15351 47933 15352
rect 54412 15352 59020 15392
rect 59060 15352 59069 15392
rect 60163 15352 60172 15392
rect 60212 15352 67660 15392
rect 67700 15352 67709 15392
rect 68131 15352 68140 15392
rect 68180 15352 68468 15392
rect 54412 15308 54452 15352
rect 54595 15308 54653 15309
rect 61219 15308 61277 15309
rect 68524 15308 68564 15436
rect 75523 15308 75581 15309
rect 42883 15268 42892 15308
rect 42932 15268 43180 15308
rect 43220 15268 45004 15308
rect 45044 15268 54452 15308
rect 54510 15268 54604 15308
rect 54644 15268 61228 15308
rect 61268 15268 61277 15308
rect 61891 15268 61900 15308
rect 61940 15268 62476 15308
rect 62516 15268 65068 15308
rect 65108 15268 65117 15308
rect 67363 15268 67372 15308
rect 67412 15268 68564 15308
rect 69667 15268 69676 15308
rect 69716 15268 70444 15308
rect 70484 15268 70493 15308
rect 75331 15268 75340 15308
rect 75380 15268 75389 15308
rect 75523 15268 75532 15308
rect 75572 15268 76492 15308
rect 76532 15268 76541 15308
rect 54595 15267 54653 15268
rect 61219 15267 61277 15268
rect 75340 15224 75380 15268
rect 75523 15267 75581 15268
rect 32035 15184 32044 15224
rect 32084 15184 33292 15224
rect 33332 15184 34828 15224
rect 34868 15184 34877 15224
rect 53443 15184 53452 15224
rect 53492 15184 54700 15224
rect 54740 15184 58636 15224
rect 58676 15184 58685 15224
rect 60748 15184 65164 15224
rect 65204 15184 65213 15224
rect 70819 15184 70828 15224
rect 70868 15184 71884 15224
rect 71924 15184 71933 15224
rect 75340 15184 75572 15224
rect 60748 15140 60788 15184
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 15103 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 15489 15140
rect 27103 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 27489 15140
rect 39103 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 39489 15140
rect 51103 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 51489 15140
rect 51811 15100 51820 15140
rect 51860 15100 56908 15140
rect 56948 15100 56957 15140
rect 58435 15100 58444 15140
rect 58484 15100 60788 15140
rect 63103 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 63489 15140
rect 75103 15100 75112 15140
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75480 15100 75489 15140
rect 75532 15056 75572 15184
rect 77923 15100 77932 15140
rect 77972 15100 78796 15140
rect 78836 15100 78845 15140
rect 60451 15016 60460 15056
rect 60500 15016 61612 15056
rect 61652 15016 63284 15056
rect 63244 14972 63284 15016
rect 75340 15016 75572 15056
rect 75340 14972 75380 15016
rect 49411 14932 49420 14972
rect 49460 14932 51724 14972
rect 51764 14932 52436 14972
rect 52483 14932 52492 14972
rect 52532 14932 53452 14972
rect 53492 14932 62860 14972
rect 62900 14932 62909 14972
rect 63235 14932 63244 14972
rect 63284 14932 63293 14972
rect 65155 14932 65164 14972
rect 65204 14932 69100 14972
rect 69140 14932 69149 14972
rect 69475 14932 69484 14972
rect 69524 14932 70924 14972
rect 70964 14932 70973 14972
rect 71107 14932 71116 14972
rect 71156 14932 73439 14972
rect 73479 14932 73488 14972
rect 75331 14932 75340 14972
rect 75380 14932 75389 14972
rect 75436 14932 75916 14972
rect 75956 14932 75965 14972
rect 0 14888 80 14908
rect 52396 14888 52436 14932
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 38659 14848 38668 14888
rect 38708 14848 39916 14888
rect 39956 14848 39965 14888
rect 51523 14848 51532 14888
rect 51572 14848 51916 14888
rect 51956 14848 51965 14888
rect 52396 14848 53300 14888
rect 54595 14848 54604 14888
rect 54644 14848 55084 14888
rect 55124 14848 55133 14888
rect 60643 14848 60652 14888
rect 60692 14848 61036 14888
rect 61076 14848 61085 14888
rect 61315 14848 61324 14888
rect 61364 14848 61804 14888
rect 61844 14848 61853 14888
rect 70147 14848 70156 14888
rect 70196 14848 71212 14888
rect 71252 14848 72076 14888
rect 72116 14848 72748 14888
rect 72788 14848 72797 14888
rect 0 14828 80 14848
rect 53260 14804 53300 14848
rect 56707 14804 56765 14805
rect 60163 14804 60221 14805
rect 60355 14804 60413 14805
rect 70723 14804 70781 14805
rect 37315 14764 37324 14804
rect 37364 14764 37708 14804
rect 37748 14764 37757 14804
rect 45667 14764 45676 14804
rect 45716 14764 46636 14804
rect 46676 14764 46828 14804
rect 46868 14764 46877 14804
rect 51619 14764 51628 14804
rect 51668 14764 53108 14804
rect 53260 14764 53836 14804
rect 53876 14764 54260 14804
rect 56622 14764 56716 14804
rect 56756 14764 56765 14804
rect 57571 14764 57580 14804
rect 57620 14764 59692 14804
rect 59732 14764 59741 14804
rect 60078 14764 60172 14804
rect 60212 14764 60221 14804
rect 60270 14764 60364 14804
rect 60404 14764 69292 14804
rect 69332 14764 69341 14804
rect 70638 14764 70732 14804
rect 70772 14764 70781 14804
rect 43459 14720 43517 14721
rect 47875 14720 47933 14721
rect 34435 14680 34444 14720
rect 34484 14680 34924 14720
rect 34964 14680 34973 14720
rect 37411 14680 37420 14720
rect 37460 14680 38284 14720
rect 38324 14680 38333 14720
rect 42211 14680 42220 14720
rect 42260 14680 42700 14720
rect 42740 14680 43084 14720
rect 43124 14680 43133 14720
rect 43267 14680 43276 14720
rect 43316 14680 43468 14720
rect 43508 14680 43517 14720
rect 45571 14680 45580 14720
rect 45620 14680 47884 14720
rect 47924 14680 47933 14720
rect 48739 14680 48748 14720
rect 48788 14680 49324 14720
rect 49364 14680 49373 14720
rect 49987 14680 49996 14720
rect 50036 14680 51340 14720
rect 51380 14680 52052 14720
rect 43459 14679 43517 14680
rect 47875 14679 47933 14680
rect 52012 14636 52052 14680
rect 53068 14636 53108 14764
rect 54220 14720 54260 14764
rect 56707 14763 56765 14764
rect 60163 14763 60221 14764
rect 60355 14763 60413 14764
rect 70723 14763 70781 14764
rect 75436 14720 75476 14932
rect 76099 14764 76108 14804
rect 76148 14764 77836 14804
rect 77876 14764 77885 14804
rect 53155 14680 53164 14720
rect 53204 14680 53452 14720
rect 53492 14680 53501 14720
rect 53635 14680 53644 14720
rect 53684 14680 54028 14720
rect 54068 14680 54077 14720
rect 54211 14680 54220 14720
rect 54260 14680 54269 14720
rect 55459 14680 55468 14720
rect 55508 14680 56044 14720
rect 56084 14680 56093 14720
rect 56899 14680 56908 14720
rect 56948 14680 58636 14720
rect 58676 14680 58685 14720
rect 61411 14680 61420 14720
rect 61460 14680 62092 14720
rect 62132 14680 62141 14720
rect 67459 14680 67468 14720
rect 67508 14680 67948 14720
rect 67988 14680 67997 14720
rect 68611 14680 68620 14720
rect 68660 14680 69100 14720
rect 69140 14680 69772 14720
rect 69812 14680 69821 14720
rect 70339 14680 70348 14720
rect 70388 14680 71116 14720
rect 71156 14680 71165 14720
rect 73430 14680 73439 14720
rect 73479 14680 74188 14720
rect 74228 14680 74237 14720
rect 75427 14680 75436 14720
rect 75476 14680 75485 14720
rect 75907 14680 75916 14720
rect 75956 14680 76396 14720
rect 76436 14680 76445 14720
rect 76867 14680 76876 14720
rect 76916 14680 77740 14720
rect 77780 14680 77789 14720
rect 55468 14636 55508 14680
rect 37027 14596 37036 14636
rect 37076 14596 38956 14636
rect 38996 14596 39005 14636
rect 45379 14596 45388 14636
rect 45428 14596 45868 14636
rect 45908 14596 45917 14636
rect 52003 14596 52012 14636
rect 52052 14596 52061 14636
rect 53068 14596 53260 14636
rect 53300 14596 55508 14636
rect 38956 14384 38996 14596
rect 52099 14512 52108 14552
rect 52148 14512 52780 14552
rect 52820 14512 54508 14552
rect 54548 14512 54557 14552
rect 51619 14468 51677 14469
rect 44803 14428 44812 14468
rect 44852 14428 45484 14468
rect 45524 14428 45533 14468
rect 50851 14428 50860 14468
rect 50900 14428 51628 14468
rect 51668 14428 53068 14468
rect 53108 14428 53117 14468
rect 53539 14428 53548 14468
rect 53588 14428 54700 14468
rect 54740 14428 54749 14468
rect 51619 14427 51677 14428
rect 56044 14384 56084 14680
rect 60835 14596 60844 14636
rect 60884 14596 64876 14636
rect 64916 14596 64925 14636
rect 65059 14596 65068 14636
rect 65108 14596 67564 14636
rect 67604 14596 68236 14636
rect 68276 14596 68285 14636
rect 70435 14596 70444 14636
rect 70484 14596 71404 14636
rect 71444 14596 72460 14636
rect 72500 14596 72509 14636
rect 75619 14596 75628 14636
rect 75668 14596 76012 14636
rect 76052 14596 76061 14636
rect 76195 14596 76204 14636
rect 76244 14596 76780 14636
rect 76820 14596 76829 14636
rect 65644 14552 65684 14596
rect 58915 14512 58924 14552
rect 58964 14512 59116 14552
rect 59156 14512 59165 14552
rect 61987 14512 61996 14552
rect 62036 14512 62380 14552
rect 62420 14512 62429 14552
rect 64771 14512 64780 14552
rect 64820 14512 65452 14552
rect 65492 14512 65501 14552
rect 65635 14512 65644 14552
rect 65684 14512 65693 14552
rect 68419 14512 68428 14552
rect 68468 14512 69484 14552
rect 69524 14512 69533 14552
rect 70915 14512 70924 14552
rect 70964 14512 72172 14552
rect 72212 14512 72221 14552
rect 73027 14512 73036 14552
rect 73076 14512 73612 14552
rect 73652 14512 73661 14552
rect 63235 14428 63244 14468
rect 63284 14428 63532 14468
rect 63572 14428 63581 14468
rect 65155 14384 65213 14385
rect 66307 14384 66365 14385
rect 72547 14384 72605 14385
rect 76867 14384 76925 14385
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 16343 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 16729 14384
rect 28343 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 28729 14384
rect 38956 14344 39340 14384
rect 39380 14344 39389 14384
rect 40343 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 40729 14384
rect 41347 14344 41356 14384
rect 41396 14344 42604 14384
rect 42644 14344 43852 14384
rect 43892 14344 45772 14384
rect 45812 14344 45821 14384
rect 46915 14344 46924 14384
rect 46964 14344 48268 14384
rect 48308 14344 48317 14384
rect 52343 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 52729 14384
rect 53923 14344 53932 14384
rect 53972 14344 54412 14384
rect 54452 14344 54461 14384
rect 56035 14344 56044 14384
rect 56084 14344 56093 14384
rect 58819 14344 58828 14384
rect 58868 14344 60692 14384
rect 64343 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 64729 14384
rect 65059 14344 65068 14384
rect 65108 14344 65164 14384
rect 65204 14344 65213 14384
rect 66222 14344 66316 14384
rect 66356 14344 66365 14384
rect 70339 14344 70348 14384
rect 70388 14344 70636 14384
rect 70676 14344 72268 14384
rect 72308 14344 72317 14384
rect 72462 14344 72556 14384
rect 72596 14344 72605 14384
rect 76343 14344 76352 14384
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76720 14344 76729 14384
rect 76867 14344 76876 14384
rect 76916 14344 77260 14384
rect 77300 14344 77309 14384
rect 60652 14300 60692 14344
rect 65155 14343 65213 14344
rect 66307 14343 66365 14344
rect 72547 14343 72605 14344
rect 76867 14343 76925 14344
rect 40771 14260 40780 14300
rect 40820 14260 42316 14300
rect 42356 14260 42365 14300
rect 44419 14260 44428 14300
rect 44468 14260 46252 14300
rect 46292 14260 47212 14300
rect 47252 14260 47261 14300
rect 48643 14260 48652 14300
rect 48692 14260 49516 14300
rect 49556 14260 49565 14300
rect 49699 14260 49708 14300
rect 49748 14260 50092 14300
rect 50132 14260 52108 14300
rect 52148 14260 52876 14300
rect 52916 14260 52925 14300
rect 53251 14260 53260 14300
rect 53300 14260 54316 14300
rect 54356 14260 54365 14300
rect 54787 14260 54796 14300
rect 54836 14260 60268 14300
rect 60308 14260 60317 14300
rect 60652 14260 63724 14300
rect 63764 14260 63773 14300
rect 77539 14260 77548 14300
rect 77588 14260 78892 14300
rect 78932 14260 78941 14300
rect 39715 14176 39724 14216
rect 39764 14176 40396 14216
rect 40436 14176 41068 14216
rect 41108 14176 41117 14216
rect 41164 14176 42220 14216
rect 42260 14176 42269 14216
rect 45187 14176 45196 14216
rect 45236 14176 46060 14216
rect 46100 14176 46348 14216
rect 46388 14176 47020 14216
rect 47060 14176 47069 14216
rect 49123 14176 49132 14216
rect 49172 14176 59788 14216
rect 59828 14176 59837 14216
rect 61315 14176 61324 14216
rect 61364 14176 61708 14216
rect 61748 14176 61757 14216
rect 66019 14176 66028 14216
rect 66068 14176 66988 14216
rect 67028 14176 72652 14216
rect 72692 14176 72701 14216
rect 72835 14176 72844 14216
rect 72884 14176 73804 14216
rect 73844 14176 74284 14216
rect 74324 14176 74333 14216
rect 75331 14176 75340 14216
rect 75380 14176 75820 14216
rect 75860 14176 75869 14216
rect 78691 14176 78700 14216
rect 78740 14176 79372 14216
rect 79412 14176 79421 14216
rect 41164 14132 41204 14176
rect 60643 14132 60701 14133
rect 61411 14132 61469 14133
rect 39907 14092 39916 14132
rect 39956 14092 40300 14132
rect 40340 14092 40349 14132
rect 40675 14092 40684 14132
rect 40724 14092 41204 14132
rect 42019 14092 42028 14132
rect 42068 14092 42892 14132
rect 42932 14092 42941 14132
rect 45091 14092 45100 14132
rect 45140 14092 46732 14132
rect 46772 14092 46781 14132
rect 48355 14092 48364 14132
rect 48404 14092 49324 14132
rect 49364 14092 49373 14132
rect 49507 14092 49516 14132
rect 49556 14092 53260 14132
rect 53300 14092 53309 14132
rect 57379 14092 57388 14132
rect 57428 14092 60652 14132
rect 60692 14092 60701 14132
rect 61027 14092 61036 14132
rect 61076 14092 61420 14132
rect 61460 14092 61469 14132
rect 62083 14092 62092 14132
rect 62132 14092 63436 14132
rect 63476 14092 63485 14132
rect 69763 14092 69772 14132
rect 69812 14092 70924 14132
rect 70964 14092 70973 14132
rect 76588 14092 78508 14132
rect 78548 14092 78988 14132
rect 79028 14092 79037 14132
rect 60643 14091 60701 14092
rect 61411 14091 61469 14092
rect 0 14048 80 14068
rect 70924 14048 70964 14092
rect 75715 14048 75773 14049
rect 76588 14048 76628 14092
rect 77347 14048 77405 14049
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 34819 14008 34828 14048
rect 34868 14008 37036 14048
rect 37076 14008 37085 14048
rect 40195 14008 40204 14048
rect 40244 14008 40588 14048
rect 40628 14008 40637 14048
rect 41251 14008 41260 14048
rect 41300 14008 45580 14048
rect 45620 14008 45629 14048
rect 46531 14008 46540 14048
rect 46580 14008 47116 14048
rect 47156 14008 47980 14048
rect 48020 14008 48029 14048
rect 48451 14008 48460 14048
rect 48500 14008 49804 14048
rect 49844 14008 49853 14048
rect 52771 14008 52780 14048
rect 52820 14008 53740 14048
rect 53780 14008 55372 14048
rect 55412 14008 56620 14048
rect 56660 14008 57964 14048
rect 58004 14008 59212 14048
rect 59252 14008 61228 14048
rect 61268 14008 62284 14048
rect 62324 14008 64108 14048
rect 64148 14008 65836 14048
rect 65876 14008 65885 14048
rect 70147 14008 70156 14048
rect 70196 14008 70540 14048
rect 70580 14008 70589 14048
rect 70924 14008 71404 14048
rect 71444 14008 71453 14048
rect 71587 14008 71596 14048
rect 71636 14008 73132 14048
rect 73172 14008 73804 14048
rect 73844 14008 74092 14048
rect 74132 14008 74141 14048
rect 75235 14008 75244 14048
rect 75284 14008 75724 14048
rect 75764 14008 75773 14048
rect 76003 14008 76012 14048
rect 76052 14008 76204 14048
rect 76244 14008 76253 14048
rect 76579 14008 76588 14048
rect 76628 14008 76637 14048
rect 77262 14008 77356 14048
rect 77396 14008 77405 14048
rect 77635 14008 77644 14048
rect 77684 14008 78124 14048
rect 78164 14008 78173 14048
rect 0 13988 80 14008
rect 45580 13964 45620 14008
rect 75715 14007 75773 14008
rect 77347 14007 77405 14008
rect 1699 13924 1708 13964
rect 1748 13924 9388 13964
rect 9428 13924 9437 13964
rect 40867 13924 40876 13964
rect 40916 13924 42796 13964
rect 42836 13924 43276 13964
rect 43316 13924 43660 13964
rect 43700 13924 43709 13964
rect 45580 13924 48940 13964
rect 48980 13924 51724 13964
rect 51764 13924 51773 13964
rect 51820 13924 57388 13964
rect 57428 13924 57437 13964
rect 58051 13924 58060 13964
rect 58100 13924 58772 13964
rect 59971 13924 59980 13964
rect 60020 13924 60556 13964
rect 60596 13924 60605 13964
rect 62371 13924 62380 13964
rect 62420 13924 63284 13964
rect 63427 13924 63436 13964
rect 63476 13924 63820 13964
rect 63860 13924 63869 13964
rect 68995 13924 69004 13964
rect 69044 13924 69868 13964
rect 69908 13924 69917 13964
rect 71203 13924 71212 13964
rect 71252 13924 71692 13964
rect 71732 13924 71741 13964
rect 72259 13924 72268 13964
rect 72308 13924 74572 13964
rect 74612 13924 74621 13964
rect 76483 13924 76492 13964
rect 76532 13924 77452 13964
rect 77492 13924 77501 13964
rect 51820 13880 51860 13924
rect 58732 13880 58772 13924
rect 63244 13880 63284 13924
rect 63523 13880 63581 13881
rect 50179 13840 50188 13880
rect 50228 13840 51860 13880
rect 51907 13840 51916 13880
rect 51956 13840 52204 13880
rect 52244 13840 53356 13880
rect 53396 13840 54508 13880
rect 54548 13840 54557 13880
rect 57667 13840 57676 13880
rect 57716 13840 58252 13880
rect 58292 13840 58301 13880
rect 58723 13840 58732 13880
rect 58772 13840 59212 13880
rect 59252 13840 59261 13880
rect 60739 13840 60748 13880
rect 60788 13840 61516 13880
rect 61556 13840 62668 13880
rect 62708 13840 62717 13880
rect 63235 13840 63244 13880
rect 63284 13840 63532 13880
rect 63572 13840 63581 13880
rect 68611 13840 68620 13880
rect 68660 13840 69964 13880
rect 70004 13840 70013 13880
rect 70531 13840 70540 13880
rect 70580 13840 70828 13880
rect 70868 13840 70877 13880
rect 51916 13796 51956 13840
rect 63523 13839 63581 13840
rect 70147 13796 70205 13797
rect 42787 13756 42796 13796
rect 42836 13756 43084 13796
rect 43124 13756 43133 13796
rect 49027 13756 49036 13796
rect 49076 13756 50380 13796
rect 50420 13756 51956 13796
rect 55747 13756 55756 13796
rect 55796 13756 56524 13796
rect 56564 13756 56573 13796
rect 59779 13756 59788 13796
rect 59828 13756 60460 13796
rect 60500 13756 60509 13796
rect 61795 13756 61804 13796
rect 61844 13756 62380 13796
rect 62420 13756 62572 13796
rect 62612 13756 62621 13796
rect 68227 13756 68236 13796
rect 68276 13756 68812 13796
rect 68852 13756 69580 13796
rect 69620 13756 69629 13796
rect 70062 13756 70156 13796
rect 70196 13756 70205 13796
rect 70147 13755 70205 13756
rect 70819 13796 70877 13797
rect 70819 13756 70828 13796
rect 70868 13756 70924 13796
rect 70964 13756 70973 13796
rect 70819 13755 70877 13756
rect 60835 13712 60893 13713
rect 56323 13672 56332 13712
rect 56372 13672 58060 13712
rect 58100 13672 58828 13712
rect 58868 13672 58877 13712
rect 58924 13672 60844 13712
rect 60884 13672 60893 13712
rect 62659 13672 62668 13712
rect 62708 13672 65932 13712
rect 65972 13672 65981 13712
rect 58924 13628 58964 13672
rect 60835 13671 60893 13672
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 15103 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 15489 13628
rect 27103 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 27489 13628
rect 39103 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 39489 13628
rect 51103 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 51489 13628
rect 53260 13588 58964 13628
rect 60163 13588 60172 13628
rect 60212 13588 60252 13628
rect 63103 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 63489 13628
rect 68131 13588 68140 13628
rect 68180 13588 68812 13628
rect 68852 13588 68861 13628
rect 70627 13588 70636 13628
rect 70676 13588 71020 13628
rect 71060 13588 71069 13628
rect 75103 13588 75112 13628
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75480 13588 75489 13628
rect 78307 13588 78316 13628
rect 78356 13588 78365 13628
rect 53260 13544 53300 13588
rect 60172 13544 60212 13588
rect 78316 13544 78356 13588
rect 49411 13504 49420 13544
rect 49460 13504 53300 13544
rect 59971 13504 59980 13544
rect 60020 13504 64876 13544
rect 64916 13504 66700 13544
rect 66740 13504 67372 13544
rect 67412 13504 67421 13544
rect 71107 13504 71116 13544
rect 71156 13504 71165 13544
rect 78220 13504 78356 13544
rect 51427 13420 51436 13460
rect 51476 13420 51820 13460
rect 51860 13420 51869 13460
rect 54691 13420 54700 13460
rect 54740 13420 55180 13460
rect 55220 13420 55564 13460
rect 55604 13420 55613 13460
rect 57187 13420 57196 13460
rect 57236 13420 59116 13460
rect 59156 13420 59165 13460
rect 59683 13420 59692 13460
rect 59732 13420 60172 13460
rect 60212 13420 60364 13460
rect 60404 13420 61516 13460
rect 61556 13420 61996 13460
rect 62036 13420 62045 13460
rect 67171 13420 67180 13460
rect 67220 13420 67468 13460
rect 67508 13420 67517 13460
rect 67555 13376 67613 13377
rect 71116 13376 71156 13504
rect 73219 13420 73228 13460
rect 73268 13420 73996 13460
rect 74036 13420 74476 13460
rect 74516 13420 74525 13460
rect 76195 13420 76204 13460
rect 76244 13420 76588 13460
rect 76628 13420 76637 13460
rect 46723 13336 46732 13376
rect 46772 13336 47020 13376
rect 47060 13336 47069 13376
rect 49795 13336 49804 13376
rect 49844 13336 50284 13376
rect 50324 13336 50333 13376
rect 60259 13336 60268 13376
rect 60308 13336 62188 13376
rect 62228 13336 62237 13376
rect 63811 13336 63820 13376
rect 63860 13336 66220 13376
rect 66260 13336 66644 13376
rect 66787 13336 66796 13376
rect 66836 13336 67276 13376
rect 67316 13336 67325 13376
rect 67470 13336 67564 13376
rect 67604 13336 67613 13376
rect 70627 13336 70636 13376
rect 70676 13336 71156 13376
rect 71299 13336 71308 13376
rect 71348 13336 72172 13376
rect 72212 13336 72221 13376
rect 74179 13336 74188 13376
rect 74228 13336 76876 13376
rect 76916 13336 76925 13376
rect 77059 13336 77068 13376
rect 77108 13336 77548 13376
rect 77588 13336 77597 13376
rect 77740 13336 77836 13376
rect 77876 13336 77885 13376
rect 66604 13292 66644 13336
rect 67555 13335 67613 13336
rect 77740 13292 77780 13336
rect 78220 13292 78260 13504
rect 78307 13420 78316 13460
rect 78356 13420 78508 13460
rect 78548 13420 78557 13460
rect 835 13252 844 13292
rect 884 13252 1516 13292
rect 1556 13252 1565 13292
rect 1699 13252 1708 13292
rect 1748 13252 11980 13292
rect 12020 13252 12029 13292
rect 39235 13252 39244 13292
rect 39284 13252 40108 13292
rect 40148 13252 41740 13292
rect 41780 13252 41789 13292
rect 46828 13252 47788 13292
rect 47828 13252 57580 13292
rect 57620 13252 57629 13292
rect 61603 13252 61612 13292
rect 61652 13252 62092 13292
rect 62132 13252 62141 13292
rect 66499 13252 66508 13292
rect 66548 13252 66557 13292
rect 66604 13252 68044 13292
rect 68084 13252 68093 13292
rect 68323 13252 68332 13292
rect 68372 13252 69004 13292
rect 69044 13252 69964 13292
rect 70004 13252 70348 13292
rect 70388 13252 70397 13292
rect 73420 13252 76012 13292
rect 76052 13252 76061 13292
rect 77155 13252 77164 13292
rect 77204 13252 77780 13292
rect 78211 13252 78220 13292
rect 78260 13252 78269 13292
rect 0 13208 80 13228
rect 46828 13208 46868 13252
rect 51619 13208 51677 13209
rect 65251 13208 65309 13209
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 38755 13168 38764 13208
rect 38804 13168 39532 13208
rect 39572 13168 39581 13208
rect 41347 13168 41356 13208
rect 41396 13168 41836 13208
rect 41876 13168 41885 13208
rect 44995 13168 45004 13208
rect 45044 13168 45292 13208
rect 45332 13168 45868 13208
rect 45908 13168 45917 13208
rect 46819 13168 46828 13208
rect 46868 13168 46877 13208
rect 47683 13168 47692 13208
rect 47732 13168 49132 13208
rect 49172 13168 49181 13208
rect 50371 13168 50380 13208
rect 50420 13168 50956 13208
rect 50996 13168 51005 13208
rect 51534 13168 51628 13208
rect 51668 13168 51677 13208
rect 53827 13168 53836 13208
rect 53876 13168 54316 13208
rect 54356 13168 54365 13208
rect 55267 13168 55276 13208
rect 55316 13168 55756 13208
rect 55796 13168 55805 13208
rect 56419 13168 56428 13208
rect 56468 13168 57292 13208
rect 57332 13168 57341 13208
rect 57955 13168 57964 13208
rect 58004 13168 58924 13208
rect 58964 13168 58973 13208
rect 59587 13168 59596 13208
rect 59636 13168 61708 13208
rect 61748 13168 61757 13208
rect 62947 13168 62956 13208
rect 62996 13168 63820 13208
rect 63860 13168 63869 13208
rect 65166 13168 65260 13208
rect 65300 13168 65309 13208
rect 66508 13208 66548 13252
rect 66508 13168 66932 13208
rect 67075 13168 67084 13208
rect 67124 13168 67660 13208
rect 67700 13168 68140 13208
rect 68180 13168 68189 13208
rect 68419 13168 68428 13208
rect 68468 13168 69868 13208
rect 69908 13168 70732 13208
rect 70772 13168 71116 13208
rect 71156 13168 71596 13208
rect 71636 13168 71645 13208
rect 71971 13168 71980 13208
rect 72020 13168 72652 13208
rect 72692 13168 72701 13208
rect 0 13148 80 13168
rect 47692 13124 47732 13168
rect 51619 13167 51677 13168
rect 54316 13124 54356 13168
rect 65251 13167 65309 13168
rect 66787 13124 66845 13125
rect 44611 13084 44620 13124
rect 44660 13084 44908 13124
rect 44948 13084 44957 13124
rect 46531 13084 46540 13124
rect 46580 13084 47732 13124
rect 51715 13084 51724 13124
rect 51764 13084 51916 13124
rect 51956 13084 51965 13124
rect 53635 13084 53644 13124
rect 53684 13084 53693 13124
rect 54316 13084 55468 13124
rect 55508 13084 55517 13124
rect 55843 13084 55852 13124
rect 55892 13084 56524 13124
rect 56564 13084 56573 13124
rect 59107 13084 59116 13124
rect 59156 13084 63628 13124
rect 63668 13084 63677 13124
rect 65347 13084 65356 13124
rect 65396 13084 65740 13124
rect 65780 13084 66412 13124
rect 66452 13084 66461 13124
rect 66702 13084 66796 13124
rect 66836 13084 66845 13124
rect 66892 13124 66932 13168
rect 73420 13124 73460 13252
rect 73795 13168 73804 13208
rect 73844 13168 75436 13208
rect 75476 13168 75956 13208
rect 77731 13168 77740 13208
rect 77780 13168 78316 13208
rect 78356 13168 78700 13208
rect 78740 13168 78749 13208
rect 75916 13124 75956 13168
rect 66892 13084 66988 13124
rect 67028 13084 67563 13124
rect 67603 13084 67612 13124
rect 68515 13084 68524 13124
rect 68564 13084 68573 13124
rect 68899 13084 68908 13124
rect 68948 13084 71404 13124
rect 71444 13084 71788 13124
rect 71828 13084 73460 13124
rect 75907 13084 75916 13124
rect 75956 13084 78124 13124
rect 78164 13084 78173 13124
rect 53644 13040 53684 13084
rect 66787 13083 66845 13084
rect 68524 13040 68564 13084
rect 835 13000 844 13040
rect 884 13000 1516 13040
rect 1556 13000 1565 13040
rect 44803 13000 44812 13040
rect 44852 13000 45484 13040
rect 45524 13000 45533 13040
rect 45859 13000 45868 13040
rect 45908 13000 46444 13040
rect 46484 13000 46493 13040
rect 50275 13000 50284 13040
rect 50324 13000 51244 13040
rect 51284 13000 55084 13040
rect 55124 13000 55700 13040
rect 55747 13000 55756 13040
rect 55796 13000 56332 13040
rect 56372 13000 56381 13040
rect 61219 13000 61228 13040
rect 61268 13000 61516 13040
rect 61556 13000 61565 13040
rect 62083 13000 62092 13040
rect 62132 13000 62668 13040
rect 62708 13000 62717 13040
rect 65892 13000 65932 13040
rect 65972 13000 65981 13040
rect 68227 13000 68236 13040
rect 68276 13000 68564 13040
rect 55660 12956 55700 13000
rect 60451 12956 60509 12957
rect 65932 12956 65972 13000
rect 67555 12956 67613 12957
rect 51715 12916 51724 12956
rect 51764 12916 52204 12956
rect 52244 12916 52253 12956
rect 55651 12916 55660 12956
rect 55700 12916 55740 12956
rect 60355 12916 60364 12956
rect 60404 12916 60460 12956
rect 60500 12916 60509 12956
rect 60643 12916 60652 12956
rect 60692 12916 63532 12956
rect 63572 12916 64780 12956
rect 64820 12916 64829 12956
rect 65539 12916 65548 12956
rect 65588 12916 65972 12956
rect 66595 12916 66604 12956
rect 66644 12916 67564 12956
rect 67604 12916 67613 12956
rect 72067 12916 72076 12956
rect 72116 12916 72460 12956
rect 72500 12916 72940 12956
rect 72980 12916 72989 12956
rect 76195 12916 76204 12956
rect 76244 12916 77260 12956
rect 77300 12916 77309 12956
rect 60451 12915 60509 12916
rect 67555 12915 67613 12916
rect 75715 12872 75773 12873
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 16343 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 16729 12872
rect 28343 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 28729 12872
rect 40343 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 40729 12872
rect 46147 12832 46156 12872
rect 46196 12832 48076 12872
rect 48116 12832 48125 12872
rect 52343 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 52729 12872
rect 62371 12832 62380 12872
rect 62420 12832 62956 12872
rect 62996 12832 63005 12872
rect 64343 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 64729 12872
rect 69379 12832 69388 12872
rect 69428 12832 75724 12872
rect 75764 12832 76244 12872
rect 76343 12832 76352 12872
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76720 12832 76729 12872
rect 75715 12831 75773 12832
rect 45379 12748 45388 12788
rect 45428 12748 45964 12788
rect 46004 12748 46013 12788
rect 48259 12748 48268 12788
rect 48308 12748 49804 12788
rect 49844 12748 49853 12788
rect 52771 12748 52780 12788
rect 52820 12748 61324 12788
rect 61364 12748 61373 12788
rect 63715 12748 63724 12788
rect 63764 12748 69196 12788
rect 69236 12748 69245 12788
rect 74851 12748 74860 12788
rect 74900 12748 75436 12788
rect 75476 12748 75485 12788
rect 76204 12704 76244 12832
rect 44035 12664 44044 12704
rect 44084 12664 44620 12704
rect 44660 12664 44669 12704
rect 48067 12664 48076 12704
rect 48116 12664 49516 12704
rect 49556 12664 49900 12704
rect 49940 12664 52588 12704
rect 52628 12664 52637 12704
rect 55555 12664 55564 12704
rect 55604 12664 56236 12704
rect 56276 12664 56285 12704
rect 59491 12664 59500 12704
rect 59540 12664 60076 12704
rect 60116 12664 60125 12704
rect 67747 12664 67756 12704
rect 67796 12664 68620 12704
rect 68660 12664 68669 12704
rect 72739 12664 72748 12704
rect 72788 12664 73460 12704
rect 73699 12664 73708 12704
rect 73748 12664 73900 12704
rect 73940 12664 75052 12704
rect 75092 12664 75101 12704
rect 76204 12664 76396 12704
rect 76436 12664 76445 12704
rect 41539 12580 41548 12620
rect 41588 12580 43948 12620
rect 43988 12580 44428 12620
rect 44468 12580 44477 12620
rect 45955 12580 45964 12620
rect 46004 12580 46013 12620
rect 48163 12580 48172 12620
rect 48212 12580 49708 12620
rect 49748 12580 49757 12620
rect 56035 12580 56044 12620
rect 56084 12580 56428 12620
rect 56468 12580 56477 12620
rect 56611 12580 56620 12620
rect 56660 12580 57196 12620
rect 57236 12580 57245 12620
rect 61891 12580 61900 12620
rect 61940 12580 62092 12620
rect 62132 12580 62141 12620
rect 66211 12580 66220 12620
rect 66260 12580 67180 12620
rect 67220 12580 67948 12620
rect 67988 12580 67997 12620
rect 69475 12580 69484 12620
rect 69524 12580 70636 12620
rect 70676 12580 70685 12620
rect 43267 12496 43276 12536
rect 43316 12496 43756 12536
rect 43796 12496 43805 12536
rect 45964 12452 46004 12580
rect 52195 12536 52253 12537
rect 46051 12496 46060 12536
rect 46100 12496 47212 12536
rect 47252 12496 48652 12536
rect 48692 12496 48701 12536
rect 49987 12496 49996 12536
rect 50036 12496 50572 12536
rect 50612 12496 50621 12536
rect 51043 12496 51052 12536
rect 51092 12496 52204 12536
rect 52244 12496 52253 12536
rect 56131 12496 56140 12536
rect 56180 12496 56716 12536
rect 56756 12496 56765 12536
rect 57091 12496 57100 12536
rect 57140 12496 58060 12536
rect 58100 12496 58109 12536
rect 59299 12496 59308 12536
rect 59348 12496 60652 12536
rect 60692 12496 60701 12536
rect 63619 12496 63628 12536
rect 63668 12496 65164 12536
rect 65204 12496 65213 12536
rect 65635 12496 65644 12536
rect 65684 12496 68428 12536
rect 68468 12496 68908 12536
rect 68948 12496 68957 12536
rect 52195 12495 52253 12496
rect 73420 12452 73460 12664
rect 76780 12536 76820 12916
rect 78211 12580 78220 12620
rect 78260 12580 78300 12620
rect 78220 12536 78260 12580
rect 76771 12496 76780 12536
rect 76820 12496 76829 12536
rect 77827 12496 77836 12536
rect 77876 12496 79372 12536
rect 79412 12496 79421 12536
rect 1699 12412 1708 12452
rect 1748 12412 10252 12452
rect 10292 12412 10301 12452
rect 45964 12412 49900 12452
rect 49940 12412 49949 12452
rect 51139 12412 51148 12452
rect 51188 12412 51628 12452
rect 51668 12412 51677 12452
rect 56803 12412 56812 12452
rect 56852 12412 64204 12452
rect 64244 12412 64253 12452
rect 64771 12412 64780 12452
rect 64820 12412 66604 12452
rect 66644 12412 66653 12452
rect 68035 12412 68044 12452
rect 68084 12412 68812 12452
rect 68852 12412 70060 12452
rect 70100 12412 70109 12452
rect 73315 12412 73324 12452
rect 73364 12412 77740 12452
rect 77780 12412 77789 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 44035 12328 44044 12368
rect 44084 12328 44428 12368
rect 44468 12328 44477 12368
rect 0 12308 80 12328
rect 45964 12284 46004 12412
rect 77347 12328 77356 12368
rect 77396 12328 77405 12368
rect 61027 12284 61085 12285
rect 43843 12244 43852 12284
rect 43892 12244 44716 12284
rect 44756 12244 46004 12284
rect 48931 12244 48940 12284
rect 48980 12244 61036 12284
rect 61076 12244 61085 12284
rect 77356 12284 77396 12328
rect 77356 12244 78124 12284
rect 78164 12244 78412 12284
rect 78452 12244 78461 12284
rect 61027 12243 61085 12244
rect 59011 12200 59069 12201
rect 64771 12200 64829 12201
rect 77347 12200 77405 12201
rect 43267 12160 43276 12200
rect 43316 12160 43468 12200
rect 43508 12160 59020 12200
rect 59060 12160 59069 12200
rect 59011 12159 59069 12160
rect 59116 12160 64780 12200
rect 64820 12160 64829 12200
rect 77262 12160 77356 12200
rect 77396 12160 77405 12200
rect 44611 12116 44669 12117
rect 59116 12116 59156 12160
rect 64771 12159 64829 12160
rect 77347 12159 77405 12160
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 15103 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 15489 12116
rect 27103 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 27489 12116
rect 39103 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 39489 12116
rect 43555 12076 43564 12116
rect 43604 12076 43700 12116
rect 44526 12076 44620 12116
rect 44660 12076 44669 12116
rect 51103 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 51489 12116
rect 58051 12076 58060 12116
rect 58100 12076 59156 12116
rect 63103 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 63489 12116
rect 75103 12076 75112 12116
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75480 12076 75489 12116
rect 43660 11780 43700 12076
rect 44611 12075 44669 12076
rect 56131 12032 56189 12033
rect 56046 11992 56140 12032
rect 56180 11992 58636 12032
rect 58676 11992 58685 12032
rect 63340 11992 66124 12032
rect 66164 11992 66173 12032
rect 56131 11991 56189 11992
rect 56035 11948 56093 11949
rect 51715 11908 51724 11948
rect 51764 11908 53740 11948
rect 53780 11908 53789 11948
rect 55950 11908 56044 11948
rect 56084 11908 56093 11948
rect 56227 11908 56236 11948
rect 56276 11908 56524 11948
rect 56564 11908 56573 11948
rect 61699 11908 61708 11948
rect 61748 11908 61788 11948
rect 56035 11907 56093 11908
rect 61708 11864 61748 11908
rect 63340 11864 63380 11992
rect 74467 11908 74476 11948
rect 74516 11908 75052 11948
rect 75092 11908 75101 11948
rect 45763 11824 45772 11864
rect 45812 11824 46924 11864
rect 46964 11824 46973 11864
rect 53260 11824 54796 11864
rect 54836 11824 54845 11864
rect 55267 11824 55276 11864
rect 55316 11824 56620 11864
rect 56660 11824 57100 11864
rect 57140 11824 57149 11864
rect 61027 11824 61036 11864
rect 61076 11824 62380 11864
rect 62420 11824 63380 11864
rect 64387 11824 64396 11864
rect 64436 11824 65548 11864
rect 65588 11824 65597 11864
rect 71971 11824 71980 11864
rect 72020 11824 72844 11864
rect 72884 11824 73132 11864
rect 73172 11824 73181 11864
rect 53260 11780 53300 11824
rect 835 11740 844 11780
rect 884 11740 1516 11780
rect 1556 11740 1565 11780
rect 1699 11740 1708 11780
rect 1748 11740 6124 11780
rect 6164 11740 6173 11780
rect 43651 11740 43660 11780
rect 43700 11740 53300 11780
rect 53347 11740 53356 11780
rect 53396 11740 55468 11780
rect 55508 11740 56428 11780
rect 56468 11740 56477 11780
rect 61699 11740 61708 11780
rect 61748 11740 61996 11780
rect 62036 11740 62188 11780
rect 62228 11740 65972 11780
rect 67459 11740 67468 11780
rect 67508 11740 67517 11780
rect 73315 11740 73324 11780
rect 73364 11740 73652 11780
rect 76003 11740 76012 11780
rect 76052 11740 76684 11780
rect 76724 11740 77452 11780
rect 77492 11740 77501 11780
rect 60163 11696 60221 11697
rect 65932 11696 65972 11740
rect 50947 11656 50956 11696
rect 50996 11656 51820 11696
rect 51860 11656 51869 11696
rect 55939 11656 55948 11696
rect 55988 11656 55997 11696
rect 56044 11656 56332 11696
rect 56372 11656 56381 11696
rect 59107 11656 59116 11696
rect 59156 11656 60172 11696
rect 60212 11656 60221 11696
rect 61411 11656 61420 11696
rect 61460 11656 63148 11696
rect 63188 11656 63197 11696
rect 64867 11656 64876 11696
rect 64916 11656 65740 11696
rect 65780 11656 65789 11696
rect 65923 11656 65932 11696
rect 65972 11656 67084 11696
rect 67124 11656 67133 11696
rect 844 11572 1420 11612
rect 1460 11572 1469 11612
rect 41251 11572 41260 11612
rect 41300 11572 42412 11612
rect 42452 11572 42461 11612
rect 45868 11572 46252 11612
rect 46292 11572 46301 11612
rect 51052 11572 51532 11612
rect 51572 11572 51581 11612
rect 0 11528 80 11548
rect 844 11528 884 11572
rect 45868 11528 45908 11572
rect 51052 11528 51092 11572
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 835 11488 844 11528
rect 884 11488 893 11528
rect 43843 11488 43852 11528
rect 43892 11488 44428 11528
rect 44468 11488 44477 11528
rect 45859 11488 45868 11528
rect 45908 11488 45917 11528
rect 51043 11488 51052 11528
rect 51092 11488 51101 11528
rect 0 11468 80 11488
rect 55948 11444 55988 11656
rect 56044 11528 56084 11656
rect 60163 11655 60221 11656
rect 67468 11612 67508 11740
rect 73612 11696 73652 11740
rect 68035 11656 68044 11696
rect 68084 11656 68332 11696
rect 68372 11656 68381 11696
rect 72547 11656 72556 11696
rect 72596 11656 73508 11696
rect 73548 11656 73557 11696
rect 73603 11656 73612 11696
rect 73652 11656 73661 11696
rect 73795 11656 73804 11696
rect 73844 11656 77644 11696
rect 77684 11656 77693 11696
rect 73804 11612 73844 11656
rect 61795 11572 61804 11612
rect 61844 11572 62284 11612
rect 62324 11572 62333 11612
rect 63331 11572 63340 11612
rect 63380 11572 63724 11612
rect 63764 11572 63773 11612
rect 66115 11572 66124 11612
rect 66164 11572 67604 11612
rect 69475 11572 69484 11612
rect 69524 11572 70252 11612
rect 70292 11572 70301 11612
rect 72451 11572 72460 11612
rect 72500 11572 73844 11612
rect 56035 11488 56044 11528
rect 56084 11488 56093 11528
rect 66211 11488 66220 11528
rect 66260 11488 66892 11528
rect 66932 11488 66941 11528
rect 67564 11444 67604 11572
rect 72067 11488 72076 11528
rect 72116 11488 72364 11528
rect 72404 11488 72413 11528
rect 55948 11404 56180 11444
rect 67555 11404 67564 11444
rect 67604 11404 67613 11444
rect 72259 11404 72268 11444
rect 72308 11404 73172 11444
rect 56140 11360 56180 11404
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 16343 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 16729 11360
rect 28343 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 28729 11360
rect 40343 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 40729 11360
rect 42691 11320 42700 11360
rect 42740 11320 43276 11360
rect 43316 11320 43325 11360
rect 52343 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 52729 11360
rect 55555 11320 55564 11360
rect 55604 11320 55948 11360
rect 55988 11320 55997 11360
rect 56131 11320 56140 11360
rect 56180 11320 56189 11360
rect 64343 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 64729 11360
rect 70435 11320 70444 11360
rect 70484 11320 72748 11360
rect 72788 11320 72797 11360
rect 73132 11276 73172 11404
rect 76343 11320 76352 11360
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76720 11320 76729 11360
rect 41443 11236 41452 11276
rect 41492 11236 44332 11276
rect 44372 11236 44381 11276
rect 47107 11236 47116 11276
rect 47156 11236 50188 11276
rect 50228 11236 50237 11276
rect 54115 11236 54124 11276
rect 54164 11236 61132 11276
rect 61172 11236 61181 11276
rect 66979 11236 66988 11276
rect 67028 11236 67468 11276
rect 67508 11236 67852 11276
rect 67892 11236 67901 11276
rect 73123 11236 73132 11276
rect 73172 11236 73181 11276
rect 63523 11192 63581 11193
rect 51619 11152 51628 11192
rect 51668 11152 52780 11192
rect 52820 11152 52829 11192
rect 55171 11152 55180 11192
rect 55220 11152 58252 11192
rect 58292 11152 58444 11192
rect 58484 11152 58493 11192
rect 59683 11152 59692 11192
rect 59732 11152 61324 11192
rect 61364 11152 61373 11192
rect 62083 11152 62092 11192
rect 62132 11152 62764 11192
rect 62804 11152 62813 11192
rect 63438 11152 63532 11192
rect 63572 11152 63581 11192
rect 64771 11152 64780 11192
rect 64820 11152 66220 11192
rect 66260 11152 66269 11192
rect 77059 11152 77068 11192
rect 77108 11152 77932 11192
rect 77972 11152 77981 11192
rect 63523 11151 63581 11152
rect 42787 11068 42796 11108
rect 42836 11068 43220 11108
rect 43267 11068 43276 11108
rect 43316 11068 43660 11108
rect 43700 11068 43709 11108
rect 44419 11068 44428 11108
rect 44468 11068 46252 11108
rect 46292 11068 46301 11108
rect 49315 11068 49324 11108
rect 49364 11068 50380 11108
rect 50420 11068 60940 11108
rect 60980 11068 60989 11108
rect 61891 11068 61900 11108
rect 61940 11068 62476 11108
rect 62516 11068 62525 11108
rect 43180 11024 43220 11068
rect 42595 10984 42604 11024
rect 42644 10984 42988 11024
rect 43028 10984 43037 11024
rect 43180 10984 43756 11024
rect 43796 10984 43805 11024
rect 45667 10984 45676 11024
rect 45716 10984 46348 11024
rect 46388 10984 46397 11024
rect 52099 10984 52108 11024
rect 52148 10984 52876 11024
rect 52916 10984 52925 11024
rect 54988 10984 55180 11024
rect 55220 10984 55229 11024
rect 55747 10984 55756 11024
rect 55796 10984 56236 11024
rect 56276 10984 56285 11024
rect 57475 10984 57484 11024
rect 57524 10984 57772 11024
rect 57812 10984 60172 11024
rect 60212 10984 60221 11024
rect 62563 10984 62572 11024
rect 62612 10984 63436 11024
rect 63476 10984 63485 11024
rect 64003 10984 64012 11024
rect 64052 10984 65932 11024
rect 65972 10984 65981 11024
rect 69955 10984 69964 11024
rect 70004 10984 71884 11024
rect 71924 10984 71933 11024
rect 74659 10984 74668 11024
rect 74708 10984 77164 11024
rect 77204 10984 77213 11024
rect 43363 10940 43421 10941
rect 43278 10900 43372 10940
rect 43412 10900 43421 10940
rect 48835 10900 48844 10940
rect 48884 10900 50284 10940
rect 50324 10900 50996 10940
rect 51715 10900 51724 10940
rect 51764 10900 52012 10940
rect 52052 10900 52061 10940
rect 52387 10900 52396 10940
rect 52436 10900 54796 10940
rect 54836 10900 54845 10940
rect 43363 10899 43421 10900
rect 50956 10856 50996 10900
rect 54988 10856 55028 10984
rect 55075 10900 55084 10940
rect 55124 10900 58636 10940
rect 58676 10900 58685 10940
rect 62083 10900 62092 10940
rect 62132 10900 62141 10940
rect 68899 10900 68908 10940
rect 68948 10900 73516 10940
rect 73556 10900 74284 10940
rect 74324 10900 78604 10940
rect 78644 10900 78653 10940
rect 56707 10856 56765 10857
rect 62092 10856 62132 10900
rect 66691 10856 66749 10857
rect 48259 10816 48268 10856
rect 48308 10816 50860 10856
rect 50900 10816 50909 10856
rect 50956 10816 55028 10856
rect 55939 10816 55948 10856
rect 55988 10816 56716 10856
rect 56756 10816 56765 10856
rect 60643 10816 60652 10856
rect 60692 10816 61900 10856
rect 61940 10816 61949 10856
rect 62092 10816 63532 10856
rect 63572 10816 63581 10856
rect 66691 10816 66700 10856
rect 66740 10816 66796 10856
rect 66836 10816 66845 10856
rect 56707 10815 56765 10816
rect 66691 10815 66749 10816
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 43363 10732 43372 10772
rect 43412 10732 44140 10772
rect 44180 10732 44189 10772
rect 51331 10732 51340 10772
rect 51380 10732 51724 10772
rect 51764 10732 51773 10772
rect 54787 10732 54796 10772
rect 54836 10732 56908 10772
rect 56948 10732 56957 10772
rect 61987 10732 61996 10772
rect 62036 10732 62284 10772
rect 62324 10732 63052 10772
rect 63092 10732 63101 10772
rect 77347 10732 77356 10772
rect 77396 10732 77740 10772
rect 77780 10732 78028 10772
rect 78068 10732 78077 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 56035 10688 56093 10689
rect 0 10648 692 10688
rect 52003 10648 52012 10688
rect 52052 10648 55948 10688
rect 55988 10648 56044 10688
rect 56084 10648 56112 10688
rect 59779 10648 59788 10688
rect 59828 10648 66124 10688
rect 66164 10648 66173 10688
rect 0 10628 80 10648
rect 56035 10647 56093 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 15103 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 15489 10604
rect 27103 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 27489 10604
rect 39103 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 39489 10604
rect 51103 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 51489 10604
rect 59587 10564 59596 10604
rect 59636 10564 59980 10604
rect 60020 10564 60556 10604
rect 60596 10564 60605 10604
rect 63103 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 63489 10604
rect 64963 10564 64972 10604
rect 65012 10564 69676 10604
rect 69716 10564 69725 10604
rect 75103 10564 75112 10604
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75480 10564 75489 10604
rect 52867 10480 52876 10520
rect 52916 10480 54124 10520
rect 54164 10480 54173 10520
rect 66403 10480 66412 10520
rect 66452 10480 69292 10520
rect 69332 10480 69341 10520
rect 70051 10480 70060 10520
rect 70100 10480 73036 10520
rect 73076 10480 73085 10520
rect 47779 10396 47788 10436
rect 47828 10396 48940 10436
rect 48980 10396 48989 10436
rect 51235 10396 51244 10436
rect 51284 10396 56236 10436
rect 56276 10396 56285 10436
rect 61123 10396 61132 10436
rect 61172 10396 64684 10436
rect 64724 10396 64733 10436
rect 68323 10396 68332 10436
rect 68372 10396 70348 10436
rect 70388 10396 70397 10436
rect 73795 10396 73804 10436
rect 73844 10396 74764 10436
rect 74804 10396 75244 10436
rect 75284 10396 75293 10436
rect 68515 10352 68573 10353
rect 835 10312 844 10352
rect 884 10312 1516 10352
rect 1556 10312 1565 10352
rect 42595 10312 42604 10352
rect 42644 10312 43276 10352
rect 43316 10312 43325 10352
rect 45091 10312 45100 10352
rect 45140 10312 45772 10352
rect 45812 10312 45821 10352
rect 53443 10312 53452 10352
rect 53492 10312 54988 10352
rect 55028 10312 55037 10352
rect 56515 10312 56524 10352
rect 56564 10312 56908 10352
rect 56948 10312 56957 10352
rect 62755 10312 62764 10352
rect 62804 10312 68236 10352
rect 68276 10312 68285 10352
rect 68430 10312 68524 10352
rect 68564 10312 68573 10352
rect 68899 10312 68908 10352
rect 68948 10312 69292 10352
rect 69332 10312 69341 10352
rect 73123 10312 73132 10352
rect 73172 10312 73324 10352
rect 73364 10312 73373 10352
rect 76675 10312 76684 10352
rect 76724 10312 78124 10352
rect 78164 10312 78173 10352
rect 68515 10311 68573 10312
rect 1699 10228 1708 10268
rect 1748 10228 3628 10268
rect 3668 10228 3677 10268
rect 43459 10228 43468 10268
rect 43508 10228 45388 10268
rect 45428 10228 45964 10268
rect 46004 10228 46013 10268
rect 50947 10228 50956 10268
rect 50996 10228 52012 10268
rect 52052 10228 52061 10268
rect 55075 10228 55084 10268
rect 55124 10228 55852 10268
rect 55892 10228 55901 10268
rect 56227 10228 56236 10268
rect 56276 10228 58444 10268
rect 58484 10228 58493 10268
rect 60163 10228 60172 10268
rect 60212 10228 60460 10268
rect 60500 10228 60509 10268
rect 64675 10228 64684 10268
rect 64724 10228 66604 10268
rect 66644 10228 66653 10268
rect 69091 10228 69100 10268
rect 69140 10228 70060 10268
rect 70100 10228 70109 10268
rect 77059 10228 77068 10268
rect 77108 10228 77932 10268
rect 77972 10228 77981 10268
rect 43075 10144 43084 10184
rect 43124 10144 43564 10184
rect 43604 10144 44044 10184
rect 44084 10144 44093 10184
rect 44227 10144 44236 10184
rect 44276 10144 44812 10184
rect 44852 10144 44861 10184
rect 44995 10144 45004 10184
rect 45044 10144 47116 10184
rect 47156 10144 47165 10184
rect 50467 10144 50476 10184
rect 50516 10144 51148 10184
rect 51188 10144 51197 10184
rect 51427 10144 51436 10184
rect 51476 10144 52204 10184
rect 52244 10144 52253 10184
rect 55459 10144 55468 10184
rect 55508 10144 56332 10184
rect 56372 10144 56381 10184
rect 58243 10144 58252 10184
rect 58292 10144 58732 10184
rect 58772 10144 59500 10184
rect 59540 10144 59549 10184
rect 61891 10144 61900 10184
rect 61940 10144 64012 10184
rect 64052 10144 64061 10184
rect 64867 10144 64876 10184
rect 64916 10144 66412 10184
rect 66452 10144 66461 10184
rect 69187 10144 69196 10184
rect 69236 10144 70252 10184
rect 70292 10144 70301 10184
rect 71683 10144 71692 10184
rect 71732 10144 76972 10184
rect 77012 10144 77021 10184
rect 47011 10100 47069 10101
rect 66499 10100 66557 10101
rect 68419 10100 68477 10101
rect 71011 10100 71069 10101
rect 75811 10100 75869 10101
rect 43843 10060 43852 10100
rect 43892 10060 46444 10100
rect 46484 10060 46636 10100
rect 46676 10060 46685 10100
rect 46926 10060 47020 10100
rect 47060 10060 47069 10100
rect 49987 10060 49996 10100
rect 50036 10060 51340 10100
rect 51380 10060 51389 10100
rect 51523 10060 51532 10100
rect 51572 10060 51916 10100
rect 51956 10060 51965 10100
rect 52963 10060 52972 10100
rect 53012 10060 54700 10100
rect 54740 10060 54749 10100
rect 55171 10060 55180 10100
rect 55220 10060 55372 10100
rect 55412 10060 55421 10100
rect 58627 10060 58636 10100
rect 58676 10060 59116 10100
rect 59156 10060 59165 10100
rect 59299 10060 59308 10100
rect 59348 10060 59636 10100
rect 60451 10060 60460 10100
rect 60500 10060 62764 10100
rect 62804 10060 63148 10100
rect 63188 10060 63197 10100
rect 66414 10060 66508 10100
rect 66548 10060 66557 10100
rect 68334 10060 68428 10100
rect 68468 10060 68477 10100
rect 70926 10060 71020 10100
rect 71060 10060 71069 10100
rect 75726 10060 75820 10100
rect 75860 10060 75869 10100
rect 47011 10059 47069 10060
rect 43363 10016 43421 10017
rect 59596 10016 59636 10060
rect 66499 10059 66557 10060
rect 68419 10059 68477 10060
rect 71011 10059 71069 10060
rect 75811 10059 75869 10060
rect 42979 9976 42988 10016
rect 43028 9976 43220 10016
rect 0 9848 80 9868
rect 43180 9848 43220 9976
rect 43363 9976 43372 10016
rect 43412 9976 46252 10016
rect 46292 9976 46301 10016
rect 54787 9976 54796 10016
rect 54836 9976 56044 10016
rect 56084 9976 56093 10016
rect 58147 9976 58156 10016
rect 58196 9976 58924 10016
rect 58964 9976 59404 10016
rect 59444 9976 59453 10016
rect 59587 9976 59596 10016
rect 59636 9976 60268 10016
rect 60308 9976 62860 10016
rect 62900 9976 64204 10016
rect 64244 9976 64253 10016
rect 64387 9976 64396 10016
rect 64436 9976 64445 10016
rect 68227 9976 68236 10016
rect 68276 9976 68524 10016
rect 68564 9976 68573 10016
rect 75331 9976 75340 10016
rect 75380 9976 76492 10016
rect 76532 9976 76541 10016
rect 77347 9976 77356 10016
rect 77396 9976 77548 10016
rect 77588 9976 77597 10016
rect 43363 9975 43421 9976
rect 56044 9932 56084 9976
rect 64396 9932 64436 9976
rect 44899 9892 44908 9932
rect 44948 9892 46636 9932
rect 46676 9892 48364 9932
rect 48404 9892 48413 9932
rect 56044 9892 59020 9932
rect 59060 9892 59069 9932
rect 64204 9892 64436 9932
rect 77059 9892 77068 9932
rect 77108 9892 77644 9932
rect 77684 9892 77693 9932
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 16343 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 16729 9848
rect 28343 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 28729 9848
rect 40343 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 40729 9848
rect 43180 9808 45772 9848
rect 45812 9808 46060 9848
rect 46100 9808 48460 9848
rect 48500 9808 48509 9848
rect 52343 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 52729 9848
rect 0 9788 80 9808
rect 48259 9724 48268 9764
rect 48308 9724 49420 9764
rect 49460 9724 49469 9764
rect 64204 9680 64244 9892
rect 64343 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 64729 9848
rect 76343 9808 76352 9848
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76720 9808 76729 9848
rect 50380 9640 52108 9680
rect 52148 9640 53836 9680
rect 53876 9640 53885 9680
rect 63523 9640 63532 9680
rect 63572 9640 64012 9680
rect 64052 9640 64061 9680
rect 64204 9640 64396 9680
rect 64436 9640 65068 9680
rect 65108 9640 65117 9680
rect 72931 9640 72940 9680
rect 72980 9640 73420 9680
rect 73460 9640 73469 9680
rect 50380 9596 50420 9640
rect 46243 9556 46252 9596
rect 46292 9556 46828 9596
rect 46868 9556 47020 9596
rect 47060 9556 48748 9596
rect 48788 9556 48797 9596
rect 49699 9556 49708 9596
rect 49748 9556 50284 9596
rect 50324 9556 50420 9596
rect 68611 9556 68620 9596
rect 68660 9556 68812 9596
rect 68852 9556 70444 9596
rect 70484 9556 70493 9596
rect 72259 9556 72268 9596
rect 72308 9556 72652 9596
rect 72692 9556 72701 9596
rect 46147 9472 46156 9512
rect 46196 9472 46540 9512
rect 46580 9472 46589 9512
rect 46723 9472 46732 9512
rect 46772 9472 47212 9512
rect 47252 9472 47788 9512
rect 47828 9472 47837 9512
rect 49027 9472 49036 9512
rect 49076 9472 51148 9512
rect 51188 9472 52012 9512
rect 52052 9472 52061 9512
rect 57091 9472 57100 9512
rect 57140 9472 58732 9512
rect 58772 9472 58781 9512
rect 63715 9472 63724 9512
rect 63764 9472 64972 9512
rect 65012 9472 65021 9512
rect 65251 9472 65260 9512
rect 65300 9472 65932 9512
rect 65972 9472 67372 9512
rect 67412 9472 69484 9512
rect 69524 9472 70540 9512
rect 70580 9472 70589 9512
rect 71491 9472 71500 9512
rect 71540 9472 71980 9512
rect 72020 9472 72029 9512
rect 72835 9472 72844 9512
rect 72884 9472 73612 9512
rect 73652 9472 73661 9512
rect 835 9388 844 9428
rect 884 9388 29452 9428
rect 29492 9388 29501 9428
rect 31747 9388 31756 9428
rect 31796 9388 45484 9428
rect 45524 9388 45772 9428
rect 45812 9388 45821 9428
rect 49507 9388 49516 9428
rect 49556 9388 56140 9428
rect 56180 9388 56189 9428
rect 60163 9388 60172 9428
rect 60212 9388 61132 9428
rect 61172 9388 61420 9428
rect 61460 9388 61469 9428
rect 72355 9388 72364 9428
rect 72404 9388 73036 9428
rect 73076 9388 73085 9428
rect 68515 9344 68573 9345
rect 44611 9304 44620 9344
rect 44660 9304 45292 9344
rect 45332 9304 45341 9344
rect 53347 9304 53356 9344
rect 53396 9304 60844 9344
rect 60884 9304 60893 9344
rect 63331 9304 63340 9344
rect 63380 9304 63820 9344
rect 63860 9304 63869 9344
rect 67651 9304 67660 9344
rect 67700 9304 68524 9344
rect 68564 9304 68573 9344
rect 68515 9303 68573 9304
rect 56323 9220 56332 9260
rect 56372 9220 57484 9260
rect 57524 9220 57533 9260
rect 73411 9220 73420 9260
rect 73460 9220 73900 9260
rect 73940 9220 73949 9260
rect 77251 9220 77260 9260
rect 77300 9220 78412 9260
rect 78452 9220 78461 9260
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 15103 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 15489 9092
rect 27103 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 27489 9092
rect 39103 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 39489 9092
rect 50755 9052 50764 9092
rect 50804 9052 50813 9092
rect 51103 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 51489 9092
rect 57859 9052 57868 9092
rect 57908 9052 58540 9092
rect 58580 9052 58589 9092
rect 59107 9052 59116 9092
rect 59156 9052 59308 9092
rect 59348 9052 59357 9092
rect 63103 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 63489 9092
rect 64387 9052 64396 9092
rect 64436 9052 64780 9092
rect 64820 9052 64829 9092
rect 75103 9052 75112 9092
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75480 9052 75489 9092
rect 0 9008 80 9028
rect 50764 9008 50804 9052
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 48355 8968 48364 9008
rect 48404 8968 49172 9008
rect 50764 8968 55700 9008
rect 68803 8968 68812 9008
rect 68852 8968 69004 9008
rect 69044 8968 69053 9008
rect 73507 8968 73516 9008
rect 73556 8968 73996 9008
rect 74036 8968 74045 9008
rect 0 8948 80 8968
rect 49132 8924 49172 8968
rect 49123 8884 49132 8924
rect 49172 8884 49181 8924
rect 50755 8884 50764 8924
rect 50804 8884 51244 8924
rect 51284 8884 51628 8924
rect 51668 8884 51677 8924
rect 44419 8800 44428 8840
rect 44468 8800 44908 8840
rect 44948 8800 47596 8840
rect 47636 8800 47645 8840
rect 49891 8800 49900 8840
rect 49940 8800 50668 8840
rect 50708 8800 50717 8840
rect 52099 8800 52108 8840
rect 52148 8800 52300 8840
rect 52340 8800 52349 8840
rect 47779 8756 47837 8757
rect 45091 8716 45100 8756
rect 45140 8716 45964 8756
rect 46004 8716 47788 8756
rect 47828 8716 47837 8756
rect 48739 8716 48748 8756
rect 48788 8716 49324 8756
rect 49364 8716 49373 8756
rect 49699 8716 49708 8756
rect 49748 8716 50188 8756
rect 50228 8716 50237 8756
rect 51619 8716 51628 8756
rect 51668 8716 52876 8756
rect 52916 8716 52925 8756
rect 45292 8672 45332 8716
rect 47779 8715 47837 8716
rect 45283 8632 45292 8672
rect 45332 8632 45372 8672
rect 45580 8632 46060 8672
rect 46100 8632 46109 8672
rect 46435 8632 46444 8672
rect 46484 8632 48940 8672
rect 48980 8632 48989 8672
rect 50851 8632 50860 8672
rect 50900 8632 52588 8672
rect 52628 8632 52637 8672
rect 54499 8632 54508 8672
rect 54548 8632 54892 8672
rect 54932 8632 54941 8672
rect 45580 8504 45620 8632
rect 45667 8548 45676 8588
rect 45716 8548 46348 8588
rect 46388 8548 46397 8588
rect 48355 8548 48364 8588
rect 48404 8548 48844 8588
rect 48884 8548 49420 8588
rect 49460 8548 49469 8588
rect 45571 8464 45580 8504
rect 45620 8464 45629 8504
rect 48643 8464 48652 8504
rect 48692 8464 49036 8504
rect 49076 8464 49085 8504
rect 51724 8420 51764 8632
rect 55660 8420 55700 8968
rect 60739 8884 60748 8924
rect 60788 8884 62188 8924
rect 62228 8884 62237 8924
rect 63811 8884 63820 8924
rect 63860 8884 64300 8924
rect 64340 8884 64349 8924
rect 65923 8884 65932 8924
rect 65972 8884 67756 8924
rect 67796 8884 67805 8924
rect 70435 8884 70444 8924
rect 70484 8884 71692 8924
rect 71732 8884 71741 8924
rect 72547 8884 72556 8924
rect 72596 8884 74572 8924
rect 74612 8884 74621 8924
rect 58627 8800 58636 8840
rect 58676 8800 59116 8840
rect 59156 8800 59165 8840
rect 63619 8800 63628 8840
rect 63668 8800 66316 8840
rect 66356 8800 66365 8840
rect 69859 8800 69868 8840
rect 69908 8800 72652 8840
rect 72692 8800 73516 8840
rect 73556 8800 73565 8840
rect 76483 8800 76492 8840
rect 76532 8800 76876 8840
rect 76916 8800 76925 8840
rect 78124 8800 78316 8840
rect 78356 8800 78365 8840
rect 78124 8756 78164 8800
rect 62659 8716 62668 8756
rect 62708 8716 62956 8756
rect 62996 8716 63005 8756
rect 63139 8716 63148 8756
rect 63188 8716 63532 8756
rect 63572 8716 63581 8756
rect 64483 8716 64492 8756
rect 64532 8716 65260 8756
rect 65300 8716 66508 8756
rect 66548 8716 66557 8756
rect 69667 8716 69676 8756
rect 69716 8716 71788 8756
rect 71828 8716 72844 8756
rect 72884 8716 72893 8756
rect 73795 8716 73804 8756
rect 73844 8716 74476 8756
rect 74516 8716 75052 8756
rect 75092 8716 75532 8756
rect 75572 8716 75581 8756
rect 76387 8716 76396 8756
rect 76436 8716 78164 8756
rect 78211 8716 78220 8756
rect 78260 8716 79276 8756
rect 79316 8716 79325 8756
rect 68995 8672 69053 8673
rect 55747 8632 55756 8672
rect 55796 8632 56044 8672
rect 56084 8632 56332 8672
rect 56372 8632 56381 8672
rect 56899 8632 56908 8672
rect 56948 8632 58252 8672
rect 58292 8632 58301 8672
rect 59020 8632 62860 8672
rect 62900 8632 64972 8672
rect 65012 8632 67468 8672
rect 67508 8632 67517 8672
rect 68899 8632 68908 8672
rect 68948 8632 69004 8672
rect 69044 8632 69053 8672
rect 70819 8632 70828 8672
rect 70868 8632 74092 8672
rect 74132 8632 76780 8672
rect 76820 8632 78124 8672
rect 78164 8632 78173 8672
rect 59020 8588 59060 8632
rect 68995 8631 69053 8632
rect 59011 8548 59020 8588
rect 59060 8548 59069 8588
rect 63907 8548 63916 8588
rect 63956 8548 64492 8588
rect 64532 8548 64541 8588
rect 65059 8548 65068 8588
rect 65108 8548 67948 8588
rect 67988 8548 67997 8588
rect 73900 8504 73940 8632
rect 63235 8464 63244 8504
rect 63284 8464 64012 8504
rect 64052 8464 64061 8504
rect 64291 8464 64300 8504
rect 64340 8464 66028 8504
rect 66068 8464 66077 8504
rect 72355 8464 72364 8504
rect 72404 8464 72652 8504
rect 72692 8464 72701 8504
rect 73891 8464 73900 8504
rect 73940 8464 73949 8504
rect 76291 8464 76300 8504
rect 76340 8464 76349 8504
rect 76675 8464 76684 8504
rect 76724 8464 77452 8504
rect 77492 8464 78028 8504
rect 78068 8464 78077 8504
rect 66019 8420 66077 8421
rect 51715 8380 51724 8420
rect 51764 8380 51773 8420
rect 55651 8380 55660 8420
rect 55700 8380 55709 8420
rect 63139 8380 63148 8420
rect 63188 8380 66028 8420
rect 66068 8380 66077 8420
rect 76300 8420 76340 8464
rect 76300 8380 77836 8420
rect 77876 8380 77885 8420
rect 66019 8379 66077 8380
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 16343 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 16729 8336
rect 28343 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 28729 8336
rect 40343 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 40729 8336
rect 52343 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 52729 8336
rect 64343 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 64729 8336
rect 65347 8296 65356 8336
rect 65396 8296 66220 8336
rect 66260 8296 66269 8336
rect 68035 8296 68044 8336
rect 68084 8296 69004 8336
rect 69044 8296 69053 8336
rect 71683 8296 71692 8336
rect 71732 8296 72268 8336
rect 72308 8296 72317 8336
rect 76343 8296 76352 8336
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76720 8296 76729 8336
rect 62083 8212 62092 8252
rect 62132 8212 66412 8252
rect 66452 8212 66461 8252
rect 68899 8212 68908 8252
rect 68948 8212 73228 8252
rect 73268 8212 77356 8252
rect 77396 8212 77405 8252
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 49603 8128 49612 8168
rect 49652 8128 50092 8168
rect 50132 8128 50284 8168
rect 50324 8128 50333 8168
rect 52579 8128 52588 8168
rect 52628 8128 53836 8168
rect 53876 8128 53885 8168
rect 54115 8128 54124 8168
rect 54164 8128 54700 8168
rect 54740 8128 54749 8168
rect 58339 8128 58348 8168
rect 58388 8128 59404 8168
rect 59444 8128 59692 8168
rect 59732 8128 59741 8168
rect 65923 8128 65932 8168
rect 65972 8128 66700 8168
rect 66740 8128 70156 8168
rect 70196 8128 70205 8168
rect 73699 8128 73708 8168
rect 73748 8128 74380 8168
rect 74420 8128 74429 8168
rect 0 8108 80 8128
rect 54787 8044 54796 8084
rect 54836 8044 56140 8084
rect 56180 8044 56189 8084
rect 59491 8044 59500 8084
rect 59540 8044 60844 8084
rect 60884 8044 61804 8084
rect 61844 8044 61853 8084
rect 62179 8044 62188 8084
rect 62228 8044 63052 8084
rect 63092 8044 63101 8084
rect 48259 7960 48268 8000
rect 48308 7960 48460 8000
rect 48500 7960 48509 8000
rect 50659 7960 50668 8000
rect 50708 7960 54316 8000
rect 54356 7960 54365 8000
rect 54883 7960 54892 8000
rect 54932 7960 55852 8000
rect 55892 7960 55901 8000
rect 56035 7960 56044 8000
rect 56084 7960 57964 8000
rect 58004 7960 58013 8000
rect 58435 7960 58444 8000
rect 58484 7960 59308 8000
rect 59348 7960 59357 8000
rect 59587 7960 59596 8000
rect 59636 7960 60556 8000
rect 60596 7960 60605 8000
rect 61315 7960 61324 8000
rect 61364 7960 62572 8000
rect 62612 7960 62621 8000
rect 66019 7960 66028 8000
rect 66068 7960 66356 8000
rect 66403 7960 66412 8000
rect 66452 7960 66796 8000
rect 66836 7960 68428 8000
rect 68468 7960 68477 8000
rect 72163 7960 72172 8000
rect 72212 7960 73708 8000
rect 73748 7960 73757 8000
rect 76675 7960 76684 8000
rect 76724 7960 78988 8000
rect 79028 7960 79037 8000
rect 66316 7916 66356 7960
rect 53059 7876 53068 7916
rect 53108 7876 53548 7916
rect 53588 7876 53597 7916
rect 54403 7876 54412 7916
rect 54452 7876 54988 7916
rect 55028 7876 55037 7916
rect 66307 7876 66316 7916
rect 66356 7876 66365 7916
rect 68035 7876 68044 7916
rect 68084 7876 68524 7916
rect 68564 7876 68573 7916
rect 56323 7832 56381 7833
rect 55555 7792 55564 7832
rect 55604 7792 56332 7832
rect 56372 7792 56381 7832
rect 69091 7792 69100 7832
rect 69140 7792 77644 7832
rect 77684 7792 77932 7832
rect 77972 7792 77981 7832
rect 56323 7791 56381 7792
rect 451 7708 460 7748
rect 500 7708 940 7748
rect 980 7708 989 7748
rect 46915 7708 46924 7748
rect 46964 7708 47596 7748
rect 47636 7708 47645 7748
rect 54211 7708 54220 7748
rect 54260 7708 55180 7748
rect 55220 7708 55468 7748
rect 55508 7708 55517 7748
rect 62275 7708 62284 7748
rect 62324 7708 63148 7748
rect 63188 7708 63197 7748
rect 68323 7708 68332 7748
rect 68372 7708 69292 7748
rect 69332 7708 71404 7748
rect 71444 7708 71453 7748
rect 71779 7708 71788 7748
rect 71828 7708 72460 7748
rect 72500 7708 72509 7748
rect 47875 7624 47884 7664
rect 47924 7624 47933 7664
rect 68131 7624 68140 7664
rect 68180 7624 68620 7664
rect 68660 7624 68669 7664
rect 47884 7580 47924 7624
rect 68995 7580 69053 7581
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 15103 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 15489 7580
rect 27103 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 27489 7580
rect 39103 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 39489 7580
rect 47884 7540 48076 7580
rect 48116 7540 48125 7580
rect 51103 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 51489 7580
rect 63103 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 63489 7580
rect 68707 7540 68716 7580
rect 68756 7540 69004 7580
rect 69044 7540 69053 7580
rect 75103 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 75489 7580
rect 68995 7539 69053 7540
rect 53443 7456 53452 7496
rect 53492 7456 53644 7496
rect 53684 7456 54604 7496
rect 54644 7456 56812 7496
rect 56852 7456 56861 7496
rect 45667 7372 45676 7412
rect 45716 7372 46828 7412
rect 46868 7372 46877 7412
rect 50371 7372 50380 7412
rect 50420 7372 50572 7412
rect 50612 7372 50621 7412
rect 52867 7372 52876 7412
rect 52916 7372 53740 7412
rect 53780 7372 54796 7412
rect 54836 7372 54845 7412
rect 65731 7372 65740 7412
rect 65780 7372 66124 7412
rect 66164 7372 66173 7412
rect 0 7328 80 7348
rect 64771 7328 64829 7329
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 53347 7288 53356 7328
rect 53396 7288 53405 7328
rect 64579 7288 64588 7328
rect 64628 7288 64780 7328
rect 64820 7288 64829 7328
rect 73027 7288 73036 7328
rect 73076 7288 73612 7328
rect 73652 7288 75764 7328
rect 0 7268 80 7288
rect 47779 7160 47837 7161
rect 53356 7160 53396 7288
rect 64771 7287 64829 7288
rect 75724 7244 75764 7288
rect 71395 7204 71404 7244
rect 71444 7204 72172 7244
rect 72212 7204 72221 7244
rect 73507 7204 73516 7244
rect 73556 7204 73996 7244
rect 74036 7204 74045 7244
rect 75715 7204 75724 7244
rect 75764 7204 76012 7244
rect 76052 7204 76061 7244
rect 47779 7120 47788 7160
rect 47828 7120 47884 7160
rect 47924 7120 47933 7160
rect 51811 7120 51820 7160
rect 51860 7120 53396 7160
rect 57091 7120 57100 7160
rect 57140 7120 59884 7160
rect 59924 7120 59933 7160
rect 61027 7120 61036 7160
rect 61076 7120 62380 7160
rect 62420 7120 63532 7160
rect 63572 7120 64780 7160
rect 64820 7120 64829 7160
rect 71875 7120 71884 7160
rect 71924 7120 72268 7160
rect 72308 7120 72748 7160
rect 72788 7120 72797 7160
rect 75619 7120 75628 7160
rect 75668 7120 76492 7160
rect 76532 7120 76541 7160
rect 76771 7120 76780 7160
rect 76820 7120 76829 7160
rect 76963 7120 76972 7160
rect 77012 7120 77356 7160
rect 77396 7120 77836 7160
rect 77876 7120 78220 7160
rect 78260 7120 78269 7160
rect 47779 7119 47837 7120
rect 76780 7076 76820 7120
rect 55267 7036 55276 7076
rect 55316 7036 56716 7076
rect 56756 7036 57868 7076
rect 57908 7036 57917 7076
rect 60643 7036 60652 7076
rect 60692 7036 61612 7076
rect 61652 7036 61661 7076
rect 62755 7036 62764 7076
rect 62804 7036 64012 7076
rect 64052 7036 64396 7076
rect 64436 7036 64445 7076
rect 65059 7036 65068 7076
rect 65108 7036 65740 7076
rect 65780 7036 65789 7076
rect 75043 7036 75052 7076
rect 75092 7036 75820 7076
rect 75860 7036 75869 7076
rect 76780 7036 77068 7076
rect 77108 7036 78124 7076
rect 78164 7036 78173 7076
rect 50947 6952 50956 6992
rect 50996 6952 52108 6992
rect 52148 6952 52588 6992
rect 52628 6952 52637 6992
rect 58819 6952 58828 6992
rect 58868 6952 60076 6992
rect 60116 6952 62668 6992
rect 62708 6952 62717 6992
rect 64195 6952 64204 6992
rect 64244 6952 64588 6992
rect 64628 6952 64637 6992
rect 76780 6908 76820 7036
rect 78019 6952 78028 6992
rect 78068 6952 78700 6992
rect 78740 6952 78749 6992
rect 56323 6868 56332 6908
rect 56372 6868 56620 6908
rect 56660 6868 57964 6908
rect 58004 6868 65260 6908
rect 65300 6868 65309 6908
rect 73795 6868 73804 6908
rect 73844 6868 74092 6908
rect 74132 6868 76820 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 16343 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 16729 6824
rect 28343 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 28729 6824
rect 40343 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 40729 6824
rect 52343 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 52729 6824
rect 64343 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 64729 6824
rect 76343 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 76729 6824
rect 50179 6700 50188 6740
rect 50228 6700 53204 6740
rect 61699 6700 61708 6740
rect 61748 6700 62092 6740
rect 62132 6700 63532 6740
rect 63572 6700 66892 6740
rect 66932 6700 66941 6740
rect 53164 6656 53204 6700
rect 52675 6616 52684 6656
rect 52724 6616 52876 6656
rect 52916 6616 52925 6656
rect 53155 6616 53164 6656
rect 53204 6616 54220 6656
rect 54260 6616 54988 6656
rect 55028 6616 55037 6656
rect 63715 6616 63724 6656
rect 63764 6616 64108 6656
rect 64148 6616 64876 6656
rect 64916 6616 64925 6656
rect 69571 6616 69580 6656
rect 69620 6616 70828 6656
rect 70868 6616 71020 6656
rect 71060 6616 71069 6656
rect 74947 6616 74956 6656
rect 74996 6616 75628 6656
rect 75668 6616 75677 6656
rect 78499 6616 78508 6656
rect 78548 6616 79468 6656
rect 79508 6616 79517 6656
rect 51715 6532 51724 6572
rect 51764 6532 53548 6572
rect 53588 6532 53597 6572
rect 55075 6532 55084 6572
rect 55124 6532 55564 6572
rect 55604 6532 55613 6572
rect 55747 6532 55756 6572
rect 55796 6532 55948 6572
rect 55988 6532 57580 6572
rect 57620 6532 57629 6572
rect 60739 6532 60748 6572
rect 60788 6532 62188 6572
rect 62228 6532 62237 6572
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 52579 6448 52588 6488
rect 52628 6448 53452 6488
rect 53492 6448 53501 6488
rect 55363 6448 55372 6488
rect 55412 6448 55660 6488
rect 55700 6448 55709 6488
rect 56803 6448 56812 6488
rect 56852 6448 58348 6488
rect 58388 6448 58397 6488
rect 60931 6448 60940 6488
rect 60980 6448 61132 6488
rect 61172 6448 61181 6488
rect 61891 6448 61900 6488
rect 61940 6448 62380 6488
rect 62420 6448 62429 6488
rect 64867 6448 64876 6488
rect 64916 6448 66604 6488
rect 66644 6448 66653 6488
rect 67939 6448 67948 6488
rect 67988 6448 68428 6488
rect 68468 6448 68477 6488
rect 69667 6448 69676 6488
rect 69716 6448 70540 6488
rect 70580 6448 70732 6488
rect 70772 6448 71308 6488
rect 71348 6448 71357 6488
rect 72931 6448 72940 6488
rect 72980 6448 75052 6488
rect 75092 6448 75101 6488
rect 0 6428 80 6448
rect 55660 6404 55700 6448
rect 50371 6364 50380 6404
rect 50420 6364 52972 6404
rect 53012 6364 53021 6404
rect 55660 6364 56908 6404
rect 56948 6364 56957 6404
rect 68803 6364 68812 6404
rect 68852 6364 70156 6404
rect 70196 6364 70444 6404
rect 70484 6364 70493 6404
rect 76771 6364 76780 6404
rect 76820 6364 77740 6404
rect 77780 6364 77789 6404
rect 52972 6320 53012 6364
rect 51907 6280 51916 6320
rect 51956 6280 52300 6320
rect 52340 6280 52349 6320
rect 52972 6280 53164 6320
rect 53204 6280 53213 6320
rect 53539 6280 53548 6320
rect 53588 6280 56044 6320
rect 56084 6280 56093 6320
rect 68131 6280 68140 6320
rect 68180 6280 69100 6320
rect 69140 6280 69149 6320
rect 70051 6280 70060 6320
rect 70100 6280 71692 6320
rect 71732 6280 71741 6320
rect 73027 6280 73036 6320
rect 73076 6280 73804 6320
rect 73844 6280 73853 6320
rect 65731 6152 65789 6153
rect 65646 6112 65740 6152
rect 65780 6112 65789 6152
rect 65731 6111 65789 6112
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 15103 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 15489 6068
rect 27103 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 27489 6068
rect 39103 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 39489 6068
rect 51103 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 51489 6068
rect 63103 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 63489 6068
rect 75103 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 75489 6068
rect 64963 5984 65021 5985
rect 59875 5944 59884 5984
rect 59924 5944 61652 5984
rect 61612 5900 61652 5944
rect 64963 5944 64972 5984
rect 65012 5944 65740 5984
rect 65780 5944 65789 5984
rect 72067 5944 72076 5984
rect 72116 5944 72460 5984
rect 72500 5944 72509 5984
rect 64963 5943 65021 5944
rect 64771 5900 64829 5901
rect 77635 5900 77693 5901
rect 60067 5860 60076 5900
rect 60116 5860 61132 5900
rect 61172 5860 61181 5900
rect 61603 5860 61612 5900
rect 61652 5860 62764 5900
rect 62804 5860 62813 5900
rect 64579 5860 64588 5900
rect 64628 5860 64780 5900
rect 64820 5860 64829 5900
rect 65347 5860 65356 5900
rect 65396 5860 65644 5900
rect 65684 5860 65693 5900
rect 77539 5860 77548 5900
rect 77588 5860 77644 5900
rect 77684 5860 77693 5900
rect 64771 5859 64829 5860
rect 77635 5859 77693 5860
rect 54211 5776 54220 5816
rect 54260 5776 56524 5816
rect 56564 5776 56573 5816
rect 58339 5776 58348 5816
rect 58388 5776 61900 5816
rect 61940 5776 61949 5816
rect 64675 5776 64684 5816
rect 64724 5776 66124 5816
rect 66164 5776 66173 5816
rect 68899 5776 68908 5816
rect 68948 5776 69388 5816
rect 69428 5776 69437 5816
rect 73219 5776 73228 5816
rect 73268 5776 74284 5816
rect 74324 5776 74333 5816
rect 74467 5776 74476 5816
rect 74516 5776 74956 5816
rect 74996 5776 75005 5816
rect 59404 5732 59444 5776
rect 76867 5732 76925 5733
rect 835 5692 844 5732
rect 884 5692 1612 5732
rect 1652 5692 1661 5732
rect 52675 5692 52684 5732
rect 52724 5692 52876 5732
rect 52916 5692 52925 5732
rect 59395 5692 59404 5732
rect 59444 5692 59453 5732
rect 64771 5692 64780 5732
rect 64820 5692 65548 5732
rect 65588 5692 65597 5732
rect 68131 5692 68140 5732
rect 68180 5692 68716 5732
rect 68756 5692 68765 5732
rect 69763 5692 69772 5732
rect 69812 5692 72172 5732
rect 72212 5692 72221 5732
rect 76003 5692 76012 5732
rect 76052 5692 76876 5732
rect 76916 5692 76925 5732
rect 77539 5692 77548 5732
rect 77588 5692 77836 5732
rect 77876 5692 77885 5732
rect 76867 5691 76925 5692
rect 0 5648 80 5668
rect 65347 5648 65405 5649
rect 77155 5648 77213 5649
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 55555 5608 55564 5648
rect 55604 5608 56236 5648
rect 56276 5608 57484 5648
rect 57524 5608 57533 5648
rect 65251 5608 65260 5648
rect 65300 5608 65356 5648
rect 65396 5608 65405 5648
rect 65635 5608 65644 5648
rect 65684 5608 66316 5648
rect 66356 5608 66365 5648
rect 68419 5608 68428 5648
rect 68468 5608 69292 5648
rect 69332 5608 70348 5648
rect 70388 5608 70397 5648
rect 71491 5608 71500 5648
rect 71540 5608 72268 5648
rect 72308 5608 72317 5648
rect 72643 5608 72652 5648
rect 72692 5608 73420 5648
rect 73460 5608 73469 5648
rect 74083 5608 74092 5648
rect 74132 5608 74380 5648
rect 74420 5608 74429 5648
rect 76963 5608 76972 5648
rect 77012 5608 77164 5648
rect 77204 5608 77213 5648
rect 77443 5608 77452 5648
rect 77492 5608 78124 5648
rect 78164 5608 78173 5648
rect 0 5588 80 5608
rect 65347 5607 65405 5608
rect 77155 5607 77213 5608
rect 68995 5564 69053 5565
rect 57955 5524 57964 5564
rect 58004 5524 59884 5564
rect 59924 5524 65452 5564
rect 65492 5524 65501 5564
rect 68323 5524 68332 5564
rect 68372 5524 68812 5564
rect 68852 5524 68861 5564
rect 68995 5524 69004 5564
rect 69044 5524 69676 5564
rect 69716 5524 69725 5564
rect 68995 5523 69053 5524
rect 58243 5440 58252 5480
rect 58292 5440 59788 5480
rect 59828 5440 59837 5480
rect 61027 5440 61036 5480
rect 61076 5440 61324 5480
rect 61364 5440 61373 5480
rect 73315 5440 73324 5480
rect 73364 5440 74572 5480
rect 74612 5440 74621 5480
rect 76483 5440 76492 5480
rect 76532 5440 77644 5480
rect 77684 5440 78316 5480
rect 78356 5440 78365 5480
rect 73987 5356 73996 5396
rect 74036 5356 76780 5396
rect 76820 5356 77548 5396
rect 77588 5356 77597 5396
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 16343 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 16729 5312
rect 28343 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 28729 5312
rect 40343 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 40729 5312
rect 52343 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 52729 5312
rect 64343 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 64729 5312
rect 76343 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 76729 5312
rect 64771 5144 64829 5145
rect 54787 5104 54796 5144
rect 54836 5104 55756 5144
rect 55796 5104 55805 5144
rect 64579 5104 64588 5144
rect 64628 5104 64780 5144
rect 64820 5104 64972 5144
rect 65012 5104 65021 5144
rect 65731 5104 65740 5144
rect 65780 5104 67756 5144
rect 67796 5104 67805 5144
rect 70147 5104 70156 5144
rect 70196 5104 70924 5144
rect 70964 5104 70973 5144
rect 64771 5103 64829 5104
rect 60547 5020 60556 5060
rect 60596 5020 60748 5060
rect 60788 5020 61420 5060
rect 61460 5020 61469 5060
rect 70531 5020 70540 5060
rect 70580 5020 72460 5060
rect 72500 5020 72509 5060
rect 77827 5020 77836 5060
rect 77876 5020 78604 5060
rect 78644 5020 78653 5060
rect 65731 4976 65789 4977
rect 45763 4936 45772 4976
rect 45812 4936 55796 4976
rect 55843 4936 55852 4976
rect 55892 4936 56236 4976
rect 56276 4936 56285 4976
rect 56995 4936 57004 4976
rect 57044 4936 58060 4976
rect 58100 4936 58109 4976
rect 59779 4936 59788 4976
rect 59828 4936 60460 4976
rect 60500 4936 60509 4976
rect 64867 4936 64876 4976
rect 64916 4936 65548 4976
rect 65588 4936 65597 4976
rect 65731 4936 65740 4976
rect 65780 4936 66796 4976
rect 66836 4936 68332 4976
rect 68372 4936 68381 4976
rect 69187 4936 69196 4976
rect 69236 4936 71020 4976
rect 71060 4936 71788 4976
rect 71828 4936 73996 4976
rect 74036 4936 74668 4976
rect 74708 4936 75820 4976
rect 75860 4936 78220 4976
rect 78260 4936 78269 4976
rect 55756 4892 55796 4936
rect 65731 4935 65789 4936
rect 52195 4852 52204 4892
rect 52244 4852 52876 4892
rect 52916 4852 53356 4892
rect 53396 4852 53405 4892
rect 54691 4852 54700 4892
rect 54740 4852 55180 4892
rect 55220 4852 55229 4892
rect 55756 4852 61804 4892
rect 61844 4852 61853 4892
rect 64963 4852 64972 4892
rect 65012 4852 65452 4892
rect 65492 4852 65836 4892
rect 65876 4852 65885 4892
rect 76963 4852 76972 4892
rect 77012 4852 77260 4892
rect 77300 4852 77309 4892
rect 0 4808 80 4828
rect 77635 4808 77693 4809
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 51715 4768 51724 4808
rect 51764 4768 52396 4808
rect 52436 4768 52445 4808
rect 52579 4768 52588 4808
rect 52628 4768 53164 4808
rect 53204 4768 54124 4808
rect 54164 4768 54173 4808
rect 56035 4768 56044 4808
rect 56084 4768 57772 4808
rect 57812 4768 57821 4808
rect 77550 4768 77644 4808
rect 77684 4768 77693 4808
rect 0 4748 80 4768
rect 77635 4767 77693 4768
rect 54211 4684 54220 4724
rect 54260 4684 54508 4724
rect 54548 4684 54557 4724
rect 71299 4684 71308 4724
rect 71348 4684 72940 4724
rect 72980 4684 73132 4724
rect 73172 4684 73181 4724
rect 61411 4600 61420 4640
rect 61460 4600 61804 4640
rect 61844 4600 61853 4640
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 15103 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 15489 4556
rect 27103 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 27489 4556
rect 39103 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 39489 4556
rect 51103 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 51489 4556
rect 63103 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 63489 4556
rect 75103 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 75489 4556
rect 68419 4432 68428 4472
rect 68468 4432 68620 4472
rect 68660 4432 68669 4472
rect 74563 4432 74572 4472
rect 74612 4432 75820 4472
rect 75860 4432 75869 4472
rect 61027 4348 61036 4388
rect 61076 4348 61420 4388
rect 61460 4348 61469 4388
rect 76867 4348 76876 4388
rect 76916 4348 77164 4388
rect 77204 4348 77213 4388
rect 53059 4264 53068 4304
rect 53108 4264 55084 4304
rect 55124 4264 55133 4304
rect 60739 4264 60748 4304
rect 60788 4264 62476 4304
rect 62516 4264 63052 4304
rect 63092 4264 63101 4304
rect 64483 4264 64492 4304
rect 64532 4264 66604 4304
rect 66644 4264 66653 4304
rect 68899 4264 68908 4304
rect 68948 4264 68957 4304
rect 69667 4264 69676 4304
rect 69716 4264 71692 4304
rect 71732 4264 71741 4304
rect 74275 4264 74284 4304
rect 74324 4264 75148 4304
rect 75188 4264 75532 4304
rect 75572 4264 75581 4304
rect 76099 4264 76108 4304
rect 76148 4264 77356 4304
rect 77396 4264 77405 4304
rect 66595 4220 66653 4221
rect 835 4180 844 4220
rect 884 4180 1420 4220
rect 1460 4180 1469 4220
rect 53827 4180 53836 4220
rect 53876 4180 54604 4220
rect 54644 4180 54653 4220
rect 56515 4180 56524 4220
rect 56564 4180 57140 4220
rect 57379 4180 57388 4220
rect 57428 4180 57964 4220
rect 58004 4180 58013 4220
rect 66115 4180 66124 4220
rect 66164 4180 66604 4220
rect 66644 4180 66653 4220
rect 68908 4220 68948 4264
rect 68908 4180 71212 4220
rect 71252 4180 71404 4220
rect 71444 4180 72076 4220
rect 72116 4180 72125 4220
rect 74947 4180 74956 4220
rect 74996 4180 75724 4220
rect 75764 4180 77068 4220
rect 77108 4180 77117 4220
rect 78115 4180 78124 4220
rect 78164 4180 79372 4220
rect 79412 4180 79421 4220
rect 57100 4136 57140 4180
rect 66595 4179 66653 4180
rect 74956 4136 74996 4180
rect 54403 4096 54412 4136
rect 54452 4096 56332 4136
rect 56372 4096 56716 4136
rect 56756 4096 56765 4136
rect 57091 4096 57100 4136
rect 57140 4096 57149 4136
rect 57283 4096 57292 4136
rect 57332 4096 57676 4136
rect 57716 4096 57725 4136
rect 60355 4096 60364 4136
rect 60404 4096 62284 4136
rect 62324 4096 62333 4136
rect 68323 4096 68332 4136
rect 68372 4096 69196 4136
rect 69236 4096 69245 4136
rect 71011 4096 71020 4136
rect 71060 4096 71500 4136
rect 71540 4096 71549 4136
rect 73123 4096 73132 4136
rect 73172 4096 74996 4136
rect 76579 4096 76588 4136
rect 76628 4096 77452 4136
rect 77492 4096 77501 4136
rect 71020 4052 71060 4096
rect 60163 4012 60172 4052
rect 60212 4012 60652 4052
rect 60692 4012 60701 4052
rect 68707 4012 68716 4052
rect 68756 4012 71060 4052
rect 72547 4012 72556 4052
rect 72596 4012 74380 4052
rect 74420 4012 74429 4052
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 52099 3928 52108 3968
rect 52148 3928 54220 3968
rect 54260 3928 56428 3968
rect 56468 3928 56477 3968
rect 60067 3928 60076 3968
rect 60116 3928 61036 3968
rect 61076 3928 62572 3968
rect 62612 3928 63628 3968
rect 63668 3928 63677 3968
rect 65155 3928 65164 3968
rect 65204 3928 65644 3968
rect 65684 3928 65693 3968
rect 71107 3928 71116 3968
rect 71156 3928 71596 3968
rect 71636 3928 71645 3968
rect 71875 3928 71884 3968
rect 71924 3928 72076 3968
rect 72116 3928 72125 3968
rect 75907 3928 75916 3968
rect 75956 3928 76300 3968
rect 76340 3928 76349 3968
rect 0 3908 80 3928
rect 76300 3884 76340 3928
rect 71779 3844 71788 3884
rect 71828 3844 72652 3884
rect 72692 3844 72701 3884
rect 76300 3844 77068 3884
rect 77108 3844 77117 3884
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 16343 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 16729 3800
rect 28343 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 28729 3800
rect 40343 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 40729 3800
rect 52343 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 52729 3800
rect 64343 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 64729 3800
rect 72259 3760 72268 3800
rect 72308 3760 73996 3800
rect 74036 3760 74045 3800
rect 76343 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 76729 3800
rect 60835 3676 60844 3716
rect 60884 3676 61516 3716
rect 61556 3676 62092 3716
rect 62132 3676 62141 3716
rect 68995 3676 69004 3716
rect 69044 3676 77644 3716
rect 77684 3676 77693 3716
rect 5155 3592 5164 3632
rect 5204 3592 7372 3632
rect 7412 3592 7421 3632
rect 65539 3592 65548 3632
rect 65588 3592 67660 3632
rect 67700 3592 68812 3632
rect 68852 3592 68861 3632
rect 71875 3592 71884 3632
rect 71924 3592 73036 3632
rect 73076 3592 73085 3632
rect 77059 3548 77117 3549
rect 60163 3508 60172 3548
rect 60212 3508 60844 3548
rect 60884 3508 60893 3548
rect 65635 3508 65644 3548
rect 65684 3508 66220 3548
rect 66260 3508 66269 3548
rect 76675 3508 76684 3548
rect 76724 3508 77068 3548
rect 77108 3508 77117 3548
rect 77059 3507 77117 3508
rect 64771 3464 64829 3465
rect 55075 3424 55084 3464
rect 55124 3424 57292 3464
rect 57332 3424 58636 3464
rect 58676 3424 58685 3464
rect 60067 3424 60076 3464
rect 60116 3424 60556 3464
rect 60596 3424 60605 3464
rect 64579 3424 64588 3464
rect 64628 3424 64780 3464
rect 64820 3424 64829 3464
rect 65923 3424 65932 3464
rect 65972 3424 66412 3464
rect 66452 3424 66461 3464
rect 76771 3424 76780 3464
rect 76820 3424 76972 3464
rect 77012 3424 78028 3464
rect 78068 3424 78077 3464
rect 64771 3423 64829 3424
rect 50179 3380 50237 3381
rect 835 3340 844 3380
rect 884 3340 2476 3380
rect 2516 3340 2525 3380
rect 50179 3340 50188 3380
rect 50228 3340 61996 3380
rect 62036 3340 69196 3380
rect 69236 3340 69245 3380
rect 50179 3339 50237 3340
rect 76771 3296 76829 3297
rect 63235 3256 63244 3296
rect 63284 3256 64492 3296
rect 64532 3256 64541 3296
rect 73123 3256 73132 3296
rect 73172 3256 73612 3296
rect 73652 3256 73661 3296
rect 76291 3256 76300 3296
rect 76340 3256 76780 3296
rect 76820 3256 76829 3296
rect 76771 3255 76829 3256
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 71587 3172 71596 3212
rect 71636 3172 72076 3212
rect 72116 3172 72940 3212
rect 72980 3172 72989 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 15103 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 15489 3044
rect 27103 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 27489 3044
rect 39103 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 39489 3044
rect 51103 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 51489 3044
rect 63103 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 63489 3044
rect 71395 3004 71404 3044
rect 71444 3004 74572 3044
rect 74612 3004 74621 3044
rect 75103 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 75489 3044
rect 61027 2960 61085 2961
rect 60942 2920 61036 2960
rect 61076 2920 61085 2960
rect 62083 2920 62092 2960
rect 62132 2920 62764 2960
rect 62804 2920 62813 2960
rect 61027 2919 61085 2920
rect 75523 2876 75581 2877
rect 56716 2836 57484 2876
rect 57524 2836 57868 2876
rect 57908 2836 57917 2876
rect 60643 2836 60652 2876
rect 60692 2836 62668 2876
rect 62708 2836 62717 2876
rect 70051 2836 70060 2876
rect 70100 2836 70924 2876
rect 70964 2836 70973 2876
rect 75043 2836 75052 2876
rect 75092 2836 75532 2876
rect 75572 2836 75581 2876
rect 56035 2752 56044 2792
rect 56084 2752 56524 2792
rect 56564 2752 56573 2792
rect 56716 2624 56756 2836
rect 75523 2835 75581 2836
rect 57091 2752 57100 2792
rect 57140 2752 58540 2792
rect 58580 2752 58589 2792
rect 61219 2752 61228 2792
rect 61268 2752 61708 2792
rect 61748 2752 62476 2792
rect 62516 2752 62525 2792
rect 72067 2752 72076 2792
rect 72116 2752 72364 2792
rect 72404 2752 72413 2792
rect 74947 2752 74956 2792
rect 74996 2752 75628 2792
rect 75668 2752 75677 2792
rect 60547 2668 60556 2708
rect 60596 2668 61516 2708
rect 61556 2668 61565 2708
rect 62563 2668 62572 2708
rect 62612 2668 63340 2708
rect 63380 2668 63389 2708
rect 64483 2668 64492 2708
rect 64532 2668 64972 2708
rect 65012 2668 65021 2708
rect 65155 2668 65164 2708
rect 65204 2668 66028 2708
rect 66068 2668 66077 2708
rect 66211 2668 66220 2708
rect 66260 2668 66796 2708
rect 66836 2668 66845 2708
rect 72739 2668 72748 2708
rect 72788 2668 74284 2708
rect 74324 2668 76972 2708
rect 77012 2668 77164 2708
rect 77204 2668 77213 2708
rect 56707 2584 56716 2624
rect 56756 2584 56765 2624
rect 57580 2584 58732 2624
rect 58772 2584 58781 2624
rect 58915 2584 58924 2624
rect 58964 2584 60748 2624
rect 60788 2584 60940 2624
rect 60980 2584 61420 2624
rect 61460 2584 61469 2624
rect 61603 2584 61612 2624
rect 61652 2584 62284 2624
rect 62324 2584 62860 2624
rect 62900 2584 62909 2624
rect 64387 2584 64396 2624
rect 64436 2584 64876 2624
rect 64916 2584 66892 2624
rect 66932 2584 67564 2624
rect 67604 2584 67613 2624
rect 68419 2584 68428 2624
rect 68468 2584 69484 2624
rect 69524 2584 69533 2624
rect 71299 2584 71308 2624
rect 71348 2584 71788 2624
rect 71828 2584 71837 2624
rect 72163 2584 72172 2624
rect 72212 2584 72844 2624
rect 72884 2584 72893 2624
rect 74083 2584 74092 2624
rect 74132 2584 74380 2624
rect 74420 2584 74429 2624
rect 75715 2584 75724 2624
rect 75764 2584 76300 2624
rect 76340 2584 76588 2624
rect 76628 2584 76637 2624
rect 77635 2584 77644 2624
rect 77684 2584 77932 2624
rect 77972 2584 78412 2624
rect 78452 2584 78461 2624
rect 57580 2540 57620 2584
rect 56323 2500 56332 2540
rect 56372 2500 57620 2540
rect 77059 2500 77068 2540
rect 77108 2500 77836 2540
rect 77876 2500 77885 2540
rect 61315 2416 61324 2456
rect 61364 2416 62188 2456
rect 62228 2416 62956 2456
rect 62996 2416 63005 2456
rect 64003 2416 64012 2456
rect 64052 2416 64588 2456
rect 64628 2416 66700 2456
rect 66740 2416 66749 2456
rect 68131 2416 68140 2456
rect 68180 2416 68812 2456
rect 68852 2416 68861 2456
rect 74083 2416 74092 2456
rect 74132 2416 76108 2456
rect 76148 2416 76157 2456
rect 76387 2416 76396 2456
rect 76436 2416 76972 2456
rect 77012 2416 77021 2456
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 16343 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 16729 2288
rect 28343 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 28729 2288
rect 40343 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 40729 2288
rect 52343 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 52729 2288
rect 64343 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 64729 2288
rect 76343 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 76729 2288
rect 0 2228 80 2248
rect 68611 2164 68620 2204
rect 68660 2164 69100 2204
rect 69140 2164 69149 2204
rect 63235 2080 63244 2120
rect 63284 2080 64780 2120
rect 64820 2080 66220 2120
rect 66260 2080 66269 2120
rect 72643 2080 72652 2120
rect 72692 2080 73996 2120
rect 74036 2080 74045 2120
rect 75811 2080 75820 2120
rect 75860 2080 76396 2120
rect 76436 2080 77452 2120
rect 77492 2080 77501 2120
rect 61027 2036 61085 2037
rect 58339 1996 58348 2036
rect 58388 1996 59116 2036
rect 59156 1996 59165 2036
rect 60259 1996 60268 2036
rect 60308 1996 61036 2036
rect 61076 1996 62764 2036
rect 62804 1996 62813 2036
rect 66787 1996 66796 2036
rect 66836 1996 67660 2036
rect 67700 1996 67709 2036
rect 69187 1996 69196 2036
rect 69236 1996 70156 2036
rect 70196 1996 71828 2036
rect 73795 1996 73804 2036
rect 73844 1996 74476 2036
rect 74516 1996 74525 2036
rect 75436 1996 77356 2036
rect 77396 1996 77405 2036
rect 61027 1995 61085 1996
rect 65731 1952 65789 1953
rect 71788 1952 71828 1996
rect 75436 1952 75476 1996
rect 59587 1912 59596 1952
rect 59636 1912 61132 1952
rect 61172 1912 61900 1952
rect 61940 1912 63628 1952
rect 63668 1912 63677 1952
rect 65347 1912 65356 1952
rect 65396 1912 65740 1952
rect 65780 1912 65789 1952
rect 66211 1912 66220 1952
rect 66260 1912 67756 1952
rect 67796 1912 68044 1952
rect 68084 1912 70060 1952
rect 70100 1912 70109 1952
rect 71779 1912 71788 1952
rect 71828 1912 71837 1952
rect 72643 1912 72652 1952
rect 72692 1912 74380 1952
rect 74420 1912 74429 1952
rect 74755 1912 74764 1952
rect 74804 1912 75436 1952
rect 75476 1912 75485 1952
rect 75619 1912 75628 1952
rect 75668 1912 75677 1952
rect 75811 1912 75820 1952
rect 75860 1912 77068 1952
rect 77108 1912 77117 1952
rect 77251 1912 77260 1952
rect 77300 1912 78220 1952
rect 78260 1912 78269 1952
rect 65731 1911 65789 1912
rect 61219 1868 61277 1869
rect 75628 1868 75668 1912
rect 61200 1828 61228 1868
rect 61268 1828 61324 1868
rect 61364 1828 71116 1868
rect 71156 1828 71165 1868
rect 74179 1828 74188 1868
rect 74228 1828 75668 1868
rect 61219 1827 61277 1828
rect 67939 1744 67948 1784
rect 67988 1744 68620 1784
rect 68660 1744 68669 1784
rect 74755 1744 74764 1784
rect 74804 1744 75532 1784
rect 75572 1744 75581 1784
rect 62755 1660 62764 1700
rect 62804 1660 63244 1700
rect 63284 1660 63293 1700
rect 66211 1660 66220 1700
rect 66260 1660 66604 1700
rect 66644 1660 67372 1700
rect 67412 1660 67421 1700
rect 68515 1660 68524 1700
rect 68564 1660 69772 1700
rect 69812 1660 69821 1700
rect 75628 1532 75668 1828
rect 76483 1576 76492 1616
rect 76532 1576 77164 1616
rect 77204 1576 77213 1616
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 15103 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 15489 1532
rect 27103 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 27489 1532
rect 39103 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 39489 1532
rect 51103 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 51489 1532
rect 58723 1492 58732 1532
rect 58772 1492 60268 1532
rect 60308 1492 60317 1532
rect 63103 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 63489 1532
rect 69571 1492 69580 1532
rect 69620 1492 71500 1532
rect 71540 1492 72460 1532
rect 72500 1492 72509 1532
rect 75103 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 75489 1532
rect 75619 1492 75628 1532
rect 75668 1492 75677 1532
rect 76099 1492 76108 1532
rect 76148 1492 76684 1532
rect 76724 1492 76733 1532
rect 71683 1408 71692 1448
rect 71732 1408 72076 1448
rect 72116 1408 72125 1448
rect 71587 1324 71596 1364
rect 71636 1324 74956 1364
rect 74996 1324 75005 1364
rect 65731 1196 65789 1197
rect 65731 1156 65740 1196
rect 65780 1156 67180 1196
rect 67220 1156 67229 1196
rect 69667 1156 69676 1196
rect 69716 1156 71212 1196
rect 71252 1156 71261 1196
rect 76579 1156 76588 1196
rect 76628 1156 79372 1196
rect 79412 1156 79421 1196
rect 65731 1155 65789 1156
rect 59875 1072 59884 1112
rect 59924 1072 61036 1112
rect 61076 1072 61085 1112
rect 66787 1072 66796 1112
rect 66836 1072 67756 1112
rect 67796 1072 67805 1112
rect 68419 1072 68428 1112
rect 68468 1072 69484 1112
rect 69524 1072 69533 1112
rect 71107 1072 71116 1112
rect 71156 1072 72844 1112
rect 72884 1072 73132 1112
rect 73172 1072 73181 1112
rect 71779 988 71788 1028
rect 71828 988 73228 1028
rect 73268 988 73277 1028
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 16343 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 16729 776
rect 28343 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 28729 776
rect 40343 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 40729 776
rect 52343 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 52729 776
rect 64343 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 64729 776
rect 76343 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 76729 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 50284 38200 50324 38240
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 66316 37108 66356 37148
rect 76204 37108 76244 37148
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 74188 36856 74228 36896
rect 74188 36520 74228 36560
rect 75628 36436 75668 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 56620 36268 56660 36308
rect 61708 36268 61748 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 61228 36016 61268 36056
rect 76684 35932 76724 35972
rect 73804 35848 73844 35888
rect 61708 35764 61748 35804
rect 61036 35680 61076 35720
rect 56620 35596 56660 35636
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 61228 35512 61268 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 61036 35260 61076 35300
rect 73804 35176 73844 35216
rect 76876 35176 76916 35216
rect 76780 35092 76820 35132
rect 61036 35008 61076 35048
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 76780 34924 76820 34964
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 77356 34252 77396 34292
rect 77932 34084 77972 34124
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 77164 33664 77204 33704
rect 77356 33412 77396 33452
rect 61228 33328 61268 33368
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55372 33244 55412 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 72844 32992 72884 33032
rect 72364 32740 72404 32780
rect 55372 32656 55412 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 73612 32488 73652 32528
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 63532 32152 63572 32192
rect 77932 32236 77972 32276
rect 72844 32068 72884 32108
rect 56428 31816 56468 31856
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 53068 31732 53108 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 72844 31648 72884 31688
rect 62668 31480 62708 31520
rect 73324 31480 73364 31520
rect 63532 31396 63572 31436
rect 61132 31312 61172 31352
rect 63916 31312 63956 31352
rect 73612 31312 73652 31352
rect 77260 31312 77300 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 61132 30556 61172 30596
rect 64012 30472 64052 30512
rect 62668 30388 62708 30428
rect 72364 30388 72404 30428
rect 51820 30304 51860 30344
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 61228 30220 61268 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 73804 30220 73844 30260
rect 74956 30220 74996 30260
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 77260 30220 77300 30260
rect 78028 30220 78068 30260
rect 53164 29884 53204 29924
rect 39916 29632 39956 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 64204 29296 64244 29336
rect 65836 29296 65876 29336
rect 39916 29044 39956 29084
rect 50380 29044 50420 29084
rect 77932 28876 77972 28916
rect 42892 28792 42932 28832
rect 71020 28792 71060 28832
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 66316 28624 66356 28664
rect 43276 28540 43316 28580
rect 65836 28540 65876 28580
rect 73324 28540 73364 28580
rect 52204 28456 52244 28496
rect 70924 28456 70964 28496
rect 50092 28204 50132 28244
rect 77260 28036 77300 28076
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 48364 27952 48404 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 53356 27952 53396 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 43372 27784 43412 27824
rect 42892 27616 42932 27656
rect 62860 27700 62900 27740
rect 73324 27532 73364 27572
rect 48364 27280 48404 27320
rect 68716 27280 68756 27320
rect 69100 27280 69140 27320
rect 69676 27280 69716 27320
rect 71308 27280 71348 27320
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 42892 27196 42932 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 52204 27196 52244 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 68812 27196 68852 27236
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 74860 27112 74900 27152
rect 40204 27028 40244 27068
rect 40108 26944 40148 26984
rect 52972 27028 53012 27068
rect 71692 26944 71732 26984
rect 58444 26860 58484 26900
rect 61612 26860 61652 26900
rect 64204 26860 64244 26900
rect 70924 26860 70964 26900
rect 40012 26692 40052 26732
rect 49132 26608 49172 26648
rect 71692 26608 71732 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 49900 26440 49940 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 52972 26440 53012 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 69772 26440 69812 26480
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 43276 26356 43316 26396
rect 69292 26272 69332 26312
rect 41068 26104 41108 26144
rect 77260 26104 77300 26144
rect 69868 25936 69908 25976
rect 43372 25852 43412 25892
rect 53356 25852 53396 25892
rect 40012 25768 40052 25808
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 42892 25600 42932 25640
rect 54508 25600 54548 25640
rect 51532 25516 51572 25556
rect 66604 25516 66644 25556
rect 51916 25432 51956 25472
rect 58732 25348 58772 25388
rect 69772 25348 69812 25388
rect 75052 25264 75092 25304
rect 40300 25180 40340 25220
rect 45580 25180 45620 25220
rect 50572 25180 50612 25220
rect 41068 25096 41108 25136
rect 50764 25096 50804 25136
rect 67564 25180 67604 25220
rect 76780 25096 76820 25136
rect 77260 25012 77300 25052
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 52780 24928 52820 24968
rect 56140 24928 56180 24968
rect 57580 24928 57620 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 51916 24508 51956 24548
rect 41356 24424 41396 24464
rect 58252 24424 58292 24464
rect 67564 24424 67604 24464
rect 69292 24424 69332 24464
rect 66604 24340 66644 24380
rect 50380 24256 50420 24296
rect 69868 24256 69908 24296
rect 75052 24256 75092 24296
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 40204 24172 40244 24212
rect 56236 24172 56276 24212
rect 56428 24172 56468 24212
rect 56620 24172 56660 24212
rect 64012 24172 64052 24212
rect 68716 24172 68756 24212
rect 62668 24088 62708 24128
rect 53068 24004 53108 24044
rect 64012 24004 64052 24044
rect 52780 23920 52820 23960
rect 55660 23920 55700 23960
rect 53164 23836 53204 23876
rect 48748 23752 48788 23792
rect 50764 23752 50804 23792
rect 53836 23752 53876 23792
rect 68812 23752 68852 23792
rect 75148 23752 75188 23792
rect 78988 23752 79028 23792
rect 50380 23668 50420 23708
rect 63916 23668 63956 23708
rect 69100 23584 69140 23624
rect 74860 23584 74900 23624
rect 77356 23584 77396 23624
rect 43372 23500 43412 23540
rect 60748 23500 60788 23540
rect 71308 23500 71348 23540
rect 76204 23500 76244 23540
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 52780 23332 52820 23372
rect 39820 23248 39860 23288
rect 57868 23248 57908 23288
rect 69676 23164 69716 23204
rect 75628 23164 75668 23204
rect 51532 23080 51572 23120
rect 51820 23080 51860 23120
rect 53452 22996 53492 23036
rect 54700 22912 54740 22952
rect 55180 23080 55220 23120
rect 62668 23080 62708 23120
rect 57100 22996 57140 23036
rect 62860 22996 62900 23036
rect 74956 22996 74996 23036
rect 78028 22996 78068 23036
rect 55180 22912 55185 22952
rect 55185 22912 55220 22952
rect 55756 22912 55796 22952
rect 57964 22912 58004 22952
rect 59020 22912 59060 22952
rect 64780 22912 64820 22952
rect 66316 22912 66356 22952
rect 53260 22828 53300 22868
rect 56236 22828 56276 22868
rect 57772 22828 57812 22868
rect 60748 22828 60788 22868
rect 66220 22828 66260 22868
rect 66604 22828 66644 22868
rect 71020 22828 71060 22868
rect 54892 22744 54895 22784
rect 54895 22744 54932 22784
rect 55564 22744 55585 22784
rect 55585 22744 55604 22784
rect 55852 22744 55892 22784
rect 57676 22744 57695 22784
rect 57695 22744 57716 22784
rect 59116 22744 59145 22784
rect 59145 22744 59156 22784
rect 60460 22744 60500 22784
rect 61900 22744 61940 22784
rect 66508 22744 66548 22784
rect 71884 22744 71924 22784
rect 76876 22744 76895 22784
rect 76895 22744 76916 22784
rect 77164 22744 77185 22784
rect 77185 22744 77204 22784
rect 77932 22744 77945 22784
rect 77945 22744 77972 22784
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43468 22492 43508 22532
rect 52396 22492 52436 22532
rect 40108 22156 40148 22196
rect 42412 22156 42452 22196
rect 51628 22156 51668 22196
rect 38860 22072 38900 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 40108 21652 40148 21692
rect 3916 21568 3956 21608
rect 4588 21568 4628 21608
rect 7372 21568 7412 21608
rect 52204 21568 52244 21608
rect 43468 21484 43508 21524
rect 51820 21484 51860 21524
rect 53068 21400 53108 21440
rect 51628 21316 51668 21356
rect 51916 21316 51956 21356
rect 52972 21316 53012 21356
rect 51724 21232 51764 21272
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 51628 21148 51668 21188
rect 52684 21148 52724 21188
rect 52300 20980 52340 21020
rect 52492 20896 52532 20936
rect 50572 20812 50612 20852
rect 52108 20728 52148 20768
rect 52780 20728 52820 20768
rect 10924 20560 10964 20600
rect 52300 20560 52340 20600
rect 52588 20560 52628 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 42796 20392 42836 20432
rect 52780 20308 52820 20348
rect 42796 20140 42836 20180
rect 40108 19972 40148 20012
rect 51916 19972 51956 20012
rect 42412 19888 42452 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 47020 19636 47060 19676
rect 37036 19468 37076 19508
rect 41356 19216 41396 19256
rect 34348 18964 34388 19004
rect 42988 18964 43028 19004
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 50380 18880 50420 18920
rect 41740 18628 41780 18668
rect 7660 18544 7700 18584
rect 32236 18544 32276 18584
rect 40876 18544 40916 18584
rect 40780 18376 40820 18416
rect 43660 18376 43700 18416
rect 34732 18292 34772 18332
rect 7564 18208 7604 18248
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 34348 18124 34388 18164
rect 47500 18376 47540 18416
rect 42988 18292 43028 18332
rect 44620 18292 44660 18332
rect 51916 18208 51956 18248
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 48940 18124 48980 18164
rect 51820 17956 51860 17996
rect 31756 17788 31796 17828
rect 40204 17788 40244 17828
rect 49804 17788 49844 17828
rect 33100 17704 33140 17744
rect 43468 17704 43508 17744
rect 7564 17536 7604 17576
rect 38284 17536 38324 17576
rect 40780 17536 40820 17576
rect 53068 17452 53108 17492
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 56140 17284 56180 17324
rect 56908 17284 56948 17324
rect 57292 17284 57295 17324
rect 57295 17284 57332 17324
rect 57580 17284 57620 17324
rect 59020 17284 59060 17324
rect 59404 17284 59444 17324
rect 59692 17284 59695 17324
rect 59695 17284 59732 17324
rect 60844 17284 60884 17324
rect 61900 17284 61940 17324
rect 63916 17284 63956 17324
rect 64780 17284 64820 17324
rect 66028 17284 66055 17324
rect 66055 17284 66068 17324
rect 66220 17284 66260 17324
rect 69100 17284 69140 17324
rect 71020 17284 71060 17324
rect 77164 17284 77185 17324
rect 77185 17284 77204 17324
rect 53260 17200 53300 17240
rect 56428 17200 56455 17240
rect 56455 17200 56468 17240
rect 56716 17200 56756 17240
rect 57388 17200 57428 17240
rect 57676 17200 57695 17240
rect 57695 17200 57716 17240
rect 58060 17200 58095 17240
rect 58095 17200 58100 17240
rect 58444 17200 58455 17240
rect 58455 17200 58484 17240
rect 58924 17200 58964 17240
rect 59212 17200 59252 17240
rect 60652 17200 60692 17240
rect 61996 17200 62036 17240
rect 65260 17200 65300 17240
rect 66508 17200 66548 17240
rect 76780 17200 76820 17240
rect 54700 17116 54740 17156
rect 65164 17116 65185 17156
rect 65185 17116 65204 17156
rect 66316 17116 66356 17156
rect 66700 17116 66740 17156
rect 68428 17116 68468 17156
rect 70156 17116 70196 17156
rect 32236 17032 32276 17072
rect 42412 17032 42452 17072
rect 43660 17032 43700 17072
rect 35308 16948 35348 16988
rect 37996 16948 38036 16988
rect 40780 16948 40820 16988
rect 40684 16780 40724 16820
rect 40876 16780 40916 16820
rect 50380 16948 50420 16988
rect 72556 17116 72596 17156
rect 75820 17116 75860 17156
rect 66796 17032 66836 17072
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 61036 16612 61076 16652
rect 47500 16528 47540 16568
rect 49804 16528 49844 16568
rect 65740 16528 65780 16568
rect 56332 16444 56372 16484
rect 60748 16360 60788 16400
rect 60940 16360 60980 16400
rect 71788 16360 71828 16400
rect 70924 16276 70964 16316
rect 60460 16192 60500 16232
rect 70828 16192 70868 16232
rect 78508 16192 78548 16232
rect 42796 16108 42836 16148
rect 71020 16108 71060 16148
rect 74860 16108 74900 16148
rect 36748 16024 36788 16064
rect 41164 16024 41204 16064
rect 51148 16024 51188 16064
rect 52204 16024 52244 16064
rect 61420 16024 61460 16064
rect 66604 15940 66644 15980
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 53164 15856 53204 15896
rect 59116 15856 59156 15896
rect 56140 15772 56180 15812
rect 53260 15688 53300 15728
rect 64108 15688 64148 15728
rect 37036 15604 37076 15644
rect 41164 15604 41204 15644
rect 53164 15604 53204 15644
rect 60556 15604 60596 15644
rect 77068 15688 77108 15728
rect 47500 15520 47540 15560
rect 47788 15520 47828 15560
rect 51148 15520 51188 15560
rect 60940 15520 60980 15560
rect 62284 15436 62324 15476
rect 64972 15436 65012 15476
rect 47884 15352 47924 15392
rect 54604 15268 54644 15308
rect 61228 15268 61268 15308
rect 75532 15268 75572 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 56716 14764 56756 14804
rect 60172 14764 60212 14804
rect 60364 14764 60404 14804
rect 70732 14764 70772 14804
rect 43468 14680 43508 14720
rect 47884 14680 47924 14720
rect 51628 14428 51668 14468
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 65164 14344 65204 14384
rect 66316 14344 66356 14384
rect 72556 14344 72596 14384
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 76876 14344 76916 14384
rect 60652 14092 60692 14132
rect 61420 14092 61460 14132
rect 75724 14008 75764 14048
rect 77356 14008 77396 14048
rect 63532 13840 63572 13880
rect 70156 13756 70196 13796
rect 70828 13756 70868 13796
rect 60844 13672 60884 13712
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 67564 13336 67604 13376
rect 51628 13168 51668 13208
rect 65260 13168 65300 13208
rect 66796 13084 66836 13124
rect 60460 12916 60500 12956
rect 67564 12916 67604 12956
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 75724 12832 75764 12872
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 52204 12496 52244 12536
rect 61036 12244 61076 12284
rect 59020 12160 59060 12200
rect 64780 12160 64820 12200
rect 77356 12160 77396 12200
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 44620 12076 44660 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 56140 11992 56180 12032
rect 56044 11908 56084 11948
rect 60172 11656 60212 11696
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 63532 11152 63572 11192
rect 43372 10900 43412 10940
rect 56716 10816 56756 10856
rect 66700 10816 66740 10856
rect 56044 10648 56084 10688
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 68524 10312 68564 10352
rect 47020 10060 47060 10100
rect 66508 10060 66548 10100
rect 68428 10060 68468 10100
rect 71020 10060 71060 10100
rect 75820 10060 75860 10100
rect 43372 9976 43412 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 68524 9304 68564 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 47788 8716 47828 8756
rect 69004 8632 69044 8672
rect 66028 8380 66068 8420
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 56332 7792 56372 7832
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 69004 7540 69044 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 64780 7288 64820 7328
rect 47788 7120 47828 7160
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 65740 6112 65780 6152
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 64972 5944 65012 5984
rect 64780 5860 64820 5900
rect 77644 5860 77684 5900
rect 76876 5692 76916 5732
rect 65356 5608 65396 5648
rect 77164 5608 77204 5648
rect 69004 5524 69044 5564
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 64780 5104 64820 5144
rect 65740 4936 65780 4976
rect 77644 4768 77684 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 66604 4180 66644 4220
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 77068 3508 77108 3548
rect 64780 3424 64820 3464
rect 50188 3340 50228 3380
rect 76780 3256 76820 3296
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 61036 2920 61076 2960
rect 75532 2836 75572 2876
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 61036 1996 61076 2036
rect 65740 1912 65780 1952
rect 61228 1828 61268 1868
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 65740 1156 65780 1196
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 50284 38240 50324 38249
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 39916 29672 39956 29681
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 39916 29084 39956 29632
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 7371 27404 7413 27413
rect 7371 27364 7372 27404
rect 7412 27364 7413 27404
rect 7371 27355 7413 27364
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3916 21608 3956 21617
rect 3916 21449 3956 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 5931 21608 5973 21617
rect 5931 21568 5932 21608
rect 5972 21568 5973 21608
rect 5931 21559 5973 21568
rect 7372 21608 7412 27355
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 39819 23708 39861 23717
rect 39819 23668 39820 23708
rect 39860 23668 39861 23708
rect 39819 23659 39861 23668
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 38859 23288 38901 23297
rect 38859 23248 38860 23288
rect 38900 23248 38901 23288
rect 38859 23239 38901 23248
rect 39820 23288 39860 23659
rect 39820 23239 39860 23248
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 38860 22112 38900 23239
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 38860 22063 38900 22072
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 7372 21559 7412 21568
rect 4588 21474 4628 21559
rect 5932 21449 5972 21559
rect 3915 21440 3957 21449
rect 3915 21400 3916 21440
rect 3956 21400 3957 21440
rect 3915 21391 3957 21400
rect 5931 21440 5973 21449
rect 5931 21400 5932 21440
rect 5972 21400 5973 21440
rect 5931 21391 5973 21400
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 10923 20768 10965 20777
rect 10923 20728 10924 20768
rect 10964 20728 10965 20768
rect 10923 20719 10965 20728
rect 10924 20600 10964 20719
rect 10924 20551 10964 20560
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 39916 20021 39956 29044
rect 42892 28832 42932 28841
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 42892 27656 42932 28792
rect 42892 27236 42932 27616
rect 40204 27068 40244 27077
rect 40108 26984 40148 26993
rect 40012 26732 40052 26741
rect 40012 25808 40052 26692
rect 40012 25759 40052 25768
rect 40108 22196 40148 26944
rect 40204 26312 40244 27028
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 40204 26272 40340 26312
rect 40300 25397 40340 26272
rect 41068 26144 41108 26153
rect 40299 25388 40341 25397
rect 40299 25348 40300 25388
rect 40340 25348 40341 25388
rect 40299 25339 40341 25348
rect 40300 25220 40340 25339
rect 40300 25171 40340 25180
rect 41068 25145 41108 26104
rect 42892 25640 42932 27196
rect 43276 28580 43316 28589
rect 43276 26396 43316 28540
rect 50092 28244 50132 28253
rect 48364 27992 48404 28001
rect 43276 26347 43316 26356
rect 43372 27824 43412 27833
rect 42892 25591 42932 25600
rect 43372 25892 43412 27784
rect 48364 27320 48404 27952
rect 48364 27271 48404 27280
rect 49899 26900 49941 26909
rect 49899 26860 49900 26900
rect 49940 26860 49941 26900
rect 49899 26851 49941 26860
rect 41067 25136 41109 25145
rect 41067 25096 41068 25136
rect 41108 25096 41109 25136
rect 41067 25087 41109 25096
rect 41068 25002 41108 25087
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 41356 24464 41396 24473
rect 40108 21692 40148 22156
rect 40108 21643 40148 21652
rect 40204 24212 40244 24221
rect 39915 20012 39957 20021
rect 39915 19972 39916 20012
rect 39956 19972 39957 20012
rect 39915 19963 39957 19972
rect 40107 20012 40149 20021
rect 40107 19972 40108 20012
rect 40148 19972 40149 20012
rect 40107 19963 40149 19972
rect 40108 19878 40148 19963
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 37036 19508 37076 19517
rect 34348 19004 34388 19013
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 7659 18584 7701 18593
rect 7659 18544 7660 18584
rect 7700 18544 7701 18584
rect 7659 18535 7701 18544
rect 32236 18584 32276 18593
rect 7660 18450 7700 18535
rect 7564 18248 7604 18257
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 7564 17585 7604 18208
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 31756 17828 31796 17837
rect 31756 17585 31796 17788
rect 7563 17576 7605 17585
rect 7563 17536 7564 17576
rect 7604 17536 7605 17576
rect 7563 17527 7605 17536
rect 31755 17576 31797 17585
rect 31755 17536 31756 17576
rect 31796 17536 31797 17576
rect 31755 17527 31797 17536
rect 7564 17442 7604 17527
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 32236 17072 32276 18544
rect 34348 18164 34388 18964
rect 34348 18115 34388 18124
rect 34732 18332 34772 18341
rect 33100 17744 33140 17753
rect 33140 17704 33236 17744
rect 33100 17676 33140 17704
rect 32236 17023 32276 17032
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 33196 15401 33236 17704
rect 34732 16997 34772 18292
rect 34731 16988 34773 16997
rect 34731 16948 34732 16988
rect 34772 16948 34773 16988
rect 34731 16939 34773 16948
rect 35308 16988 35348 16997
rect 35308 16829 35348 16948
rect 35307 16820 35349 16829
rect 35307 16780 35308 16820
rect 35348 16780 35349 16820
rect 35307 16771 35349 16780
rect 36748 16064 36788 16073
rect 33195 15392 33237 15401
rect 33195 15352 33196 15392
rect 33236 15352 33237 15392
rect 33195 15343 33237 15352
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 36748 14981 36788 16024
rect 37036 15644 37076 19468
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 40204 17828 40244 24172
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 41356 19256 41396 24424
rect 43372 23540 43412 25852
rect 49132 26648 49172 26657
rect 45579 25304 45621 25313
rect 45579 25264 45580 25304
rect 45620 25264 45621 25304
rect 45579 25255 45621 25264
rect 45580 25220 45620 25255
rect 49132 25229 49172 26608
rect 49900 26480 49940 26851
rect 45580 25169 45620 25180
rect 49131 25220 49173 25229
rect 49131 25180 49132 25220
rect 49172 25180 49173 25220
rect 49131 25171 49173 25180
rect 48747 23792 48789 23801
rect 48747 23752 48748 23792
rect 48788 23752 48789 23792
rect 48747 23743 48789 23752
rect 48748 23658 48788 23743
rect 43467 23624 43509 23633
rect 43467 23584 43468 23624
rect 43508 23584 43509 23624
rect 43467 23575 43509 23584
rect 43372 23491 43412 23500
rect 43468 22532 43508 23575
rect 42412 22196 42452 22205
rect 42412 19928 42452 22156
rect 43468 21524 43508 22492
rect 43468 21475 43508 21484
rect 42796 20432 42836 20441
rect 42796 20180 42836 20392
rect 42796 20131 42836 20140
rect 42412 19879 42452 19888
rect 47020 19676 47060 19685
rect 41739 19508 41781 19517
rect 41739 19468 41740 19508
rect 41780 19468 41781 19508
rect 41739 19459 41781 19468
rect 41356 19207 41396 19216
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 41740 18668 41780 19459
rect 41835 19424 41877 19433
rect 41835 19384 41836 19424
rect 41876 19384 41877 19424
rect 41835 19375 41877 19384
rect 41740 18619 41780 18628
rect 41836 18593 41876 19375
rect 42988 19004 43028 19013
rect 40876 18584 40916 18593
rect 40204 17779 40244 17788
rect 40780 18416 40820 18425
rect 38284 17576 38324 17585
rect 37996 16988 38036 16999
rect 37996 16913 38036 16948
rect 37995 16904 38037 16913
rect 37995 16864 37996 16904
rect 38036 16864 38037 16904
rect 37995 16855 38037 16864
rect 38284 16493 38324 17536
rect 40780 17576 40820 18376
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 40780 17240 40820 17536
rect 40684 17200 40820 17240
rect 40684 16820 40724 17200
rect 40684 16771 40724 16780
rect 40780 16988 40820 16997
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 38283 16484 38325 16493
rect 38283 16444 38284 16484
rect 38324 16444 38325 16484
rect 38283 16435 38325 16444
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 37036 15595 37076 15604
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 36747 14972 36789 14981
rect 36747 14932 36748 14972
rect 36788 14932 36789 14972
rect 36747 14923 36789 14932
rect 40780 14897 40820 16948
rect 40876 16820 40916 18544
rect 41835 18584 41877 18593
rect 41835 18544 41836 18584
rect 41876 18544 41877 18584
rect 41835 18535 41877 18544
rect 42988 18332 43028 18964
rect 42988 18283 43028 18292
rect 43660 18416 43700 18425
rect 43468 17744 43508 17753
rect 42411 17072 42453 17081
rect 42411 17032 42412 17072
rect 42452 17032 42453 17072
rect 42411 17023 42453 17032
rect 42412 16938 42452 17023
rect 40876 15821 40916 16780
rect 42795 16148 42837 16157
rect 42795 16108 42796 16148
rect 42836 16108 42837 16148
rect 42795 16099 42837 16108
rect 41163 16064 41205 16073
rect 41163 16024 41164 16064
rect 41204 16024 41205 16064
rect 41163 16015 41205 16024
rect 40875 15812 40917 15821
rect 40875 15772 40876 15812
rect 40916 15772 40917 15812
rect 40875 15763 40917 15772
rect 41164 15644 41204 16015
rect 42796 16014 42836 16099
rect 41164 15595 41204 15604
rect 40779 14888 40821 14897
rect 40779 14848 40780 14888
rect 40820 14848 40821 14888
rect 40779 14839 40821 14848
rect 43468 14720 43508 17704
rect 43660 17072 43700 18376
rect 43660 17023 43700 17032
rect 44620 18332 44660 18341
rect 43468 14671 43508 14680
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 44620 12116 44660 18292
rect 44620 12067 44660 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 43372 10940 43412 10949
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 43372 10016 43412 10900
rect 47020 10100 47060 19636
rect 47500 18416 47540 18425
rect 47500 16568 47540 18376
rect 47500 15560 47540 16528
rect 48940 18164 48980 18173
rect 48940 15737 48980 18124
rect 49804 17828 49844 17837
rect 49804 16568 49844 17788
rect 49804 16519 49844 16528
rect 48939 15728 48981 15737
rect 48939 15688 48940 15728
rect 48980 15688 48981 15728
rect 48939 15679 48981 15688
rect 47787 15644 47829 15653
rect 47787 15604 47788 15644
rect 47828 15604 47829 15644
rect 47787 15595 47829 15604
rect 47500 15511 47540 15520
rect 47788 15560 47828 15595
rect 47788 15509 47828 15520
rect 47884 15392 47924 15403
rect 47884 15317 47924 15352
rect 47883 15308 47925 15317
rect 47883 15268 47884 15308
rect 47924 15268 47925 15308
rect 47883 15259 47925 15268
rect 47884 14720 47924 15259
rect 49900 14813 49940 26440
rect 49995 25388 50037 25397
rect 49995 25348 49996 25388
rect 50036 25348 50037 25388
rect 49995 25339 50037 25348
rect 49899 14804 49941 14813
rect 49899 14764 49900 14804
rect 49940 14764 49941 14804
rect 49899 14755 49941 14764
rect 47884 14671 47924 14680
rect 49996 14225 50036 25339
rect 50092 14729 50132 28204
rect 50187 26984 50229 26993
rect 50187 26944 50188 26984
rect 50228 26944 50229 26984
rect 50187 26935 50229 26944
rect 50091 14720 50133 14729
rect 50091 14680 50092 14720
rect 50132 14680 50133 14720
rect 50091 14671 50133 14680
rect 49995 14216 50037 14225
rect 49995 14176 49996 14216
rect 50036 14176 50037 14216
rect 49995 14167 50037 14176
rect 47020 10051 47060 10060
rect 43372 9967 43412 9976
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 47788 8756 47828 8765
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 47788 7160 47828 8716
rect 47788 7111 47828 7120
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 50188 3380 50228 26935
rect 50284 15569 50324 38200
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 66316 37148 66356 37157
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 56620 36308 56660 36317
rect 56620 35636 56660 36268
rect 61708 36308 61748 36317
rect 61228 36056 61268 36065
rect 56620 35587 56660 35596
rect 61036 35720 61076 35729
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 61036 35300 61076 35680
rect 61228 35552 61268 36016
rect 61708 35804 61748 36268
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 61708 35755 61748 35764
rect 61228 35503 61268 35512
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 61036 35048 61076 35260
rect 61036 34999 61076 35008
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 61228 33368 61268 33377
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 55372 33284 55412 33293
rect 55372 32696 55412 33244
rect 55372 32647 55412 32656
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 56428 31856 56468 31865
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 53068 31772 53108 31781
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 51820 30344 51860 30353
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 50380 29084 50420 29093
rect 50380 24296 50420 29044
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 51532 25556 51572 25565
rect 50380 24247 50420 24256
rect 50572 25220 50612 25229
rect 50380 23708 50420 23717
rect 50380 21533 50420 23668
rect 50379 21524 50421 21533
rect 50379 21484 50380 21524
rect 50420 21484 50421 21524
rect 50379 21475 50421 21484
rect 50572 20852 50612 25180
rect 50764 25136 50804 25145
rect 50764 23792 50804 25096
rect 50764 23743 50804 23752
rect 51532 23120 51572 25516
rect 51627 24632 51669 24641
rect 51627 24592 51628 24632
rect 51668 24592 51669 24632
rect 51627 24583 51669 24592
rect 51532 23071 51572 23080
rect 51628 22196 51668 24583
rect 51723 24548 51765 24557
rect 51723 24508 51724 24548
rect 51764 24508 51765 24548
rect 51723 24499 51765 24508
rect 51628 22147 51668 22156
rect 50572 20803 50612 20812
rect 51628 21356 51668 21365
rect 51628 21188 51668 21316
rect 51724 21272 51764 24499
rect 51820 23969 51860 30304
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 52204 28496 52244 28505
rect 52204 27236 52244 28456
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 52204 27187 52244 27196
rect 52972 27068 53012 27077
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 52972 26480 53012 27028
rect 52972 26431 53012 26440
rect 51916 25472 51956 25481
rect 51916 24809 51956 25432
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 52780 24968 52820 24977
rect 51915 24800 51957 24809
rect 51915 24760 51916 24800
rect 51956 24760 51957 24800
rect 51915 24751 51957 24760
rect 51916 24548 51956 24751
rect 52107 24716 52149 24725
rect 52107 24676 52108 24716
rect 52148 24676 52149 24716
rect 52107 24667 52149 24676
rect 51916 24499 51956 24508
rect 51819 23960 51861 23969
rect 51819 23920 51820 23960
rect 51860 23920 51861 23960
rect 51819 23911 51861 23920
rect 51820 23120 51860 23911
rect 51820 23071 51860 23080
rect 51819 22784 51861 22793
rect 51819 22744 51820 22784
rect 51860 22744 51861 22784
rect 51819 22735 51861 22744
rect 51820 21524 51860 22735
rect 51820 21475 51860 21484
rect 51724 21223 51764 21232
rect 51916 21356 51956 21365
rect 51628 19517 51668 21148
rect 51916 20777 51956 21316
rect 51915 20768 51957 20777
rect 51915 20728 51916 20768
rect 51956 20728 51957 20768
rect 51915 20719 51957 20728
rect 52108 20768 52148 24667
rect 52780 23960 52820 24928
rect 52780 23911 52820 23920
rect 53068 24044 53108 31732
rect 53068 23885 53108 24004
rect 53164 29924 53204 29933
rect 53067 23876 53109 23885
rect 53067 23836 53068 23876
rect 53108 23836 53109 23876
rect 53067 23827 53109 23836
rect 53164 23876 53204 29884
rect 53356 27992 53396 28001
rect 53356 25892 53396 27952
rect 55659 27404 55701 27413
rect 55659 27364 55660 27404
rect 55700 27364 55701 27404
rect 55659 27355 55701 27364
rect 53356 25843 53396 25852
rect 53164 23827 53204 23836
rect 54508 25640 54548 25649
rect 53836 23792 53876 23801
rect 52587 23456 52629 23465
rect 52587 23416 52588 23456
rect 52628 23416 52629 23456
rect 52587 23407 52629 23416
rect 53739 23456 53781 23465
rect 53739 23416 53740 23456
rect 53780 23416 53781 23456
rect 53739 23407 53781 23416
rect 52203 23204 52245 23213
rect 52203 23164 52204 23204
rect 52244 23164 52245 23204
rect 52203 23155 52245 23164
rect 52204 21608 52244 23155
rect 52299 23120 52341 23129
rect 52299 23080 52300 23120
rect 52340 23080 52341 23120
rect 52299 23071 52341 23080
rect 52204 21559 52244 21568
rect 52300 21020 52340 23071
rect 52395 22868 52437 22877
rect 52395 22828 52396 22868
rect 52436 22828 52437 22868
rect 52395 22819 52437 22828
rect 52396 22532 52436 22819
rect 52396 22483 52436 22492
rect 52491 21608 52533 21617
rect 52491 21568 52492 21608
rect 52532 21568 52533 21608
rect 52491 21559 52533 21568
rect 52300 20971 52340 20980
rect 52492 20936 52532 21559
rect 52492 20887 52532 20896
rect 52108 20719 52148 20728
rect 52300 20600 52340 20609
rect 51915 20012 51957 20021
rect 51915 19972 51916 20012
rect 51956 19972 52052 20012
rect 51915 19963 51957 19972
rect 51916 19878 51956 19963
rect 51627 19508 51669 19517
rect 51627 19468 51628 19508
rect 51668 19468 51669 19508
rect 51627 19459 51669 19468
rect 50380 18920 50420 18929
rect 50380 16988 50420 18880
rect 51916 18248 51956 18257
rect 51820 17996 51860 18005
rect 51820 17249 51860 17956
rect 51819 17240 51861 17249
rect 51819 17200 51820 17240
rect 51860 17200 51861 17240
rect 51819 17191 51861 17200
rect 51916 17165 51956 18208
rect 51915 17156 51957 17165
rect 51915 17116 51916 17156
rect 51956 17116 51957 17156
rect 51915 17107 51957 17116
rect 50380 16939 50420 16948
rect 51148 16064 51188 16075
rect 51148 15989 51188 16024
rect 51147 15980 51189 15989
rect 51147 15940 51148 15980
rect 51188 15940 51189 15980
rect 51147 15931 51189 15940
rect 50283 15560 50325 15569
rect 50283 15520 50284 15560
rect 50324 15520 50325 15560
rect 50283 15511 50325 15520
rect 51148 15560 51188 15931
rect 52012 15821 52052 19972
rect 52300 19433 52340 20560
rect 52588 20600 52628 23407
rect 52683 23372 52725 23381
rect 52683 23332 52684 23372
rect 52724 23332 52725 23372
rect 52683 23323 52725 23332
rect 52780 23372 52820 23381
rect 52684 21188 52724 23323
rect 52684 21139 52724 21148
rect 52588 20551 52628 20560
rect 52780 20768 52820 23332
rect 53740 23297 53780 23407
rect 53739 23288 53781 23297
rect 53739 23248 53740 23288
rect 53780 23248 53781 23288
rect 53739 23239 53781 23248
rect 53836 23204 53876 23752
rect 54508 23213 54548 25600
rect 54891 24548 54933 24557
rect 54891 24508 54892 24548
rect 54932 24508 54933 24548
rect 54891 24499 54933 24508
rect 54219 23204 54261 23213
rect 53836 23164 54220 23204
rect 54260 23164 54261 23204
rect 54219 23155 54261 23164
rect 54507 23204 54549 23213
rect 54507 23164 54508 23204
rect 54548 23164 54549 23204
rect 54507 23155 54549 23164
rect 52875 23036 52917 23045
rect 52875 22996 52876 23036
rect 52916 22996 52917 23036
rect 52875 22987 52917 22996
rect 53451 23036 53493 23045
rect 53451 22996 53452 23036
rect 53492 22996 53493 23036
rect 53451 22987 53493 22996
rect 53643 23036 53685 23045
rect 53643 22996 53644 23036
rect 53684 22996 53685 23036
rect 53643 22987 53685 22996
rect 52876 21617 52916 22987
rect 52971 22952 53013 22961
rect 52971 22912 52972 22952
rect 53012 22912 53013 22952
rect 52971 22903 53013 22912
rect 52875 21608 52917 21617
rect 52875 21568 52876 21608
rect 52916 21568 52917 21608
rect 52875 21559 52917 21568
rect 52972 21356 53012 22903
rect 53452 22902 53492 22987
rect 53260 22868 53300 22877
rect 53068 22828 53260 22868
rect 53068 21440 53108 22828
rect 53260 22819 53300 22828
rect 53355 22784 53397 22793
rect 53644 22784 53684 22987
rect 54699 22952 54741 22961
rect 54699 22912 54700 22952
rect 54740 22912 54741 22952
rect 54699 22903 54741 22912
rect 54700 22818 54740 22903
rect 53355 22744 53356 22784
rect 53396 22744 53684 22784
rect 54892 22784 54932 24499
rect 55660 23960 55700 27355
rect 56139 24968 56181 24977
rect 56139 24928 56140 24968
rect 56180 24928 56181 24968
rect 56139 24919 56181 24928
rect 56140 24834 56180 24919
rect 55755 24716 55797 24725
rect 55755 24676 55756 24716
rect 55796 24676 55797 24716
rect 55755 24667 55797 24676
rect 55660 23911 55700 23920
rect 55563 23372 55605 23381
rect 55563 23332 55564 23372
rect 55604 23332 55605 23372
rect 55563 23323 55605 23332
rect 55179 23288 55221 23297
rect 55179 23248 55180 23288
rect 55220 23248 55221 23288
rect 55179 23239 55221 23248
rect 55083 23120 55125 23129
rect 55083 23080 55084 23120
rect 55124 23080 55125 23120
rect 55083 23071 55125 23080
rect 55180 23120 55220 23239
rect 55180 23071 55220 23080
rect 55084 22952 55124 23071
rect 55180 22952 55220 22961
rect 55084 22912 55180 22952
rect 55180 22903 55220 22912
rect 53355 22735 53397 22744
rect 54892 22735 54932 22744
rect 55564 22784 55604 23323
rect 55756 22952 55796 24667
rect 56235 24212 56277 24221
rect 56235 24172 56236 24212
rect 56276 24172 56277 24212
rect 56235 24163 56277 24172
rect 56428 24212 56468 31816
rect 61132 31352 61172 31361
rect 61132 30596 61172 31312
rect 61132 30547 61172 30556
rect 61228 30260 61268 33328
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 63532 32192 63572 32201
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 61228 30211 61268 30220
rect 62668 31520 62708 31529
rect 62668 30428 62708 31480
rect 63532 31436 63572 32152
rect 63532 31387 63572 31396
rect 61611 26984 61653 26993
rect 61611 26944 61612 26984
rect 61652 26944 61653 26984
rect 61611 26935 61653 26944
rect 58443 26900 58485 26909
rect 58443 26860 58444 26900
rect 58484 26860 58485 26900
rect 58443 26851 58485 26860
rect 61612 26900 61652 26935
rect 58444 26766 58484 26851
rect 61612 26849 61652 26860
rect 58731 25388 58773 25397
rect 58731 25348 58732 25388
rect 58772 25348 58773 25388
rect 58731 25339 58773 25348
rect 58732 25254 58772 25339
rect 59115 25304 59157 25313
rect 59115 25264 59116 25304
rect 59156 25264 59157 25304
rect 59115 25255 59157 25264
rect 57963 25136 58005 25145
rect 57963 25096 57964 25136
rect 58004 25096 58005 25136
rect 57963 25087 58005 25096
rect 57579 24968 57621 24977
rect 57579 24928 57580 24968
rect 57620 24928 57621 24968
rect 57579 24919 57621 24928
rect 57580 24834 57620 24919
rect 57771 24632 57813 24641
rect 57771 24592 57772 24632
rect 57812 24592 57813 24632
rect 57771 24583 57813 24592
rect 56236 24078 56276 24163
rect 56428 23549 56468 24172
rect 56619 24212 56661 24221
rect 56619 24172 56620 24212
rect 56660 24172 56661 24212
rect 56619 24163 56661 24172
rect 56620 24078 56660 24163
rect 57675 23708 57717 23717
rect 57675 23668 57676 23708
rect 57716 23668 57717 23708
rect 57675 23659 57717 23668
rect 55851 23540 55893 23549
rect 55851 23500 55852 23540
rect 55892 23500 55893 23540
rect 55851 23491 55893 23500
rect 56427 23540 56469 23549
rect 56427 23500 56428 23540
rect 56468 23500 56469 23540
rect 56427 23491 56469 23500
rect 55756 22903 55796 22912
rect 55564 22735 55604 22744
rect 55852 22784 55892 23491
rect 56235 23456 56277 23465
rect 56235 23416 56236 23456
rect 56276 23416 56277 23456
rect 56235 23407 56277 23416
rect 56236 22868 56276 23407
rect 57100 23036 57140 23045
rect 57100 22877 57140 22996
rect 56236 22819 56276 22828
rect 57099 22868 57141 22877
rect 57099 22828 57100 22868
rect 57140 22828 57141 22868
rect 57099 22819 57141 22828
rect 55852 22735 55892 22744
rect 57676 22784 57716 23659
rect 57772 22868 57812 24583
rect 57867 23708 57909 23717
rect 57867 23668 57868 23708
rect 57908 23668 57909 23708
rect 57867 23659 57909 23668
rect 57868 23288 57908 23659
rect 57868 23239 57908 23248
rect 57964 22952 58004 25087
rect 58252 24464 58292 24473
rect 58252 23717 58292 24424
rect 58251 23708 58293 23717
rect 58251 23668 58252 23708
rect 58292 23668 58293 23708
rect 58251 23659 58293 23668
rect 59019 23624 59061 23633
rect 59019 23584 59020 23624
rect 59060 23584 59061 23624
rect 59019 23575 59061 23584
rect 57964 22903 58004 22912
rect 59020 22952 59060 23575
rect 59020 22903 59060 22912
rect 57772 22819 57812 22828
rect 57676 22735 57716 22744
rect 59116 22784 59156 25255
rect 61899 25220 61941 25229
rect 61899 25180 61900 25220
rect 61940 25180 61941 25220
rect 61899 25171 61941 25180
rect 60459 23792 60501 23801
rect 60459 23752 60460 23792
rect 60500 23752 60501 23792
rect 60459 23743 60501 23752
rect 59116 22735 59156 22744
rect 60460 22784 60500 23743
rect 60748 23540 60788 23549
rect 60748 23045 60788 23500
rect 60747 23036 60789 23045
rect 60747 22996 60748 23036
rect 60788 22996 60789 23036
rect 60747 22987 60789 22996
rect 60748 22868 60788 22987
rect 60748 22819 60788 22828
rect 60460 22735 60500 22744
rect 61900 22784 61940 25171
rect 62668 24128 62708 30388
rect 63916 31352 63956 31361
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 62668 23120 62708 24088
rect 62668 23071 62708 23080
rect 62860 27740 62900 27749
rect 62860 23036 62900 27700
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 63916 23708 63956 31312
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 64012 30512 64052 30521
rect 64012 24212 64052 30472
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 64204 29336 64244 29345
rect 64204 26900 64244 29296
rect 65836 29336 65876 29345
rect 65836 28580 65876 29296
rect 66316 28664 66356 37108
rect 76204 37148 76244 37157
rect 74188 36896 74228 36905
rect 74188 36560 74228 36856
rect 74188 36511 74228 36520
rect 75628 36476 75668 36485
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 73804 35888 73844 35897
rect 73804 35216 73844 35848
rect 72844 33032 72884 33041
rect 72364 32780 72404 32789
rect 72364 30428 72404 32740
rect 72844 32108 72884 32992
rect 72844 31688 72884 32068
rect 72844 31639 72884 31648
rect 73612 32528 73652 32537
rect 72364 30379 72404 30388
rect 73324 31520 73364 31529
rect 66316 28615 66356 28624
rect 71020 28832 71060 28841
rect 65836 28531 65876 28540
rect 70924 28496 70964 28505
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 64204 26851 64244 26860
rect 68716 27320 68756 27329
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 66604 25556 66644 25565
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 66604 24380 66644 25516
rect 67564 25220 67604 25229
rect 67564 24464 67604 25180
rect 67564 24415 67604 24424
rect 66604 24331 66644 24340
rect 64012 24044 64052 24172
rect 68716 24212 68756 27280
rect 69100 27320 69140 27329
rect 68716 24163 68756 24172
rect 68812 27236 68852 27245
rect 64012 23995 64052 24004
rect 64779 23960 64821 23969
rect 64779 23920 64780 23960
rect 64820 23920 64821 23960
rect 64779 23911 64821 23920
rect 63916 23659 63956 23668
rect 62860 22987 62900 22996
rect 64780 22952 64820 23911
rect 66507 23876 66549 23885
rect 66507 23836 66508 23876
rect 66548 23836 66549 23876
rect 66507 23827 66549 23836
rect 66315 23540 66357 23549
rect 66315 23500 66316 23540
rect 66356 23500 66357 23540
rect 66315 23491 66357 23500
rect 66219 23204 66261 23213
rect 66219 23164 66220 23204
rect 66260 23164 66261 23204
rect 66219 23155 66261 23164
rect 64780 22903 64820 22912
rect 66220 22868 66260 23155
rect 66316 22952 66356 23491
rect 66316 22903 66356 22912
rect 66220 22819 66260 22828
rect 61900 22735 61940 22744
rect 66508 22784 66548 23827
rect 68812 23792 68852 27196
rect 68812 23743 68852 23752
rect 66603 23708 66645 23717
rect 66603 23668 66604 23708
rect 66644 23668 66645 23708
rect 66603 23659 66645 23668
rect 66604 22868 66644 23659
rect 69100 23624 69140 27280
rect 69676 27320 69716 27329
rect 69292 26312 69332 26321
rect 69292 24464 69332 26272
rect 69292 24415 69332 24424
rect 69100 23575 69140 23584
rect 69676 23204 69716 27280
rect 70924 26900 70964 28456
rect 70924 26851 70964 26860
rect 69772 26480 69812 26489
rect 69772 25388 69812 26440
rect 69772 25339 69812 25348
rect 69868 25976 69908 25985
rect 69868 24296 69908 25936
rect 69868 24247 69908 24256
rect 69676 23155 69716 23164
rect 66604 22819 66644 22828
rect 71020 22868 71060 28792
rect 73324 28580 73364 31480
rect 73612 31352 73652 32488
rect 73612 31303 73652 31312
rect 73804 30260 73844 35176
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 75112 33284 75480 33293
rect 75152 33244 75194 33284
rect 75234 33244 75276 33284
rect 75316 33244 75358 33284
rect 75398 33244 75440 33284
rect 75112 33235 75480 33244
rect 75112 31772 75480 31781
rect 75152 31732 75194 31772
rect 75234 31732 75276 31772
rect 75316 31732 75358 31772
rect 75398 31732 75440 31772
rect 75112 31723 75480 31732
rect 73804 30211 73844 30220
rect 74956 30260 74996 30269
rect 73324 27572 73364 28540
rect 73324 27523 73364 27532
rect 71308 27320 71348 27329
rect 71308 23540 71348 27280
rect 74860 27152 74900 27161
rect 71692 26984 71732 26993
rect 71692 26648 71732 26944
rect 71692 26599 71732 26608
rect 74860 23624 74900 27112
rect 74860 23575 74900 23584
rect 71308 23491 71348 23500
rect 74956 23036 74996 30220
rect 75112 30260 75480 30269
rect 75152 30220 75194 30260
rect 75234 30220 75276 30260
rect 75316 30220 75358 30260
rect 75398 30220 75440 30260
rect 75112 30211 75480 30220
rect 75112 28748 75480 28757
rect 75152 28708 75194 28748
rect 75234 28708 75276 28748
rect 75316 28708 75358 28748
rect 75398 28708 75440 28748
rect 75112 28699 75480 28708
rect 75112 27236 75480 27245
rect 75152 27196 75194 27236
rect 75234 27196 75276 27236
rect 75316 27196 75358 27236
rect 75398 27196 75440 27236
rect 75112 27187 75480 27196
rect 75112 25724 75480 25733
rect 75152 25684 75194 25724
rect 75234 25684 75276 25724
rect 75316 25684 75358 25724
rect 75398 25684 75440 25724
rect 75112 25675 75480 25684
rect 75052 25304 75092 25313
rect 75052 24296 75092 25264
rect 75052 24247 75092 24256
rect 75148 23792 75188 23801
rect 75148 23129 75188 23752
rect 75628 23204 75668 36436
rect 76204 23540 76244 37108
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 76684 35972 76724 35981
rect 76724 35932 76820 35972
rect 76684 35923 76724 35932
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 76780 35132 76820 35932
rect 76780 35083 76820 35092
rect 76876 35216 76916 35225
rect 76780 34964 76820 34973
rect 76352 34040 76720 34049
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 76352 32528 76720 32537
rect 76392 32488 76434 32528
rect 76474 32488 76516 32528
rect 76556 32488 76598 32528
rect 76638 32488 76680 32528
rect 76352 32479 76720 32488
rect 76352 31016 76720 31025
rect 76392 30976 76434 31016
rect 76474 30976 76516 31016
rect 76556 30976 76598 31016
rect 76638 30976 76680 31016
rect 76352 30967 76720 30976
rect 76352 29504 76720 29513
rect 76392 29464 76434 29504
rect 76474 29464 76516 29504
rect 76556 29464 76598 29504
rect 76638 29464 76680 29504
rect 76352 29455 76720 29464
rect 76352 27992 76720 28001
rect 76392 27952 76434 27992
rect 76474 27952 76516 27992
rect 76556 27952 76598 27992
rect 76638 27952 76680 27992
rect 76352 27943 76720 27952
rect 76352 26480 76720 26489
rect 76392 26440 76434 26480
rect 76474 26440 76516 26480
rect 76556 26440 76598 26480
rect 76638 26440 76680 26480
rect 76352 26431 76720 26440
rect 76780 25136 76820 34924
rect 76780 25087 76820 25096
rect 76352 24968 76720 24977
rect 76392 24928 76434 24968
rect 76474 24928 76516 24968
rect 76556 24928 76598 24968
rect 76638 24928 76680 24968
rect 76352 24919 76720 24928
rect 76204 23491 76244 23500
rect 75628 23155 75668 23164
rect 75147 23120 75189 23129
rect 75147 23080 75148 23120
rect 75188 23080 75189 23120
rect 75147 23071 75189 23080
rect 74956 22987 74996 22996
rect 71020 22819 71060 22828
rect 71884 22793 71924 22878
rect 66508 22735 66548 22744
rect 71883 22784 71925 22793
rect 71883 22744 71884 22784
rect 71924 22744 71925 22784
rect 71883 22735 71925 22744
rect 76876 22784 76916 35176
rect 77356 34292 77396 34301
rect 76876 22735 76916 22744
rect 77164 33704 77204 33713
rect 77164 22784 77204 33664
rect 77356 33452 77396 34252
rect 77260 31352 77300 31361
rect 77260 30260 77300 31312
rect 77260 30211 77300 30220
rect 77260 28076 77300 28085
rect 77260 26144 77300 28036
rect 77260 25052 77300 26104
rect 77260 25003 77300 25012
rect 77356 23624 77396 33412
rect 77932 34124 77972 34133
rect 77932 32276 77972 34084
rect 77932 32227 77972 32236
rect 78028 30260 78068 30269
rect 77356 23575 77396 23584
rect 77932 28916 77972 28925
rect 77164 22735 77204 22744
rect 77932 22784 77972 28876
rect 78028 23036 78068 30220
rect 78987 24800 79029 24809
rect 78987 24760 78988 24800
rect 79028 24760 79029 24800
rect 78987 24751 79029 24760
rect 78988 23801 79028 24751
rect 78987 23792 79029 23801
rect 78987 23752 78988 23792
rect 79028 23752 79029 23792
rect 78987 23743 79029 23752
rect 78988 23658 79028 23743
rect 78028 22987 78068 22996
rect 77932 22735 77972 22744
rect 53068 21391 53108 21400
rect 52972 21307 53012 21316
rect 52780 20348 52820 20728
rect 52780 20299 52820 20308
rect 52299 19424 52341 19433
rect 52299 19384 52300 19424
rect 52340 19384 52341 19424
rect 52299 19375 52341 19384
rect 53068 17492 53108 17501
rect 53068 17240 53108 17452
rect 56140 17324 56180 17333
rect 53260 17240 53300 17249
rect 53068 17200 53260 17240
rect 53260 17191 53300 17200
rect 56140 17165 56180 17284
rect 56908 17324 56948 17333
rect 56428 17240 56468 17249
rect 54700 17156 54740 17165
rect 54700 16913 54740 17116
rect 56139 17156 56181 17165
rect 56139 17116 56140 17156
rect 56180 17116 56181 17156
rect 56139 17107 56181 17116
rect 56331 17156 56373 17165
rect 56331 17116 56332 17156
rect 56372 17116 56373 17156
rect 56331 17107 56373 17116
rect 54699 16904 54741 16913
rect 54699 16864 54700 16904
rect 54740 16864 54741 16904
rect 54699 16855 54741 16864
rect 56332 16484 56372 17107
rect 52204 16064 52244 16073
rect 52204 15905 52244 16024
rect 52203 15896 52245 15905
rect 52203 15856 52204 15896
rect 52244 15856 52245 15896
rect 52203 15847 52245 15856
rect 53164 15896 53204 15905
rect 52011 15812 52053 15821
rect 52011 15772 52012 15812
rect 52052 15772 52053 15812
rect 52011 15763 52053 15772
rect 51148 15511 51188 15520
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 51628 14468 51668 14477
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 51628 13208 51668 14428
rect 51628 13159 51668 13168
rect 52204 12536 52244 15847
rect 53164 15644 53204 15856
rect 56140 15812 56180 15821
rect 53259 15728 53301 15737
rect 53259 15688 53260 15728
rect 53300 15688 53301 15728
rect 53259 15679 53301 15688
rect 53164 15595 53204 15604
rect 53260 15594 53300 15679
rect 54603 15560 54645 15569
rect 54603 15520 54604 15560
rect 54644 15520 54645 15560
rect 54603 15511 54645 15520
rect 54604 15308 54644 15511
rect 54604 15259 54644 15268
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 52204 12487 52244 12496
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 56140 12032 56180 15772
rect 56140 11983 56180 11992
rect 56044 11948 56084 11957
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 56044 10688 56084 11908
rect 56044 10639 56084 10648
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 56332 7832 56372 16444
rect 56428 15485 56468 17200
rect 56716 17240 56756 17249
rect 56716 16493 56756 17200
rect 56811 17240 56853 17249
rect 56908 17240 56948 17284
rect 56811 17200 56812 17240
rect 56852 17200 56948 17240
rect 57292 17324 57332 17333
rect 56811 17191 56853 17200
rect 57292 16997 57332 17284
rect 57580 17324 57620 17333
rect 57388 17240 57428 17249
rect 57291 16988 57333 16997
rect 57291 16948 57292 16988
rect 57332 16948 57333 16988
rect 57291 16939 57333 16948
rect 57388 16829 57428 17200
rect 57580 17081 57620 17284
rect 59020 17324 59060 17333
rect 57676 17240 57716 17249
rect 57579 17072 57621 17081
rect 57579 17032 57580 17072
rect 57620 17032 57621 17072
rect 57579 17023 57621 17032
rect 57387 16820 57429 16829
rect 57387 16780 57388 16820
rect 57428 16780 57429 16820
rect 57387 16771 57429 16780
rect 56715 16484 56757 16493
rect 56715 16444 56716 16484
rect 56756 16444 56757 16484
rect 56715 16435 56757 16444
rect 56427 15476 56469 15485
rect 56427 15436 56428 15476
rect 56468 15436 56469 15476
rect 56427 15427 56469 15436
rect 57676 15401 57716 17200
rect 58060 17240 58100 17249
rect 57675 15392 57717 15401
rect 57675 15352 57676 15392
rect 57716 15352 57717 15392
rect 57675 15343 57717 15352
rect 58060 14981 58100 17200
rect 58444 17240 58484 17249
rect 58059 14972 58101 14981
rect 58059 14932 58060 14972
rect 58100 14932 58101 14972
rect 58059 14923 58101 14932
rect 58444 14897 58484 17200
rect 58924 17240 58964 17249
rect 58924 16073 58964 17200
rect 59020 16157 59060 17284
rect 59404 17324 59444 17333
rect 59212 17240 59252 17249
rect 59019 16148 59061 16157
rect 59019 16108 59020 16148
rect 59060 16108 59061 16148
rect 59019 16099 59061 16108
rect 58923 16064 58965 16073
rect 58923 16024 58924 16064
rect 58964 16024 58965 16064
rect 58923 16015 58965 16024
rect 59116 15896 59156 15905
rect 58443 14888 58485 14897
rect 58443 14848 58444 14888
rect 58484 14848 58485 14888
rect 58443 14839 58485 14848
rect 56716 14804 56756 14813
rect 56716 10856 56756 14764
rect 59116 14225 59156 15856
rect 59115 14216 59157 14225
rect 59115 14176 59116 14216
rect 59156 14176 59157 14216
rect 59115 14167 59157 14176
rect 59020 12200 59060 12209
rect 59212 12200 59252 17200
rect 59404 15653 59444 17284
rect 59692 17324 59732 17333
rect 59403 15644 59445 15653
rect 59403 15604 59404 15644
rect 59444 15604 59445 15644
rect 59403 15595 59445 15604
rect 59692 15317 59732 17284
rect 60844 17324 60884 17333
rect 60652 17240 60692 17249
rect 60459 16904 60501 16913
rect 60459 16864 60460 16904
rect 60500 16864 60501 16904
rect 60459 16855 60501 16864
rect 60460 16232 60500 16855
rect 59691 15308 59733 15317
rect 59691 15268 59692 15308
rect 59732 15268 59733 15308
rect 59691 15259 59733 15268
rect 59060 12160 59252 12200
rect 60172 14804 60212 14813
rect 59020 12151 59060 12160
rect 60172 11696 60212 14764
rect 60363 14804 60405 14813
rect 60363 14764 60364 14804
rect 60404 14764 60405 14804
rect 60363 14755 60405 14764
rect 60364 14670 60404 14755
rect 60460 12956 60500 16192
rect 60555 15728 60597 15737
rect 60555 15688 60556 15728
rect 60596 15688 60597 15728
rect 60555 15679 60597 15688
rect 60556 15644 60596 15679
rect 60556 15593 60596 15604
rect 60652 14132 60692 17200
rect 60748 16400 60788 16409
rect 60748 16325 60788 16360
rect 60747 16316 60789 16325
rect 60747 16276 60748 16316
rect 60788 16276 60789 16316
rect 60747 16267 60789 16276
rect 60748 15821 60788 16267
rect 60747 15812 60789 15821
rect 60747 15772 60748 15812
rect 60788 15772 60789 15812
rect 60747 15763 60789 15772
rect 60652 14083 60692 14092
rect 60844 13712 60884 17284
rect 61900 17324 61940 17333
rect 61036 16652 61076 16661
rect 60940 16400 60980 16409
rect 60940 15560 60980 16360
rect 60940 15511 60980 15520
rect 60844 13663 60884 13672
rect 60460 12907 60500 12916
rect 61036 12284 61076 16612
rect 61420 16064 61460 16073
rect 61036 12235 61076 12244
rect 61228 15308 61268 15317
rect 60172 11647 60212 11656
rect 56716 10807 56756 10816
rect 56332 7783 56372 7792
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 50188 3331 50228 3340
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 61036 2960 61076 2969
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 61036 2036 61076 2920
rect 61036 1987 61076 1996
rect 61228 1868 61268 15268
rect 61420 14132 61460 16024
rect 61900 15905 61940 17284
rect 63916 17324 63956 17333
rect 61996 17240 62036 17249
rect 61996 15989 62036 17200
rect 63916 17165 63956 17284
rect 64780 17324 64820 17333
rect 63915 17156 63957 17165
rect 63915 17116 63916 17156
rect 63956 17116 63957 17156
rect 63915 17107 63957 17116
rect 61995 15980 62037 15989
rect 61995 15940 61996 15980
rect 62036 15940 62037 15980
rect 61995 15931 62037 15940
rect 61899 15896 61941 15905
rect 61899 15856 61900 15896
rect 61940 15856 61941 15896
rect 61899 15847 61941 15856
rect 64107 15728 64149 15737
rect 64107 15688 64108 15728
rect 64148 15688 64149 15728
rect 64107 15679 64149 15688
rect 64108 15594 64148 15679
rect 61899 15476 61941 15485
rect 61899 15436 61900 15476
rect 61940 15436 61941 15476
rect 61899 15427 61941 15436
rect 62283 15476 62325 15485
rect 62283 15436 62284 15476
rect 62324 15436 62325 15476
rect 62283 15427 62325 15436
rect 61900 14729 61940 15427
rect 62284 15342 62324 15427
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 61899 14720 61941 14729
rect 61899 14680 61900 14720
rect 61940 14680 61941 14720
rect 61899 14671 61941 14680
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 61420 14083 61460 14092
rect 63532 13880 63572 13889
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 63532 11192 63572 13840
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 64780 12200 64820 17284
rect 66028 17324 66068 17333
rect 65260 17240 65300 17249
rect 65164 17156 65204 17165
rect 64780 12151 64820 12160
rect 64972 15476 65012 15485
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 63532 11143 63572 11152
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 64780 7328 64820 7337
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 64780 5900 64820 7288
rect 64972 5984 65012 15436
rect 65164 14384 65204 17116
rect 65164 14335 65204 14344
rect 65260 13208 65300 17200
rect 65355 16568 65397 16577
rect 65355 16528 65356 16568
rect 65396 16528 65397 16568
rect 65355 16519 65397 16528
rect 65739 16568 65781 16577
rect 65739 16528 65740 16568
rect 65780 16528 65781 16568
rect 65739 16519 65781 16528
rect 65260 13159 65300 13168
rect 64972 5935 65012 5944
rect 64780 5851 64820 5860
rect 65356 5648 65396 16519
rect 65740 16434 65780 16519
rect 66028 8420 66068 17284
rect 66220 17324 66260 17333
rect 66220 16913 66260 17284
rect 69100 17324 69140 17333
rect 66508 17240 66548 17249
rect 66316 17156 66356 17165
rect 66219 16904 66261 16913
rect 66219 16864 66220 16904
rect 66260 16864 66261 16904
rect 66219 16855 66261 16864
rect 66316 14384 66356 17116
rect 66316 14335 66356 14344
rect 66508 10100 66548 17200
rect 66700 17156 66740 17165
rect 66508 10051 66548 10060
rect 66604 15980 66644 15989
rect 66028 8371 66068 8380
rect 65356 5599 65396 5608
rect 65740 6152 65780 6161
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 64780 5144 64820 5153
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 64780 3464 64820 5104
rect 64780 3415 64820 3424
rect 65740 4976 65780 6112
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 61228 1819 61268 1828
rect 65740 1952 65780 4936
rect 66604 4220 66644 15940
rect 66700 10856 66740 17116
rect 68428 17156 68468 17165
rect 66796 17072 66836 17081
rect 66796 13124 66836 17032
rect 66796 13075 66836 13084
rect 67564 13376 67604 13385
rect 67564 12956 67604 13336
rect 67564 12907 67604 12916
rect 66700 10807 66740 10816
rect 68428 10100 68468 17116
rect 69100 16577 69140 17284
rect 71020 17324 71060 17333
rect 70156 17156 70196 17165
rect 69099 16568 69141 16577
rect 69099 16528 69100 16568
rect 69140 16528 69141 16568
rect 69099 16519 69141 16528
rect 70156 13796 70196 17116
rect 70923 16316 70965 16325
rect 70923 16276 70924 16316
rect 70964 16276 70965 16316
rect 70923 16267 70965 16276
rect 70828 16232 70868 16241
rect 70731 15476 70773 15485
rect 70731 15436 70732 15476
rect 70772 15436 70773 15476
rect 70731 15427 70773 15436
rect 70732 14804 70772 15427
rect 70732 14755 70772 14764
rect 70156 13747 70196 13756
rect 70828 13796 70868 16192
rect 70924 16182 70964 16267
rect 70828 13747 70868 13756
rect 71020 16148 71060 17284
rect 77164 17324 77204 17333
rect 74859 17240 74901 17249
rect 74859 17200 74860 17240
rect 74900 17200 74901 17240
rect 74859 17191 74901 17200
rect 76780 17240 76820 17249
rect 72556 17156 72596 17165
rect 71787 16400 71829 16409
rect 71787 16360 71788 16400
rect 71828 16360 71829 16400
rect 71787 16351 71829 16360
rect 71788 16266 71828 16351
rect 68428 10051 68468 10060
rect 68524 10352 68564 10361
rect 68524 9344 68564 10312
rect 71020 10100 71060 16108
rect 72556 14384 72596 17116
rect 74860 16148 74900 17191
rect 74860 16099 74900 16108
rect 75820 17156 75860 17165
rect 75532 15308 75572 15317
rect 75112 15140 75480 15149
rect 75152 15100 75194 15140
rect 75234 15100 75276 15140
rect 75316 15100 75358 15140
rect 75398 15100 75440 15140
rect 75112 15091 75480 15100
rect 72556 14335 72596 14344
rect 75112 13628 75480 13637
rect 75152 13588 75194 13628
rect 75234 13588 75276 13628
rect 75316 13588 75358 13628
rect 75398 13588 75440 13628
rect 75112 13579 75480 13588
rect 75112 12116 75480 12125
rect 75152 12076 75194 12116
rect 75234 12076 75276 12116
rect 75316 12076 75358 12116
rect 75398 12076 75440 12116
rect 75112 12067 75480 12076
rect 75112 10604 75480 10613
rect 75152 10564 75194 10604
rect 75234 10564 75276 10604
rect 75316 10564 75358 10604
rect 75398 10564 75440 10604
rect 75112 10555 75480 10564
rect 71020 10051 71060 10060
rect 68524 9295 68564 9304
rect 75112 9092 75480 9101
rect 75152 9052 75194 9092
rect 75234 9052 75276 9092
rect 75316 9052 75358 9092
rect 75398 9052 75440 9092
rect 75112 9043 75480 9052
rect 69004 8672 69044 8681
rect 69004 7580 69044 8632
rect 69004 5564 69044 7540
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 69004 5515 69044 5524
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 66604 4171 66644 4180
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 75532 2876 75572 15268
rect 75724 14048 75764 14057
rect 75724 12872 75764 14008
rect 75724 12823 75764 12832
rect 75820 10100 75860 17116
rect 76352 14384 76720 14393
rect 76392 14344 76434 14384
rect 76474 14344 76516 14384
rect 76556 14344 76598 14384
rect 76638 14344 76680 14384
rect 76352 14335 76720 14344
rect 76352 12872 76720 12881
rect 76392 12832 76434 12872
rect 76474 12832 76516 12872
rect 76556 12832 76598 12872
rect 76638 12832 76680 12872
rect 76352 12823 76720 12832
rect 76352 11360 76720 11369
rect 76392 11320 76434 11360
rect 76474 11320 76516 11360
rect 76556 11320 76598 11360
rect 76638 11320 76680 11360
rect 76352 11311 76720 11320
rect 75820 10051 75860 10060
rect 76352 9848 76720 9857
rect 76392 9808 76434 9848
rect 76474 9808 76516 9848
rect 76556 9808 76598 9848
rect 76638 9808 76680 9848
rect 76352 9799 76720 9808
rect 76352 8336 76720 8345
rect 76392 8296 76434 8336
rect 76474 8296 76516 8336
rect 76556 8296 76598 8336
rect 76638 8296 76680 8336
rect 76352 8287 76720 8296
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 76780 3296 76820 17200
rect 77068 15728 77108 15737
rect 76876 14384 76916 14393
rect 76876 5732 76916 14344
rect 76876 5683 76916 5692
rect 77068 3548 77108 15688
rect 77164 5648 77204 17284
rect 78507 16232 78549 16241
rect 78507 16192 78508 16232
rect 78548 16192 78549 16232
rect 78507 16183 78549 16192
rect 78508 16098 78548 16183
rect 77356 14048 77396 14057
rect 77356 12200 77396 14008
rect 77356 12151 77396 12160
rect 77164 5599 77204 5608
rect 77644 5900 77684 5909
rect 77644 4808 77684 5860
rect 77644 4759 77684 4768
rect 77068 3499 77108 3508
rect 76780 3247 76820 3256
rect 75532 2827 75572 2836
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 65740 1196 65780 1912
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 65740 1147 65780 1156
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 7372 27364 7412 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4588 21568 4628 21608
rect 5932 21568 5972 21608
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 39820 23668 39860 23708
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 38860 23248 38900 23288
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 3916 21400 3956 21440
rect 5932 21400 5972 21440
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 10924 20728 10964 20768
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 40300 25348 40340 25388
rect 49900 26860 49940 26900
rect 41068 25096 41108 25136
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 39916 19972 39956 20012
rect 40108 19972 40148 20012
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 7660 18544 7700 18584
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 7564 17536 7604 17576
rect 31756 17536 31796 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 34732 16948 34772 16988
rect 35308 16780 35348 16820
rect 33196 15352 33236 15392
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 45580 25264 45620 25304
rect 49132 25180 49172 25220
rect 48748 23752 48788 23792
rect 43468 23584 43508 23624
rect 41740 19468 41780 19508
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 41836 19384 41876 19424
rect 37996 16864 38036 16904
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 38284 16444 38324 16484
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 36748 14932 36788 14972
rect 41836 18544 41876 18584
rect 42412 17032 42452 17072
rect 42796 16108 42836 16148
rect 41164 16024 41204 16064
rect 40876 15772 40916 15812
rect 40780 14848 40820 14888
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 48940 15688 48980 15728
rect 47788 15604 47828 15644
rect 47884 15268 47924 15308
rect 49996 25348 50036 25388
rect 49900 14764 49940 14804
rect 50188 26944 50228 26984
rect 50092 14680 50132 14720
rect 49996 14176 50036 14216
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 50380 21484 50420 21524
rect 51628 24592 51668 24632
rect 51724 24508 51764 24548
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 51916 24760 51956 24800
rect 52108 24676 52148 24716
rect 51820 23920 51860 23960
rect 51820 22744 51860 22784
rect 51916 20728 51956 20768
rect 53068 23836 53108 23876
rect 55660 27364 55700 27404
rect 52588 23416 52628 23456
rect 53740 23416 53780 23456
rect 52204 23164 52244 23204
rect 52300 23080 52340 23120
rect 52396 22828 52436 22868
rect 52492 21568 52532 21608
rect 51916 19972 51956 20012
rect 51628 19468 51668 19508
rect 51820 17200 51860 17240
rect 51916 17116 51956 17156
rect 51148 15940 51188 15980
rect 50284 15520 50324 15560
rect 52684 23332 52724 23372
rect 53740 23248 53780 23288
rect 54892 24508 54932 24548
rect 54220 23164 54260 23204
rect 54508 23164 54548 23204
rect 52876 22996 52916 23036
rect 53452 22996 53492 23036
rect 53644 22996 53684 23036
rect 52972 22912 53012 22952
rect 52876 21568 52916 21608
rect 54700 22912 54740 22952
rect 53356 22744 53396 22784
rect 56140 24928 56180 24968
rect 55756 24676 55796 24716
rect 55564 23332 55604 23372
rect 55180 23248 55220 23288
rect 55084 23080 55124 23120
rect 56236 24172 56276 24212
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 61612 26944 61652 26984
rect 58444 26860 58484 26900
rect 58732 25348 58772 25388
rect 59116 25264 59156 25304
rect 57964 25096 58004 25136
rect 57580 24928 57620 24968
rect 57772 24592 57812 24632
rect 56620 24172 56660 24212
rect 57676 23668 57716 23708
rect 55852 23500 55892 23540
rect 56428 23500 56468 23540
rect 56236 23416 56276 23456
rect 57100 22828 57140 22868
rect 57868 23668 57908 23708
rect 58252 23668 58292 23708
rect 59020 23584 59060 23624
rect 61900 25180 61940 25220
rect 60460 23752 60500 23792
rect 60748 22996 60788 23036
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 64780 23920 64820 23960
rect 66508 23836 66548 23876
rect 66316 23500 66356 23540
rect 66220 23164 66260 23204
rect 66604 23668 66644 23708
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 75112 33244 75152 33284
rect 75194 33244 75234 33284
rect 75276 33244 75316 33284
rect 75358 33244 75398 33284
rect 75440 33244 75480 33284
rect 75112 31732 75152 31772
rect 75194 31732 75234 31772
rect 75276 31732 75316 31772
rect 75358 31732 75398 31772
rect 75440 31732 75480 31772
rect 75112 30220 75152 30260
rect 75194 30220 75234 30260
rect 75276 30220 75316 30260
rect 75358 30220 75398 30260
rect 75440 30220 75480 30260
rect 75112 28708 75152 28748
rect 75194 28708 75234 28748
rect 75276 28708 75316 28748
rect 75358 28708 75398 28748
rect 75440 28708 75480 28748
rect 75112 27196 75152 27236
rect 75194 27196 75234 27236
rect 75276 27196 75316 27236
rect 75358 27196 75398 27236
rect 75440 27196 75480 27236
rect 75112 25684 75152 25724
rect 75194 25684 75234 25724
rect 75276 25684 75316 25724
rect 75358 25684 75398 25724
rect 75440 25684 75480 25724
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 76352 32488 76392 32528
rect 76434 32488 76474 32528
rect 76516 32488 76556 32528
rect 76598 32488 76638 32528
rect 76680 32488 76720 32528
rect 76352 30976 76392 31016
rect 76434 30976 76474 31016
rect 76516 30976 76556 31016
rect 76598 30976 76638 31016
rect 76680 30976 76720 31016
rect 76352 29464 76392 29504
rect 76434 29464 76474 29504
rect 76516 29464 76556 29504
rect 76598 29464 76638 29504
rect 76680 29464 76720 29504
rect 76352 27952 76392 27992
rect 76434 27952 76474 27992
rect 76516 27952 76556 27992
rect 76598 27952 76638 27992
rect 76680 27952 76720 27992
rect 76352 26440 76392 26480
rect 76434 26440 76474 26480
rect 76516 26440 76556 26480
rect 76598 26440 76638 26480
rect 76680 26440 76720 26480
rect 76352 24928 76392 24968
rect 76434 24928 76474 24968
rect 76516 24928 76556 24968
rect 76598 24928 76638 24968
rect 76680 24928 76720 24968
rect 75148 23080 75188 23120
rect 71884 22744 71924 22784
rect 78988 24760 79028 24800
rect 78988 23752 79028 23792
rect 52300 19384 52340 19424
rect 56140 17116 56180 17156
rect 56332 17116 56372 17156
rect 54700 16864 54740 16904
rect 52204 15856 52244 15896
rect 52012 15772 52052 15812
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 53260 15688 53300 15728
rect 54604 15520 54644 15560
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56812 17200 56852 17240
rect 57292 16948 57332 16988
rect 57580 17032 57620 17072
rect 57388 16780 57428 16820
rect 56716 16444 56756 16484
rect 56428 15436 56468 15476
rect 57676 15352 57716 15392
rect 58060 14932 58100 14972
rect 59020 16108 59060 16148
rect 58924 16024 58964 16064
rect 58444 14848 58484 14888
rect 59116 14176 59156 14216
rect 59404 15604 59444 15644
rect 60460 16864 60500 16904
rect 59692 15268 59732 15308
rect 60364 14764 60404 14804
rect 60556 15688 60596 15728
rect 60748 16276 60788 16316
rect 60748 15772 60788 15812
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 63916 17116 63956 17156
rect 61996 15940 62036 15980
rect 61900 15856 61940 15896
rect 64108 15688 64148 15728
rect 61900 15436 61940 15476
rect 62284 15436 62324 15476
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 61900 14680 61940 14720
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 65356 16528 65396 16568
rect 65740 16528 65780 16568
rect 66220 16864 66260 16904
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 69100 16528 69140 16568
rect 70924 16276 70964 16316
rect 70732 15436 70772 15476
rect 74860 17200 74900 17240
rect 71788 16360 71828 16400
rect 75112 15100 75152 15140
rect 75194 15100 75234 15140
rect 75276 15100 75316 15140
rect 75358 15100 75398 15140
rect 75440 15100 75480 15140
rect 75112 13588 75152 13628
rect 75194 13588 75234 13628
rect 75276 13588 75316 13628
rect 75358 13588 75398 13628
rect 75440 13588 75480 13628
rect 75112 12076 75152 12116
rect 75194 12076 75234 12116
rect 75276 12076 75316 12116
rect 75358 12076 75398 12116
rect 75440 12076 75480 12116
rect 75112 10564 75152 10604
rect 75194 10564 75234 10604
rect 75276 10564 75316 10604
rect 75358 10564 75398 10604
rect 75440 10564 75480 10604
rect 75112 9052 75152 9092
rect 75194 9052 75234 9092
rect 75276 9052 75316 9092
rect 75358 9052 75398 9092
rect 75440 9052 75480 9092
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 76352 14344 76392 14384
rect 76434 14344 76474 14384
rect 76516 14344 76556 14384
rect 76598 14344 76638 14384
rect 76680 14344 76720 14384
rect 76352 12832 76392 12872
rect 76434 12832 76474 12872
rect 76516 12832 76556 12872
rect 76598 12832 76638 12872
rect 76680 12832 76720 12872
rect 76352 11320 76392 11360
rect 76434 11320 76474 11360
rect 76516 11320 76556 11360
rect 76598 11320 76638 11360
rect 76680 11320 76720 11360
rect 76352 9808 76392 9848
rect 76434 9808 76474 9848
rect 76516 9808 76556 9848
rect 76598 9808 76638 9848
rect 76680 9808 76720 9848
rect 76352 8296 76392 8336
rect 76434 8296 76474 8336
rect 76516 8296 76556 8336
rect 76598 8296 76638 8336
rect 76680 8296 76720 8336
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 78508 16192 78548 16232
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
<< metal5 >>
rect 4343 38576 4390 38618
rect 4514 38576 4558 38618
rect 4682 38576 4729 38618
rect 4343 38536 4352 38576
rect 4514 38536 4516 38576
rect 4556 38536 4558 38576
rect 4720 38536 4729 38576
rect 4343 38494 4390 38536
rect 4514 38494 4558 38536
rect 4682 38494 4729 38536
rect 16343 38576 16390 38618
rect 16514 38576 16558 38618
rect 16682 38576 16729 38618
rect 16343 38536 16352 38576
rect 16514 38536 16516 38576
rect 16556 38536 16558 38576
rect 16720 38536 16729 38576
rect 16343 38494 16390 38536
rect 16514 38494 16558 38536
rect 16682 38494 16729 38536
rect 28343 38576 28390 38618
rect 28514 38576 28558 38618
rect 28682 38576 28729 38618
rect 28343 38536 28352 38576
rect 28514 38536 28516 38576
rect 28556 38536 28558 38576
rect 28720 38536 28729 38576
rect 28343 38494 28390 38536
rect 28514 38494 28558 38536
rect 28682 38494 28729 38536
rect 40343 38576 40390 38618
rect 40514 38576 40558 38618
rect 40682 38576 40729 38618
rect 40343 38536 40352 38576
rect 40514 38536 40516 38576
rect 40556 38536 40558 38576
rect 40720 38536 40729 38576
rect 40343 38494 40390 38536
rect 40514 38494 40558 38536
rect 40682 38494 40729 38536
rect 52343 38576 52390 38618
rect 52514 38576 52558 38618
rect 52682 38576 52729 38618
rect 52343 38536 52352 38576
rect 52514 38536 52516 38576
rect 52556 38536 52558 38576
rect 52720 38536 52729 38576
rect 52343 38494 52390 38536
rect 52514 38494 52558 38536
rect 52682 38494 52729 38536
rect 64343 38576 64390 38618
rect 64514 38576 64558 38618
rect 64682 38576 64729 38618
rect 64343 38536 64352 38576
rect 64514 38536 64516 38576
rect 64556 38536 64558 38576
rect 64720 38536 64729 38576
rect 64343 38494 64390 38536
rect 64514 38494 64558 38536
rect 64682 38494 64729 38536
rect 76343 38576 76390 38618
rect 76514 38576 76558 38618
rect 76682 38576 76729 38618
rect 76343 38536 76352 38576
rect 76514 38536 76516 38576
rect 76556 38536 76558 38576
rect 76720 38536 76729 38576
rect 76343 38494 76390 38536
rect 76514 38494 76558 38536
rect 76682 38494 76729 38536
rect 3103 37820 3150 37862
rect 3274 37820 3318 37862
rect 3442 37820 3489 37862
rect 3103 37780 3112 37820
rect 3274 37780 3276 37820
rect 3316 37780 3318 37820
rect 3480 37780 3489 37820
rect 3103 37738 3150 37780
rect 3274 37738 3318 37780
rect 3442 37738 3489 37780
rect 15103 37820 15150 37862
rect 15274 37820 15318 37862
rect 15442 37820 15489 37862
rect 15103 37780 15112 37820
rect 15274 37780 15276 37820
rect 15316 37780 15318 37820
rect 15480 37780 15489 37820
rect 15103 37738 15150 37780
rect 15274 37738 15318 37780
rect 15442 37738 15489 37780
rect 27103 37820 27150 37862
rect 27274 37820 27318 37862
rect 27442 37820 27489 37862
rect 27103 37780 27112 37820
rect 27274 37780 27276 37820
rect 27316 37780 27318 37820
rect 27480 37780 27489 37820
rect 27103 37738 27150 37780
rect 27274 37738 27318 37780
rect 27442 37738 27489 37780
rect 39103 37820 39150 37862
rect 39274 37820 39318 37862
rect 39442 37820 39489 37862
rect 39103 37780 39112 37820
rect 39274 37780 39276 37820
rect 39316 37780 39318 37820
rect 39480 37780 39489 37820
rect 39103 37738 39150 37780
rect 39274 37738 39318 37780
rect 39442 37738 39489 37780
rect 51103 37820 51150 37862
rect 51274 37820 51318 37862
rect 51442 37820 51489 37862
rect 51103 37780 51112 37820
rect 51274 37780 51276 37820
rect 51316 37780 51318 37820
rect 51480 37780 51489 37820
rect 51103 37738 51150 37780
rect 51274 37738 51318 37780
rect 51442 37738 51489 37780
rect 63103 37820 63150 37862
rect 63274 37820 63318 37862
rect 63442 37820 63489 37862
rect 63103 37780 63112 37820
rect 63274 37780 63276 37820
rect 63316 37780 63318 37820
rect 63480 37780 63489 37820
rect 63103 37738 63150 37780
rect 63274 37738 63318 37780
rect 63442 37738 63489 37780
rect 75103 37820 75150 37862
rect 75274 37820 75318 37862
rect 75442 37820 75489 37862
rect 75103 37780 75112 37820
rect 75274 37780 75276 37820
rect 75316 37780 75318 37820
rect 75480 37780 75489 37820
rect 75103 37738 75150 37780
rect 75274 37738 75318 37780
rect 75442 37738 75489 37780
rect 4343 37064 4390 37106
rect 4514 37064 4558 37106
rect 4682 37064 4729 37106
rect 4343 37024 4352 37064
rect 4514 37024 4516 37064
rect 4556 37024 4558 37064
rect 4720 37024 4729 37064
rect 4343 36982 4390 37024
rect 4514 36982 4558 37024
rect 4682 36982 4729 37024
rect 16343 37064 16390 37106
rect 16514 37064 16558 37106
rect 16682 37064 16729 37106
rect 16343 37024 16352 37064
rect 16514 37024 16516 37064
rect 16556 37024 16558 37064
rect 16720 37024 16729 37064
rect 16343 36982 16390 37024
rect 16514 36982 16558 37024
rect 16682 36982 16729 37024
rect 28343 37064 28390 37106
rect 28514 37064 28558 37106
rect 28682 37064 28729 37106
rect 28343 37024 28352 37064
rect 28514 37024 28516 37064
rect 28556 37024 28558 37064
rect 28720 37024 28729 37064
rect 28343 36982 28390 37024
rect 28514 36982 28558 37024
rect 28682 36982 28729 37024
rect 40343 37064 40390 37106
rect 40514 37064 40558 37106
rect 40682 37064 40729 37106
rect 40343 37024 40352 37064
rect 40514 37024 40516 37064
rect 40556 37024 40558 37064
rect 40720 37024 40729 37064
rect 40343 36982 40390 37024
rect 40514 36982 40558 37024
rect 40682 36982 40729 37024
rect 52343 37064 52390 37106
rect 52514 37064 52558 37106
rect 52682 37064 52729 37106
rect 52343 37024 52352 37064
rect 52514 37024 52516 37064
rect 52556 37024 52558 37064
rect 52720 37024 52729 37064
rect 52343 36982 52390 37024
rect 52514 36982 52558 37024
rect 52682 36982 52729 37024
rect 64343 37064 64390 37106
rect 64514 37064 64558 37106
rect 64682 37064 64729 37106
rect 64343 37024 64352 37064
rect 64514 37024 64516 37064
rect 64556 37024 64558 37064
rect 64720 37024 64729 37064
rect 64343 36982 64390 37024
rect 64514 36982 64558 37024
rect 64682 36982 64729 37024
rect 76343 37064 76390 37106
rect 76514 37064 76558 37106
rect 76682 37064 76729 37106
rect 76343 37024 76352 37064
rect 76514 37024 76516 37064
rect 76556 37024 76558 37064
rect 76720 37024 76729 37064
rect 76343 36982 76390 37024
rect 76514 36982 76558 37024
rect 76682 36982 76729 37024
rect 3103 36308 3150 36350
rect 3274 36308 3318 36350
rect 3442 36308 3489 36350
rect 3103 36268 3112 36308
rect 3274 36268 3276 36308
rect 3316 36268 3318 36308
rect 3480 36268 3489 36308
rect 3103 36226 3150 36268
rect 3274 36226 3318 36268
rect 3442 36226 3489 36268
rect 15103 36308 15150 36350
rect 15274 36308 15318 36350
rect 15442 36308 15489 36350
rect 15103 36268 15112 36308
rect 15274 36268 15276 36308
rect 15316 36268 15318 36308
rect 15480 36268 15489 36308
rect 15103 36226 15150 36268
rect 15274 36226 15318 36268
rect 15442 36226 15489 36268
rect 27103 36308 27150 36350
rect 27274 36308 27318 36350
rect 27442 36308 27489 36350
rect 27103 36268 27112 36308
rect 27274 36268 27276 36308
rect 27316 36268 27318 36308
rect 27480 36268 27489 36308
rect 27103 36226 27150 36268
rect 27274 36226 27318 36268
rect 27442 36226 27489 36268
rect 39103 36308 39150 36350
rect 39274 36308 39318 36350
rect 39442 36308 39489 36350
rect 39103 36268 39112 36308
rect 39274 36268 39276 36308
rect 39316 36268 39318 36308
rect 39480 36268 39489 36308
rect 39103 36226 39150 36268
rect 39274 36226 39318 36268
rect 39442 36226 39489 36268
rect 51103 36308 51150 36350
rect 51274 36308 51318 36350
rect 51442 36308 51489 36350
rect 51103 36268 51112 36308
rect 51274 36268 51276 36308
rect 51316 36268 51318 36308
rect 51480 36268 51489 36308
rect 51103 36226 51150 36268
rect 51274 36226 51318 36268
rect 51442 36226 51489 36268
rect 63103 36308 63150 36350
rect 63274 36308 63318 36350
rect 63442 36308 63489 36350
rect 63103 36268 63112 36308
rect 63274 36268 63276 36308
rect 63316 36268 63318 36308
rect 63480 36268 63489 36308
rect 63103 36226 63150 36268
rect 63274 36226 63318 36268
rect 63442 36226 63489 36268
rect 75103 36308 75150 36350
rect 75274 36308 75318 36350
rect 75442 36308 75489 36350
rect 75103 36268 75112 36308
rect 75274 36268 75276 36308
rect 75316 36268 75318 36308
rect 75480 36268 75489 36308
rect 75103 36226 75150 36268
rect 75274 36226 75318 36268
rect 75442 36226 75489 36268
rect 4343 35552 4390 35594
rect 4514 35552 4558 35594
rect 4682 35552 4729 35594
rect 4343 35512 4352 35552
rect 4514 35512 4516 35552
rect 4556 35512 4558 35552
rect 4720 35512 4729 35552
rect 4343 35470 4390 35512
rect 4514 35470 4558 35512
rect 4682 35470 4729 35512
rect 16343 35552 16390 35594
rect 16514 35552 16558 35594
rect 16682 35552 16729 35594
rect 16343 35512 16352 35552
rect 16514 35512 16516 35552
rect 16556 35512 16558 35552
rect 16720 35512 16729 35552
rect 16343 35470 16390 35512
rect 16514 35470 16558 35512
rect 16682 35470 16729 35512
rect 28343 35552 28390 35594
rect 28514 35552 28558 35594
rect 28682 35552 28729 35594
rect 28343 35512 28352 35552
rect 28514 35512 28516 35552
rect 28556 35512 28558 35552
rect 28720 35512 28729 35552
rect 28343 35470 28390 35512
rect 28514 35470 28558 35512
rect 28682 35470 28729 35512
rect 40343 35552 40390 35594
rect 40514 35552 40558 35594
rect 40682 35552 40729 35594
rect 40343 35512 40352 35552
rect 40514 35512 40516 35552
rect 40556 35512 40558 35552
rect 40720 35512 40729 35552
rect 40343 35470 40390 35512
rect 40514 35470 40558 35512
rect 40682 35470 40729 35512
rect 52343 35552 52390 35594
rect 52514 35552 52558 35594
rect 52682 35552 52729 35594
rect 52343 35512 52352 35552
rect 52514 35512 52516 35552
rect 52556 35512 52558 35552
rect 52720 35512 52729 35552
rect 52343 35470 52390 35512
rect 52514 35470 52558 35512
rect 52682 35470 52729 35512
rect 64343 35552 64390 35594
rect 64514 35552 64558 35594
rect 64682 35552 64729 35594
rect 64343 35512 64352 35552
rect 64514 35512 64516 35552
rect 64556 35512 64558 35552
rect 64720 35512 64729 35552
rect 64343 35470 64390 35512
rect 64514 35470 64558 35512
rect 64682 35470 64729 35512
rect 76343 35552 76390 35594
rect 76514 35552 76558 35594
rect 76682 35552 76729 35594
rect 76343 35512 76352 35552
rect 76514 35512 76516 35552
rect 76556 35512 76558 35552
rect 76720 35512 76729 35552
rect 76343 35470 76390 35512
rect 76514 35470 76558 35512
rect 76682 35470 76729 35512
rect 3103 34796 3150 34838
rect 3274 34796 3318 34838
rect 3442 34796 3489 34838
rect 3103 34756 3112 34796
rect 3274 34756 3276 34796
rect 3316 34756 3318 34796
rect 3480 34756 3489 34796
rect 3103 34714 3150 34756
rect 3274 34714 3318 34756
rect 3442 34714 3489 34756
rect 15103 34796 15150 34838
rect 15274 34796 15318 34838
rect 15442 34796 15489 34838
rect 15103 34756 15112 34796
rect 15274 34756 15276 34796
rect 15316 34756 15318 34796
rect 15480 34756 15489 34796
rect 15103 34714 15150 34756
rect 15274 34714 15318 34756
rect 15442 34714 15489 34756
rect 27103 34796 27150 34838
rect 27274 34796 27318 34838
rect 27442 34796 27489 34838
rect 27103 34756 27112 34796
rect 27274 34756 27276 34796
rect 27316 34756 27318 34796
rect 27480 34756 27489 34796
rect 27103 34714 27150 34756
rect 27274 34714 27318 34756
rect 27442 34714 27489 34756
rect 39103 34796 39150 34838
rect 39274 34796 39318 34838
rect 39442 34796 39489 34838
rect 39103 34756 39112 34796
rect 39274 34756 39276 34796
rect 39316 34756 39318 34796
rect 39480 34756 39489 34796
rect 39103 34714 39150 34756
rect 39274 34714 39318 34756
rect 39442 34714 39489 34756
rect 51103 34796 51150 34838
rect 51274 34796 51318 34838
rect 51442 34796 51489 34838
rect 51103 34756 51112 34796
rect 51274 34756 51276 34796
rect 51316 34756 51318 34796
rect 51480 34756 51489 34796
rect 51103 34714 51150 34756
rect 51274 34714 51318 34756
rect 51442 34714 51489 34756
rect 63103 34796 63150 34838
rect 63274 34796 63318 34838
rect 63442 34796 63489 34838
rect 63103 34756 63112 34796
rect 63274 34756 63276 34796
rect 63316 34756 63318 34796
rect 63480 34756 63489 34796
rect 63103 34714 63150 34756
rect 63274 34714 63318 34756
rect 63442 34714 63489 34756
rect 75103 34796 75150 34838
rect 75274 34796 75318 34838
rect 75442 34796 75489 34838
rect 75103 34756 75112 34796
rect 75274 34756 75276 34796
rect 75316 34756 75318 34796
rect 75480 34756 75489 34796
rect 75103 34714 75150 34756
rect 75274 34714 75318 34756
rect 75442 34714 75489 34756
rect 4343 34040 4390 34082
rect 4514 34040 4558 34082
rect 4682 34040 4729 34082
rect 4343 34000 4352 34040
rect 4514 34000 4516 34040
rect 4556 34000 4558 34040
rect 4720 34000 4729 34040
rect 4343 33958 4390 34000
rect 4514 33958 4558 34000
rect 4682 33958 4729 34000
rect 16343 34040 16390 34082
rect 16514 34040 16558 34082
rect 16682 34040 16729 34082
rect 16343 34000 16352 34040
rect 16514 34000 16516 34040
rect 16556 34000 16558 34040
rect 16720 34000 16729 34040
rect 16343 33958 16390 34000
rect 16514 33958 16558 34000
rect 16682 33958 16729 34000
rect 28343 34040 28390 34082
rect 28514 34040 28558 34082
rect 28682 34040 28729 34082
rect 28343 34000 28352 34040
rect 28514 34000 28516 34040
rect 28556 34000 28558 34040
rect 28720 34000 28729 34040
rect 28343 33958 28390 34000
rect 28514 33958 28558 34000
rect 28682 33958 28729 34000
rect 40343 34040 40390 34082
rect 40514 34040 40558 34082
rect 40682 34040 40729 34082
rect 40343 34000 40352 34040
rect 40514 34000 40516 34040
rect 40556 34000 40558 34040
rect 40720 34000 40729 34040
rect 40343 33958 40390 34000
rect 40514 33958 40558 34000
rect 40682 33958 40729 34000
rect 52343 34040 52390 34082
rect 52514 34040 52558 34082
rect 52682 34040 52729 34082
rect 52343 34000 52352 34040
rect 52514 34000 52516 34040
rect 52556 34000 52558 34040
rect 52720 34000 52729 34040
rect 52343 33958 52390 34000
rect 52514 33958 52558 34000
rect 52682 33958 52729 34000
rect 64343 34040 64390 34082
rect 64514 34040 64558 34082
rect 64682 34040 64729 34082
rect 64343 34000 64352 34040
rect 64514 34000 64516 34040
rect 64556 34000 64558 34040
rect 64720 34000 64729 34040
rect 64343 33958 64390 34000
rect 64514 33958 64558 34000
rect 64682 33958 64729 34000
rect 76343 34040 76390 34082
rect 76514 34040 76558 34082
rect 76682 34040 76729 34082
rect 76343 34000 76352 34040
rect 76514 34000 76516 34040
rect 76556 34000 76558 34040
rect 76720 34000 76729 34040
rect 76343 33958 76390 34000
rect 76514 33958 76558 34000
rect 76682 33958 76729 34000
rect 3103 33284 3150 33326
rect 3274 33284 3318 33326
rect 3442 33284 3489 33326
rect 3103 33244 3112 33284
rect 3274 33244 3276 33284
rect 3316 33244 3318 33284
rect 3480 33244 3489 33284
rect 3103 33202 3150 33244
rect 3274 33202 3318 33244
rect 3442 33202 3489 33244
rect 15103 33284 15150 33326
rect 15274 33284 15318 33326
rect 15442 33284 15489 33326
rect 15103 33244 15112 33284
rect 15274 33244 15276 33284
rect 15316 33244 15318 33284
rect 15480 33244 15489 33284
rect 15103 33202 15150 33244
rect 15274 33202 15318 33244
rect 15442 33202 15489 33244
rect 27103 33284 27150 33326
rect 27274 33284 27318 33326
rect 27442 33284 27489 33326
rect 27103 33244 27112 33284
rect 27274 33244 27276 33284
rect 27316 33244 27318 33284
rect 27480 33244 27489 33284
rect 27103 33202 27150 33244
rect 27274 33202 27318 33244
rect 27442 33202 27489 33244
rect 39103 33284 39150 33326
rect 39274 33284 39318 33326
rect 39442 33284 39489 33326
rect 39103 33244 39112 33284
rect 39274 33244 39276 33284
rect 39316 33244 39318 33284
rect 39480 33244 39489 33284
rect 39103 33202 39150 33244
rect 39274 33202 39318 33244
rect 39442 33202 39489 33244
rect 51103 33284 51150 33326
rect 51274 33284 51318 33326
rect 51442 33284 51489 33326
rect 51103 33244 51112 33284
rect 51274 33244 51276 33284
rect 51316 33244 51318 33284
rect 51480 33244 51489 33284
rect 51103 33202 51150 33244
rect 51274 33202 51318 33244
rect 51442 33202 51489 33244
rect 63103 33284 63150 33326
rect 63274 33284 63318 33326
rect 63442 33284 63489 33326
rect 63103 33244 63112 33284
rect 63274 33244 63276 33284
rect 63316 33244 63318 33284
rect 63480 33244 63489 33284
rect 63103 33202 63150 33244
rect 63274 33202 63318 33244
rect 63442 33202 63489 33244
rect 75103 33284 75150 33326
rect 75274 33284 75318 33326
rect 75442 33284 75489 33326
rect 75103 33244 75112 33284
rect 75274 33244 75276 33284
rect 75316 33244 75318 33284
rect 75480 33244 75489 33284
rect 75103 33202 75150 33244
rect 75274 33202 75318 33244
rect 75442 33202 75489 33244
rect 4343 32528 4390 32570
rect 4514 32528 4558 32570
rect 4682 32528 4729 32570
rect 4343 32488 4352 32528
rect 4514 32488 4516 32528
rect 4556 32488 4558 32528
rect 4720 32488 4729 32528
rect 4343 32446 4390 32488
rect 4514 32446 4558 32488
rect 4682 32446 4729 32488
rect 16343 32528 16390 32570
rect 16514 32528 16558 32570
rect 16682 32528 16729 32570
rect 16343 32488 16352 32528
rect 16514 32488 16516 32528
rect 16556 32488 16558 32528
rect 16720 32488 16729 32528
rect 16343 32446 16390 32488
rect 16514 32446 16558 32488
rect 16682 32446 16729 32488
rect 28343 32528 28390 32570
rect 28514 32528 28558 32570
rect 28682 32528 28729 32570
rect 28343 32488 28352 32528
rect 28514 32488 28516 32528
rect 28556 32488 28558 32528
rect 28720 32488 28729 32528
rect 28343 32446 28390 32488
rect 28514 32446 28558 32488
rect 28682 32446 28729 32488
rect 40343 32528 40390 32570
rect 40514 32528 40558 32570
rect 40682 32528 40729 32570
rect 40343 32488 40352 32528
rect 40514 32488 40516 32528
rect 40556 32488 40558 32528
rect 40720 32488 40729 32528
rect 40343 32446 40390 32488
rect 40514 32446 40558 32488
rect 40682 32446 40729 32488
rect 52343 32528 52390 32570
rect 52514 32528 52558 32570
rect 52682 32528 52729 32570
rect 52343 32488 52352 32528
rect 52514 32488 52516 32528
rect 52556 32488 52558 32528
rect 52720 32488 52729 32528
rect 52343 32446 52390 32488
rect 52514 32446 52558 32488
rect 52682 32446 52729 32488
rect 64343 32528 64390 32570
rect 64514 32528 64558 32570
rect 64682 32528 64729 32570
rect 64343 32488 64352 32528
rect 64514 32488 64516 32528
rect 64556 32488 64558 32528
rect 64720 32488 64729 32528
rect 64343 32446 64390 32488
rect 64514 32446 64558 32488
rect 64682 32446 64729 32488
rect 76343 32528 76390 32570
rect 76514 32528 76558 32570
rect 76682 32528 76729 32570
rect 76343 32488 76352 32528
rect 76514 32488 76516 32528
rect 76556 32488 76558 32528
rect 76720 32488 76729 32528
rect 76343 32446 76390 32488
rect 76514 32446 76558 32488
rect 76682 32446 76729 32488
rect 3103 31772 3150 31814
rect 3274 31772 3318 31814
rect 3442 31772 3489 31814
rect 3103 31732 3112 31772
rect 3274 31732 3276 31772
rect 3316 31732 3318 31772
rect 3480 31732 3489 31772
rect 3103 31690 3150 31732
rect 3274 31690 3318 31732
rect 3442 31690 3489 31732
rect 15103 31772 15150 31814
rect 15274 31772 15318 31814
rect 15442 31772 15489 31814
rect 15103 31732 15112 31772
rect 15274 31732 15276 31772
rect 15316 31732 15318 31772
rect 15480 31732 15489 31772
rect 15103 31690 15150 31732
rect 15274 31690 15318 31732
rect 15442 31690 15489 31732
rect 27103 31772 27150 31814
rect 27274 31772 27318 31814
rect 27442 31772 27489 31814
rect 27103 31732 27112 31772
rect 27274 31732 27276 31772
rect 27316 31732 27318 31772
rect 27480 31732 27489 31772
rect 27103 31690 27150 31732
rect 27274 31690 27318 31732
rect 27442 31690 27489 31732
rect 39103 31772 39150 31814
rect 39274 31772 39318 31814
rect 39442 31772 39489 31814
rect 39103 31732 39112 31772
rect 39274 31732 39276 31772
rect 39316 31732 39318 31772
rect 39480 31732 39489 31772
rect 39103 31690 39150 31732
rect 39274 31690 39318 31732
rect 39442 31690 39489 31732
rect 51103 31772 51150 31814
rect 51274 31772 51318 31814
rect 51442 31772 51489 31814
rect 51103 31732 51112 31772
rect 51274 31732 51276 31772
rect 51316 31732 51318 31772
rect 51480 31732 51489 31772
rect 51103 31690 51150 31732
rect 51274 31690 51318 31732
rect 51442 31690 51489 31732
rect 63103 31772 63150 31814
rect 63274 31772 63318 31814
rect 63442 31772 63489 31814
rect 63103 31732 63112 31772
rect 63274 31732 63276 31772
rect 63316 31732 63318 31772
rect 63480 31732 63489 31772
rect 63103 31690 63150 31732
rect 63274 31690 63318 31732
rect 63442 31690 63489 31732
rect 75103 31772 75150 31814
rect 75274 31772 75318 31814
rect 75442 31772 75489 31814
rect 75103 31732 75112 31772
rect 75274 31732 75276 31772
rect 75316 31732 75318 31772
rect 75480 31732 75489 31772
rect 75103 31690 75150 31732
rect 75274 31690 75318 31732
rect 75442 31690 75489 31732
rect 4343 31016 4390 31058
rect 4514 31016 4558 31058
rect 4682 31016 4729 31058
rect 4343 30976 4352 31016
rect 4514 30976 4516 31016
rect 4556 30976 4558 31016
rect 4720 30976 4729 31016
rect 4343 30934 4390 30976
rect 4514 30934 4558 30976
rect 4682 30934 4729 30976
rect 16343 31016 16390 31058
rect 16514 31016 16558 31058
rect 16682 31016 16729 31058
rect 16343 30976 16352 31016
rect 16514 30976 16516 31016
rect 16556 30976 16558 31016
rect 16720 30976 16729 31016
rect 16343 30934 16390 30976
rect 16514 30934 16558 30976
rect 16682 30934 16729 30976
rect 28343 31016 28390 31058
rect 28514 31016 28558 31058
rect 28682 31016 28729 31058
rect 28343 30976 28352 31016
rect 28514 30976 28516 31016
rect 28556 30976 28558 31016
rect 28720 30976 28729 31016
rect 28343 30934 28390 30976
rect 28514 30934 28558 30976
rect 28682 30934 28729 30976
rect 40343 31016 40390 31058
rect 40514 31016 40558 31058
rect 40682 31016 40729 31058
rect 40343 30976 40352 31016
rect 40514 30976 40516 31016
rect 40556 30976 40558 31016
rect 40720 30976 40729 31016
rect 40343 30934 40390 30976
rect 40514 30934 40558 30976
rect 40682 30934 40729 30976
rect 52343 31016 52390 31058
rect 52514 31016 52558 31058
rect 52682 31016 52729 31058
rect 52343 30976 52352 31016
rect 52514 30976 52516 31016
rect 52556 30976 52558 31016
rect 52720 30976 52729 31016
rect 52343 30934 52390 30976
rect 52514 30934 52558 30976
rect 52682 30934 52729 30976
rect 64343 31016 64390 31058
rect 64514 31016 64558 31058
rect 64682 31016 64729 31058
rect 64343 30976 64352 31016
rect 64514 30976 64516 31016
rect 64556 30976 64558 31016
rect 64720 30976 64729 31016
rect 64343 30934 64390 30976
rect 64514 30934 64558 30976
rect 64682 30934 64729 30976
rect 76343 31016 76390 31058
rect 76514 31016 76558 31058
rect 76682 31016 76729 31058
rect 76343 30976 76352 31016
rect 76514 30976 76516 31016
rect 76556 30976 76558 31016
rect 76720 30976 76729 31016
rect 76343 30934 76390 30976
rect 76514 30934 76558 30976
rect 76682 30934 76729 30976
rect 3103 30260 3150 30302
rect 3274 30260 3318 30302
rect 3442 30260 3489 30302
rect 3103 30220 3112 30260
rect 3274 30220 3276 30260
rect 3316 30220 3318 30260
rect 3480 30220 3489 30260
rect 3103 30178 3150 30220
rect 3274 30178 3318 30220
rect 3442 30178 3489 30220
rect 15103 30260 15150 30302
rect 15274 30260 15318 30302
rect 15442 30260 15489 30302
rect 15103 30220 15112 30260
rect 15274 30220 15276 30260
rect 15316 30220 15318 30260
rect 15480 30220 15489 30260
rect 15103 30178 15150 30220
rect 15274 30178 15318 30220
rect 15442 30178 15489 30220
rect 27103 30260 27150 30302
rect 27274 30260 27318 30302
rect 27442 30260 27489 30302
rect 27103 30220 27112 30260
rect 27274 30220 27276 30260
rect 27316 30220 27318 30260
rect 27480 30220 27489 30260
rect 27103 30178 27150 30220
rect 27274 30178 27318 30220
rect 27442 30178 27489 30220
rect 39103 30260 39150 30302
rect 39274 30260 39318 30302
rect 39442 30260 39489 30302
rect 39103 30220 39112 30260
rect 39274 30220 39276 30260
rect 39316 30220 39318 30260
rect 39480 30220 39489 30260
rect 39103 30178 39150 30220
rect 39274 30178 39318 30220
rect 39442 30178 39489 30220
rect 51103 30260 51150 30302
rect 51274 30260 51318 30302
rect 51442 30260 51489 30302
rect 51103 30220 51112 30260
rect 51274 30220 51276 30260
rect 51316 30220 51318 30260
rect 51480 30220 51489 30260
rect 51103 30178 51150 30220
rect 51274 30178 51318 30220
rect 51442 30178 51489 30220
rect 63103 30260 63150 30302
rect 63274 30260 63318 30302
rect 63442 30260 63489 30302
rect 63103 30220 63112 30260
rect 63274 30220 63276 30260
rect 63316 30220 63318 30260
rect 63480 30220 63489 30260
rect 63103 30178 63150 30220
rect 63274 30178 63318 30220
rect 63442 30178 63489 30220
rect 75103 30260 75150 30302
rect 75274 30260 75318 30302
rect 75442 30260 75489 30302
rect 75103 30220 75112 30260
rect 75274 30220 75276 30260
rect 75316 30220 75318 30260
rect 75480 30220 75489 30260
rect 75103 30178 75150 30220
rect 75274 30178 75318 30220
rect 75442 30178 75489 30220
rect 4343 29504 4390 29546
rect 4514 29504 4558 29546
rect 4682 29504 4729 29546
rect 4343 29464 4352 29504
rect 4514 29464 4516 29504
rect 4556 29464 4558 29504
rect 4720 29464 4729 29504
rect 4343 29422 4390 29464
rect 4514 29422 4558 29464
rect 4682 29422 4729 29464
rect 16343 29504 16390 29546
rect 16514 29504 16558 29546
rect 16682 29504 16729 29546
rect 16343 29464 16352 29504
rect 16514 29464 16516 29504
rect 16556 29464 16558 29504
rect 16720 29464 16729 29504
rect 16343 29422 16390 29464
rect 16514 29422 16558 29464
rect 16682 29422 16729 29464
rect 28343 29504 28390 29546
rect 28514 29504 28558 29546
rect 28682 29504 28729 29546
rect 28343 29464 28352 29504
rect 28514 29464 28516 29504
rect 28556 29464 28558 29504
rect 28720 29464 28729 29504
rect 28343 29422 28390 29464
rect 28514 29422 28558 29464
rect 28682 29422 28729 29464
rect 40343 29504 40390 29546
rect 40514 29504 40558 29546
rect 40682 29504 40729 29546
rect 40343 29464 40352 29504
rect 40514 29464 40516 29504
rect 40556 29464 40558 29504
rect 40720 29464 40729 29504
rect 40343 29422 40390 29464
rect 40514 29422 40558 29464
rect 40682 29422 40729 29464
rect 52343 29504 52390 29546
rect 52514 29504 52558 29546
rect 52682 29504 52729 29546
rect 52343 29464 52352 29504
rect 52514 29464 52516 29504
rect 52556 29464 52558 29504
rect 52720 29464 52729 29504
rect 52343 29422 52390 29464
rect 52514 29422 52558 29464
rect 52682 29422 52729 29464
rect 64343 29504 64390 29546
rect 64514 29504 64558 29546
rect 64682 29504 64729 29546
rect 64343 29464 64352 29504
rect 64514 29464 64516 29504
rect 64556 29464 64558 29504
rect 64720 29464 64729 29504
rect 64343 29422 64390 29464
rect 64514 29422 64558 29464
rect 64682 29422 64729 29464
rect 76343 29504 76390 29546
rect 76514 29504 76558 29546
rect 76682 29504 76729 29546
rect 76343 29464 76352 29504
rect 76514 29464 76516 29504
rect 76556 29464 76558 29504
rect 76720 29464 76729 29504
rect 76343 29422 76390 29464
rect 76514 29422 76558 29464
rect 76682 29422 76729 29464
rect 3103 28748 3150 28790
rect 3274 28748 3318 28790
rect 3442 28748 3489 28790
rect 3103 28708 3112 28748
rect 3274 28708 3276 28748
rect 3316 28708 3318 28748
rect 3480 28708 3489 28748
rect 3103 28666 3150 28708
rect 3274 28666 3318 28708
rect 3442 28666 3489 28708
rect 15103 28748 15150 28790
rect 15274 28748 15318 28790
rect 15442 28748 15489 28790
rect 15103 28708 15112 28748
rect 15274 28708 15276 28748
rect 15316 28708 15318 28748
rect 15480 28708 15489 28748
rect 15103 28666 15150 28708
rect 15274 28666 15318 28708
rect 15442 28666 15489 28708
rect 27103 28748 27150 28790
rect 27274 28748 27318 28790
rect 27442 28748 27489 28790
rect 27103 28708 27112 28748
rect 27274 28708 27276 28748
rect 27316 28708 27318 28748
rect 27480 28708 27489 28748
rect 27103 28666 27150 28708
rect 27274 28666 27318 28708
rect 27442 28666 27489 28708
rect 39103 28748 39150 28790
rect 39274 28748 39318 28790
rect 39442 28748 39489 28790
rect 39103 28708 39112 28748
rect 39274 28708 39276 28748
rect 39316 28708 39318 28748
rect 39480 28708 39489 28748
rect 39103 28666 39150 28708
rect 39274 28666 39318 28708
rect 39442 28666 39489 28708
rect 51103 28748 51150 28790
rect 51274 28748 51318 28790
rect 51442 28748 51489 28790
rect 51103 28708 51112 28748
rect 51274 28708 51276 28748
rect 51316 28708 51318 28748
rect 51480 28708 51489 28748
rect 51103 28666 51150 28708
rect 51274 28666 51318 28708
rect 51442 28666 51489 28708
rect 63103 28748 63150 28790
rect 63274 28748 63318 28790
rect 63442 28748 63489 28790
rect 63103 28708 63112 28748
rect 63274 28708 63276 28748
rect 63316 28708 63318 28748
rect 63480 28708 63489 28748
rect 63103 28666 63150 28708
rect 63274 28666 63318 28708
rect 63442 28666 63489 28708
rect 75103 28748 75150 28790
rect 75274 28748 75318 28790
rect 75442 28748 75489 28790
rect 75103 28708 75112 28748
rect 75274 28708 75276 28748
rect 75316 28708 75318 28748
rect 75480 28708 75489 28748
rect 75103 28666 75150 28708
rect 75274 28666 75318 28708
rect 75442 28666 75489 28708
rect 4343 27992 4390 28034
rect 4514 27992 4558 28034
rect 4682 27992 4729 28034
rect 4343 27952 4352 27992
rect 4514 27952 4516 27992
rect 4556 27952 4558 27992
rect 4720 27952 4729 27992
rect 4343 27910 4390 27952
rect 4514 27910 4558 27952
rect 4682 27910 4729 27952
rect 16343 27992 16390 28034
rect 16514 27992 16558 28034
rect 16682 27992 16729 28034
rect 16343 27952 16352 27992
rect 16514 27952 16516 27992
rect 16556 27952 16558 27992
rect 16720 27952 16729 27992
rect 16343 27910 16390 27952
rect 16514 27910 16558 27952
rect 16682 27910 16729 27952
rect 28343 27992 28390 28034
rect 28514 27992 28558 28034
rect 28682 27992 28729 28034
rect 28343 27952 28352 27992
rect 28514 27952 28516 27992
rect 28556 27952 28558 27992
rect 28720 27952 28729 27992
rect 28343 27910 28390 27952
rect 28514 27910 28558 27952
rect 28682 27910 28729 27952
rect 40343 27992 40390 28034
rect 40514 27992 40558 28034
rect 40682 27992 40729 28034
rect 40343 27952 40352 27992
rect 40514 27952 40516 27992
rect 40556 27952 40558 27992
rect 40720 27952 40729 27992
rect 40343 27910 40390 27952
rect 40514 27910 40558 27952
rect 40682 27910 40729 27952
rect 52343 27992 52390 28034
rect 52514 27992 52558 28034
rect 52682 27992 52729 28034
rect 52343 27952 52352 27992
rect 52514 27952 52516 27992
rect 52556 27952 52558 27992
rect 52720 27952 52729 27992
rect 52343 27910 52390 27952
rect 52514 27910 52558 27952
rect 52682 27910 52729 27952
rect 64343 27992 64390 28034
rect 64514 27992 64558 28034
rect 64682 27992 64729 28034
rect 64343 27952 64352 27992
rect 64514 27952 64516 27992
rect 64556 27952 64558 27992
rect 64720 27952 64729 27992
rect 64343 27910 64390 27952
rect 64514 27910 64558 27952
rect 64682 27910 64729 27952
rect 76343 27992 76390 28034
rect 76514 27992 76558 28034
rect 76682 27992 76729 28034
rect 76343 27952 76352 27992
rect 76514 27952 76516 27992
rect 76556 27952 76558 27992
rect 76720 27952 76729 27992
rect 76343 27910 76390 27952
rect 76514 27910 76558 27952
rect 76682 27910 76729 27952
rect 7363 27364 7372 27404
rect 7412 27364 55660 27404
rect 55700 27364 55709 27404
rect 3103 27236 3150 27278
rect 3274 27236 3318 27278
rect 3442 27236 3489 27278
rect 3103 27196 3112 27236
rect 3274 27196 3276 27236
rect 3316 27196 3318 27236
rect 3480 27196 3489 27236
rect 3103 27154 3150 27196
rect 3274 27154 3318 27196
rect 3442 27154 3489 27196
rect 15103 27236 15150 27278
rect 15274 27236 15318 27278
rect 15442 27236 15489 27278
rect 15103 27196 15112 27236
rect 15274 27196 15276 27236
rect 15316 27196 15318 27236
rect 15480 27196 15489 27236
rect 15103 27154 15150 27196
rect 15274 27154 15318 27196
rect 15442 27154 15489 27196
rect 27103 27236 27150 27278
rect 27274 27236 27318 27278
rect 27442 27236 27489 27278
rect 27103 27196 27112 27236
rect 27274 27196 27276 27236
rect 27316 27196 27318 27236
rect 27480 27196 27489 27236
rect 27103 27154 27150 27196
rect 27274 27154 27318 27196
rect 27442 27154 27489 27196
rect 39103 27236 39150 27278
rect 39274 27236 39318 27278
rect 39442 27236 39489 27278
rect 39103 27196 39112 27236
rect 39274 27196 39276 27236
rect 39316 27196 39318 27236
rect 39480 27196 39489 27236
rect 39103 27154 39150 27196
rect 39274 27154 39318 27196
rect 39442 27154 39489 27196
rect 51103 27236 51150 27278
rect 51274 27236 51318 27278
rect 51442 27236 51489 27278
rect 51103 27196 51112 27236
rect 51274 27196 51276 27236
rect 51316 27196 51318 27236
rect 51480 27196 51489 27236
rect 51103 27154 51150 27196
rect 51274 27154 51318 27196
rect 51442 27154 51489 27196
rect 63103 27236 63150 27278
rect 63274 27236 63318 27278
rect 63442 27236 63489 27278
rect 63103 27196 63112 27236
rect 63274 27196 63276 27236
rect 63316 27196 63318 27236
rect 63480 27196 63489 27236
rect 63103 27154 63150 27196
rect 63274 27154 63318 27196
rect 63442 27154 63489 27196
rect 75103 27236 75150 27278
rect 75274 27236 75318 27278
rect 75442 27236 75489 27278
rect 75103 27196 75112 27236
rect 75274 27196 75276 27236
rect 75316 27196 75318 27236
rect 75480 27196 75489 27236
rect 75103 27154 75150 27196
rect 75274 27154 75318 27196
rect 75442 27154 75489 27196
rect 50179 26944 50188 26984
rect 50228 26944 61612 26984
rect 61652 26944 61661 26984
rect 49891 26860 49900 26900
rect 49940 26860 58444 26900
rect 58484 26860 58493 26900
rect 4343 26480 4390 26522
rect 4514 26480 4558 26522
rect 4682 26480 4729 26522
rect 4343 26440 4352 26480
rect 4514 26440 4516 26480
rect 4556 26440 4558 26480
rect 4720 26440 4729 26480
rect 4343 26398 4390 26440
rect 4514 26398 4558 26440
rect 4682 26398 4729 26440
rect 16343 26480 16390 26522
rect 16514 26480 16558 26522
rect 16682 26480 16729 26522
rect 16343 26440 16352 26480
rect 16514 26440 16516 26480
rect 16556 26440 16558 26480
rect 16720 26440 16729 26480
rect 16343 26398 16390 26440
rect 16514 26398 16558 26440
rect 16682 26398 16729 26440
rect 28343 26480 28390 26522
rect 28514 26480 28558 26522
rect 28682 26480 28729 26522
rect 28343 26440 28352 26480
rect 28514 26440 28516 26480
rect 28556 26440 28558 26480
rect 28720 26440 28729 26480
rect 28343 26398 28390 26440
rect 28514 26398 28558 26440
rect 28682 26398 28729 26440
rect 40343 26480 40390 26522
rect 40514 26480 40558 26522
rect 40682 26480 40729 26522
rect 40343 26440 40352 26480
rect 40514 26440 40516 26480
rect 40556 26440 40558 26480
rect 40720 26440 40729 26480
rect 40343 26398 40390 26440
rect 40514 26398 40558 26440
rect 40682 26398 40729 26440
rect 52343 26480 52390 26522
rect 52514 26480 52558 26522
rect 52682 26480 52729 26522
rect 52343 26440 52352 26480
rect 52514 26440 52516 26480
rect 52556 26440 52558 26480
rect 52720 26440 52729 26480
rect 52343 26398 52390 26440
rect 52514 26398 52558 26440
rect 52682 26398 52729 26440
rect 64343 26480 64390 26522
rect 64514 26480 64558 26522
rect 64682 26480 64729 26522
rect 64343 26440 64352 26480
rect 64514 26440 64516 26480
rect 64556 26440 64558 26480
rect 64720 26440 64729 26480
rect 64343 26398 64390 26440
rect 64514 26398 64558 26440
rect 64682 26398 64729 26440
rect 76343 26480 76390 26522
rect 76514 26480 76558 26522
rect 76682 26480 76729 26522
rect 76343 26440 76352 26480
rect 76514 26440 76516 26480
rect 76556 26440 76558 26480
rect 76720 26440 76729 26480
rect 76343 26398 76390 26440
rect 76514 26398 76558 26440
rect 76682 26398 76729 26440
rect 3103 25724 3150 25766
rect 3274 25724 3318 25766
rect 3442 25724 3489 25766
rect 3103 25684 3112 25724
rect 3274 25684 3276 25724
rect 3316 25684 3318 25724
rect 3480 25684 3489 25724
rect 3103 25642 3150 25684
rect 3274 25642 3318 25684
rect 3442 25642 3489 25684
rect 15103 25724 15150 25766
rect 15274 25724 15318 25766
rect 15442 25724 15489 25766
rect 15103 25684 15112 25724
rect 15274 25684 15276 25724
rect 15316 25684 15318 25724
rect 15480 25684 15489 25724
rect 15103 25642 15150 25684
rect 15274 25642 15318 25684
rect 15442 25642 15489 25684
rect 27103 25724 27150 25766
rect 27274 25724 27318 25766
rect 27442 25724 27489 25766
rect 27103 25684 27112 25724
rect 27274 25684 27276 25724
rect 27316 25684 27318 25724
rect 27480 25684 27489 25724
rect 27103 25642 27150 25684
rect 27274 25642 27318 25684
rect 27442 25642 27489 25684
rect 39103 25724 39150 25766
rect 39274 25724 39318 25766
rect 39442 25724 39489 25766
rect 39103 25684 39112 25724
rect 39274 25684 39276 25724
rect 39316 25684 39318 25724
rect 39480 25684 39489 25724
rect 39103 25642 39150 25684
rect 39274 25642 39318 25684
rect 39442 25642 39489 25684
rect 51103 25724 51150 25766
rect 51274 25724 51318 25766
rect 51442 25724 51489 25766
rect 51103 25684 51112 25724
rect 51274 25684 51276 25724
rect 51316 25684 51318 25724
rect 51480 25684 51489 25724
rect 51103 25642 51150 25684
rect 51274 25642 51318 25684
rect 51442 25642 51489 25684
rect 63103 25724 63150 25766
rect 63274 25724 63318 25766
rect 63442 25724 63489 25766
rect 63103 25684 63112 25724
rect 63274 25684 63276 25724
rect 63316 25684 63318 25724
rect 63480 25684 63489 25724
rect 63103 25642 63150 25684
rect 63274 25642 63318 25684
rect 63442 25642 63489 25684
rect 75103 25724 75150 25766
rect 75274 25724 75318 25766
rect 75442 25724 75489 25766
rect 75103 25684 75112 25724
rect 75274 25684 75276 25724
rect 75316 25684 75318 25724
rect 75480 25684 75489 25724
rect 75103 25642 75150 25684
rect 75274 25642 75318 25684
rect 75442 25642 75489 25684
rect 40291 25348 40300 25388
rect 40340 25348 49996 25388
rect 50036 25348 58732 25388
rect 58772 25348 58781 25388
rect 45571 25264 45580 25304
rect 45620 25264 59116 25304
rect 59156 25264 59165 25304
rect 49123 25180 49132 25220
rect 49172 25180 61900 25220
rect 61940 25180 61949 25220
rect 41059 25096 41068 25136
rect 41108 25096 57964 25136
rect 58004 25096 58013 25136
rect 4343 24968 4390 25010
rect 4514 24968 4558 25010
rect 4682 24968 4729 25010
rect 4343 24928 4352 24968
rect 4514 24928 4516 24968
rect 4556 24928 4558 24968
rect 4720 24928 4729 24968
rect 4343 24886 4390 24928
rect 4514 24886 4558 24928
rect 4682 24886 4729 24928
rect 16343 24968 16390 25010
rect 16514 24968 16558 25010
rect 16682 24968 16729 25010
rect 16343 24928 16352 24968
rect 16514 24928 16516 24968
rect 16556 24928 16558 24968
rect 16720 24928 16729 24968
rect 16343 24886 16390 24928
rect 16514 24886 16558 24928
rect 16682 24886 16729 24928
rect 28343 24968 28390 25010
rect 28514 24968 28558 25010
rect 28682 24968 28729 25010
rect 28343 24928 28352 24968
rect 28514 24928 28516 24968
rect 28556 24928 28558 24968
rect 28720 24928 28729 24968
rect 28343 24886 28390 24928
rect 28514 24886 28558 24928
rect 28682 24886 28729 24928
rect 40343 24968 40390 25010
rect 40514 24968 40558 25010
rect 40682 24968 40729 25010
rect 40343 24928 40352 24968
rect 40514 24928 40516 24968
rect 40556 24928 40558 24968
rect 40720 24928 40729 24968
rect 40343 24886 40390 24928
rect 40514 24886 40558 24928
rect 40682 24886 40729 24928
rect 52343 24968 52390 25010
rect 52514 24968 52558 25010
rect 52682 24968 52729 25010
rect 64343 24968 64390 25010
rect 64514 24968 64558 25010
rect 64682 24968 64729 25010
rect 52343 24928 52352 24968
rect 52514 24928 52516 24968
rect 52556 24928 52558 24968
rect 52720 24928 52729 24968
rect 56131 24928 56140 24968
rect 56180 24928 57580 24968
rect 57620 24928 57629 24968
rect 64343 24928 64352 24968
rect 64514 24928 64516 24968
rect 64556 24928 64558 24968
rect 64720 24928 64729 24968
rect 52343 24886 52390 24928
rect 52514 24886 52558 24928
rect 52682 24886 52729 24928
rect 64343 24886 64390 24928
rect 64514 24886 64558 24928
rect 64682 24886 64729 24928
rect 76343 24968 76390 25010
rect 76514 24968 76558 25010
rect 76682 24968 76729 25010
rect 76343 24928 76352 24968
rect 76514 24928 76516 24968
rect 76556 24928 76558 24968
rect 76720 24928 76729 24968
rect 76343 24886 76390 24928
rect 76514 24886 76558 24928
rect 76682 24886 76729 24928
rect 51907 24760 51916 24800
rect 51956 24760 78988 24800
rect 79028 24760 79037 24800
rect 52099 24676 52108 24716
rect 52148 24676 55756 24716
rect 55796 24676 55805 24716
rect 51619 24592 51628 24632
rect 51668 24592 57772 24632
rect 57812 24592 57821 24632
rect 51715 24508 51724 24548
rect 51764 24508 54892 24548
rect 54932 24508 54941 24548
rect 3103 24212 3150 24254
rect 3274 24212 3318 24254
rect 3442 24212 3489 24254
rect 3103 24172 3112 24212
rect 3274 24172 3276 24212
rect 3316 24172 3318 24212
rect 3480 24172 3489 24212
rect 3103 24130 3150 24172
rect 3274 24130 3318 24172
rect 3442 24130 3489 24172
rect 15103 24212 15150 24254
rect 15274 24212 15318 24254
rect 15442 24212 15489 24254
rect 15103 24172 15112 24212
rect 15274 24172 15276 24212
rect 15316 24172 15318 24212
rect 15480 24172 15489 24212
rect 15103 24130 15150 24172
rect 15274 24130 15318 24172
rect 15442 24130 15489 24172
rect 27103 24212 27150 24254
rect 27274 24212 27318 24254
rect 27442 24212 27489 24254
rect 27103 24172 27112 24212
rect 27274 24172 27276 24212
rect 27316 24172 27318 24212
rect 27480 24172 27489 24212
rect 27103 24130 27150 24172
rect 27274 24130 27318 24172
rect 27442 24130 27489 24172
rect 39103 24212 39150 24254
rect 39274 24212 39318 24254
rect 39442 24212 39489 24254
rect 39103 24172 39112 24212
rect 39274 24172 39276 24212
rect 39316 24172 39318 24212
rect 39480 24172 39489 24212
rect 56227 24172 56236 24212
rect 56276 24172 56620 24212
rect 56660 24172 56669 24212
rect 39103 24130 39150 24172
rect 39274 24130 39318 24172
rect 39442 24130 39489 24172
rect 51811 23920 51820 23960
rect 51860 23920 64780 23960
rect 64820 23920 64829 23960
rect 53059 23836 53068 23876
rect 53108 23836 66508 23876
rect 66548 23836 66557 23876
rect 48739 23752 48748 23792
rect 48788 23752 60460 23792
rect 60500 23752 60509 23792
rect 78822 23752 78988 23792
rect 79028 23752 79037 23792
rect 39811 23668 39820 23708
rect 39860 23668 57676 23708
rect 57716 23668 57725 23708
rect 57859 23668 57868 23708
rect 57908 23668 58252 23708
rect 58292 23668 66604 23708
rect 66644 23668 66653 23708
rect 43459 23584 43468 23624
rect 43508 23584 59020 23624
rect 59060 23584 59069 23624
rect 53452 23500 55852 23540
rect 55892 23500 55901 23540
rect 56419 23500 56428 23540
rect 56468 23500 66316 23540
rect 66356 23500 66365 23540
rect 4343 23456 4390 23498
rect 4514 23456 4558 23498
rect 4682 23456 4729 23498
rect 4343 23416 4352 23456
rect 4514 23416 4516 23456
rect 4556 23416 4558 23456
rect 4720 23416 4729 23456
rect 4343 23374 4390 23416
rect 4514 23374 4558 23416
rect 4682 23374 4729 23416
rect 16343 23456 16390 23498
rect 16514 23456 16558 23498
rect 16682 23456 16729 23498
rect 16343 23416 16352 23456
rect 16514 23416 16516 23456
rect 16556 23416 16558 23456
rect 16720 23416 16729 23456
rect 16343 23374 16390 23416
rect 16514 23374 16558 23416
rect 16682 23374 16729 23416
rect 28343 23456 28390 23498
rect 28514 23456 28558 23498
rect 28682 23456 28729 23498
rect 28343 23416 28352 23456
rect 28514 23416 28516 23456
rect 28556 23416 28558 23456
rect 28720 23416 28729 23456
rect 28343 23374 28390 23416
rect 28514 23374 28558 23416
rect 28682 23374 28729 23416
rect 40343 23456 40390 23498
rect 40514 23456 40558 23498
rect 40682 23456 40729 23498
rect 53452 23456 53492 23500
rect 40343 23416 40352 23456
rect 40514 23416 40516 23456
rect 40556 23416 40558 23456
rect 40720 23416 40729 23456
rect 52579 23416 52588 23456
rect 52628 23416 53492 23456
rect 53731 23416 53740 23456
rect 53780 23416 56236 23456
rect 56276 23416 56285 23456
rect 40343 23374 40390 23416
rect 40514 23374 40558 23416
rect 40682 23374 40729 23416
rect 52675 23332 52684 23372
rect 52724 23332 55564 23372
rect 55604 23332 55613 23372
rect 38851 23248 38860 23288
rect 38900 23248 53740 23288
rect 53780 23248 53789 23288
rect 54116 23248 55180 23288
rect 55220 23248 55229 23288
rect 54116 23204 54156 23248
rect 52195 23164 52204 23204
rect 52244 23164 54156 23204
rect 54211 23164 54220 23204
rect 54260 23164 54508 23204
rect 54548 23164 66220 23204
rect 66260 23164 66269 23204
rect 52291 23080 52300 23120
rect 52340 23080 55084 23120
rect 55124 23080 55133 23120
rect 74262 23080 75148 23120
rect 75188 23080 75197 23120
rect 52867 22996 52876 23036
rect 52916 22996 53452 23036
rect 53492 22996 53501 23036
rect 53635 22996 53644 23036
rect 53684 22996 60748 23036
rect 60788 22996 60797 23036
rect 52963 22912 52972 22952
rect 53012 22912 54700 22952
rect 54740 22912 54749 22952
rect 52387 22828 52396 22868
rect 52436 22828 57100 22868
rect 57140 22828 57149 22868
rect 51811 22744 51820 22784
rect 51860 22744 53356 22784
rect 53396 22744 53405 22784
rect 3103 22700 3150 22742
rect 3274 22700 3318 22742
rect 3442 22700 3489 22742
rect 3103 22660 3112 22700
rect 3274 22660 3276 22700
rect 3316 22660 3318 22700
rect 3480 22660 3489 22700
rect 3103 22618 3150 22660
rect 3274 22618 3318 22660
rect 3442 22618 3489 22660
rect 15103 22700 15150 22742
rect 15274 22700 15318 22742
rect 15442 22700 15489 22742
rect 15103 22660 15112 22700
rect 15274 22660 15276 22700
rect 15316 22660 15318 22700
rect 15480 22660 15489 22700
rect 15103 22618 15150 22660
rect 15274 22618 15318 22660
rect 15442 22618 15489 22660
rect 27103 22700 27150 22742
rect 27274 22700 27318 22742
rect 27442 22700 27489 22742
rect 27103 22660 27112 22700
rect 27274 22660 27276 22700
rect 27316 22660 27318 22700
rect 27480 22660 27489 22700
rect 27103 22618 27150 22660
rect 27274 22618 27318 22660
rect 27442 22618 27489 22660
rect 39103 22700 39150 22742
rect 39274 22700 39318 22742
rect 39442 22700 39489 22742
rect 39103 22660 39112 22700
rect 39274 22660 39276 22700
rect 39316 22660 39318 22700
rect 39480 22660 39489 22700
rect 39103 22618 39150 22660
rect 39274 22618 39318 22660
rect 39442 22618 39489 22660
rect 64316 22541 64756 22652
rect 64316 22417 64390 22541
rect 64514 22417 64558 22541
rect 64682 22417 64756 22541
rect 64316 22373 64756 22417
rect 64316 22249 64390 22373
rect 64514 22249 64558 22373
rect 64682 22249 64756 22373
rect 64316 22205 64756 22249
rect 64316 22081 64390 22205
rect 64514 22081 64558 22205
rect 64682 22081 64756 22205
rect 64316 22037 64756 22081
rect 4343 21944 4390 21986
rect 4514 21944 4558 21986
rect 4682 21944 4729 21986
rect 4343 21904 4352 21944
rect 4514 21904 4516 21944
rect 4556 21904 4558 21944
rect 4720 21904 4729 21944
rect 4343 21862 4390 21904
rect 4514 21862 4558 21904
rect 4682 21862 4729 21904
rect 16343 21944 16390 21986
rect 16514 21944 16558 21986
rect 16682 21944 16729 21986
rect 16343 21904 16352 21944
rect 16514 21904 16516 21944
rect 16556 21904 16558 21944
rect 16720 21904 16729 21944
rect 16343 21862 16390 21904
rect 16514 21862 16558 21904
rect 16682 21862 16729 21904
rect 28343 21944 28390 21986
rect 28514 21944 28558 21986
rect 28682 21944 28729 21986
rect 28343 21904 28352 21944
rect 28514 21904 28516 21944
rect 28556 21904 28558 21944
rect 28720 21904 28729 21944
rect 28343 21862 28390 21904
rect 28514 21862 28558 21904
rect 28682 21862 28729 21904
rect 40343 21944 40390 21986
rect 40514 21944 40558 21986
rect 40682 21944 40729 21986
rect 40343 21904 40352 21944
rect 40514 21904 40516 21944
rect 40556 21904 40558 21944
rect 40720 21904 40729 21944
rect 40343 21862 40390 21904
rect 40514 21862 40558 21904
rect 40682 21862 40729 21904
rect 64316 21913 64390 22037
rect 64514 21913 64558 22037
rect 64682 21913 64756 22037
rect 64316 21869 64756 21913
rect 64316 21745 64390 21869
rect 64514 21745 64558 21869
rect 64682 21745 64756 21869
rect 64316 21701 64756 21745
rect 4579 21568 4588 21608
rect 4628 21568 5820 21608
rect 5923 21568 5932 21608
rect 5972 21568 52492 21608
rect 52532 21568 52876 21608
rect 52916 21568 52925 21608
rect 64316 21577 64390 21701
rect 64514 21577 64558 21701
rect 64682 21577 64756 21701
rect 5780 21524 5820 21568
rect 64316 21533 64756 21577
rect 5780 21484 50380 21524
rect 50420 21484 50429 21524
rect 3907 21400 3916 21440
rect 3956 21400 5932 21440
rect 5972 21400 5981 21440
rect 64316 21409 64390 21533
rect 64514 21409 64558 21533
rect 64682 21409 64756 21533
rect 64316 21365 64756 21409
rect 64316 21241 64390 21365
rect 64514 21241 64558 21365
rect 64682 21241 64756 21365
rect 3103 21188 3150 21230
rect 3274 21188 3318 21230
rect 3442 21188 3489 21230
rect 3103 21148 3112 21188
rect 3274 21148 3276 21188
rect 3316 21148 3318 21188
rect 3480 21148 3489 21188
rect 3103 21106 3150 21148
rect 3274 21106 3318 21148
rect 3442 21106 3489 21148
rect 15103 21188 15150 21230
rect 15274 21188 15318 21230
rect 15442 21188 15489 21230
rect 15103 21148 15112 21188
rect 15274 21148 15276 21188
rect 15316 21148 15318 21188
rect 15480 21148 15489 21188
rect 15103 21106 15150 21148
rect 15274 21106 15318 21148
rect 15442 21106 15489 21148
rect 27103 21188 27150 21230
rect 27274 21188 27318 21230
rect 27442 21188 27489 21230
rect 27103 21148 27112 21188
rect 27274 21148 27276 21188
rect 27316 21148 27318 21188
rect 27480 21148 27489 21188
rect 27103 21106 27150 21148
rect 27274 21106 27318 21148
rect 27442 21106 27489 21148
rect 39103 21188 39150 21230
rect 39274 21188 39318 21230
rect 39442 21188 39489 21230
rect 39103 21148 39112 21188
rect 39274 21148 39276 21188
rect 39316 21148 39318 21188
rect 39480 21148 39489 21188
rect 39103 21106 39150 21148
rect 39274 21106 39318 21148
rect 39442 21106 39489 21148
rect 64316 21197 64756 21241
rect 64316 21073 64390 21197
rect 64514 21073 64558 21197
rect 64682 21073 64756 21197
rect 64316 21029 64756 21073
rect 64316 20905 64390 21029
rect 64514 20905 64558 21029
rect 64682 20905 64756 21029
rect 64316 20861 64756 20905
rect 10915 20728 10924 20768
rect 10964 20728 51916 20768
rect 51956 20728 51965 20768
rect 64316 20737 64390 20861
rect 64514 20737 64558 20861
rect 64682 20737 64756 20861
rect 64316 20693 64756 20737
rect 64316 20569 64390 20693
rect 64514 20569 64558 20693
rect 64682 20569 64756 20693
rect 64316 20525 64756 20569
rect 4343 20432 4390 20474
rect 4514 20432 4558 20474
rect 4682 20432 4729 20474
rect 4343 20392 4352 20432
rect 4514 20392 4516 20432
rect 4556 20392 4558 20432
rect 4720 20392 4729 20432
rect 4343 20350 4390 20392
rect 4514 20350 4558 20392
rect 4682 20350 4729 20392
rect 16343 20432 16390 20474
rect 16514 20432 16558 20474
rect 16682 20432 16729 20474
rect 16343 20392 16352 20432
rect 16514 20392 16516 20432
rect 16556 20392 16558 20432
rect 16720 20392 16729 20432
rect 16343 20350 16390 20392
rect 16514 20350 16558 20392
rect 16682 20350 16729 20392
rect 28343 20432 28390 20474
rect 28514 20432 28558 20474
rect 28682 20432 28729 20474
rect 28343 20392 28352 20432
rect 28514 20392 28516 20432
rect 28556 20392 28558 20432
rect 28720 20392 28729 20432
rect 28343 20350 28390 20392
rect 28514 20350 28558 20392
rect 28682 20350 28729 20392
rect 40343 20432 40390 20474
rect 40514 20432 40558 20474
rect 40682 20432 40729 20474
rect 40343 20392 40352 20432
rect 40514 20392 40516 20432
rect 40556 20392 40558 20432
rect 40720 20392 40729 20432
rect 40343 20350 40390 20392
rect 40514 20350 40558 20392
rect 40682 20350 40729 20392
rect 64316 20401 64390 20525
rect 64514 20401 64558 20525
rect 64682 20401 64756 20525
rect 64316 20290 64756 20401
rect 76316 22541 76756 22652
rect 76316 22417 76390 22541
rect 76514 22417 76558 22541
rect 76682 22417 76756 22541
rect 76316 22373 76756 22417
rect 76316 22249 76390 22373
rect 76514 22249 76558 22373
rect 76682 22249 76756 22373
rect 76316 22205 76756 22249
rect 76316 22081 76390 22205
rect 76514 22081 76558 22205
rect 76682 22081 76756 22205
rect 76316 22037 76756 22081
rect 76316 21913 76390 22037
rect 76514 21913 76558 22037
rect 76682 21913 76756 22037
rect 76316 21869 76756 21913
rect 76316 21745 76390 21869
rect 76514 21745 76558 21869
rect 76682 21745 76756 21869
rect 76316 21701 76756 21745
rect 76316 21577 76390 21701
rect 76514 21577 76558 21701
rect 76682 21577 76756 21701
rect 76316 21533 76756 21577
rect 76316 21409 76390 21533
rect 76514 21409 76558 21533
rect 76682 21409 76756 21533
rect 76316 21365 76756 21409
rect 76316 21241 76390 21365
rect 76514 21241 76558 21365
rect 76682 21241 76756 21365
rect 76316 21197 76756 21241
rect 76316 21073 76390 21197
rect 76514 21073 76558 21197
rect 76682 21073 76756 21197
rect 76316 21029 76756 21073
rect 76316 20905 76390 21029
rect 76514 20905 76558 21029
rect 76682 20905 76756 21029
rect 76316 20861 76756 20905
rect 76316 20737 76390 20861
rect 76514 20737 76558 20861
rect 76682 20737 76756 20861
rect 76316 20693 76756 20737
rect 76316 20569 76390 20693
rect 76514 20569 76558 20693
rect 76682 20569 76756 20693
rect 76316 20525 76756 20569
rect 76316 20401 76390 20525
rect 76514 20401 76558 20525
rect 76682 20401 76756 20525
rect 76316 20290 76756 20401
rect 39907 19972 39916 20012
rect 39956 19972 40108 20012
rect 40148 19972 51916 20012
rect 51956 19972 51965 20012
rect 3103 19676 3150 19718
rect 3274 19676 3318 19718
rect 3442 19676 3489 19718
rect 3103 19636 3112 19676
rect 3274 19636 3276 19676
rect 3316 19636 3318 19676
rect 3480 19636 3489 19676
rect 3103 19594 3150 19636
rect 3274 19594 3318 19636
rect 3442 19594 3489 19636
rect 15103 19676 15150 19718
rect 15274 19676 15318 19718
rect 15442 19676 15489 19718
rect 15103 19636 15112 19676
rect 15274 19636 15276 19676
rect 15316 19636 15318 19676
rect 15480 19636 15489 19676
rect 15103 19594 15150 19636
rect 15274 19594 15318 19636
rect 15442 19594 15489 19636
rect 27103 19676 27150 19718
rect 27274 19676 27318 19718
rect 27442 19676 27489 19718
rect 27103 19636 27112 19676
rect 27274 19636 27276 19676
rect 27316 19636 27318 19676
rect 27480 19636 27489 19676
rect 27103 19594 27150 19636
rect 27274 19594 27318 19636
rect 27442 19594 27489 19636
rect 39103 19676 39150 19718
rect 39274 19676 39318 19718
rect 39442 19676 39489 19718
rect 39103 19636 39112 19676
rect 39274 19636 39276 19676
rect 39316 19636 39318 19676
rect 39480 19636 39489 19676
rect 39103 19594 39150 19636
rect 39274 19594 39318 19636
rect 39442 19594 39489 19636
rect 63076 19665 63516 19776
rect 63076 19541 63150 19665
rect 63274 19541 63318 19665
rect 63442 19541 63516 19665
rect 41731 19468 41740 19508
rect 41780 19468 51628 19508
rect 51668 19468 51677 19508
rect 63076 19497 63516 19541
rect 41827 19384 41836 19424
rect 41876 19384 52300 19424
rect 52340 19384 52349 19424
rect 63076 19373 63150 19497
rect 63274 19373 63318 19497
rect 63442 19373 63516 19497
rect 63076 19329 63516 19373
rect 63076 19205 63150 19329
rect 63274 19205 63318 19329
rect 63442 19205 63516 19329
rect 63076 19161 63516 19205
rect 63076 19037 63150 19161
rect 63274 19037 63318 19161
rect 63442 19037 63516 19161
rect 63076 18993 63516 19037
rect 4343 18920 4390 18962
rect 4514 18920 4558 18962
rect 4682 18920 4729 18962
rect 4343 18880 4352 18920
rect 4514 18880 4516 18920
rect 4556 18880 4558 18920
rect 4720 18880 4729 18920
rect 4343 18838 4390 18880
rect 4514 18838 4558 18880
rect 4682 18838 4729 18880
rect 16343 18920 16390 18962
rect 16514 18920 16558 18962
rect 16682 18920 16729 18962
rect 16343 18880 16352 18920
rect 16514 18880 16516 18920
rect 16556 18880 16558 18920
rect 16720 18880 16729 18920
rect 16343 18838 16390 18880
rect 16514 18838 16558 18880
rect 16682 18838 16729 18880
rect 28343 18920 28390 18962
rect 28514 18920 28558 18962
rect 28682 18920 28729 18962
rect 28343 18880 28352 18920
rect 28514 18880 28516 18920
rect 28556 18880 28558 18920
rect 28720 18880 28729 18920
rect 28343 18838 28390 18880
rect 28514 18838 28558 18880
rect 28682 18838 28729 18880
rect 40343 18920 40390 18962
rect 40514 18920 40558 18962
rect 40682 18920 40729 18962
rect 40343 18880 40352 18920
rect 40514 18880 40516 18920
rect 40556 18880 40558 18920
rect 40720 18880 40729 18920
rect 40343 18838 40390 18880
rect 40514 18838 40558 18880
rect 40682 18838 40729 18880
rect 63076 18869 63150 18993
rect 63274 18869 63318 18993
rect 63442 18869 63516 18993
rect 63076 18825 63516 18869
rect 63076 18701 63150 18825
rect 63274 18701 63318 18825
rect 63442 18701 63516 18825
rect 63076 18657 63516 18701
rect 7651 18544 7660 18584
rect 7700 18544 41836 18584
rect 41876 18544 41885 18584
rect 63076 18533 63150 18657
rect 63274 18533 63318 18657
rect 63442 18533 63516 18657
rect 63076 18489 63516 18533
rect 63076 18365 63150 18489
rect 63274 18365 63318 18489
rect 63442 18365 63516 18489
rect 63076 18321 63516 18365
rect 3103 18164 3150 18206
rect 3274 18164 3318 18206
rect 3442 18164 3489 18206
rect 3103 18124 3112 18164
rect 3274 18124 3276 18164
rect 3316 18124 3318 18164
rect 3480 18124 3489 18164
rect 3103 18082 3150 18124
rect 3274 18082 3318 18124
rect 3442 18082 3489 18124
rect 15103 18164 15150 18206
rect 15274 18164 15318 18206
rect 15442 18164 15489 18206
rect 15103 18124 15112 18164
rect 15274 18124 15276 18164
rect 15316 18124 15318 18164
rect 15480 18124 15489 18164
rect 15103 18082 15150 18124
rect 15274 18082 15318 18124
rect 15442 18082 15489 18124
rect 27103 18164 27150 18206
rect 27274 18164 27318 18206
rect 27442 18164 27489 18206
rect 27103 18124 27112 18164
rect 27274 18124 27276 18164
rect 27316 18124 27318 18164
rect 27480 18124 27489 18164
rect 27103 18082 27150 18124
rect 27274 18082 27318 18124
rect 27442 18082 27489 18124
rect 39103 18164 39150 18206
rect 39274 18164 39318 18206
rect 39442 18164 39489 18206
rect 39103 18124 39112 18164
rect 39274 18124 39276 18164
rect 39316 18124 39318 18164
rect 39480 18124 39489 18164
rect 39103 18082 39150 18124
rect 39274 18082 39318 18124
rect 39442 18082 39489 18124
rect 63076 18197 63150 18321
rect 63274 18197 63318 18321
rect 63442 18197 63516 18321
rect 63076 18153 63516 18197
rect 63076 18029 63150 18153
rect 63274 18029 63318 18153
rect 63442 18029 63516 18153
rect 63076 17985 63516 18029
rect 63076 17861 63150 17985
rect 63274 17861 63318 17985
rect 63442 17861 63516 17985
rect 63076 17817 63516 17861
rect 63076 17693 63150 17817
rect 63274 17693 63318 17817
rect 63442 17693 63516 17817
rect 63076 17649 63516 17693
rect 7555 17536 7564 17576
rect 7604 17536 31756 17576
rect 31796 17536 31805 17576
rect 63076 17525 63150 17649
rect 63274 17525 63318 17649
rect 63442 17525 63516 17649
rect 4343 17408 4390 17450
rect 4514 17408 4558 17450
rect 4682 17408 4729 17450
rect 4343 17368 4352 17408
rect 4514 17368 4516 17408
rect 4556 17368 4558 17408
rect 4720 17368 4729 17408
rect 4343 17326 4390 17368
rect 4514 17326 4558 17368
rect 4682 17326 4729 17368
rect 16343 17408 16390 17450
rect 16514 17408 16558 17450
rect 16682 17408 16729 17450
rect 16343 17368 16352 17408
rect 16514 17368 16516 17408
rect 16556 17368 16558 17408
rect 16720 17368 16729 17408
rect 16343 17326 16390 17368
rect 16514 17326 16558 17368
rect 16682 17326 16729 17368
rect 28343 17408 28390 17450
rect 28514 17408 28558 17450
rect 28682 17408 28729 17450
rect 28343 17368 28352 17408
rect 28514 17368 28516 17408
rect 28556 17368 28558 17408
rect 28720 17368 28729 17408
rect 28343 17326 28390 17368
rect 28514 17326 28558 17368
rect 28682 17326 28729 17368
rect 40343 17408 40390 17450
rect 40514 17408 40558 17450
rect 40682 17408 40729 17450
rect 63076 17414 63516 17525
rect 75076 19665 75516 19776
rect 75076 19541 75150 19665
rect 75274 19541 75318 19665
rect 75442 19541 75516 19665
rect 75076 19497 75516 19541
rect 75076 19373 75150 19497
rect 75274 19373 75318 19497
rect 75442 19373 75516 19497
rect 75076 19329 75516 19373
rect 75076 19205 75150 19329
rect 75274 19205 75318 19329
rect 75442 19205 75516 19329
rect 75076 19161 75516 19205
rect 75076 19037 75150 19161
rect 75274 19037 75318 19161
rect 75442 19037 75516 19161
rect 75076 18993 75516 19037
rect 75076 18869 75150 18993
rect 75274 18869 75318 18993
rect 75442 18869 75516 18993
rect 75076 18825 75516 18869
rect 75076 18701 75150 18825
rect 75274 18701 75318 18825
rect 75442 18701 75516 18825
rect 75076 18657 75516 18701
rect 75076 18533 75150 18657
rect 75274 18533 75318 18657
rect 75442 18533 75516 18657
rect 75076 18489 75516 18533
rect 75076 18365 75150 18489
rect 75274 18365 75318 18489
rect 75442 18365 75516 18489
rect 75076 18321 75516 18365
rect 75076 18197 75150 18321
rect 75274 18197 75318 18321
rect 75442 18197 75516 18321
rect 75076 18153 75516 18197
rect 75076 18029 75150 18153
rect 75274 18029 75318 18153
rect 75442 18029 75516 18153
rect 75076 17985 75516 18029
rect 75076 17861 75150 17985
rect 75274 17861 75318 17985
rect 75442 17861 75516 17985
rect 75076 17817 75516 17861
rect 75076 17693 75150 17817
rect 75274 17693 75318 17817
rect 75442 17693 75516 17817
rect 75076 17649 75516 17693
rect 75076 17525 75150 17649
rect 75274 17525 75318 17649
rect 75442 17525 75516 17649
rect 75076 17414 75516 17525
rect 40343 17368 40352 17408
rect 40514 17368 40516 17408
rect 40556 17368 40558 17408
rect 40720 17368 40729 17408
rect 40343 17326 40390 17368
rect 40514 17326 40558 17368
rect 40682 17326 40729 17368
rect 51811 17200 51820 17240
rect 51860 17200 56812 17240
rect 56852 17200 56861 17240
rect 74262 17200 74860 17240
rect 74900 17200 74909 17240
rect 51907 17116 51916 17156
rect 51956 17116 56140 17156
rect 56180 17116 56189 17156
rect 56323 17116 56332 17156
rect 56372 17116 63916 17156
rect 63956 17116 63965 17156
rect 42403 17032 42412 17072
rect 42452 17032 57580 17072
rect 57620 17032 57629 17072
rect 34723 16948 34732 16988
rect 34772 16948 57292 16988
rect 57332 16948 57341 16988
rect 37987 16864 37996 16904
rect 38036 16864 54700 16904
rect 54740 16864 54749 16904
rect 60451 16864 60460 16904
rect 60500 16864 66220 16904
rect 66260 16864 66269 16904
rect 35299 16780 35308 16820
rect 35348 16780 57388 16820
rect 57428 16780 57437 16820
rect 3103 16652 3150 16694
rect 3274 16652 3318 16694
rect 3442 16652 3489 16694
rect 3103 16612 3112 16652
rect 3274 16612 3276 16652
rect 3316 16612 3318 16652
rect 3480 16612 3489 16652
rect 3103 16570 3150 16612
rect 3274 16570 3318 16612
rect 3442 16570 3489 16612
rect 15103 16652 15150 16694
rect 15274 16652 15318 16694
rect 15442 16652 15489 16694
rect 15103 16612 15112 16652
rect 15274 16612 15276 16652
rect 15316 16612 15318 16652
rect 15480 16612 15489 16652
rect 15103 16570 15150 16612
rect 15274 16570 15318 16612
rect 15442 16570 15489 16612
rect 27103 16652 27150 16694
rect 27274 16652 27318 16694
rect 27442 16652 27489 16694
rect 27103 16612 27112 16652
rect 27274 16612 27276 16652
rect 27316 16612 27318 16652
rect 27480 16612 27489 16652
rect 27103 16570 27150 16612
rect 27274 16570 27318 16612
rect 27442 16570 27489 16612
rect 39103 16652 39150 16694
rect 39274 16652 39318 16694
rect 39442 16652 39489 16694
rect 39103 16612 39112 16652
rect 39274 16612 39276 16652
rect 39316 16612 39318 16652
rect 39480 16612 39489 16652
rect 39103 16570 39150 16612
rect 39274 16570 39318 16612
rect 39442 16570 39489 16612
rect 65347 16528 65356 16568
rect 65396 16528 65740 16568
rect 65780 16528 69100 16568
rect 69140 16528 69149 16568
rect 38275 16444 38284 16484
rect 38324 16444 56716 16484
rect 56756 16444 56765 16484
rect 71779 16360 71788 16400
rect 71828 16360 71858 16400
rect 60739 16276 60748 16316
rect 60788 16276 70924 16316
rect 70964 16276 70973 16316
rect 78499 16192 78508 16232
rect 78548 16192 78698 16232
rect 42787 16108 42796 16148
rect 42836 16108 59020 16148
rect 59060 16108 59069 16148
rect 41155 16024 41164 16064
rect 41204 16024 58924 16064
rect 58964 16024 58973 16064
rect 51139 15940 51148 15980
rect 51188 15940 61996 15980
rect 62036 15940 62045 15980
rect 4343 15896 4390 15938
rect 4514 15896 4558 15938
rect 4682 15896 4729 15938
rect 4343 15856 4352 15896
rect 4514 15856 4516 15896
rect 4556 15856 4558 15896
rect 4720 15856 4729 15896
rect 4343 15814 4390 15856
rect 4514 15814 4558 15856
rect 4682 15814 4729 15856
rect 16343 15896 16390 15938
rect 16514 15896 16558 15938
rect 16682 15896 16729 15938
rect 16343 15856 16352 15896
rect 16514 15856 16516 15896
rect 16556 15856 16558 15896
rect 16720 15856 16729 15896
rect 16343 15814 16390 15856
rect 16514 15814 16558 15856
rect 16682 15814 16729 15856
rect 28343 15896 28390 15938
rect 28514 15896 28558 15938
rect 28682 15896 28729 15938
rect 28343 15856 28352 15896
rect 28514 15856 28516 15896
rect 28556 15856 28558 15896
rect 28720 15856 28729 15896
rect 28343 15814 28390 15856
rect 28514 15814 28558 15856
rect 28682 15814 28729 15856
rect 40343 15896 40390 15938
rect 40514 15896 40558 15938
rect 40682 15896 40729 15938
rect 40343 15856 40352 15896
rect 40514 15856 40516 15896
rect 40556 15856 40558 15896
rect 40720 15856 40729 15896
rect 52195 15856 52204 15896
rect 52244 15856 61900 15896
rect 61940 15856 61949 15896
rect 40343 15814 40390 15856
rect 40514 15814 40558 15856
rect 40682 15814 40729 15856
rect 40867 15772 40876 15812
rect 40916 15772 43220 15812
rect 52003 15772 52012 15812
rect 52052 15772 60748 15812
rect 60788 15772 60797 15812
rect 43180 15476 43220 15772
rect 48931 15688 48940 15728
rect 48980 15688 53260 15728
rect 53300 15688 53309 15728
rect 60547 15688 60556 15728
rect 60596 15688 64108 15728
rect 64148 15688 64157 15728
rect 47779 15604 47788 15644
rect 47828 15604 59404 15644
rect 59444 15604 59453 15644
rect 50275 15520 50284 15560
rect 50324 15520 54604 15560
rect 54644 15520 54653 15560
rect 43180 15436 56428 15476
rect 56468 15436 56477 15476
rect 61891 15436 61900 15476
rect 61940 15436 62284 15476
rect 62324 15436 70732 15476
rect 70772 15436 70781 15476
rect 33187 15352 33196 15392
rect 33236 15352 57676 15392
rect 57716 15352 57725 15392
rect 47875 15268 47884 15308
rect 47924 15268 59692 15308
rect 59732 15268 59741 15308
rect 3103 15140 3150 15182
rect 3274 15140 3318 15182
rect 3442 15140 3489 15182
rect 3103 15100 3112 15140
rect 3274 15100 3276 15140
rect 3316 15100 3318 15140
rect 3480 15100 3489 15140
rect 3103 15058 3150 15100
rect 3274 15058 3318 15100
rect 3442 15058 3489 15100
rect 15103 15140 15150 15182
rect 15274 15140 15318 15182
rect 15442 15140 15489 15182
rect 15103 15100 15112 15140
rect 15274 15100 15276 15140
rect 15316 15100 15318 15140
rect 15480 15100 15489 15140
rect 15103 15058 15150 15100
rect 15274 15058 15318 15100
rect 15442 15058 15489 15100
rect 27103 15140 27150 15182
rect 27274 15140 27318 15182
rect 27442 15140 27489 15182
rect 27103 15100 27112 15140
rect 27274 15100 27276 15140
rect 27316 15100 27318 15140
rect 27480 15100 27489 15140
rect 27103 15058 27150 15100
rect 27274 15058 27318 15100
rect 27442 15058 27489 15100
rect 39103 15140 39150 15182
rect 39274 15140 39318 15182
rect 39442 15140 39489 15182
rect 39103 15100 39112 15140
rect 39274 15100 39276 15140
rect 39316 15100 39318 15140
rect 39480 15100 39489 15140
rect 39103 15058 39150 15100
rect 39274 15058 39318 15100
rect 39442 15058 39489 15100
rect 51103 15140 51150 15182
rect 51274 15140 51318 15182
rect 51442 15140 51489 15182
rect 51103 15100 51112 15140
rect 51274 15100 51276 15140
rect 51316 15100 51318 15140
rect 51480 15100 51489 15140
rect 51103 15058 51150 15100
rect 51274 15058 51318 15100
rect 51442 15058 51489 15100
rect 63103 15140 63150 15182
rect 63274 15140 63318 15182
rect 63442 15140 63489 15182
rect 63103 15100 63112 15140
rect 63274 15100 63276 15140
rect 63316 15100 63318 15140
rect 63480 15100 63489 15140
rect 63103 15058 63150 15100
rect 63274 15058 63318 15100
rect 63442 15058 63489 15100
rect 75103 15140 75150 15182
rect 75274 15140 75318 15182
rect 75442 15140 75489 15182
rect 75103 15100 75112 15140
rect 75274 15100 75276 15140
rect 75316 15100 75318 15140
rect 75480 15100 75489 15140
rect 75103 15058 75150 15100
rect 75274 15058 75318 15100
rect 75442 15058 75489 15100
rect 36739 14932 36748 14972
rect 36788 14932 58060 14972
rect 58100 14932 58109 14972
rect 40771 14848 40780 14888
rect 40820 14848 58444 14888
rect 58484 14848 58493 14888
rect 49891 14764 49900 14804
rect 49940 14764 60364 14804
rect 60404 14764 60413 14804
rect 50083 14680 50092 14720
rect 50132 14680 61900 14720
rect 61940 14680 61949 14720
rect 4343 14384 4390 14426
rect 4514 14384 4558 14426
rect 4682 14384 4729 14426
rect 4343 14344 4352 14384
rect 4514 14344 4516 14384
rect 4556 14344 4558 14384
rect 4720 14344 4729 14384
rect 4343 14302 4390 14344
rect 4514 14302 4558 14344
rect 4682 14302 4729 14344
rect 16343 14384 16390 14426
rect 16514 14384 16558 14426
rect 16682 14384 16729 14426
rect 16343 14344 16352 14384
rect 16514 14344 16516 14384
rect 16556 14344 16558 14384
rect 16720 14344 16729 14384
rect 16343 14302 16390 14344
rect 16514 14302 16558 14344
rect 16682 14302 16729 14344
rect 28343 14384 28390 14426
rect 28514 14384 28558 14426
rect 28682 14384 28729 14426
rect 28343 14344 28352 14384
rect 28514 14344 28516 14384
rect 28556 14344 28558 14384
rect 28720 14344 28729 14384
rect 28343 14302 28390 14344
rect 28514 14302 28558 14344
rect 28682 14302 28729 14344
rect 40343 14384 40390 14426
rect 40514 14384 40558 14426
rect 40682 14384 40729 14426
rect 40343 14344 40352 14384
rect 40514 14344 40516 14384
rect 40556 14344 40558 14384
rect 40720 14344 40729 14384
rect 40343 14302 40390 14344
rect 40514 14302 40558 14344
rect 40682 14302 40729 14344
rect 52343 14384 52390 14426
rect 52514 14384 52558 14426
rect 52682 14384 52729 14426
rect 52343 14344 52352 14384
rect 52514 14344 52516 14384
rect 52556 14344 52558 14384
rect 52720 14344 52729 14384
rect 52343 14302 52390 14344
rect 52514 14302 52558 14344
rect 52682 14302 52729 14344
rect 64343 14384 64390 14426
rect 64514 14384 64558 14426
rect 64682 14384 64729 14426
rect 64343 14344 64352 14384
rect 64514 14344 64516 14384
rect 64556 14344 64558 14384
rect 64720 14344 64729 14384
rect 64343 14302 64390 14344
rect 64514 14302 64558 14344
rect 64682 14302 64729 14344
rect 76343 14384 76390 14426
rect 76514 14384 76558 14426
rect 76682 14384 76729 14426
rect 76343 14344 76352 14384
rect 76514 14344 76516 14384
rect 76556 14344 76558 14384
rect 76720 14344 76729 14384
rect 76343 14302 76390 14344
rect 76514 14302 76558 14344
rect 76682 14302 76729 14344
rect 49987 14176 49996 14216
rect 50036 14176 59116 14216
rect 59156 14176 59165 14216
rect 3103 13628 3150 13670
rect 3274 13628 3318 13670
rect 3442 13628 3489 13670
rect 3103 13588 3112 13628
rect 3274 13588 3276 13628
rect 3316 13588 3318 13628
rect 3480 13588 3489 13628
rect 3103 13546 3150 13588
rect 3274 13546 3318 13588
rect 3442 13546 3489 13588
rect 15103 13628 15150 13670
rect 15274 13628 15318 13670
rect 15442 13628 15489 13670
rect 15103 13588 15112 13628
rect 15274 13588 15276 13628
rect 15316 13588 15318 13628
rect 15480 13588 15489 13628
rect 15103 13546 15150 13588
rect 15274 13546 15318 13588
rect 15442 13546 15489 13588
rect 27103 13628 27150 13670
rect 27274 13628 27318 13670
rect 27442 13628 27489 13670
rect 27103 13588 27112 13628
rect 27274 13588 27276 13628
rect 27316 13588 27318 13628
rect 27480 13588 27489 13628
rect 27103 13546 27150 13588
rect 27274 13546 27318 13588
rect 27442 13546 27489 13588
rect 39103 13628 39150 13670
rect 39274 13628 39318 13670
rect 39442 13628 39489 13670
rect 39103 13588 39112 13628
rect 39274 13588 39276 13628
rect 39316 13588 39318 13628
rect 39480 13588 39489 13628
rect 39103 13546 39150 13588
rect 39274 13546 39318 13588
rect 39442 13546 39489 13588
rect 51103 13628 51150 13670
rect 51274 13628 51318 13670
rect 51442 13628 51489 13670
rect 51103 13588 51112 13628
rect 51274 13588 51276 13628
rect 51316 13588 51318 13628
rect 51480 13588 51489 13628
rect 51103 13546 51150 13588
rect 51274 13546 51318 13588
rect 51442 13546 51489 13588
rect 63103 13628 63150 13670
rect 63274 13628 63318 13670
rect 63442 13628 63489 13670
rect 63103 13588 63112 13628
rect 63274 13588 63276 13628
rect 63316 13588 63318 13628
rect 63480 13588 63489 13628
rect 63103 13546 63150 13588
rect 63274 13546 63318 13588
rect 63442 13546 63489 13588
rect 75103 13628 75150 13670
rect 75274 13628 75318 13670
rect 75442 13628 75489 13670
rect 75103 13588 75112 13628
rect 75274 13588 75276 13628
rect 75316 13588 75318 13628
rect 75480 13588 75489 13628
rect 75103 13546 75150 13588
rect 75274 13546 75318 13588
rect 75442 13546 75489 13588
rect 4343 12872 4390 12914
rect 4514 12872 4558 12914
rect 4682 12872 4729 12914
rect 4343 12832 4352 12872
rect 4514 12832 4516 12872
rect 4556 12832 4558 12872
rect 4720 12832 4729 12872
rect 4343 12790 4390 12832
rect 4514 12790 4558 12832
rect 4682 12790 4729 12832
rect 16343 12872 16390 12914
rect 16514 12872 16558 12914
rect 16682 12872 16729 12914
rect 16343 12832 16352 12872
rect 16514 12832 16516 12872
rect 16556 12832 16558 12872
rect 16720 12832 16729 12872
rect 16343 12790 16390 12832
rect 16514 12790 16558 12832
rect 16682 12790 16729 12832
rect 28343 12872 28390 12914
rect 28514 12872 28558 12914
rect 28682 12872 28729 12914
rect 28343 12832 28352 12872
rect 28514 12832 28516 12872
rect 28556 12832 28558 12872
rect 28720 12832 28729 12872
rect 28343 12790 28390 12832
rect 28514 12790 28558 12832
rect 28682 12790 28729 12832
rect 40343 12872 40390 12914
rect 40514 12872 40558 12914
rect 40682 12872 40729 12914
rect 40343 12832 40352 12872
rect 40514 12832 40516 12872
rect 40556 12832 40558 12872
rect 40720 12832 40729 12872
rect 40343 12790 40390 12832
rect 40514 12790 40558 12832
rect 40682 12790 40729 12832
rect 52343 12872 52390 12914
rect 52514 12872 52558 12914
rect 52682 12872 52729 12914
rect 52343 12832 52352 12872
rect 52514 12832 52516 12872
rect 52556 12832 52558 12872
rect 52720 12832 52729 12872
rect 52343 12790 52390 12832
rect 52514 12790 52558 12832
rect 52682 12790 52729 12832
rect 64343 12872 64390 12914
rect 64514 12872 64558 12914
rect 64682 12872 64729 12914
rect 64343 12832 64352 12872
rect 64514 12832 64516 12872
rect 64556 12832 64558 12872
rect 64720 12832 64729 12872
rect 64343 12790 64390 12832
rect 64514 12790 64558 12832
rect 64682 12790 64729 12832
rect 76343 12872 76390 12914
rect 76514 12872 76558 12914
rect 76682 12872 76729 12914
rect 76343 12832 76352 12872
rect 76514 12832 76516 12872
rect 76556 12832 76558 12872
rect 76720 12832 76729 12872
rect 76343 12790 76390 12832
rect 76514 12790 76558 12832
rect 76682 12790 76729 12832
rect 3103 12116 3150 12158
rect 3274 12116 3318 12158
rect 3442 12116 3489 12158
rect 3103 12076 3112 12116
rect 3274 12076 3276 12116
rect 3316 12076 3318 12116
rect 3480 12076 3489 12116
rect 3103 12034 3150 12076
rect 3274 12034 3318 12076
rect 3442 12034 3489 12076
rect 15103 12116 15150 12158
rect 15274 12116 15318 12158
rect 15442 12116 15489 12158
rect 15103 12076 15112 12116
rect 15274 12076 15276 12116
rect 15316 12076 15318 12116
rect 15480 12076 15489 12116
rect 15103 12034 15150 12076
rect 15274 12034 15318 12076
rect 15442 12034 15489 12076
rect 27103 12116 27150 12158
rect 27274 12116 27318 12158
rect 27442 12116 27489 12158
rect 27103 12076 27112 12116
rect 27274 12076 27276 12116
rect 27316 12076 27318 12116
rect 27480 12076 27489 12116
rect 27103 12034 27150 12076
rect 27274 12034 27318 12076
rect 27442 12034 27489 12076
rect 39103 12116 39150 12158
rect 39274 12116 39318 12158
rect 39442 12116 39489 12158
rect 39103 12076 39112 12116
rect 39274 12076 39276 12116
rect 39316 12076 39318 12116
rect 39480 12076 39489 12116
rect 39103 12034 39150 12076
rect 39274 12034 39318 12076
rect 39442 12034 39489 12076
rect 51103 12116 51150 12158
rect 51274 12116 51318 12158
rect 51442 12116 51489 12158
rect 51103 12076 51112 12116
rect 51274 12076 51276 12116
rect 51316 12076 51318 12116
rect 51480 12076 51489 12116
rect 51103 12034 51150 12076
rect 51274 12034 51318 12076
rect 51442 12034 51489 12076
rect 63103 12116 63150 12158
rect 63274 12116 63318 12158
rect 63442 12116 63489 12158
rect 63103 12076 63112 12116
rect 63274 12076 63276 12116
rect 63316 12076 63318 12116
rect 63480 12076 63489 12116
rect 63103 12034 63150 12076
rect 63274 12034 63318 12076
rect 63442 12034 63489 12076
rect 75103 12116 75150 12158
rect 75274 12116 75318 12158
rect 75442 12116 75489 12158
rect 75103 12076 75112 12116
rect 75274 12076 75276 12116
rect 75316 12076 75318 12116
rect 75480 12076 75489 12116
rect 75103 12034 75150 12076
rect 75274 12034 75318 12076
rect 75442 12034 75489 12076
rect 4343 11360 4390 11402
rect 4514 11360 4558 11402
rect 4682 11360 4729 11402
rect 4343 11320 4352 11360
rect 4514 11320 4516 11360
rect 4556 11320 4558 11360
rect 4720 11320 4729 11360
rect 4343 11278 4390 11320
rect 4514 11278 4558 11320
rect 4682 11278 4729 11320
rect 16343 11360 16390 11402
rect 16514 11360 16558 11402
rect 16682 11360 16729 11402
rect 16343 11320 16352 11360
rect 16514 11320 16516 11360
rect 16556 11320 16558 11360
rect 16720 11320 16729 11360
rect 16343 11278 16390 11320
rect 16514 11278 16558 11320
rect 16682 11278 16729 11320
rect 28343 11360 28390 11402
rect 28514 11360 28558 11402
rect 28682 11360 28729 11402
rect 28343 11320 28352 11360
rect 28514 11320 28516 11360
rect 28556 11320 28558 11360
rect 28720 11320 28729 11360
rect 28343 11278 28390 11320
rect 28514 11278 28558 11320
rect 28682 11278 28729 11320
rect 40343 11360 40390 11402
rect 40514 11360 40558 11402
rect 40682 11360 40729 11402
rect 40343 11320 40352 11360
rect 40514 11320 40516 11360
rect 40556 11320 40558 11360
rect 40720 11320 40729 11360
rect 40343 11278 40390 11320
rect 40514 11278 40558 11320
rect 40682 11278 40729 11320
rect 52343 11360 52390 11402
rect 52514 11360 52558 11402
rect 52682 11360 52729 11402
rect 52343 11320 52352 11360
rect 52514 11320 52516 11360
rect 52556 11320 52558 11360
rect 52720 11320 52729 11360
rect 52343 11278 52390 11320
rect 52514 11278 52558 11320
rect 52682 11278 52729 11320
rect 64343 11360 64390 11402
rect 64514 11360 64558 11402
rect 64682 11360 64729 11402
rect 64343 11320 64352 11360
rect 64514 11320 64516 11360
rect 64556 11320 64558 11360
rect 64720 11320 64729 11360
rect 64343 11278 64390 11320
rect 64514 11278 64558 11320
rect 64682 11278 64729 11320
rect 76343 11360 76390 11402
rect 76514 11360 76558 11402
rect 76682 11360 76729 11402
rect 76343 11320 76352 11360
rect 76514 11320 76516 11360
rect 76556 11320 76558 11360
rect 76720 11320 76729 11360
rect 76343 11278 76390 11320
rect 76514 11278 76558 11320
rect 76682 11278 76729 11320
rect 3103 10604 3150 10646
rect 3274 10604 3318 10646
rect 3442 10604 3489 10646
rect 3103 10564 3112 10604
rect 3274 10564 3276 10604
rect 3316 10564 3318 10604
rect 3480 10564 3489 10604
rect 3103 10522 3150 10564
rect 3274 10522 3318 10564
rect 3442 10522 3489 10564
rect 15103 10604 15150 10646
rect 15274 10604 15318 10646
rect 15442 10604 15489 10646
rect 15103 10564 15112 10604
rect 15274 10564 15276 10604
rect 15316 10564 15318 10604
rect 15480 10564 15489 10604
rect 15103 10522 15150 10564
rect 15274 10522 15318 10564
rect 15442 10522 15489 10564
rect 27103 10604 27150 10646
rect 27274 10604 27318 10646
rect 27442 10604 27489 10646
rect 27103 10564 27112 10604
rect 27274 10564 27276 10604
rect 27316 10564 27318 10604
rect 27480 10564 27489 10604
rect 27103 10522 27150 10564
rect 27274 10522 27318 10564
rect 27442 10522 27489 10564
rect 39103 10604 39150 10646
rect 39274 10604 39318 10646
rect 39442 10604 39489 10646
rect 39103 10564 39112 10604
rect 39274 10564 39276 10604
rect 39316 10564 39318 10604
rect 39480 10564 39489 10604
rect 39103 10522 39150 10564
rect 39274 10522 39318 10564
rect 39442 10522 39489 10564
rect 51103 10604 51150 10646
rect 51274 10604 51318 10646
rect 51442 10604 51489 10646
rect 51103 10564 51112 10604
rect 51274 10564 51276 10604
rect 51316 10564 51318 10604
rect 51480 10564 51489 10604
rect 51103 10522 51150 10564
rect 51274 10522 51318 10564
rect 51442 10522 51489 10564
rect 63103 10604 63150 10646
rect 63274 10604 63318 10646
rect 63442 10604 63489 10646
rect 63103 10564 63112 10604
rect 63274 10564 63276 10604
rect 63316 10564 63318 10604
rect 63480 10564 63489 10604
rect 63103 10522 63150 10564
rect 63274 10522 63318 10564
rect 63442 10522 63489 10564
rect 75103 10604 75150 10646
rect 75274 10604 75318 10646
rect 75442 10604 75489 10646
rect 75103 10564 75112 10604
rect 75274 10564 75276 10604
rect 75316 10564 75318 10604
rect 75480 10564 75489 10604
rect 75103 10522 75150 10564
rect 75274 10522 75318 10564
rect 75442 10522 75489 10564
rect 4343 9848 4390 9890
rect 4514 9848 4558 9890
rect 4682 9848 4729 9890
rect 4343 9808 4352 9848
rect 4514 9808 4516 9848
rect 4556 9808 4558 9848
rect 4720 9808 4729 9848
rect 4343 9766 4390 9808
rect 4514 9766 4558 9808
rect 4682 9766 4729 9808
rect 16343 9848 16390 9890
rect 16514 9848 16558 9890
rect 16682 9848 16729 9890
rect 16343 9808 16352 9848
rect 16514 9808 16516 9848
rect 16556 9808 16558 9848
rect 16720 9808 16729 9848
rect 16343 9766 16390 9808
rect 16514 9766 16558 9808
rect 16682 9766 16729 9808
rect 28343 9848 28390 9890
rect 28514 9848 28558 9890
rect 28682 9848 28729 9890
rect 28343 9808 28352 9848
rect 28514 9808 28516 9848
rect 28556 9808 28558 9848
rect 28720 9808 28729 9848
rect 28343 9766 28390 9808
rect 28514 9766 28558 9808
rect 28682 9766 28729 9808
rect 40343 9848 40390 9890
rect 40514 9848 40558 9890
rect 40682 9848 40729 9890
rect 40343 9808 40352 9848
rect 40514 9808 40516 9848
rect 40556 9808 40558 9848
rect 40720 9808 40729 9848
rect 40343 9766 40390 9808
rect 40514 9766 40558 9808
rect 40682 9766 40729 9808
rect 52343 9848 52390 9890
rect 52514 9848 52558 9890
rect 52682 9848 52729 9890
rect 52343 9808 52352 9848
rect 52514 9808 52516 9848
rect 52556 9808 52558 9848
rect 52720 9808 52729 9848
rect 52343 9766 52390 9808
rect 52514 9766 52558 9808
rect 52682 9766 52729 9808
rect 64343 9848 64390 9890
rect 64514 9848 64558 9890
rect 64682 9848 64729 9890
rect 64343 9808 64352 9848
rect 64514 9808 64516 9848
rect 64556 9808 64558 9848
rect 64720 9808 64729 9848
rect 64343 9766 64390 9808
rect 64514 9766 64558 9808
rect 64682 9766 64729 9808
rect 76343 9848 76390 9890
rect 76514 9848 76558 9890
rect 76682 9848 76729 9890
rect 76343 9808 76352 9848
rect 76514 9808 76516 9848
rect 76556 9808 76558 9848
rect 76720 9808 76729 9848
rect 76343 9766 76390 9808
rect 76514 9766 76558 9808
rect 76682 9766 76729 9808
rect 3103 9092 3150 9134
rect 3274 9092 3318 9134
rect 3442 9092 3489 9134
rect 3103 9052 3112 9092
rect 3274 9052 3276 9092
rect 3316 9052 3318 9092
rect 3480 9052 3489 9092
rect 3103 9010 3150 9052
rect 3274 9010 3318 9052
rect 3442 9010 3489 9052
rect 15103 9092 15150 9134
rect 15274 9092 15318 9134
rect 15442 9092 15489 9134
rect 15103 9052 15112 9092
rect 15274 9052 15276 9092
rect 15316 9052 15318 9092
rect 15480 9052 15489 9092
rect 15103 9010 15150 9052
rect 15274 9010 15318 9052
rect 15442 9010 15489 9052
rect 27103 9092 27150 9134
rect 27274 9092 27318 9134
rect 27442 9092 27489 9134
rect 27103 9052 27112 9092
rect 27274 9052 27276 9092
rect 27316 9052 27318 9092
rect 27480 9052 27489 9092
rect 27103 9010 27150 9052
rect 27274 9010 27318 9052
rect 27442 9010 27489 9052
rect 39103 9092 39150 9134
rect 39274 9092 39318 9134
rect 39442 9092 39489 9134
rect 39103 9052 39112 9092
rect 39274 9052 39276 9092
rect 39316 9052 39318 9092
rect 39480 9052 39489 9092
rect 39103 9010 39150 9052
rect 39274 9010 39318 9052
rect 39442 9010 39489 9052
rect 51103 9092 51150 9134
rect 51274 9092 51318 9134
rect 51442 9092 51489 9134
rect 51103 9052 51112 9092
rect 51274 9052 51276 9092
rect 51316 9052 51318 9092
rect 51480 9052 51489 9092
rect 51103 9010 51150 9052
rect 51274 9010 51318 9052
rect 51442 9010 51489 9052
rect 63103 9092 63150 9134
rect 63274 9092 63318 9134
rect 63442 9092 63489 9134
rect 63103 9052 63112 9092
rect 63274 9052 63276 9092
rect 63316 9052 63318 9092
rect 63480 9052 63489 9092
rect 63103 9010 63150 9052
rect 63274 9010 63318 9052
rect 63442 9010 63489 9052
rect 75103 9092 75150 9134
rect 75274 9092 75318 9134
rect 75442 9092 75489 9134
rect 75103 9052 75112 9092
rect 75274 9052 75276 9092
rect 75316 9052 75318 9092
rect 75480 9052 75489 9092
rect 75103 9010 75150 9052
rect 75274 9010 75318 9052
rect 75442 9010 75489 9052
rect 4343 8336 4390 8378
rect 4514 8336 4558 8378
rect 4682 8336 4729 8378
rect 4343 8296 4352 8336
rect 4514 8296 4516 8336
rect 4556 8296 4558 8336
rect 4720 8296 4729 8336
rect 4343 8254 4390 8296
rect 4514 8254 4558 8296
rect 4682 8254 4729 8296
rect 16343 8336 16390 8378
rect 16514 8336 16558 8378
rect 16682 8336 16729 8378
rect 16343 8296 16352 8336
rect 16514 8296 16516 8336
rect 16556 8296 16558 8336
rect 16720 8296 16729 8336
rect 16343 8254 16390 8296
rect 16514 8254 16558 8296
rect 16682 8254 16729 8296
rect 28343 8336 28390 8378
rect 28514 8336 28558 8378
rect 28682 8336 28729 8378
rect 28343 8296 28352 8336
rect 28514 8296 28516 8336
rect 28556 8296 28558 8336
rect 28720 8296 28729 8336
rect 28343 8254 28390 8296
rect 28514 8254 28558 8296
rect 28682 8254 28729 8296
rect 40343 8336 40390 8378
rect 40514 8336 40558 8378
rect 40682 8336 40729 8378
rect 40343 8296 40352 8336
rect 40514 8296 40516 8336
rect 40556 8296 40558 8336
rect 40720 8296 40729 8336
rect 40343 8254 40390 8296
rect 40514 8254 40558 8296
rect 40682 8254 40729 8296
rect 52343 8336 52390 8378
rect 52514 8336 52558 8378
rect 52682 8336 52729 8378
rect 52343 8296 52352 8336
rect 52514 8296 52516 8336
rect 52556 8296 52558 8336
rect 52720 8296 52729 8336
rect 52343 8254 52390 8296
rect 52514 8254 52558 8296
rect 52682 8254 52729 8296
rect 64343 8336 64390 8378
rect 64514 8336 64558 8378
rect 64682 8336 64729 8378
rect 64343 8296 64352 8336
rect 64514 8296 64516 8336
rect 64556 8296 64558 8336
rect 64720 8296 64729 8336
rect 64343 8254 64390 8296
rect 64514 8254 64558 8296
rect 64682 8254 64729 8296
rect 76343 8336 76390 8378
rect 76514 8336 76558 8378
rect 76682 8336 76729 8378
rect 76343 8296 76352 8336
rect 76514 8296 76516 8336
rect 76556 8296 76558 8336
rect 76720 8296 76729 8336
rect 76343 8254 76390 8296
rect 76514 8254 76558 8296
rect 76682 8254 76729 8296
rect 3103 7580 3150 7622
rect 3274 7580 3318 7622
rect 3442 7580 3489 7622
rect 3103 7540 3112 7580
rect 3274 7540 3276 7580
rect 3316 7540 3318 7580
rect 3480 7540 3489 7580
rect 3103 7498 3150 7540
rect 3274 7498 3318 7540
rect 3442 7498 3489 7540
rect 15103 7580 15150 7622
rect 15274 7580 15318 7622
rect 15442 7580 15489 7622
rect 15103 7540 15112 7580
rect 15274 7540 15276 7580
rect 15316 7540 15318 7580
rect 15480 7540 15489 7580
rect 15103 7498 15150 7540
rect 15274 7498 15318 7540
rect 15442 7498 15489 7540
rect 27103 7580 27150 7622
rect 27274 7580 27318 7622
rect 27442 7580 27489 7622
rect 27103 7540 27112 7580
rect 27274 7540 27276 7580
rect 27316 7540 27318 7580
rect 27480 7540 27489 7580
rect 27103 7498 27150 7540
rect 27274 7498 27318 7540
rect 27442 7498 27489 7540
rect 39103 7580 39150 7622
rect 39274 7580 39318 7622
rect 39442 7580 39489 7622
rect 39103 7540 39112 7580
rect 39274 7540 39276 7580
rect 39316 7540 39318 7580
rect 39480 7540 39489 7580
rect 39103 7498 39150 7540
rect 39274 7498 39318 7540
rect 39442 7498 39489 7540
rect 51103 7580 51150 7622
rect 51274 7580 51318 7622
rect 51442 7580 51489 7622
rect 51103 7540 51112 7580
rect 51274 7540 51276 7580
rect 51316 7540 51318 7580
rect 51480 7540 51489 7580
rect 51103 7498 51150 7540
rect 51274 7498 51318 7540
rect 51442 7498 51489 7540
rect 63103 7580 63150 7622
rect 63274 7580 63318 7622
rect 63442 7580 63489 7622
rect 63103 7540 63112 7580
rect 63274 7540 63276 7580
rect 63316 7540 63318 7580
rect 63480 7540 63489 7580
rect 63103 7498 63150 7540
rect 63274 7498 63318 7540
rect 63442 7498 63489 7540
rect 75103 7580 75150 7622
rect 75274 7580 75318 7622
rect 75442 7580 75489 7622
rect 75103 7540 75112 7580
rect 75274 7540 75276 7580
rect 75316 7540 75318 7580
rect 75480 7540 75489 7580
rect 75103 7498 75150 7540
rect 75274 7498 75318 7540
rect 75442 7498 75489 7540
rect 4343 6824 4390 6866
rect 4514 6824 4558 6866
rect 4682 6824 4729 6866
rect 4343 6784 4352 6824
rect 4514 6784 4516 6824
rect 4556 6784 4558 6824
rect 4720 6784 4729 6824
rect 4343 6742 4390 6784
rect 4514 6742 4558 6784
rect 4682 6742 4729 6784
rect 16343 6824 16390 6866
rect 16514 6824 16558 6866
rect 16682 6824 16729 6866
rect 16343 6784 16352 6824
rect 16514 6784 16516 6824
rect 16556 6784 16558 6824
rect 16720 6784 16729 6824
rect 16343 6742 16390 6784
rect 16514 6742 16558 6784
rect 16682 6742 16729 6784
rect 28343 6824 28390 6866
rect 28514 6824 28558 6866
rect 28682 6824 28729 6866
rect 28343 6784 28352 6824
rect 28514 6784 28516 6824
rect 28556 6784 28558 6824
rect 28720 6784 28729 6824
rect 28343 6742 28390 6784
rect 28514 6742 28558 6784
rect 28682 6742 28729 6784
rect 40343 6824 40390 6866
rect 40514 6824 40558 6866
rect 40682 6824 40729 6866
rect 40343 6784 40352 6824
rect 40514 6784 40516 6824
rect 40556 6784 40558 6824
rect 40720 6784 40729 6824
rect 40343 6742 40390 6784
rect 40514 6742 40558 6784
rect 40682 6742 40729 6784
rect 52343 6824 52390 6866
rect 52514 6824 52558 6866
rect 52682 6824 52729 6866
rect 52343 6784 52352 6824
rect 52514 6784 52516 6824
rect 52556 6784 52558 6824
rect 52720 6784 52729 6824
rect 52343 6742 52390 6784
rect 52514 6742 52558 6784
rect 52682 6742 52729 6784
rect 64343 6824 64390 6866
rect 64514 6824 64558 6866
rect 64682 6824 64729 6866
rect 64343 6784 64352 6824
rect 64514 6784 64516 6824
rect 64556 6784 64558 6824
rect 64720 6784 64729 6824
rect 64343 6742 64390 6784
rect 64514 6742 64558 6784
rect 64682 6742 64729 6784
rect 76343 6824 76390 6866
rect 76514 6824 76558 6866
rect 76682 6824 76729 6866
rect 76343 6784 76352 6824
rect 76514 6784 76516 6824
rect 76556 6784 76558 6824
rect 76720 6784 76729 6824
rect 76343 6742 76390 6784
rect 76514 6742 76558 6784
rect 76682 6742 76729 6784
rect 3103 6068 3150 6110
rect 3274 6068 3318 6110
rect 3442 6068 3489 6110
rect 3103 6028 3112 6068
rect 3274 6028 3276 6068
rect 3316 6028 3318 6068
rect 3480 6028 3489 6068
rect 3103 5986 3150 6028
rect 3274 5986 3318 6028
rect 3442 5986 3489 6028
rect 15103 6068 15150 6110
rect 15274 6068 15318 6110
rect 15442 6068 15489 6110
rect 15103 6028 15112 6068
rect 15274 6028 15276 6068
rect 15316 6028 15318 6068
rect 15480 6028 15489 6068
rect 15103 5986 15150 6028
rect 15274 5986 15318 6028
rect 15442 5986 15489 6028
rect 27103 6068 27150 6110
rect 27274 6068 27318 6110
rect 27442 6068 27489 6110
rect 27103 6028 27112 6068
rect 27274 6028 27276 6068
rect 27316 6028 27318 6068
rect 27480 6028 27489 6068
rect 27103 5986 27150 6028
rect 27274 5986 27318 6028
rect 27442 5986 27489 6028
rect 39103 6068 39150 6110
rect 39274 6068 39318 6110
rect 39442 6068 39489 6110
rect 39103 6028 39112 6068
rect 39274 6028 39276 6068
rect 39316 6028 39318 6068
rect 39480 6028 39489 6068
rect 39103 5986 39150 6028
rect 39274 5986 39318 6028
rect 39442 5986 39489 6028
rect 51103 6068 51150 6110
rect 51274 6068 51318 6110
rect 51442 6068 51489 6110
rect 51103 6028 51112 6068
rect 51274 6028 51276 6068
rect 51316 6028 51318 6068
rect 51480 6028 51489 6068
rect 51103 5986 51150 6028
rect 51274 5986 51318 6028
rect 51442 5986 51489 6028
rect 63103 6068 63150 6110
rect 63274 6068 63318 6110
rect 63442 6068 63489 6110
rect 63103 6028 63112 6068
rect 63274 6028 63276 6068
rect 63316 6028 63318 6068
rect 63480 6028 63489 6068
rect 63103 5986 63150 6028
rect 63274 5986 63318 6028
rect 63442 5986 63489 6028
rect 75103 6068 75150 6110
rect 75274 6068 75318 6110
rect 75442 6068 75489 6110
rect 75103 6028 75112 6068
rect 75274 6028 75276 6068
rect 75316 6028 75318 6068
rect 75480 6028 75489 6068
rect 75103 5986 75150 6028
rect 75274 5986 75318 6028
rect 75442 5986 75489 6028
rect 4343 5312 4390 5354
rect 4514 5312 4558 5354
rect 4682 5312 4729 5354
rect 4343 5272 4352 5312
rect 4514 5272 4516 5312
rect 4556 5272 4558 5312
rect 4720 5272 4729 5312
rect 4343 5230 4390 5272
rect 4514 5230 4558 5272
rect 4682 5230 4729 5272
rect 16343 5312 16390 5354
rect 16514 5312 16558 5354
rect 16682 5312 16729 5354
rect 16343 5272 16352 5312
rect 16514 5272 16516 5312
rect 16556 5272 16558 5312
rect 16720 5272 16729 5312
rect 16343 5230 16390 5272
rect 16514 5230 16558 5272
rect 16682 5230 16729 5272
rect 28343 5312 28390 5354
rect 28514 5312 28558 5354
rect 28682 5312 28729 5354
rect 28343 5272 28352 5312
rect 28514 5272 28516 5312
rect 28556 5272 28558 5312
rect 28720 5272 28729 5312
rect 28343 5230 28390 5272
rect 28514 5230 28558 5272
rect 28682 5230 28729 5272
rect 40343 5312 40390 5354
rect 40514 5312 40558 5354
rect 40682 5312 40729 5354
rect 40343 5272 40352 5312
rect 40514 5272 40516 5312
rect 40556 5272 40558 5312
rect 40720 5272 40729 5312
rect 40343 5230 40390 5272
rect 40514 5230 40558 5272
rect 40682 5230 40729 5272
rect 52343 5312 52390 5354
rect 52514 5312 52558 5354
rect 52682 5312 52729 5354
rect 52343 5272 52352 5312
rect 52514 5272 52516 5312
rect 52556 5272 52558 5312
rect 52720 5272 52729 5312
rect 52343 5230 52390 5272
rect 52514 5230 52558 5272
rect 52682 5230 52729 5272
rect 64343 5312 64390 5354
rect 64514 5312 64558 5354
rect 64682 5312 64729 5354
rect 64343 5272 64352 5312
rect 64514 5272 64516 5312
rect 64556 5272 64558 5312
rect 64720 5272 64729 5312
rect 64343 5230 64390 5272
rect 64514 5230 64558 5272
rect 64682 5230 64729 5272
rect 76343 5312 76390 5354
rect 76514 5312 76558 5354
rect 76682 5312 76729 5354
rect 76343 5272 76352 5312
rect 76514 5272 76516 5312
rect 76556 5272 76558 5312
rect 76720 5272 76729 5312
rect 76343 5230 76390 5272
rect 76514 5230 76558 5272
rect 76682 5230 76729 5272
rect 3103 4556 3150 4598
rect 3274 4556 3318 4598
rect 3442 4556 3489 4598
rect 3103 4516 3112 4556
rect 3274 4516 3276 4556
rect 3316 4516 3318 4556
rect 3480 4516 3489 4556
rect 3103 4474 3150 4516
rect 3274 4474 3318 4516
rect 3442 4474 3489 4516
rect 15103 4556 15150 4598
rect 15274 4556 15318 4598
rect 15442 4556 15489 4598
rect 15103 4516 15112 4556
rect 15274 4516 15276 4556
rect 15316 4516 15318 4556
rect 15480 4516 15489 4556
rect 15103 4474 15150 4516
rect 15274 4474 15318 4516
rect 15442 4474 15489 4516
rect 27103 4556 27150 4598
rect 27274 4556 27318 4598
rect 27442 4556 27489 4598
rect 27103 4516 27112 4556
rect 27274 4516 27276 4556
rect 27316 4516 27318 4556
rect 27480 4516 27489 4556
rect 27103 4474 27150 4516
rect 27274 4474 27318 4516
rect 27442 4474 27489 4516
rect 39103 4556 39150 4598
rect 39274 4556 39318 4598
rect 39442 4556 39489 4598
rect 39103 4516 39112 4556
rect 39274 4516 39276 4556
rect 39316 4516 39318 4556
rect 39480 4516 39489 4556
rect 39103 4474 39150 4516
rect 39274 4474 39318 4516
rect 39442 4474 39489 4516
rect 51103 4556 51150 4598
rect 51274 4556 51318 4598
rect 51442 4556 51489 4598
rect 51103 4516 51112 4556
rect 51274 4516 51276 4556
rect 51316 4516 51318 4556
rect 51480 4516 51489 4556
rect 51103 4474 51150 4516
rect 51274 4474 51318 4516
rect 51442 4474 51489 4516
rect 63103 4556 63150 4598
rect 63274 4556 63318 4598
rect 63442 4556 63489 4598
rect 63103 4516 63112 4556
rect 63274 4516 63276 4556
rect 63316 4516 63318 4556
rect 63480 4516 63489 4556
rect 63103 4474 63150 4516
rect 63274 4474 63318 4516
rect 63442 4474 63489 4516
rect 75103 4556 75150 4598
rect 75274 4556 75318 4598
rect 75442 4556 75489 4598
rect 75103 4516 75112 4556
rect 75274 4516 75276 4556
rect 75316 4516 75318 4556
rect 75480 4516 75489 4556
rect 75103 4474 75150 4516
rect 75274 4474 75318 4516
rect 75442 4474 75489 4516
rect 4343 3800 4390 3842
rect 4514 3800 4558 3842
rect 4682 3800 4729 3842
rect 4343 3760 4352 3800
rect 4514 3760 4516 3800
rect 4556 3760 4558 3800
rect 4720 3760 4729 3800
rect 4343 3718 4390 3760
rect 4514 3718 4558 3760
rect 4682 3718 4729 3760
rect 16343 3800 16390 3842
rect 16514 3800 16558 3842
rect 16682 3800 16729 3842
rect 16343 3760 16352 3800
rect 16514 3760 16516 3800
rect 16556 3760 16558 3800
rect 16720 3760 16729 3800
rect 16343 3718 16390 3760
rect 16514 3718 16558 3760
rect 16682 3718 16729 3760
rect 28343 3800 28390 3842
rect 28514 3800 28558 3842
rect 28682 3800 28729 3842
rect 28343 3760 28352 3800
rect 28514 3760 28516 3800
rect 28556 3760 28558 3800
rect 28720 3760 28729 3800
rect 28343 3718 28390 3760
rect 28514 3718 28558 3760
rect 28682 3718 28729 3760
rect 40343 3800 40390 3842
rect 40514 3800 40558 3842
rect 40682 3800 40729 3842
rect 40343 3760 40352 3800
rect 40514 3760 40516 3800
rect 40556 3760 40558 3800
rect 40720 3760 40729 3800
rect 40343 3718 40390 3760
rect 40514 3718 40558 3760
rect 40682 3718 40729 3760
rect 52343 3800 52390 3842
rect 52514 3800 52558 3842
rect 52682 3800 52729 3842
rect 52343 3760 52352 3800
rect 52514 3760 52516 3800
rect 52556 3760 52558 3800
rect 52720 3760 52729 3800
rect 52343 3718 52390 3760
rect 52514 3718 52558 3760
rect 52682 3718 52729 3760
rect 64343 3800 64390 3842
rect 64514 3800 64558 3842
rect 64682 3800 64729 3842
rect 64343 3760 64352 3800
rect 64514 3760 64516 3800
rect 64556 3760 64558 3800
rect 64720 3760 64729 3800
rect 64343 3718 64390 3760
rect 64514 3718 64558 3760
rect 64682 3718 64729 3760
rect 76343 3800 76390 3842
rect 76514 3800 76558 3842
rect 76682 3800 76729 3842
rect 76343 3760 76352 3800
rect 76514 3760 76516 3800
rect 76556 3760 76558 3800
rect 76720 3760 76729 3800
rect 76343 3718 76390 3760
rect 76514 3718 76558 3760
rect 76682 3718 76729 3760
rect 3103 3044 3150 3086
rect 3274 3044 3318 3086
rect 3442 3044 3489 3086
rect 3103 3004 3112 3044
rect 3274 3004 3276 3044
rect 3316 3004 3318 3044
rect 3480 3004 3489 3044
rect 3103 2962 3150 3004
rect 3274 2962 3318 3004
rect 3442 2962 3489 3004
rect 15103 3044 15150 3086
rect 15274 3044 15318 3086
rect 15442 3044 15489 3086
rect 15103 3004 15112 3044
rect 15274 3004 15276 3044
rect 15316 3004 15318 3044
rect 15480 3004 15489 3044
rect 15103 2962 15150 3004
rect 15274 2962 15318 3004
rect 15442 2962 15489 3004
rect 27103 3044 27150 3086
rect 27274 3044 27318 3086
rect 27442 3044 27489 3086
rect 27103 3004 27112 3044
rect 27274 3004 27276 3044
rect 27316 3004 27318 3044
rect 27480 3004 27489 3044
rect 27103 2962 27150 3004
rect 27274 2962 27318 3004
rect 27442 2962 27489 3004
rect 39103 3044 39150 3086
rect 39274 3044 39318 3086
rect 39442 3044 39489 3086
rect 39103 3004 39112 3044
rect 39274 3004 39276 3044
rect 39316 3004 39318 3044
rect 39480 3004 39489 3044
rect 39103 2962 39150 3004
rect 39274 2962 39318 3004
rect 39442 2962 39489 3004
rect 51103 3044 51150 3086
rect 51274 3044 51318 3086
rect 51442 3044 51489 3086
rect 51103 3004 51112 3044
rect 51274 3004 51276 3044
rect 51316 3004 51318 3044
rect 51480 3004 51489 3044
rect 51103 2962 51150 3004
rect 51274 2962 51318 3004
rect 51442 2962 51489 3004
rect 63103 3044 63150 3086
rect 63274 3044 63318 3086
rect 63442 3044 63489 3086
rect 63103 3004 63112 3044
rect 63274 3004 63276 3044
rect 63316 3004 63318 3044
rect 63480 3004 63489 3044
rect 63103 2962 63150 3004
rect 63274 2962 63318 3004
rect 63442 2962 63489 3004
rect 75103 3044 75150 3086
rect 75274 3044 75318 3086
rect 75442 3044 75489 3086
rect 75103 3004 75112 3044
rect 75274 3004 75276 3044
rect 75316 3004 75318 3044
rect 75480 3004 75489 3044
rect 75103 2962 75150 3004
rect 75274 2962 75318 3004
rect 75442 2962 75489 3004
rect 4343 2288 4390 2330
rect 4514 2288 4558 2330
rect 4682 2288 4729 2330
rect 4343 2248 4352 2288
rect 4514 2248 4516 2288
rect 4556 2248 4558 2288
rect 4720 2248 4729 2288
rect 4343 2206 4390 2248
rect 4514 2206 4558 2248
rect 4682 2206 4729 2248
rect 16343 2288 16390 2330
rect 16514 2288 16558 2330
rect 16682 2288 16729 2330
rect 16343 2248 16352 2288
rect 16514 2248 16516 2288
rect 16556 2248 16558 2288
rect 16720 2248 16729 2288
rect 16343 2206 16390 2248
rect 16514 2206 16558 2248
rect 16682 2206 16729 2248
rect 28343 2288 28390 2330
rect 28514 2288 28558 2330
rect 28682 2288 28729 2330
rect 28343 2248 28352 2288
rect 28514 2248 28516 2288
rect 28556 2248 28558 2288
rect 28720 2248 28729 2288
rect 28343 2206 28390 2248
rect 28514 2206 28558 2248
rect 28682 2206 28729 2248
rect 40343 2288 40390 2330
rect 40514 2288 40558 2330
rect 40682 2288 40729 2330
rect 40343 2248 40352 2288
rect 40514 2248 40516 2288
rect 40556 2248 40558 2288
rect 40720 2248 40729 2288
rect 40343 2206 40390 2248
rect 40514 2206 40558 2248
rect 40682 2206 40729 2248
rect 52343 2288 52390 2330
rect 52514 2288 52558 2330
rect 52682 2288 52729 2330
rect 52343 2248 52352 2288
rect 52514 2248 52516 2288
rect 52556 2248 52558 2288
rect 52720 2248 52729 2288
rect 52343 2206 52390 2248
rect 52514 2206 52558 2248
rect 52682 2206 52729 2248
rect 64343 2288 64390 2330
rect 64514 2288 64558 2330
rect 64682 2288 64729 2330
rect 64343 2248 64352 2288
rect 64514 2248 64516 2288
rect 64556 2248 64558 2288
rect 64720 2248 64729 2288
rect 64343 2206 64390 2248
rect 64514 2206 64558 2248
rect 64682 2206 64729 2248
rect 76343 2288 76390 2330
rect 76514 2288 76558 2330
rect 76682 2288 76729 2330
rect 76343 2248 76352 2288
rect 76514 2248 76516 2288
rect 76556 2248 76558 2288
rect 76720 2248 76729 2288
rect 76343 2206 76390 2248
rect 76514 2206 76558 2248
rect 76682 2206 76729 2248
rect 3103 1532 3150 1574
rect 3274 1532 3318 1574
rect 3442 1532 3489 1574
rect 3103 1492 3112 1532
rect 3274 1492 3276 1532
rect 3316 1492 3318 1532
rect 3480 1492 3489 1532
rect 3103 1450 3150 1492
rect 3274 1450 3318 1492
rect 3442 1450 3489 1492
rect 15103 1532 15150 1574
rect 15274 1532 15318 1574
rect 15442 1532 15489 1574
rect 15103 1492 15112 1532
rect 15274 1492 15276 1532
rect 15316 1492 15318 1532
rect 15480 1492 15489 1532
rect 15103 1450 15150 1492
rect 15274 1450 15318 1492
rect 15442 1450 15489 1492
rect 27103 1532 27150 1574
rect 27274 1532 27318 1574
rect 27442 1532 27489 1574
rect 27103 1492 27112 1532
rect 27274 1492 27276 1532
rect 27316 1492 27318 1532
rect 27480 1492 27489 1532
rect 27103 1450 27150 1492
rect 27274 1450 27318 1492
rect 27442 1450 27489 1492
rect 39103 1532 39150 1574
rect 39274 1532 39318 1574
rect 39442 1532 39489 1574
rect 39103 1492 39112 1532
rect 39274 1492 39276 1532
rect 39316 1492 39318 1532
rect 39480 1492 39489 1532
rect 39103 1450 39150 1492
rect 39274 1450 39318 1492
rect 39442 1450 39489 1492
rect 51103 1532 51150 1574
rect 51274 1532 51318 1574
rect 51442 1532 51489 1574
rect 51103 1492 51112 1532
rect 51274 1492 51276 1532
rect 51316 1492 51318 1532
rect 51480 1492 51489 1532
rect 51103 1450 51150 1492
rect 51274 1450 51318 1492
rect 51442 1450 51489 1492
rect 63103 1532 63150 1574
rect 63274 1532 63318 1574
rect 63442 1532 63489 1574
rect 63103 1492 63112 1532
rect 63274 1492 63276 1532
rect 63316 1492 63318 1532
rect 63480 1492 63489 1532
rect 63103 1450 63150 1492
rect 63274 1450 63318 1492
rect 63442 1450 63489 1492
rect 75103 1532 75150 1574
rect 75274 1532 75318 1574
rect 75442 1532 75489 1574
rect 75103 1492 75112 1532
rect 75274 1492 75276 1532
rect 75316 1492 75318 1532
rect 75480 1492 75489 1532
rect 75103 1450 75150 1492
rect 75274 1450 75318 1492
rect 75442 1450 75489 1492
rect 4343 776 4390 818
rect 4514 776 4558 818
rect 4682 776 4729 818
rect 4343 736 4352 776
rect 4514 736 4516 776
rect 4556 736 4558 776
rect 4720 736 4729 776
rect 4343 694 4390 736
rect 4514 694 4558 736
rect 4682 694 4729 736
rect 16343 776 16390 818
rect 16514 776 16558 818
rect 16682 776 16729 818
rect 16343 736 16352 776
rect 16514 736 16516 776
rect 16556 736 16558 776
rect 16720 736 16729 776
rect 16343 694 16390 736
rect 16514 694 16558 736
rect 16682 694 16729 736
rect 28343 776 28390 818
rect 28514 776 28558 818
rect 28682 776 28729 818
rect 28343 736 28352 776
rect 28514 736 28516 776
rect 28556 736 28558 776
rect 28720 736 28729 776
rect 28343 694 28390 736
rect 28514 694 28558 736
rect 28682 694 28729 736
rect 40343 776 40390 818
rect 40514 776 40558 818
rect 40682 776 40729 818
rect 40343 736 40352 776
rect 40514 736 40516 776
rect 40556 736 40558 776
rect 40720 736 40729 776
rect 40343 694 40390 736
rect 40514 694 40558 736
rect 40682 694 40729 736
rect 52343 776 52390 818
rect 52514 776 52558 818
rect 52682 776 52729 818
rect 52343 736 52352 776
rect 52514 736 52516 776
rect 52556 736 52558 776
rect 52720 736 52729 776
rect 52343 694 52390 736
rect 52514 694 52558 736
rect 52682 694 52729 736
rect 64343 776 64390 818
rect 64514 776 64558 818
rect 64682 776 64729 818
rect 64343 736 64352 776
rect 64514 736 64516 776
rect 64556 736 64558 776
rect 64720 736 64729 776
rect 64343 694 64390 736
rect 64514 694 64558 736
rect 64682 694 64729 736
rect 76343 776 76390 818
rect 76514 776 76558 818
rect 76682 776 76729 818
rect 76343 736 76352 776
rect 76514 736 76516 776
rect 76556 736 76558 776
rect 76720 736 76729 776
rect 76343 694 76390 736
rect 76514 694 76558 736
rect 76682 694 76729 736
<< via5 >>
rect 4390 38576 4514 38618
rect 4558 38576 4682 38618
rect 4390 38536 4392 38576
rect 4392 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4514 38576
rect 4558 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4680 38576
rect 4680 38536 4682 38576
rect 4390 38494 4514 38536
rect 4558 38494 4682 38536
rect 16390 38576 16514 38618
rect 16558 38576 16682 38618
rect 16390 38536 16392 38576
rect 16392 38536 16434 38576
rect 16434 38536 16474 38576
rect 16474 38536 16514 38576
rect 16558 38536 16598 38576
rect 16598 38536 16638 38576
rect 16638 38536 16680 38576
rect 16680 38536 16682 38576
rect 16390 38494 16514 38536
rect 16558 38494 16682 38536
rect 28390 38576 28514 38618
rect 28558 38576 28682 38618
rect 28390 38536 28392 38576
rect 28392 38536 28434 38576
rect 28434 38536 28474 38576
rect 28474 38536 28514 38576
rect 28558 38536 28598 38576
rect 28598 38536 28638 38576
rect 28638 38536 28680 38576
rect 28680 38536 28682 38576
rect 28390 38494 28514 38536
rect 28558 38494 28682 38536
rect 40390 38576 40514 38618
rect 40558 38576 40682 38618
rect 40390 38536 40392 38576
rect 40392 38536 40434 38576
rect 40434 38536 40474 38576
rect 40474 38536 40514 38576
rect 40558 38536 40598 38576
rect 40598 38536 40638 38576
rect 40638 38536 40680 38576
rect 40680 38536 40682 38576
rect 40390 38494 40514 38536
rect 40558 38494 40682 38536
rect 52390 38576 52514 38618
rect 52558 38576 52682 38618
rect 52390 38536 52392 38576
rect 52392 38536 52434 38576
rect 52434 38536 52474 38576
rect 52474 38536 52514 38576
rect 52558 38536 52598 38576
rect 52598 38536 52638 38576
rect 52638 38536 52680 38576
rect 52680 38536 52682 38576
rect 52390 38494 52514 38536
rect 52558 38494 52682 38536
rect 64390 38576 64514 38618
rect 64558 38576 64682 38618
rect 64390 38536 64392 38576
rect 64392 38536 64434 38576
rect 64434 38536 64474 38576
rect 64474 38536 64514 38576
rect 64558 38536 64598 38576
rect 64598 38536 64638 38576
rect 64638 38536 64680 38576
rect 64680 38536 64682 38576
rect 64390 38494 64514 38536
rect 64558 38494 64682 38536
rect 76390 38576 76514 38618
rect 76558 38576 76682 38618
rect 76390 38536 76392 38576
rect 76392 38536 76434 38576
rect 76434 38536 76474 38576
rect 76474 38536 76514 38576
rect 76558 38536 76598 38576
rect 76598 38536 76638 38576
rect 76638 38536 76680 38576
rect 76680 38536 76682 38576
rect 76390 38494 76514 38536
rect 76558 38494 76682 38536
rect 3150 37820 3274 37862
rect 3318 37820 3442 37862
rect 3150 37780 3152 37820
rect 3152 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3274 37820
rect 3318 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3440 37820
rect 3440 37780 3442 37820
rect 3150 37738 3274 37780
rect 3318 37738 3442 37780
rect 15150 37820 15274 37862
rect 15318 37820 15442 37862
rect 15150 37780 15152 37820
rect 15152 37780 15194 37820
rect 15194 37780 15234 37820
rect 15234 37780 15274 37820
rect 15318 37780 15358 37820
rect 15358 37780 15398 37820
rect 15398 37780 15440 37820
rect 15440 37780 15442 37820
rect 15150 37738 15274 37780
rect 15318 37738 15442 37780
rect 27150 37820 27274 37862
rect 27318 37820 27442 37862
rect 27150 37780 27152 37820
rect 27152 37780 27194 37820
rect 27194 37780 27234 37820
rect 27234 37780 27274 37820
rect 27318 37780 27358 37820
rect 27358 37780 27398 37820
rect 27398 37780 27440 37820
rect 27440 37780 27442 37820
rect 27150 37738 27274 37780
rect 27318 37738 27442 37780
rect 39150 37820 39274 37862
rect 39318 37820 39442 37862
rect 39150 37780 39152 37820
rect 39152 37780 39194 37820
rect 39194 37780 39234 37820
rect 39234 37780 39274 37820
rect 39318 37780 39358 37820
rect 39358 37780 39398 37820
rect 39398 37780 39440 37820
rect 39440 37780 39442 37820
rect 39150 37738 39274 37780
rect 39318 37738 39442 37780
rect 51150 37820 51274 37862
rect 51318 37820 51442 37862
rect 51150 37780 51152 37820
rect 51152 37780 51194 37820
rect 51194 37780 51234 37820
rect 51234 37780 51274 37820
rect 51318 37780 51358 37820
rect 51358 37780 51398 37820
rect 51398 37780 51440 37820
rect 51440 37780 51442 37820
rect 51150 37738 51274 37780
rect 51318 37738 51442 37780
rect 63150 37820 63274 37862
rect 63318 37820 63442 37862
rect 63150 37780 63152 37820
rect 63152 37780 63194 37820
rect 63194 37780 63234 37820
rect 63234 37780 63274 37820
rect 63318 37780 63358 37820
rect 63358 37780 63398 37820
rect 63398 37780 63440 37820
rect 63440 37780 63442 37820
rect 63150 37738 63274 37780
rect 63318 37738 63442 37780
rect 75150 37820 75274 37862
rect 75318 37820 75442 37862
rect 75150 37780 75152 37820
rect 75152 37780 75194 37820
rect 75194 37780 75234 37820
rect 75234 37780 75274 37820
rect 75318 37780 75358 37820
rect 75358 37780 75398 37820
rect 75398 37780 75440 37820
rect 75440 37780 75442 37820
rect 75150 37738 75274 37780
rect 75318 37738 75442 37780
rect 4390 37064 4514 37106
rect 4558 37064 4682 37106
rect 4390 37024 4392 37064
rect 4392 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4514 37064
rect 4558 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4680 37064
rect 4680 37024 4682 37064
rect 4390 36982 4514 37024
rect 4558 36982 4682 37024
rect 16390 37064 16514 37106
rect 16558 37064 16682 37106
rect 16390 37024 16392 37064
rect 16392 37024 16434 37064
rect 16434 37024 16474 37064
rect 16474 37024 16514 37064
rect 16558 37024 16598 37064
rect 16598 37024 16638 37064
rect 16638 37024 16680 37064
rect 16680 37024 16682 37064
rect 16390 36982 16514 37024
rect 16558 36982 16682 37024
rect 28390 37064 28514 37106
rect 28558 37064 28682 37106
rect 28390 37024 28392 37064
rect 28392 37024 28434 37064
rect 28434 37024 28474 37064
rect 28474 37024 28514 37064
rect 28558 37024 28598 37064
rect 28598 37024 28638 37064
rect 28638 37024 28680 37064
rect 28680 37024 28682 37064
rect 28390 36982 28514 37024
rect 28558 36982 28682 37024
rect 40390 37064 40514 37106
rect 40558 37064 40682 37106
rect 40390 37024 40392 37064
rect 40392 37024 40434 37064
rect 40434 37024 40474 37064
rect 40474 37024 40514 37064
rect 40558 37024 40598 37064
rect 40598 37024 40638 37064
rect 40638 37024 40680 37064
rect 40680 37024 40682 37064
rect 40390 36982 40514 37024
rect 40558 36982 40682 37024
rect 52390 37064 52514 37106
rect 52558 37064 52682 37106
rect 52390 37024 52392 37064
rect 52392 37024 52434 37064
rect 52434 37024 52474 37064
rect 52474 37024 52514 37064
rect 52558 37024 52598 37064
rect 52598 37024 52638 37064
rect 52638 37024 52680 37064
rect 52680 37024 52682 37064
rect 52390 36982 52514 37024
rect 52558 36982 52682 37024
rect 64390 37064 64514 37106
rect 64558 37064 64682 37106
rect 64390 37024 64392 37064
rect 64392 37024 64434 37064
rect 64434 37024 64474 37064
rect 64474 37024 64514 37064
rect 64558 37024 64598 37064
rect 64598 37024 64638 37064
rect 64638 37024 64680 37064
rect 64680 37024 64682 37064
rect 64390 36982 64514 37024
rect 64558 36982 64682 37024
rect 76390 37064 76514 37106
rect 76558 37064 76682 37106
rect 76390 37024 76392 37064
rect 76392 37024 76434 37064
rect 76434 37024 76474 37064
rect 76474 37024 76514 37064
rect 76558 37024 76598 37064
rect 76598 37024 76638 37064
rect 76638 37024 76680 37064
rect 76680 37024 76682 37064
rect 76390 36982 76514 37024
rect 76558 36982 76682 37024
rect 3150 36308 3274 36350
rect 3318 36308 3442 36350
rect 3150 36268 3152 36308
rect 3152 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3274 36308
rect 3318 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3440 36308
rect 3440 36268 3442 36308
rect 3150 36226 3274 36268
rect 3318 36226 3442 36268
rect 15150 36308 15274 36350
rect 15318 36308 15442 36350
rect 15150 36268 15152 36308
rect 15152 36268 15194 36308
rect 15194 36268 15234 36308
rect 15234 36268 15274 36308
rect 15318 36268 15358 36308
rect 15358 36268 15398 36308
rect 15398 36268 15440 36308
rect 15440 36268 15442 36308
rect 15150 36226 15274 36268
rect 15318 36226 15442 36268
rect 27150 36308 27274 36350
rect 27318 36308 27442 36350
rect 27150 36268 27152 36308
rect 27152 36268 27194 36308
rect 27194 36268 27234 36308
rect 27234 36268 27274 36308
rect 27318 36268 27358 36308
rect 27358 36268 27398 36308
rect 27398 36268 27440 36308
rect 27440 36268 27442 36308
rect 27150 36226 27274 36268
rect 27318 36226 27442 36268
rect 39150 36308 39274 36350
rect 39318 36308 39442 36350
rect 39150 36268 39152 36308
rect 39152 36268 39194 36308
rect 39194 36268 39234 36308
rect 39234 36268 39274 36308
rect 39318 36268 39358 36308
rect 39358 36268 39398 36308
rect 39398 36268 39440 36308
rect 39440 36268 39442 36308
rect 39150 36226 39274 36268
rect 39318 36226 39442 36268
rect 51150 36308 51274 36350
rect 51318 36308 51442 36350
rect 51150 36268 51152 36308
rect 51152 36268 51194 36308
rect 51194 36268 51234 36308
rect 51234 36268 51274 36308
rect 51318 36268 51358 36308
rect 51358 36268 51398 36308
rect 51398 36268 51440 36308
rect 51440 36268 51442 36308
rect 51150 36226 51274 36268
rect 51318 36226 51442 36268
rect 63150 36308 63274 36350
rect 63318 36308 63442 36350
rect 63150 36268 63152 36308
rect 63152 36268 63194 36308
rect 63194 36268 63234 36308
rect 63234 36268 63274 36308
rect 63318 36268 63358 36308
rect 63358 36268 63398 36308
rect 63398 36268 63440 36308
rect 63440 36268 63442 36308
rect 63150 36226 63274 36268
rect 63318 36226 63442 36268
rect 75150 36308 75274 36350
rect 75318 36308 75442 36350
rect 75150 36268 75152 36308
rect 75152 36268 75194 36308
rect 75194 36268 75234 36308
rect 75234 36268 75274 36308
rect 75318 36268 75358 36308
rect 75358 36268 75398 36308
rect 75398 36268 75440 36308
rect 75440 36268 75442 36308
rect 75150 36226 75274 36268
rect 75318 36226 75442 36268
rect 4390 35552 4514 35594
rect 4558 35552 4682 35594
rect 4390 35512 4392 35552
rect 4392 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4514 35552
rect 4558 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4680 35552
rect 4680 35512 4682 35552
rect 4390 35470 4514 35512
rect 4558 35470 4682 35512
rect 16390 35552 16514 35594
rect 16558 35552 16682 35594
rect 16390 35512 16392 35552
rect 16392 35512 16434 35552
rect 16434 35512 16474 35552
rect 16474 35512 16514 35552
rect 16558 35512 16598 35552
rect 16598 35512 16638 35552
rect 16638 35512 16680 35552
rect 16680 35512 16682 35552
rect 16390 35470 16514 35512
rect 16558 35470 16682 35512
rect 28390 35552 28514 35594
rect 28558 35552 28682 35594
rect 28390 35512 28392 35552
rect 28392 35512 28434 35552
rect 28434 35512 28474 35552
rect 28474 35512 28514 35552
rect 28558 35512 28598 35552
rect 28598 35512 28638 35552
rect 28638 35512 28680 35552
rect 28680 35512 28682 35552
rect 28390 35470 28514 35512
rect 28558 35470 28682 35512
rect 40390 35552 40514 35594
rect 40558 35552 40682 35594
rect 40390 35512 40392 35552
rect 40392 35512 40434 35552
rect 40434 35512 40474 35552
rect 40474 35512 40514 35552
rect 40558 35512 40598 35552
rect 40598 35512 40638 35552
rect 40638 35512 40680 35552
rect 40680 35512 40682 35552
rect 40390 35470 40514 35512
rect 40558 35470 40682 35512
rect 52390 35552 52514 35594
rect 52558 35552 52682 35594
rect 52390 35512 52392 35552
rect 52392 35512 52434 35552
rect 52434 35512 52474 35552
rect 52474 35512 52514 35552
rect 52558 35512 52598 35552
rect 52598 35512 52638 35552
rect 52638 35512 52680 35552
rect 52680 35512 52682 35552
rect 52390 35470 52514 35512
rect 52558 35470 52682 35512
rect 64390 35552 64514 35594
rect 64558 35552 64682 35594
rect 64390 35512 64392 35552
rect 64392 35512 64434 35552
rect 64434 35512 64474 35552
rect 64474 35512 64514 35552
rect 64558 35512 64598 35552
rect 64598 35512 64638 35552
rect 64638 35512 64680 35552
rect 64680 35512 64682 35552
rect 64390 35470 64514 35512
rect 64558 35470 64682 35512
rect 76390 35552 76514 35594
rect 76558 35552 76682 35594
rect 76390 35512 76392 35552
rect 76392 35512 76434 35552
rect 76434 35512 76474 35552
rect 76474 35512 76514 35552
rect 76558 35512 76598 35552
rect 76598 35512 76638 35552
rect 76638 35512 76680 35552
rect 76680 35512 76682 35552
rect 76390 35470 76514 35512
rect 76558 35470 76682 35512
rect 3150 34796 3274 34838
rect 3318 34796 3442 34838
rect 3150 34756 3152 34796
rect 3152 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3274 34796
rect 3318 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3440 34796
rect 3440 34756 3442 34796
rect 3150 34714 3274 34756
rect 3318 34714 3442 34756
rect 15150 34796 15274 34838
rect 15318 34796 15442 34838
rect 15150 34756 15152 34796
rect 15152 34756 15194 34796
rect 15194 34756 15234 34796
rect 15234 34756 15274 34796
rect 15318 34756 15358 34796
rect 15358 34756 15398 34796
rect 15398 34756 15440 34796
rect 15440 34756 15442 34796
rect 15150 34714 15274 34756
rect 15318 34714 15442 34756
rect 27150 34796 27274 34838
rect 27318 34796 27442 34838
rect 27150 34756 27152 34796
rect 27152 34756 27194 34796
rect 27194 34756 27234 34796
rect 27234 34756 27274 34796
rect 27318 34756 27358 34796
rect 27358 34756 27398 34796
rect 27398 34756 27440 34796
rect 27440 34756 27442 34796
rect 27150 34714 27274 34756
rect 27318 34714 27442 34756
rect 39150 34796 39274 34838
rect 39318 34796 39442 34838
rect 39150 34756 39152 34796
rect 39152 34756 39194 34796
rect 39194 34756 39234 34796
rect 39234 34756 39274 34796
rect 39318 34756 39358 34796
rect 39358 34756 39398 34796
rect 39398 34756 39440 34796
rect 39440 34756 39442 34796
rect 39150 34714 39274 34756
rect 39318 34714 39442 34756
rect 51150 34796 51274 34838
rect 51318 34796 51442 34838
rect 51150 34756 51152 34796
rect 51152 34756 51194 34796
rect 51194 34756 51234 34796
rect 51234 34756 51274 34796
rect 51318 34756 51358 34796
rect 51358 34756 51398 34796
rect 51398 34756 51440 34796
rect 51440 34756 51442 34796
rect 51150 34714 51274 34756
rect 51318 34714 51442 34756
rect 63150 34796 63274 34838
rect 63318 34796 63442 34838
rect 63150 34756 63152 34796
rect 63152 34756 63194 34796
rect 63194 34756 63234 34796
rect 63234 34756 63274 34796
rect 63318 34756 63358 34796
rect 63358 34756 63398 34796
rect 63398 34756 63440 34796
rect 63440 34756 63442 34796
rect 63150 34714 63274 34756
rect 63318 34714 63442 34756
rect 75150 34796 75274 34838
rect 75318 34796 75442 34838
rect 75150 34756 75152 34796
rect 75152 34756 75194 34796
rect 75194 34756 75234 34796
rect 75234 34756 75274 34796
rect 75318 34756 75358 34796
rect 75358 34756 75398 34796
rect 75398 34756 75440 34796
rect 75440 34756 75442 34796
rect 75150 34714 75274 34756
rect 75318 34714 75442 34756
rect 4390 34040 4514 34082
rect 4558 34040 4682 34082
rect 4390 34000 4392 34040
rect 4392 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4514 34040
rect 4558 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4680 34040
rect 4680 34000 4682 34040
rect 4390 33958 4514 34000
rect 4558 33958 4682 34000
rect 16390 34040 16514 34082
rect 16558 34040 16682 34082
rect 16390 34000 16392 34040
rect 16392 34000 16434 34040
rect 16434 34000 16474 34040
rect 16474 34000 16514 34040
rect 16558 34000 16598 34040
rect 16598 34000 16638 34040
rect 16638 34000 16680 34040
rect 16680 34000 16682 34040
rect 16390 33958 16514 34000
rect 16558 33958 16682 34000
rect 28390 34040 28514 34082
rect 28558 34040 28682 34082
rect 28390 34000 28392 34040
rect 28392 34000 28434 34040
rect 28434 34000 28474 34040
rect 28474 34000 28514 34040
rect 28558 34000 28598 34040
rect 28598 34000 28638 34040
rect 28638 34000 28680 34040
rect 28680 34000 28682 34040
rect 28390 33958 28514 34000
rect 28558 33958 28682 34000
rect 40390 34040 40514 34082
rect 40558 34040 40682 34082
rect 40390 34000 40392 34040
rect 40392 34000 40434 34040
rect 40434 34000 40474 34040
rect 40474 34000 40514 34040
rect 40558 34000 40598 34040
rect 40598 34000 40638 34040
rect 40638 34000 40680 34040
rect 40680 34000 40682 34040
rect 40390 33958 40514 34000
rect 40558 33958 40682 34000
rect 52390 34040 52514 34082
rect 52558 34040 52682 34082
rect 52390 34000 52392 34040
rect 52392 34000 52434 34040
rect 52434 34000 52474 34040
rect 52474 34000 52514 34040
rect 52558 34000 52598 34040
rect 52598 34000 52638 34040
rect 52638 34000 52680 34040
rect 52680 34000 52682 34040
rect 52390 33958 52514 34000
rect 52558 33958 52682 34000
rect 64390 34040 64514 34082
rect 64558 34040 64682 34082
rect 64390 34000 64392 34040
rect 64392 34000 64434 34040
rect 64434 34000 64474 34040
rect 64474 34000 64514 34040
rect 64558 34000 64598 34040
rect 64598 34000 64638 34040
rect 64638 34000 64680 34040
rect 64680 34000 64682 34040
rect 64390 33958 64514 34000
rect 64558 33958 64682 34000
rect 76390 34040 76514 34082
rect 76558 34040 76682 34082
rect 76390 34000 76392 34040
rect 76392 34000 76434 34040
rect 76434 34000 76474 34040
rect 76474 34000 76514 34040
rect 76558 34000 76598 34040
rect 76598 34000 76638 34040
rect 76638 34000 76680 34040
rect 76680 34000 76682 34040
rect 76390 33958 76514 34000
rect 76558 33958 76682 34000
rect 3150 33284 3274 33326
rect 3318 33284 3442 33326
rect 3150 33244 3152 33284
rect 3152 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3274 33284
rect 3318 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3440 33284
rect 3440 33244 3442 33284
rect 3150 33202 3274 33244
rect 3318 33202 3442 33244
rect 15150 33284 15274 33326
rect 15318 33284 15442 33326
rect 15150 33244 15152 33284
rect 15152 33244 15194 33284
rect 15194 33244 15234 33284
rect 15234 33244 15274 33284
rect 15318 33244 15358 33284
rect 15358 33244 15398 33284
rect 15398 33244 15440 33284
rect 15440 33244 15442 33284
rect 15150 33202 15274 33244
rect 15318 33202 15442 33244
rect 27150 33284 27274 33326
rect 27318 33284 27442 33326
rect 27150 33244 27152 33284
rect 27152 33244 27194 33284
rect 27194 33244 27234 33284
rect 27234 33244 27274 33284
rect 27318 33244 27358 33284
rect 27358 33244 27398 33284
rect 27398 33244 27440 33284
rect 27440 33244 27442 33284
rect 27150 33202 27274 33244
rect 27318 33202 27442 33244
rect 39150 33284 39274 33326
rect 39318 33284 39442 33326
rect 39150 33244 39152 33284
rect 39152 33244 39194 33284
rect 39194 33244 39234 33284
rect 39234 33244 39274 33284
rect 39318 33244 39358 33284
rect 39358 33244 39398 33284
rect 39398 33244 39440 33284
rect 39440 33244 39442 33284
rect 39150 33202 39274 33244
rect 39318 33202 39442 33244
rect 51150 33284 51274 33326
rect 51318 33284 51442 33326
rect 51150 33244 51152 33284
rect 51152 33244 51194 33284
rect 51194 33244 51234 33284
rect 51234 33244 51274 33284
rect 51318 33244 51358 33284
rect 51358 33244 51398 33284
rect 51398 33244 51440 33284
rect 51440 33244 51442 33284
rect 51150 33202 51274 33244
rect 51318 33202 51442 33244
rect 63150 33284 63274 33326
rect 63318 33284 63442 33326
rect 63150 33244 63152 33284
rect 63152 33244 63194 33284
rect 63194 33244 63234 33284
rect 63234 33244 63274 33284
rect 63318 33244 63358 33284
rect 63358 33244 63398 33284
rect 63398 33244 63440 33284
rect 63440 33244 63442 33284
rect 63150 33202 63274 33244
rect 63318 33202 63442 33244
rect 75150 33284 75274 33326
rect 75318 33284 75442 33326
rect 75150 33244 75152 33284
rect 75152 33244 75194 33284
rect 75194 33244 75234 33284
rect 75234 33244 75274 33284
rect 75318 33244 75358 33284
rect 75358 33244 75398 33284
rect 75398 33244 75440 33284
rect 75440 33244 75442 33284
rect 75150 33202 75274 33244
rect 75318 33202 75442 33244
rect 4390 32528 4514 32570
rect 4558 32528 4682 32570
rect 4390 32488 4392 32528
rect 4392 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4514 32528
rect 4558 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4680 32528
rect 4680 32488 4682 32528
rect 4390 32446 4514 32488
rect 4558 32446 4682 32488
rect 16390 32528 16514 32570
rect 16558 32528 16682 32570
rect 16390 32488 16392 32528
rect 16392 32488 16434 32528
rect 16434 32488 16474 32528
rect 16474 32488 16514 32528
rect 16558 32488 16598 32528
rect 16598 32488 16638 32528
rect 16638 32488 16680 32528
rect 16680 32488 16682 32528
rect 16390 32446 16514 32488
rect 16558 32446 16682 32488
rect 28390 32528 28514 32570
rect 28558 32528 28682 32570
rect 28390 32488 28392 32528
rect 28392 32488 28434 32528
rect 28434 32488 28474 32528
rect 28474 32488 28514 32528
rect 28558 32488 28598 32528
rect 28598 32488 28638 32528
rect 28638 32488 28680 32528
rect 28680 32488 28682 32528
rect 28390 32446 28514 32488
rect 28558 32446 28682 32488
rect 40390 32528 40514 32570
rect 40558 32528 40682 32570
rect 40390 32488 40392 32528
rect 40392 32488 40434 32528
rect 40434 32488 40474 32528
rect 40474 32488 40514 32528
rect 40558 32488 40598 32528
rect 40598 32488 40638 32528
rect 40638 32488 40680 32528
rect 40680 32488 40682 32528
rect 40390 32446 40514 32488
rect 40558 32446 40682 32488
rect 52390 32528 52514 32570
rect 52558 32528 52682 32570
rect 52390 32488 52392 32528
rect 52392 32488 52434 32528
rect 52434 32488 52474 32528
rect 52474 32488 52514 32528
rect 52558 32488 52598 32528
rect 52598 32488 52638 32528
rect 52638 32488 52680 32528
rect 52680 32488 52682 32528
rect 52390 32446 52514 32488
rect 52558 32446 52682 32488
rect 64390 32528 64514 32570
rect 64558 32528 64682 32570
rect 64390 32488 64392 32528
rect 64392 32488 64434 32528
rect 64434 32488 64474 32528
rect 64474 32488 64514 32528
rect 64558 32488 64598 32528
rect 64598 32488 64638 32528
rect 64638 32488 64680 32528
rect 64680 32488 64682 32528
rect 64390 32446 64514 32488
rect 64558 32446 64682 32488
rect 76390 32528 76514 32570
rect 76558 32528 76682 32570
rect 76390 32488 76392 32528
rect 76392 32488 76434 32528
rect 76434 32488 76474 32528
rect 76474 32488 76514 32528
rect 76558 32488 76598 32528
rect 76598 32488 76638 32528
rect 76638 32488 76680 32528
rect 76680 32488 76682 32528
rect 76390 32446 76514 32488
rect 76558 32446 76682 32488
rect 3150 31772 3274 31814
rect 3318 31772 3442 31814
rect 3150 31732 3152 31772
rect 3152 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3274 31772
rect 3318 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3440 31772
rect 3440 31732 3442 31772
rect 3150 31690 3274 31732
rect 3318 31690 3442 31732
rect 15150 31772 15274 31814
rect 15318 31772 15442 31814
rect 15150 31732 15152 31772
rect 15152 31732 15194 31772
rect 15194 31732 15234 31772
rect 15234 31732 15274 31772
rect 15318 31732 15358 31772
rect 15358 31732 15398 31772
rect 15398 31732 15440 31772
rect 15440 31732 15442 31772
rect 15150 31690 15274 31732
rect 15318 31690 15442 31732
rect 27150 31772 27274 31814
rect 27318 31772 27442 31814
rect 27150 31732 27152 31772
rect 27152 31732 27194 31772
rect 27194 31732 27234 31772
rect 27234 31732 27274 31772
rect 27318 31732 27358 31772
rect 27358 31732 27398 31772
rect 27398 31732 27440 31772
rect 27440 31732 27442 31772
rect 27150 31690 27274 31732
rect 27318 31690 27442 31732
rect 39150 31772 39274 31814
rect 39318 31772 39442 31814
rect 39150 31732 39152 31772
rect 39152 31732 39194 31772
rect 39194 31732 39234 31772
rect 39234 31732 39274 31772
rect 39318 31732 39358 31772
rect 39358 31732 39398 31772
rect 39398 31732 39440 31772
rect 39440 31732 39442 31772
rect 39150 31690 39274 31732
rect 39318 31690 39442 31732
rect 51150 31772 51274 31814
rect 51318 31772 51442 31814
rect 51150 31732 51152 31772
rect 51152 31732 51194 31772
rect 51194 31732 51234 31772
rect 51234 31732 51274 31772
rect 51318 31732 51358 31772
rect 51358 31732 51398 31772
rect 51398 31732 51440 31772
rect 51440 31732 51442 31772
rect 51150 31690 51274 31732
rect 51318 31690 51442 31732
rect 63150 31772 63274 31814
rect 63318 31772 63442 31814
rect 63150 31732 63152 31772
rect 63152 31732 63194 31772
rect 63194 31732 63234 31772
rect 63234 31732 63274 31772
rect 63318 31732 63358 31772
rect 63358 31732 63398 31772
rect 63398 31732 63440 31772
rect 63440 31732 63442 31772
rect 63150 31690 63274 31732
rect 63318 31690 63442 31732
rect 75150 31772 75274 31814
rect 75318 31772 75442 31814
rect 75150 31732 75152 31772
rect 75152 31732 75194 31772
rect 75194 31732 75234 31772
rect 75234 31732 75274 31772
rect 75318 31732 75358 31772
rect 75358 31732 75398 31772
rect 75398 31732 75440 31772
rect 75440 31732 75442 31772
rect 75150 31690 75274 31732
rect 75318 31690 75442 31732
rect 4390 31016 4514 31058
rect 4558 31016 4682 31058
rect 4390 30976 4392 31016
rect 4392 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4514 31016
rect 4558 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4680 31016
rect 4680 30976 4682 31016
rect 4390 30934 4514 30976
rect 4558 30934 4682 30976
rect 16390 31016 16514 31058
rect 16558 31016 16682 31058
rect 16390 30976 16392 31016
rect 16392 30976 16434 31016
rect 16434 30976 16474 31016
rect 16474 30976 16514 31016
rect 16558 30976 16598 31016
rect 16598 30976 16638 31016
rect 16638 30976 16680 31016
rect 16680 30976 16682 31016
rect 16390 30934 16514 30976
rect 16558 30934 16682 30976
rect 28390 31016 28514 31058
rect 28558 31016 28682 31058
rect 28390 30976 28392 31016
rect 28392 30976 28434 31016
rect 28434 30976 28474 31016
rect 28474 30976 28514 31016
rect 28558 30976 28598 31016
rect 28598 30976 28638 31016
rect 28638 30976 28680 31016
rect 28680 30976 28682 31016
rect 28390 30934 28514 30976
rect 28558 30934 28682 30976
rect 40390 31016 40514 31058
rect 40558 31016 40682 31058
rect 40390 30976 40392 31016
rect 40392 30976 40434 31016
rect 40434 30976 40474 31016
rect 40474 30976 40514 31016
rect 40558 30976 40598 31016
rect 40598 30976 40638 31016
rect 40638 30976 40680 31016
rect 40680 30976 40682 31016
rect 40390 30934 40514 30976
rect 40558 30934 40682 30976
rect 52390 31016 52514 31058
rect 52558 31016 52682 31058
rect 52390 30976 52392 31016
rect 52392 30976 52434 31016
rect 52434 30976 52474 31016
rect 52474 30976 52514 31016
rect 52558 30976 52598 31016
rect 52598 30976 52638 31016
rect 52638 30976 52680 31016
rect 52680 30976 52682 31016
rect 52390 30934 52514 30976
rect 52558 30934 52682 30976
rect 64390 31016 64514 31058
rect 64558 31016 64682 31058
rect 64390 30976 64392 31016
rect 64392 30976 64434 31016
rect 64434 30976 64474 31016
rect 64474 30976 64514 31016
rect 64558 30976 64598 31016
rect 64598 30976 64638 31016
rect 64638 30976 64680 31016
rect 64680 30976 64682 31016
rect 64390 30934 64514 30976
rect 64558 30934 64682 30976
rect 76390 31016 76514 31058
rect 76558 31016 76682 31058
rect 76390 30976 76392 31016
rect 76392 30976 76434 31016
rect 76434 30976 76474 31016
rect 76474 30976 76514 31016
rect 76558 30976 76598 31016
rect 76598 30976 76638 31016
rect 76638 30976 76680 31016
rect 76680 30976 76682 31016
rect 76390 30934 76514 30976
rect 76558 30934 76682 30976
rect 3150 30260 3274 30302
rect 3318 30260 3442 30302
rect 3150 30220 3152 30260
rect 3152 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3274 30260
rect 3318 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3440 30260
rect 3440 30220 3442 30260
rect 3150 30178 3274 30220
rect 3318 30178 3442 30220
rect 15150 30260 15274 30302
rect 15318 30260 15442 30302
rect 15150 30220 15152 30260
rect 15152 30220 15194 30260
rect 15194 30220 15234 30260
rect 15234 30220 15274 30260
rect 15318 30220 15358 30260
rect 15358 30220 15398 30260
rect 15398 30220 15440 30260
rect 15440 30220 15442 30260
rect 15150 30178 15274 30220
rect 15318 30178 15442 30220
rect 27150 30260 27274 30302
rect 27318 30260 27442 30302
rect 27150 30220 27152 30260
rect 27152 30220 27194 30260
rect 27194 30220 27234 30260
rect 27234 30220 27274 30260
rect 27318 30220 27358 30260
rect 27358 30220 27398 30260
rect 27398 30220 27440 30260
rect 27440 30220 27442 30260
rect 27150 30178 27274 30220
rect 27318 30178 27442 30220
rect 39150 30260 39274 30302
rect 39318 30260 39442 30302
rect 39150 30220 39152 30260
rect 39152 30220 39194 30260
rect 39194 30220 39234 30260
rect 39234 30220 39274 30260
rect 39318 30220 39358 30260
rect 39358 30220 39398 30260
rect 39398 30220 39440 30260
rect 39440 30220 39442 30260
rect 39150 30178 39274 30220
rect 39318 30178 39442 30220
rect 51150 30260 51274 30302
rect 51318 30260 51442 30302
rect 51150 30220 51152 30260
rect 51152 30220 51194 30260
rect 51194 30220 51234 30260
rect 51234 30220 51274 30260
rect 51318 30220 51358 30260
rect 51358 30220 51398 30260
rect 51398 30220 51440 30260
rect 51440 30220 51442 30260
rect 51150 30178 51274 30220
rect 51318 30178 51442 30220
rect 63150 30260 63274 30302
rect 63318 30260 63442 30302
rect 63150 30220 63152 30260
rect 63152 30220 63194 30260
rect 63194 30220 63234 30260
rect 63234 30220 63274 30260
rect 63318 30220 63358 30260
rect 63358 30220 63398 30260
rect 63398 30220 63440 30260
rect 63440 30220 63442 30260
rect 63150 30178 63274 30220
rect 63318 30178 63442 30220
rect 75150 30260 75274 30302
rect 75318 30260 75442 30302
rect 75150 30220 75152 30260
rect 75152 30220 75194 30260
rect 75194 30220 75234 30260
rect 75234 30220 75274 30260
rect 75318 30220 75358 30260
rect 75358 30220 75398 30260
rect 75398 30220 75440 30260
rect 75440 30220 75442 30260
rect 75150 30178 75274 30220
rect 75318 30178 75442 30220
rect 4390 29504 4514 29546
rect 4558 29504 4682 29546
rect 4390 29464 4392 29504
rect 4392 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4514 29504
rect 4558 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4680 29504
rect 4680 29464 4682 29504
rect 4390 29422 4514 29464
rect 4558 29422 4682 29464
rect 16390 29504 16514 29546
rect 16558 29504 16682 29546
rect 16390 29464 16392 29504
rect 16392 29464 16434 29504
rect 16434 29464 16474 29504
rect 16474 29464 16514 29504
rect 16558 29464 16598 29504
rect 16598 29464 16638 29504
rect 16638 29464 16680 29504
rect 16680 29464 16682 29504
rect 16390 29422 16514 29464
rect 16558 29422 16682 29464
rect 28390 29504 28514 29546
rect 28558 29504 28682 29546
rect 28390 29464 28392 29504
rect 28392 29464 28434 29504
rect 28434 29464 28474 29504
rect 28474 29464 28514 29504
rect 28558 29464 28598 29504
rect 28598 29464 28638 29504
rect 28638 29464 28680 29504
rect 28680 29464 28682 29504
rect 28390 29422 28514 29464
rect 28558 29422 28682 29464
rect 40390 29504 40514 29546
rect 40558 29504 40682 29546
rect 40390 29464 40392 29504
rect 40392 29464 40434 29504
rect 40434 29464 40474 29504
rect 40474 29464 40514 29504
rect 40558 29464 40598 29504
rect 40598 29464 40638 29504
rect 40638 29464 40680 29504
rect 40680 29464 40682 29504
rect 40390 29422 40514 29464
rect 40558 29422 40682 29464
rect 52390 29504 52514 29546
rect 52558 29504 52682 29546
rect 52390 29464 52392 29504
rect 52392 29464 52434 29504
rect 52434 29464 52474 29504
rect 52474 29464 52514 29504
rect 52558 29464 52598 29504
rect 52598 29464 52638 29504
rect 52638 29464 52680 29504
rect 52680 29464 52682 29504
rect 52390 29422 52514 29464
rect 52558 29422 52682 29464
rect 64390 29504 64514 29546
rect 64558 29504 64682 29546
rect 64390 29464 64392 29504
rect 64392 29464 64434 29504
rect 64434 29464 64474 29504
rect 64474 29464 64514 29504
rect 64558 29464 64598 29504
rect 64598 29464 64638 29504
rect 64638 29464 64680 29504
rect 64680 29464 64682 29504
rect 64390 29422 64514 29464
rect 64558 29422 64682 29464
rect 76390 29504 76514 29546
rect 76558 29504 76682 29546
rect 76390 29464 76392 29504
rect 76392 29464 76434 29504
rect 76434 29464 76474 29504
rect 76474 29464 76514 29504
rect 76558 29464 76598 29504
rect 76598 29464 76638 29504
rect 76638 29464 76680 29504
rect 76680 29464 76682 29504
rect 76390 29422 76514 29464
rect 76558 29422 76682 29464
rect 3150 28748 3274 28790
rect 3318 28748 3442 28790
rect 3150 28708 3152 28748
rect 3152 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3274 28748
rect 3318 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3440 28748
rect 3440 28708 3442 28748
rect 3150 28666 3274 28708
rect 3318 28666 3442 28708
rect 15150 28748 15274 28790
rect 15318 28748 15442 28790
rect 15150 28708 15152 28748
rect 15152 28708 15194 28748
rect 15194 28708 15234 28748
rect 15234 28708 15274 28748
rect 15318 28708 15358 28748
rect 15358 28708 15398 28748
rect 15398 28708 15440 28748
rect 15440 28708 15442 28748
rect 15150 28666 15274 28708
rect 15318 28666 15442 28708
rect 27150 28748 27274 28790
rect 27318 28748 27442 28790
rect 27150 28708 27152 28748
rect 27152 28708 27194 28748
rect 27194 28708 27234 28748
rect 27234 28708 27274 28748
rect 27318 28708 27358 28748
rect 27358 28708 27398 28748
rect 27398 28708 27440 28748
rect 27440 28708 27442 28748
rect 27150 28666 27274 28708
rect 27318 28666 27442 28708
rect 39150 28748 39274 28790
rect 39318 28748 39442 28790
rect 39150 28708 39152 28748
rect 39152 28708 39194 28748
rect 39194 28708 39234 28748
rect 39234 28708 39274 28748
rect 39318 28708 39358 28748
rect 39358 28708 39398 28748
rect 39398 28708 39440 28748
rect 39440 28708 39442 28748
rect 39150 28666 39274 28708
rect 39318 28666 39442 28708
rect 51150 28748 51274 28790
rect 51318 28748 51442 28790
rect 51150 28708 51152 28748
rect 51152 28708 51194 28748
rect 51194 28708 51234 28748
rect 51234 28708 51274 28748
rect 51318 28708 51358 28748
rect 51358 28708 51398 28748
rect 51398 28708 51440 28748
rect 51440 28708 51442 28748
rect 51150 28666 51274 28708
rect 51318 28666 51442 28708
rect 63150 28748 63274 28790
rect 63318 28748 63442 28790
rect 63150 28708 63152 28748
rect 63152 28708 63194 28748
rect 63194 28708 63234 28748
rect 63234 28708 63274 28748
rect 63318 28708 63358 28748
rect 63358 28708 63398 28748
rect 63398 28708 63440 28748
rect 63440 28708 63442 28748
rect 63150 28666 63274 28708
rect 63318 28666 63442 28708
rect 75150 28748 75274 28790
rect 75318 28748 75442 28790
rect 75150 28708 75152 28748
rect 75152 28708 75194 28748
rect 75194 28708 75234 28748
rect 75234 28708 75274 28748
rect 75318 28708 75358 28748
rect 75358 28708 75398 28748
rect 75398 28708 75440 28748
rect 75440 28708 75442 28748
rect 75150 28666 75274 28708
rect 75318 28666 75442 28708
rect 4390 27992 4514 28034
rect 4558 27992 4682 28034
rect 4390 27952 4392 27992
rect 4392 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4514 27992
rect 4558 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4680 27992
rect 4680 27952 4682 27992
rect 4390 27910 4514 27952
rect 4558 27910 4682 27952
rect 16390 27992 16514 28034
rect 16558 27992 16682 28034
rect 16390 27952 16392 27992
rect 16392 27952 16434 27992
rect 16434 27952 16474 27992
rect 16474 27952 16514 27992
rect 16558 27952 16598 27992
rect 16598 27952 16638 27992
rect 16638 27952 16680 27992
rect 16680 27952 16682 27992
rect 16390 27910 16514 27952
rect 16558 27910 16682 27952
rect 28390 27992 28514 28034
rect 28558 27992 28682 28034
rect 28390 27952 28392 27992
rect 28392 27952 28434 27992
rect 28434 27952 28474 27992
rect 28474 27952 28514 27992
rect 28558 27952 28598 27992
rect 28598 27952 28638 27992
rect 28638 27952 28680 27992
rect 28680 27952 28682 27992
rect 28390 27910 28514 27952
rect 28558 27910 28682 27952
rect 40390 27992 40514 28034
rect 40558 27992 40682 28034
rect 40390 27952 40392 27992
rect 40392 27952 40434 27992
rect 40434 27952 40474 27992
rect 40474 27952 40514 27992
rect 40558 27952 40598 27992
rect 40598 27952 40638 27992
rect 40638 27952 40680 27992
rect 40680 27952 40682 27992
rect 40390 27910 40514 27952
rect 40558 27910 40682 27952
rect 52390 27992 52514 28034
rect 52558 27992 52682 28034
rect 52390 27952 52392 27992
rect 52392 27952 52434 27992
rect 52434 27952 52474 27992
rect 52474 27952 52514 27992
rect 52558 27952 52598 27992
rect 52598 27952 52638 27992
rect 52638 27952 52680 27992
rect 52680 27952 52682 27992
rect 52390 27910 52514 27952
rect 52558 27910 52682 27952
rect 64390 27992 64514 28034
rect 64558 27992 64682 28034
rect 64390 27952 64392 27992
rect 64392 27952 64434 27992
rect 64434 27952 64474 27992
rect 64474 27952 64514 27992
rect 64558 27952 64598 27992
rect 64598 27952 64638 27992
rect 64638 27952 64680 27992
rect 64680 27952 64682 27992
rect 64390 27910 64514 27952
rect 64558 27910 64682 27952
rect 76390 27992 76514 28034
rect 76558 27992 76682 28034
rect 76390 27952 76392 27992
rect 76392 27952 76434 27992
rect 76434 27952 76474 27992
rect 76474 27952 76514 27992
rect 76558 27952 76598 27992
rect 76598 27952 76638 27992
rect 76638 27952 76680 27992
rect 76680 27952 76682 27992
rect 76390 27910 76514 27952
rect 76558 27910 76682 27952
rect 3150 27236 3274 27278
rect 3318 27236 3442 27278
rect 3150 27196 3152 27236
rect 3152 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3274 27236
rect 3318 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3440 27236
rect 3440 27196 3442 27236
rect 3150 27154 3274 27196
rect 3318 27154 3442 27196
rect 15150 27236 15274 27278
rect 15318 27236 15442 27278
rect 15150 27196 15152 27236
rect 15152 27196 15194 27236
rect 15194 27196 15234 27236
rect 15234 27196 15274 27236
rect 15318 27196 15358 27236
rect 15358 27196 15398 27236
rect 15398 27196 15440 27236
rect 15440 27196 15442 27236
rect 15150 27154 15274 27196
rect 15318 27154 15442 27196
rect 27150 27236 27274 27278
rect 27318 27236 27442 27278
rect 27150 27196 27152 27236
rect 27152 27196 27194 27236
rect 27194 27196 27234 27236
rect 27234 27196 27274 27236
rect 27318 27196 27358 27236
rect 27358 27196 27398 27236
rect 27398 27196 27440 27236
rect 27440 27196 27442 27236
rect 27150 27154 27274 27196
rect 27318 27154 27442 27196
rect 39150 27236 39274 27278
rect 39318 27236 39442 27278
rect 39150 27196 39152 27236
rect 39152 27196 39194 27236
rect 39194 27196 39234 27236
rect 39234 27196 39274 27236
rect 39318 27196 39358 27236
rect 39358 27196 39398 27236
rect 39398 27196 39440 27236
rect 39440 27196 39442 27236
rect 39150 27154 39274 27196
rect 39318 27154 39442 27196
rect 51150 27236 51274 27278
rect 51318 27236 51442 27278
rect 51150 27196 51152 27236
rect 51152 27196 51194 27236
rect 51194 27196 51234 27236
rect 51234 27196 51274 27236
rect 51318 27196 51358 27236
rect 51358 27196 51398 27236
rect 51398 27196 51440 27236
rect 51440 27196 51442 27236
rect 51150 27154 51274 27196
rect 51318 27154 51442 27196
rect 63150 27236 63274 27278
rect 63318 27236 63442 27278
rect 63150 27196 63152 27236
rect 63152 27196 63194 27236
rect 63194 27196 63234 27236
rect 63234 27196 63274 27236
rect 63318 27196 63358 27236
rect 63358 27196 63398 27236
rect 63398 27196 63440 27236
rect 63440 27196 63442 27236
rect 63150 27154 63274 27196
rect 63318 27154 63442 27196
rect 75150 27236 75274 27278
rect 75318 27236 75442 27278
rect 75150 27196 75152 27236
rect 75152 27196 75194 27236
rect 75194 27196 75234 27236
rect 75234 27196 75274 27236
rect 75318 27196 75358 27236
rect 75358 27196 75398 27236
rect 75398 27196 75440 27236
rect 75440 27196 75442 27236
rect 75150 27154 75274 27196
rect 75318 27154 75442 27196
rect 4390 26480 4514 26522
rect 4558 26480 4682 26522
rect 4390 26440 4392 26480
rect 4392 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4514 26480
rect 4558 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4680 26480
rect 4680 26440 4682 26480
rect 4390 26398 4514 26440
rect 4558 26398 4682 26440
rect 16390 26480 16514 26522
rect 16558 26480 16682 26522
rect 16390 26440 16392 26480
rect 16392 26440 16434 26480
rect 16434 26440 16474 26480
rect 16474 26440 16514 26480
rect 16558 26440 16598 26480
rect 16598 26440 16638 26480
rect 16638 26440 16680 26480
rect 16680 26440 16682 26480
rect 16390 26398 16514 26440
rect 16558 26398 16682 26440
rect 28390 26480 28514 26522
rect 28558 26480 28682 26522
rect 28390 26440 28392 26480
rect 28392 26440 28434 26480
rect 28434 26440 28474 26480
rect 28474 26440 28514 26480
rect 28558 26440 28598 26480
rect 28598 26440 28638 26480
rect 28638 26440 28680 26480
rect 28680 26440 28682 26480
rect 28390 26398 28514 26440
rect 28558 26398 28682 26440
rect 40390 26480 40514 26522
rect 40558 26480 40682 26522
rect 40390 26440 40392 26480
rect 40392 26440 40434 26480
rect 40434 26440 40474 26480
rect 40474 26440 40514 26480
rect 40558 26440 40598 26480
rect 40598 26440 40638 26480
rect 40638 26440 40680 26480
rect 40680 26440 40682 26480
rect 40390 26398 40514 26440
rect 40558 26398 40682 26440
rect 52390 26480 52514 26522
rect 52558 26480 52682 26522
rect 52390 26440 52392 26480
rect 52392 26440 52434 26480
rect 52434 26440 52474 26480
rect 52474 26440 52514 26480
rect 52558 26440 52598 26480
rect 52598 26440 52638 26480
rect 52638 26440 52680 26480
rect 52680 26440 52682 26480
rect 52390 26398 52514 26440
rect 52558 26398 52682 26440
rect 64390 26480 64514 26522
rect 64558 26480 64682 26522
rect 64390 26440 64392 26480
rect 64392 26440 64434 26480
rect 64434 26440 64474 26480
rect 64474 26440 64514 26480
rect 64558 26440 64598 26480
rect 64598 26440 64638 26480
rect 64638 26440 64680 26480
rect 64680 26440 64682 26480
rect 64390 26398 64514 26440
rect 64558 26398 64682 26440
rect 76390 26480 76514 26522
rect 76558 26480 76682 26522
rect 76390 26440 76392 26480
rect 76392 26440 76434 26480
rect 76434 26440 76474 26480
rect 76474 26440 76514 26480
rect 76558 26440 76598 26480
rect 76598 26440 76638 26480
rect 76638 26440 76680 26480
rect 76680 26440 76682 26480
rect 76390 26398 76514 26440
rect 76558 26398 76682 26440
rect 3150 25724 3274 25766
rect 3318 25724 3442 25766
rect 3150 25684 3152 25724
rect 3152 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3274 25724
rect 3318 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3440 25724
rect 3440 25684 3442 25724
rect 3150 25642 3274 25684
rect 3318 25642 3442 25684
rect 15150 25724 15274 25766
rect 15318 25724 15442 25766
rect 15150 25684 15152 25724
rect 15152 25684 15194 25724
rect 15194 25684 15234 25724
rect 15234 25684 15274 25724
rect 15318 25684 15358 25724
rect 15358 25684 15398 25724
rect 15398 25684 15440 25724
rect 15440 25684 15442 25724
rect 15150 25642 15274 25684
rect 15318 25642 15442 25684
rect 27150 25724 27274 25766
rect 27318 25724 27442 25766
rect 27150 25684 27152 25724
rect 27152 25684 27194 25724
rect 27194 25684 27234 25724
rect 27234 25684 27274 25724
rect 27318 25684 27358 25724
rect 27358 25684 27398 25724
rect 27398 25684 27440 25724
rect 27440 25684 27442 25724
rect 27150 25642 27274 25684
rect 27318 25642 27442 25684
rect 39150 25724 39274 25766
rect 39318 25724 39442 25766
rect 39150 25684 39152 25724
rect 39152 25684 39194 25724
rect 39194 25684 39234 25724
rect 39234 25684 39274 25724
rect 39318 25684 39358 25724
rect 39358 25684 39398 25724
rect 39398 25684 39440 25724
rect 39440 25684 39442 25724
rect 39150 25642 39274 25684
rect 39318 25642 39442 25684
rect 51150 25724 51274 25766
rect 51318 25724 51442 25766
rect 51150 25684 51152 25724
rect 51152 25684 51194 25724
rect 51194 25684 51234 25724
rect 51234 25684 51274 25724
rect 51318 25684 51358 25724
rect 51358 25684 51398 25724
rect 51398 25684 51440 25724
rect 51440 25684 51442 25724
rect 51150 25642 51274 25684
rect 51318 25642 51442 25684
rect 63150 25724 63274 25766
rect 63318 25724 63442 25766
rect 63150 25684 63152 25724
rect 63152 25684 63194 25724
rect 63194 25684 63234 25724
rect 63234 25684 63274 25724
rect 63318 25684 63358 25724
rect 63358 25684 63398 25724
rect 63398 25684 63440 25724
rect 63440 25684 63442 25724
rect 63150 25642 63274 25684
rect 63318 25642 63442 25684
rect 75150 25724 75274 25766
rect 75318 25724 75442 25766
rect 75150 25684 75152 25724
rect 75152 25684 75194 25724
rect 75194 25684 75234 25724
rect 75234 25684 75274 25724
rect 75318 25684 75358 25724
rect 75358 25684 75398 25724
rect 75398 25684 75440 25724
rect 75440 25684 75442 25724
rect 75150 25642 75274 25684
rect 75318 25642 75442 25684
rect 4390 24968 4514 25010
rect 4558 24968 4682 25010
rect 4390 24928 4392 24968
rect 4392 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4514 24968
rect 4558 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4680 24968
rect 4680 24928 4682 24968
rect 4390 24886 4514 24928
rect 4558 24886 4682 24928
rect 16390 24968 16514 25010
rect 16558 24968 16682 25010
rect 16390 24928 16392 24968
rect 16392 24928 16434 24968
rect 16434 24928 16474 24968
rect 16474 24928 16514 24968
rect 16558 24928 16598 24968
rect 16598 24928 16638 24968
rect 16638 24928 16680 24968
rect 16680 24928 16682 24968
rect 16390 24886 16514 24928
rect 16558 24886 16682 24928
rect 28390 24968 28514 25010
rect 28558 24968 28682 25010
rect 28390 24928 28392 24968
rect 28392 24928 28434 24968
rect 28434 24928 28474 24968
rect 28474 24928 28514 24968
rect 28558 24928 28598 24968
rect 28598 24928 28638 24968
rect 28638 24928 28680 24968
rect 28680 24928 28682 24968
rect 28390 24886 28514 24928
rect 28558 24886 28682 24928
rect 40390 24968 40514 25010
rect 40558 24968 40682 25010
rect 40390 24928 40392 24968
rect 40392 24928 40434 24968
rect 40434 24928 40474 24968
rect 40474 24928 40514 24968
rect 40558 24928 40598 24968
rect 40598 24928 40638 24968
rect 40638 24928 40680 24968
rect 40680 24928 40682 24968
rect 40390 24886 40514 24928
rect 40558 24886 40682 24928
rect 52390 24968 52514 25010
rect 52558 24968 52682 25010
rect 64390 24968 64514 25010
rect 64558 24968 64682 25010
rect 52390 24928 52392 24968
rect 52392 24928 52434 24968
rect 52434 24928 52474 24968
rect 52474 24928 52514 24968
rect 52558 24928 52598 24968
rect 52598 24928 52638 24968
rect 52638 24928 52680 24968
rect 52680 24928 52682 24968
rect 64390 24928 64392 24968
rect 64392 24928 64434 24968
rect 64434 24928 64474 24968
rect 64474 24928 64514 24968
rect 64558 24928 64598 24968
rect 64598 24928 64638 24968
rect 64638 24928 64680 24968
rect 64680 24928 64682 24968
rect 52390 24886 52514 24928
rect 52558 24886 52682 24928
rect 64390 24886 64514 24928
rect 64558 24886 64682 24928
rect 76390 24968 76514 25010
rect 76558 24968 76682 25010
rect 76390 24928 76392 24968
rect 76392 24928 76434 24968
rect 76434 24928 76474 24968
rect 76474 24928 76514 24968
rect 76558 24928 76598 24968
rect 76598 24928 76638 24968
rect 76638 24928 76680 24968
rect 76680 24928 76682 24968
rect 76390 24886 76514 24928
rect 76558 24886 76682 24928
rect 3150 24212 3274 24254
rect 3318 24212 3442 24254
rect 3150 24172 3152 24212
rect 3152 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3274 24212
rect 3318 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3440 24212
rect 3440 24172 3442 24212
rect 3150 24130 3274 24172
rect 3318 24130 3442 24172
rect 15150 24212 15274 24254
rect 15318 24212 15442 24254
rect 15150 24172 15152 24212
rect 15152 24172 15194 24212
rect 15194 24172 15234 24212
rect 15234 24172 15274 24212
rect 15318 24172 15358 24212
rect 15358 24172 15398 24212
rect 15398 24172 15440 24212
rect 15440 24172 15442 24212
rect 15150 24130 15274 24172
rect 15318 24130 15442 24172
rect 27150 24212 27274 24254
rect 27318 24212 27442 24254
rect 27150 24172 27152 24212
rect 27152 24172 27194 24212
rect 27194 24172 27234 24212
rect 27234 24172 27274 24212
rect 27318 24172 27358 24212
rect 27358 24172 27398 24212
rect 27398 24172 27440 24212
rect 27440 24172 27442 24212
rect 27150 24130 27274 24172
rect 27318 24130 27442 24172
rect 39150 24212 39274 24254
rect 39318 24212 39442 24254
rect 39150 24172 39152 24212
rect 39152 24172 39194 24212
rect 39194 24172 39234 24212
rect 39234 24172 39274 24212
rect 39318 24172 39358 24212
rect 39358 24172 39398 24212
rect 39398 24172 39440 24212
rect 39440 24172 39442 24212
rect 39150 24130 39274 24172
rect 39318 24130 39442 24172
rect 78698 23710 78822 23834
rect 4390 23456 4514 23498
rect 4558 23456 4682 23498
rect 4390 23416 4392 23456
rect 4392 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4514 23456
rect 4558 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4680 23456
rect 4680 23416 4682 23456
rect 4390 23374 4514 23416
rect 4558 23374 4682 23416
rect 16390 23456 16514 23498
rect 16558 23456 16682 23498
rect 16390 23416 16392 23456
rect 16392 23416 16434 23456
rect 16434 23416 16474 23456
rect 16474 23416 16514 23456
rect 16558 23416 16598 23456
rect 16598 23416 16638 23456
rect 16638 23416 16680 23456
rect 16680 23416 16682 23456
rect 16390 23374 16514 23416
rect 16558 23374 16682 23416
rect 28390 23456 28514 23498
rect 28558 23456 28682 23498
rect 28390 23416 28392 23456
rect 28392 23416 28434 23456
rect 28434 23416 28474 23456
rect 28474 23416 28514 23456
rect 28558 23416 28598 23456
rect 28598 23416 28638 23456
rect 28638 23416 28680 23456
rect 28680 23416 28682 23456
rect 28390 23374 28514 23416
rect 28558 23374 28682 23416
rect 40390 23456 40514 23498
rect 40558 23456 40682 23498
rect 40390 23416 40392 23456
rect 40392 23416 40434 23456
rect 40434 23416 40474 23456
rect 40474 23416 40514 23456
rect 40558 23416 40598 23456
rect 40598 23416 40638 23456
rect 40638 23416 40680 23456
rect 40680 23416 40682 23456
rect 40390 23374 40514 23416
rect 40558 23374 40682 23416
rect 74138 23038 74262 23162
rect 71858 22784 71982 22826
rect 71858 22744 71884 22784
rect 71884 22744 71924 22784
rect 71924 22744 71982 22784
rect 3150 22700 3274 22742
rect 3318 22700 3442 22742
rect 3150 22660 3152 22700
rect 3152 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3274 22700
rect 3318 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3440 22700
rect 3440 22660 3442 22700
rect 3150 22618 3274 22660
rect 3318 22618 3442 22660
rect 15150 22700 15274 22742
rect 15318 22700 15442 22742
rect 15150 22660 15152 22700
rect 15152 22660 15194 22700
rect 15194 22660 15234 22700
rect 15234 22660 15274 22700
rect 15318 22660 15358 22700
rect 15358 22660 15398 22700
rect 15398 22660 15440 22700
rect 15440 22660 15442 22700
rect 15150 22618 15274 22660
rect 15318 22618 15442 22660
rect 27150 22700 27274 22742
rect 27318 22700 27442 22742
rect 27150 22660 27152 22700
rect 27152 22660 27194 22700
rect 27194 22660 27234 22700
rect 27234 22660 27274 22700
rect 27318 22660 27358 22700
rect 27358 22660 27398 22700
rect 27398 22660 27440 22700
rect 27440 22660 27442 22700
rect 27150 22618 27274 22660
rect 27318 22618 27442 22660
rect 39150 22700 39274 22742
rect 39318 22700 39442 22742
rect 71858 22702 71982 22744
rect 39150 22660 39152 22700
rect 39152 22660 39194 22700
rect 39194 22660 39234 22700
rect 39234 22660 39274 22700
rect 39318 22660 39358 22700
rect 39358 22660 39398 22700
rect 39398 22660 39440 22700
rect 39440 22660 39442 22700
rect 39150 22618 39274 22660
rect 39318 22618 39442 22660
rect 64390 22417 64514 22541
rect 64558 22417 64682 22541
rect 64390 22249 64514 22373
rect 64558 22249 64682 22373
rect 64390 22081 64514 22205
rect 64558 22081 64682 22205
rect 4390 21944 4514 21986
rect 4558 21944 4682 21986
rect 4390 21904 4392 21944
rect 4392 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4514 21944
rect 4558 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4680 21944
rect 4680 21904 4682 21944
rect 4390 21862 4514 21904
rect 4558 21862 4682 21904
rect 16390 21944 16514 21986
rect 16558 21944 16682 21986
rect 16390 21904 16392 21944
rect 16392 21904 16434 21944
rect 16434 21904 16474 21944
rect 16474 21904 16514 21944
rect 16558 21904 16598 21944
rect 16598 21904 16638 21944
rect 16638 21904 16680 21944
rect 16680 21904 16682 21944
rect 16390 21862 16514 21904
rect 16558 21862 16682 21904
rect 28390 21944 28514 21986
rect 28558 21944 28682 21986
rect 28390 21904 28392 21944
rect 28392 21904 28434 21944
rect 28434 21904 28474 21944
rect 28474 21904 28514 21944
rect 28558 21904 28598 21944
rect 28598 21904 28638 21944
rect 28638 21904 28680 21944
rect 28680 21904 28682 21944
rect 28390 21862 28514 21904
rect 28558 21862 28682 21904
rect 40390 21944 40514 21986
rect 40558 21944 40682 21986
rect 40390 21904 40392 21944
rect 40392 21904 40434 21944
rect 40434 21904 40474 21944
rect 40474 21904 40514 21944
rect 40558 21904 40598 21944
rect 40598 21904 40638 21944
rect 40638 21904 40680 21944
rect 40680 21904 40682 21944
rect 40390 21862 40514 21904
rect 40558 21862 40682 21904
rect 64390 21913 64514 22037
rect 64558 21913 64682 22037
rect 64390 21745 64514 21869
rect 64558 21745 64682 21869
rect 64390 21577 64514 21701
rect 64558 21577 64682 21701
rect 64390 21409 64514 21533
rect 64558 21409 64682 21533
rect 64390 21241 64514 21365
rect 64558 21241 64682 21365
rect 3150 21188 3274 21230
rect 3318 21188 3442 21230
rect 3150 21148 3152 21188
rect 3152 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3274 21188
rect 3318 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3440 21188
rect 3440 21148 3442 21188
rect 3150 21106 3274 21148
rect 3318 21106 3442 21148
rect 15150 21188 15274 21230
rect 15318 21188 15442 21230
rect 15150 21148 15152 21188
rect 15152 21148 15194 21188
rect 15194 21148 15234 21188
rect 15234 21148 15274 21188
rect 15318 21148 15358 21188
rect 15358 21148 15398 21188
rect 15398 21148 15440 21188
rect 15440 21148 15442 21188
rect 15150 21106 15274 21148
rect 15318 21106 15442 21148
rect 27150 21188 27274 21230
rect 27318 21188 27442 21230
rect 27150 21148 27152 21188
rect 27152 21148 27194 21188
rect 27194 21148 27234 21188
rect 27234 21148 27274 21188
rect 27318 21148 27358 21188
rect 27358 21148 27398 21188
rect 27398 21148 27440 21188
rect 27440 21148 27442 21188
rect 27150 21106 27274 21148
rect 27318 21106 27442 21148
rect 39150 21188 39274 21230
rect 39318 21188 39442 21230
rect 39150 21148 39152 21188
rect 39152 21148 39194 21188
rect 39194 21148 39234 21188
rect 39234 21148 39274 21188
rect 39318 21148 39358 21188
rect 39358 21148 39398 21188
rect 39398 21148 39440 21188
rect 39440 21148 39442 21188
rect 39150 21106 39274 21148
rect 39318 21106 39442 21148
rect 64390 21073 64514 21197
rect 64558 21073 64682 21197
rect 64390 20905 64514 21029
rect 64558 20905 64682 21029
rect 64390 20737 64514 20861
rect 64558 20737 64682 20861
rect 64390 20569 64514 20693
rect 64558 20569 64682 20693
rect 4390 20432 4514 20474
rect 4558 20432 4682 20474
rect 4390 20392 4392 20432
rect 4392 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4514 20432
rect 4558 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4680 20432
rect 4680 20392 4682 20432
rect 4390 20350 4514 20392
rect 4558 20350 4682 20392
rect 16390 20432 16514 20474
rect 16558 20432 16682 20474
rect 16390 20392 16392 20432
rect 16392 20392 16434 20432
rect 16434 20392 16474 20432
rect 16474 20392 16514 20432
rect 16558 20392 16598 20432
rect 16598 20392 16638 20432
rect 16638 20392 16680 20432
rect 16680 20392 16682 20432
rect 16390 20350 16514 20392
rect 16558 20350 16682 20392
rect 28390 20432 28514 20474
rect 28558 20432 28682 20474
rect 28390 20392 28392 20432
rect 28392 20392 28434 20432
rect 28434 20392 28474 20432
rect 28474 20392 28514 20432
rect 28558 20392 28598 20432
rect 28598 20392 28638 20432
rect 28638 20392 28680 20432
rect 28680 20392 28682 20432
rect 28390 20350 28514 20392
rect 28558 20350 28682 20392
rect 40390 20432 40514 20474
rect 40558 20432 40682 20474
rect 40390 20392 40392 20432
rect 40392 20392 40434 20432
rect 40434 20392 40474 20432
rect 40474 20392 40514 20432
rect 40558 20392 40598 20432
rect 40598 20392 40638 20432
rect 40638 20392 40680 20432
rect 40680 20392 40682 20432
rect 40390 20350 40514 20392
rect 40558 20350 40682 20392
rect 64390 20401 64514 20525
rect 64558 20401 64682 20525
rect 76390 22417 76514 22541
rect 76558 22417 76682 22541
rect 76390 22249 76514 22373
rect 76558 22249 76682 22373
rect 76390 22081 76514 22205
rect 76558 22081 76682 22205
rect 76390 21913 76514 22037
rect 76558 21913 76682 22037
rect 76390 21745 76514 21869
rect 76558 21745 76682 21869
rect 76390 21577 76514 21701
rect 76558 21577 76682 21701
rect 76390 21409 76514 21533
rect 76558 21409 76682 21533
rect 76390 21241 76514 21365
rect 76558 21241 76682 21365
rect 76390 21073 76514 21197
rect 76558 21073 76682 21197
rect 76390 20905 76514 21029
rect 76558 20905 76682 21029
rect 76390 20737 76514 20861
rect 76558 20737 76682 20861
rect 76390 20569 76514 20693
rect 76558 20569 76682 20693
rect 76390 20401 76514 20525
rect 76558 20401 76682 20525
rect 3150 19676 3274 19718
rect 3318 19676 3442 19718
rect 3150 19636 3152 19676
rect 3152 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3274 19676
rect 3318 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3440 19676
rect 3440 19636 3442 19676
rect 3150 19594 3274 19636
rect 3318 19594 3442 19636
rect 15150 19676 15274 19718
rect 15318 19676 15442 19718
rect 15150 19636 15152 19676
rect 15152 19636 15194 19676
rect 15194 19636 15234 19676
rect 15234 19636 15274 19676
rect 15318 19636 15358 19676
rect 15358 19636 15398 19676
rect 15398 19636 15440 19676
rect 15440 19636 15442 19676
rect 15150 19594 15274 19636
rect 15318 19594 15442 19636
rect 27150 19676 27274 19718
rect 27318 19676 27442 19718
rect 27150 19636 27152 19676
rect 27152 19636 27194 19676
rect 27194 19636 27234 19676
rect 27234 19636 27274 19676
rect 27318 19636 27358 19676
rect 27358 19636 27398 19676
rect 27398 19636 27440 19676
rect 27440 19636 27442 19676
rect 27150 19594 27274 19636
rect 27318 19594 27442 19636
rect 39150 19676 39274 19718
rect 39318 19676 39442 19718
rect 39150 19636 39152 19676
rect 39152 19636 39194 19676
rect 39194 19636 39234 19676
rect 39234 19636 39274 19676
rect 39318 19636 39358 19676
rect 39358 19636 39398 19676
rect 39398 19636 39440 19676
rect 39440 19636 39442 19676
rect 39150 19594 39274 19636
rect 39318 19594 39442 19636
rect 63150 19541 63274 19665
rect 63318 19541 63442 19665
rect 63150 19373 63274 19497
rect 63318 19373 63442 19497
rect 63150 19205 63274 19329
rect 63318 19205 63442 19329
rect 63150 19037 63274 19161
rect 63318 19037 63442 19161
rect 4390 18920 4514 18962
rect 4558 18920 4682 18962
rect 4390 18880 4392 18920
rect 4392 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4514 18920
rect 4558 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4680 18920
rect 4680 18880 4682 18920
rect 4390 18838 4514 18880
rect 4558 18838 4682 18880
rect 16390 18920 16514 18962
rect 16558 18920 16682 18962
rect 16390 18880 16392 18920
rect 16392 18880 16434 18920
rect 16434 18880 16474 18920
rect 16474 18880 16514 18920
rect 16558 18880 16598 18920
rect 16598 18880 16638 18920
rect 16638 18880 16680 18920
rect 16680 18880 16682 18920
rect 16390 18838 16514 18880
rect 16558 18838 16682 18880
rect 28390 18920 28514 18962
rect 28558 18920 28682 18962
rect 28390 18880 28392 18920
rect 28392 18880 28434 18920
rect 28434 18880 28474 18920
rect 28474 18880 28514 18920
rect 28558 18880 28598 18920
rect 28598 18880 28638 18920
rect 28638 18880 28680 18920
rect 28680 18880 28682 18920
rect 28390 18838 28514 18880
rect 28558 18838 28682 18880
rect 40390 18920 40514 18962
rect 40558 18920 40682 18962
rect 40390 18880 40392 18920
rect 40392 18880 40434 18920
rect 40434 18880 40474 18920
rect 40474 18880 40514 18920
rect 40558 18880 40598 18920
rect 40598 18880 40638 18920
rect 40638 18880 40680 18920
rect 40680 18880 40682 18920
rect 40390 18838 40514 18880
rect 40558 18838 40682 18880
rect 63150 18869 63274 18993
rect 63318 18869 63442 18993
rect 63150 18701 63274 18825
rect 63318 18701 63442 18825
rect 63150 18533 63274 18657
rect 63318 18533 63442 18657
rect 63150 18365 63274 18489
rect 63318 18365 63442 18489
rect 3150 18164 3274 18206
rect 3318 18164 3442 18206
rect 3150 18124 3152 18164
rect 3152 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3274 18164
rect 3318 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3440 18164
rect 3440 18124 3442 18164
rect 3150 18082 3274 18124
rect 3318 18082 3442 18124
rect 15150 18164 15274 18206
rect 15318 18164 15442 18206
rect 15150 18124 15152 18164
rect 15152 18124 15194 18164
rect 15194 18124 15234 18164
rect 15234 18124 15274 18164
rect 15318 18124 15358 18164
rect 15358 18124 15398 18164
rect 15398 18124 15440 18164
rect 15440 18124 15442 18164
rect 15150 18082 15274 18124
rect 15318 18082 15442 18124
rect 27150 18164 27274 18206
rect 27318 18164 27442 18206
rect 27150 18124 27152 18164
rect 27152 18124 27194 18164
rect 27194 18124 27234 18164
rect 27234 18124 27274 18164
rect 27318 18124 27358 18164
rect 27358 18124 27398 18164
rect 27398 18124 27440 18164
rect 27440 18124 27442 18164
rect 27150 18082 27274 18124
rect 27318 18082 27442 18124
rect 39150 18164 39274 18206
rect 39318 18164 39442 18206
rect 39150 18124 39152 18164
rect 39152 18124 39194 18164
rect 39194 18124 39234 18164
rect 39234 18124 39274 18164
rect 39318 18124 39358 18164
rect 39358 18124 39398 18164
rect 39398 18124 39440 18164
rect 39440 18124 39442 18164
rect 39150 18082 39274 18124
rect 39318 18082 39442 18124
rect 63150 18197 63274 18321
rect 63318 18197 63442 18321
rect 63150 18029 63274 18153
rect 63318 18029 63442 18153
rect 63150 17861 63274 17985
rect 63318 17861 63442 17985
rect 63150 17693 63274 17817
rect 63318 17693 63442 17817
rect 63150 17525 63274 17649
rect 63318 17525 63442 17649
rect 4390 17408 4514 17450
rect 4558 17408 4682 17450
rect 4390 17368 4392 17408
rect 4392 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4514 17408
rect 4558 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4680 17408
rect 4680 17368 4682 17408
rect 4390 17326 4514 17368
rect 4558 17326 4682 17368
rect 16390 17408 16514 17450
rect 16558 17408 16682 17450
rect 16390 17368 16392 17408
rect 16392 17368 16434 17408
rect 16434 17368 16474 17408
rect 16474 17368 16514 17408
rect 16558 17368 16598 17408
rect 16598 17368 16638 17408
rect 16638 17368 16680 17408
rect 16680 17368 16682 17408
rect 16390 17326 16514 17368
rect 16558 17326 16682 17368
rect 28390 17408 28514 17450
rect 28558 17408 28682 17450
rect 28390 17368 28392 17408
rect 28392 17368 28434 17408
rect 28434 17368 28474 17408
rect 28474 17368 28514 17408
rect 28558 17368 28598 17408
rect 28598 17368 28638 17408
rect 28638 17368 28680 17408
rect 28680 17368 28682 17408
rect 28390 17326 28514 17368
rect 28558 17326 28682 17368
rect 40390 17408 40514 17450
rect 40558 17408 40682 17450
rect 75150 19541 75274 19665
rect 75318 19541 75442 19665
rect 75150 19373 75274 19497
rect 75318 19373 75442 19497
rect 75150 19205 75274 19329
rect 75318 19205 75442 19329
rect 75150 19037 75274 19161
rect 75318 19037 75442 19161
rect 75150 18869 75274 18993
rect 75318 18869 75442 18993
rect 75150 18701 75274 18825
rect 75318 18701 75442 18825
rect 75150 18533 75274 18657
rect 75318 18533 75442 18657
rect 75150 18365 75274 18489
rect 75318 18365 75442 18489
rect 75150 18197 75274 18321
rect 75318 18197 75442 18321
rect 75150 18029 75274 18153
rect 75318 18029 75442 18153
rect 75150 17861 75274 17985
rect 75318 17861 75442 17985
rect 75150 17693 75274 17817
rect 75318 17693 75442 17817
rect 75150 17525 75274 17649
rect 75318 17525 75442 17649
rect 40390 17368 40392 17408
rect 40392 17368 40434 17408
rect 40434 17368 40474 17408
rect 40474 17368 40514 17408
rect 40558 17368 40598 17408
rect 40598 17368 40638 17408
rect 40638 17368 40680 17408
rect 40680 17368 40682 17408
rect 40390 17326 40514 17368
rect 40558 17326 40682 17368
rect 74138 17158 74262 17282
rect 3150 16652 3274 16694
rect 3318 16652 3442 16694
rect 3150 16612 3152 16652
rect 3152 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3274 16652
rect 3318 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3440 16652
rect 3440 16612 3442 16652
rect 3150 16570 3274 16612
rect 3318 16570 3442 16612
rect 15150 16652 15274 16694
rect 15318 16652 15442 16694
rect 15150 16612 15152 16652
rect 15152 16612 15194 16652
rect 15194 16612 15234 16652
rect 15234 16612 15274 16652
rect 15318 16612 15358 16652
rect 15358 16612 15398 16652
rect 15398 16612 15440 16652
rect 15440 16612 15442 16652
rect 15150 16570 15274 16612
rect 15318 16570 15442 16612
rect 27150 16652 27274 16694
rect 27318 16652 27442 16694
rect 27150 16612 27152 16652
rect 27152 16612 27194 16652
rect 27194 16612 27234 16652
rect 27234 16612 27274 16652
rect 27318 16612 27358 16652
rect 27358 16612 27398 16652
rect 27398 16612 27440 16652
rect 27440 16612 27442 16652
rect 27150 16570 27274 16612
rect 27318 16570 27442 16612
rect 39150 16652 39274 16694
rect 39318 16652 39442 16694
rect 39150 16612 39152 16652
rect 39152 16612 39194 16652
rect 39194 16612 39234 16652
rect 39234 16612 39274 16652
rect 39318 16612 39358 16652
rect 39358 16612 39398 16652
rect 39398 16612 39440 16652
rect 39440 16612 39442 16652
rect 39150 16570 39274 16612
rect 39318 16570 39442 16612
rect 71858 16318 71982 16442
rect 78698 16150 78822 16274
rect 4390 15896 4514 15938
rect 4558 15896 4682 15938
rect 4390 15856 4392 15896
rect 4392 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4514 15896
rect 4558 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4680 15896
rect 4680 15856 4682 15896
rect 4390 15814 4514 15856
rect 4558 15814 4682 15856
rect 16390 15896 16514 15938
rect 16558 15896 16682 15938
rect 16390 15856 16392 15896
rect 16392 15856 16434 15896
rect 16434 15856 16474 15896
rect 16474 15856 16514 15896
rect 16558 15856 16598 15896
rect 16598 15856 16638 15896
rect 16638 15856 16680 15896
rect 16680 15856 16682 15896
rect 16390 15814 16514 15856
rect 16558 15814 16682 15856
rect 28390 15896 28514 15938
rect 28558 15896 28682 15938
rect 28390 15856 28392 15896
rect 28392 15856 28434 15896
rect 28434 15856 28474 15896
rect 28474 15856 28514 15896
rect 28558 15856 28598 15896
rect 28598 15856 28638 15896
rect 28638 15856 28680 15896
rect 28680 15856 28682 15896
rect 28390 15814 28514 15856
rect 28558 15814 28682 15856
rect 40390 15896 40514 15938
rect 40558 15896 40682 15938
rect 40390 15856 40392 15896
rect 40392 15856 40434 15896
rect 40434 15856 40474 15896
rect 40474 15856 40514 15896
rect 40558 15856 40598 15896
rect 40598 15856 40638 15896
rect 40638 15856 40680 15896
rect 40680 15856 40682 15896
rect 40390 15814 40514 15856
rect 40558 15814 40682 15856
rect 3150 15140 3274 15182
rect 3318 15140 3442 15182
rect 3150 15100 3152 15140
rect 3152 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3274 15140
rect 3318 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3440 15140
rect 3440 15100 3442 15140
rect 3150 15058 3274 15100
rect 3318 15058 3442 15100
rect 15150 15140 15274 15182
rect 15318 15140 15442 15182
rect 15150 15100 15152 15140
rect 15152 15100 15194 15140
rect 15194 15100 15234 15140
rect 15234 15100 15274 15140
rect 15318 15100 15358 15140
rect 15358 15100 15398 15140
rect 15398 15100 15440 15140
rect 15440 15100 15442 15140
rect 15150 15058 15274 15100
rect 15318 15058 15442 15100
rect 27150 15140 27274 15182
rect 27318 15140 27442 15182
rect 27150 15100 27152 15140
rect 27152 15100 27194 15140
rect 27194 15100 27234 15140
rect 27234 15100 27274 15140
rect 27318 15100 27358 15140
rect 27358 15100 27398 15140
rect 27398 15100 27440 15140
rect 27440 15100 27442 15140
rect 27150 15058 27274 15100
rect 27318 15058 27442 15100
rect 39150 15140 39274 15182
rect 39318 15140 39442 15182
rect 39150 15100 39152 15140
rect 39152 15100 39194 15140
rect 39194 15100 39234 15140
rect 39234 15100 39274 15140
rect 39318 15100 39358 15140
rect 39358 15100 39398 15140
rect 39398 15100 39440 15140
rect 39440 15100 39442 15140
rect 39150 15058 39274 15100
rect 39318 15058 39442 15100
rect 51150 15140 51274 15182
rect 51318 15140 51442 15182
rect 51150 15100 51152 15140
rect 51152 15100 51194 15140
rect 51194 15100 51234 15140
rect 51234 15100 51274 15140
rect 51318 15100 51358 15140
rect 51358 15100 51398 15140
rect 51398 15100 51440 15140
rect 51440 15100 51442 15140
rect 51150 15058 51274 15100
rect 51318 15058 51442 15100
rect 63150 15140 63274 15182
rect 63318 15140 63442 15182
rect 63150 15100 63152 15140
rect 63152 15100 63194 15140
rect 63194 15100 63234 15140
rect 63234 15100 63274 15140
rect 63318 15100 63358 15140
rect 63358 15100 63398 15140
rect 63398 15100 63440 15140
rect 63440 15100 63442 15140
rect 63150 15058 63274 15100
rect 63318 15058 63442 15100
rect 75150 15140 75274 15182
rect 75318 15140 75442 15182
rect 75150 15100 75152 15140
rect 75152 15100 75194 15140
rect 75194 15100 75234 15140
rect 75234 15100 75274 15140
rect 75318 15100 75358 15140
rect 75358 15100 75398 15140
rect 75398 15100 75440 15140
rect 75440 15100 75442 15140
rect 75150 15058 75274 15100
rect 75318 15058 75442 15100
rect 4390 14384 4514 14426
rect 4558 14384 4682 14426
rect 4390 14344 4392 14384
rect 4392 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4514 14384
rect 4558 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4680 14384
rect 4680 14344 4682 14384
rect 4390 14302 4514 14344
rect 4558 14302 4682 14344
rect 16390 14384 16514 14426
rect 16558 14384 16682 14426
rect 16390 14344 16392 14384
rect 16392 14344 16434 14384
rect 16434 14344 16474 14384
rect 16474 14344 16514 14384
rect 16558 14344 16598 14384
rect 16598 14344 16638 14384
rect 16638 14344 16680 14384
rect 16680 14344 16682 14384
rect 16390 14302 16514 14344
rect 16558 14302 16682 14344
rect 28390 14384 28514 14426
rect 28558 14384 28682 14426
rect 28390 14344 28392 14384
rect 28392 14344 28434 14384
rect 28434 14344 28474 14384
rect 28474 14344 28514 14384
rect 28558 14344 28598 14384
rect 28598 14344 28638 14384
rect 28638 14344 28680 14384
rect 28680 14344 28682 14384
rect 28390 14302 28514 14344
rect 28558 14302 28682 14344
rect 40390 14384 40514 14426
rect 40558 14384 40682 14426
rect 40390 14344 40392 14384
rect 40392 14344 40434 14384
rect 40434 14344 40474 14384
rect 40474 14344 40514 14384
rect 40558 14344 40598 14384
rect 40598 14344 40638 14384
rect 40638 14344 40680 14384
rect 40680 14344 40682 14384
rect 40390 14302 40514 14344
rect 40558 14302 40682 14344
rect 52390 14384 52514 14426
rect 52558 14384 52682 14426
rect 52390 14344 52392 14384
rect 52392 14344 52434 14384
rect 52434 14344 52474 14384
rect 52474 14344 52514 14384
rect 52558 14344 52598 14384
rect 52598 14344 52638 14384
rect 52638 14344 52680 14384
rect 52680 14344 52682 14384
rect 52390 14302 52514 14344
rect 52558 14302 52682 14344
rect 64390 14384 64514 14426
rect 64558 14384 64682 14426
rect 64390 14344 64392 14384
rect 64392 14344 64434 14384
rect 64434 14344 64474 14384
rect 64474 14344 64514 14384
rect 64558 14344 64598 14384
rect 64598 14344 64638 14384
rect 64638 14344 64680 14384
rect 64680 14344 64682 14384
rect 64390 14302 64514 14344
rect 64558 14302 64682 14344
rect 76390 14384 76514 14426
rect 76558 14384 76682 14426
rect 76390 14344 76392 14384
rect 76392 14344 76434 14384
rect 76434 14344 76474 14384
rect 76474 14344 76514 14384
rect 76558 14344 76598 14384
rect 76598 14344 76638 14384
rect 76638 14344 76680 14384
rect 76680 14344 76682 14384
rect 76390 14302 76514 14344
rect 76558 14302 76682 14344
rect 3150 13628 3274 13670
rect 3318 13628 3442 13670
rect 3150 13588 3152 13628
rect 3152 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3274 13628
rect 3318 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3440 13628
rect 3440 13588 3442 13628
rect 3150 13546 3274 13588
rect 3318 13546 3442 13588
rect 15150 13628 15274 13670
rect 15318 13628 15442 13670
rect 15150 13588 15152 13628
rect 15152 13588 15194 13628
rect 15194 13588 15234 13628
rect 15234 13588 15274 13628
rect 15318 13588 15358 13628
rect 15358 13588 15398 13628
rect 15398 13588 15440 13628
rect 15440 13588 15442 13628
rect 15150 13546 15274 13588
rect 15318 13546 15442 13588
rect 27150 13628 27274 13670
rect 27318 13628 27442 13670
rect 27150 13588 27152 13628
rect 27152 13588 27194 13628
rect 27194 13588 27234 13628
rect 27234 13588 27274 13628
rect 27318 13588 27358 13628
rect 27358 13588 27398 13628
rect 27398 13588 27440 13628
rect 27440 13588 27442 13628
rect 27150 13546 27274 13588
rect 27318 13546 27442 13588
rect 39150 13628 39274 13670
rect 39318 13628 39442 13670
rect 39150 13588 39152 13628
rect 39152 13588 39194 13628
rect 39194 13588 39234 13628
rect 39234 13588 39274 13628
rect 39318 13588 39358 13628
rect 39358 13588 39398 13628
rect 39398 13588 39440 13628
rect 39440 13588 39442 13628
rect 39150 13546 39274 13588
rect 39318 13546 39442 13588
rect 51150 13628 51274 13670
rect 51318 13628 51442 13670
rect 51150 13588 51152 13628
rect 51152 13588 51194 13628
rect 51194 13588 51234 13628
rect 51234 13588 51274 13628
rect 51318 13588 51358 13628
rect 51358 13588 51398 13628
rect 51398 13588 51440 13628
rect 51440 13588 51442 13628
rect 51150 13546 51274 13588
rect 51318 13546 51442 13588
rect 63150 13628 63274 13670
rect 63318 13628 63442 13670
rect 63150 13588 63152 13628
rect 63152 13588 63194 13628
rect 63194 13588 63234 13628
rect 63234 13588 63274 13628
rect 63318 13588 63358 13628
rect 63358 13588 63398 13628
rect 63398 13588 63440 13628
rect 63440 13588 63442 13628
rect 63150 13546 63274 13588
rect 63318 13546 63442 13588
rect 75150 13628 75274 13670
rect 75318 13628 75442 13670
rect 75150 13588 75152 13628
rect 75152 13588 75194 13628
rect 75194 13588 75234 13628
rect 75234 13588 75274 13628
rect 75318 13588 75358 13628
rect 75358 13588 75398 13628
rect 75398 13588 75440 13628
rect 75440 13588 75442 13628
rect 75150 13546 75274 13588
rect 75318 13546 75442 13588
rect 4390 12872 4514 12914
rect 4558 12872 4682 12914
rect 4390 12832 4392 12872
rect 4392 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4514 12872
rect 4558 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4680 12872
rect 4680 12832 4682 12872
rect 4390 12790 4514 12832
rect 4558 12790 4682 12832
rect 16390 12872 16514 12914
rect 16558 12872 16682 12914
rect 16390 12832 16392 12872
rect 16392 12832 16434 12872
rect 16434 12832 16474 12872
rect 16474 12832 16514 12872
rect 16558 12832 16598 12872
rect 16598 12832 16638 12872
rect 16638 12832 16680 12872
rect 16680 12832 16682 12872
rect 16390 12790 16514 12832
rect 16558 12790 16682 12832
rect 28390 12872 28514 12914
rect 28558 12872 28682 12914
rect 28390 12832 28392 12872
rect 28392 12832 28434 12872
rect 28434 12832 28474 12872
rect 28474 12832 28514 12872
rect 28558 12832 28598 12872
rect 28598 12832 28638 12872
rect 28638 12832 28680 12872
rect 28680 12832 28682 12872
rect 28390 12790 28514 12832
rect 28558 12790 28682 12832
rect 40390 12872 40514 12914
rect 40558 12872 40682 12914
rect 40390 12832 40392 12872
rect 40392 12832 40434 12872
rect 40434 12832 40474 12872
rect 40474 12832 40514 12872
rect 40558 12832 40598 12872
rect 40598 12832 40638 12872
rect 40638 12832 40680 12872
rect 40680 12832 40682 12872
rect 40390 12790 40514 12832
rect 40558 12790 40682 12832
rect 52390 12872 52514 12914
rect 52558 12872 52682 12914
rect 52390 12832 52392 12872
rect 52392 12832 52434 12872
rect 52434 12832 52474 12872
rect 52474 12832 52514 12872
rect 52558 12832 52598 12872
rect 52598 12832 52638 12872
rect 52638 12832 52680 12872
rect 52680 12832 52682 12872
rect 52390 12790 52514 12832
rect 52558 12790 52682 12832
rect 64390 12872 64514 12914
rect 64558 12872 64682 12914
rect 64390 12832 64392 12872
rect 64392 12832 64434 12872
rect 64434 12832 64474 12872
rect 64474 12832 64514 12872
rect 64558 12832 64598 12872
rect 64598 12832 64638 12872
rect 64638 12832 64680 12872
rect 64680 12832 64682 12872
rect 64390 12790 64514 12832
rect 64558 12790 64682 12832
rect 76390 12872 76514 12914
rect 76558 12872 76682 12914
rect 76390 12832 76392 12872
rect 76392 12832 76434 12872
rect 76434 12832 76474 12872
rect 76474 12832 76514 12872
rect 76558 12832 76598 12872
rect 76598 12832 76638 12872
rect 76638 12832 76680 12872
rect 76680 12832 76682 12872
rect 76390 12790 76514 12832
rect 76558 12790 76682 12832
rect 3150 12116 3274 12158
rect 3318 12116 3442 12158
rect 3150 12076 3152 12116
rect 3152 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3274 12116
rect 3318 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3440 12116
rect 3440 12076 3442 12116
rect 3150 12034 3274 12076
rect 3318 12034 3442 12076
rect 15150 12116 15274 12158
rect 15318 12116 15442 12158
rect 15150 12076 15152 12116
rect 15152 12076 15194 12116
rect 15194 12076 15234 12116
rect 15234 12076 15274 12116
rect 15318 12076 15358 12116
rect 15358 12076 15398 12116
rect 15398 12076 15440 12116
rect 15440 12076 15442 12116
rect 15150 12034 15274 12076
rect 15318 12034 15442 12076
rect 27150 12116 27274 12158
rect 27318 12116 27442 12158
rect 27150 12076 27152 12116
rect 27152 12076 27194 12116
rect 27194 12076 27234 12116
rect 27234 12076 27274 12116
rect 27318 12076 27358 12116
rect 27358 12076 27398 12116
rect 27398 12076 27440 12116
rect 27440 12076 27442 12116
rect 27150 12034 27274 12076
rect 27318 12034 27442 12076
rect 39150 12116 39274 12158
rect 39318 12116 39442 12158
rect 39150 12076 39152 12116
rect 39152 12076 39194 12116
rect 39194 12076 39234 12116
rect 39234 12076 39274 12116
rect 39318 12076 39358 12116
rect 39358 12076 39398 12116
rect 39398 12076 39440 12116
rect 39440 12076 39442 12116
rect 39150 12034 39274 12076
rect 39318 12034 39442 12076
rect 51150 12116 51274 12158
rect 51318 12116 51442 12158
rect 51150 12076 51152 12116
rect 51152 12076 51194 12116
rect 51194 12076 51234 12116
rect 51234 12076 51274 12116
rect 51318 12076 51358 12116
rect 51358 12076 51398 12116
rect 51398 12076 51440 12116
rect 51440 12076 51442 12116
rect 51150 12034 51274 12076
rect 51318 12034 51442 12076
rect 63150 12116 63274 12158
rect 63318 12116 63442 12158
rect 63150 12076 63152 12116
rect 63152 12076 63194 12116
rect 63194 12076 63234 12116
rect 63234 12076 63274 12116
rect 63318 12076 63358 12116
rect 63358 12076 63398 12116
rect 63398 12076 63440 12116
rect 63440 12076 63442 12116
rect 63150 12034 63274 12076
rect 63318 12034 63442 12076
rect 75150 12116 75274 12158
rect 75318 12116 75442 12158
rect 75150 12076 75152 12116
rect 75152 12076 75194 12116
rect 75194 12076 75234 12116
rect 75234 12076 75274 12116
rect 75318 12076 75358 12116
rect 75358 12076 75398 12116
rect 75398 12076 75440 12116
rect 75440 12076 75442 12116
rect 75150 12034 75274 12076
rect 75318 12034 75442 12076
rect 4390 11360 4514 11402
rect 4558 11360 4682 11402
rect 4390 11320 4392 11360
rect 4392 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4514 11360
rect 4558 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4680 11360
rect 4680 11320 4682 11360
rect 4390 11278 4514 11320
rect 4558 11278 4682 11320
rect 16390 11360 16514 11402
rect 16558 11360 16682 11402
rect 16390 11320 16392 11360
rect 16392 11320 16434 11360
rect 16434 11320 16474 11360
rect 16474 11320 16514 11360
rect 16558 11320 16598 11360
rect 16598 11320 16638 11360
rect 16638 11320 16680 11360
rect 16680 11320 16682 11360
rect 16390 11278 16514 11320
rect 16558 11278 16682 11320
rect 28390 11360 28514 11402
rect 28558 11360 28682 11402
rect 28390 11320 28392 11360
rect 28392 11320 28434 11360
rect 28434 11320 28474 11360
rect 28474 11320 28514 11360
rect 28558 11320 28598 11360
rect 28598 11320 28638 11360
rect 28638 11320 28680 11360
rect 28680 11320 28682 11360
rect 28390 11278 28514 11320
rect 28558 11278 28682 11320
rect 40390 11360 40514 11402
rect 40558 11360 40682 11402
rect 40390 11320 40392 11360
rect 40392 11320 40434 11360
rect 40434 11320 40474 11360
rect 40474 11320 40514 11360
rect 40558 11320 40598 11360
rect 40598 11320 40638 11360
rect 40638 11320 40680 11360
rect 40680 11320 40682 11360
rect 40390 11278 40514 11320
rect 40558 11278 40682 11320
rect 52390 11360 52514 11402
rect 52558 11360 52682 11402
rect 52390 11320 52392 11360
rect 52392 11320 52434 11360
rect 52434 11320 52474 11360
rect 52474 11320 52514 11360
rect 52558 11320 52598 11360
rect 52598 11320 52638 11360
rect 52638 11320 52680 11360
rect 52680 11320 52682 11360
rect 52390 11278 52514 11320
rect 52558 11278 52682 11320
rect 64390 11360 64514 11402
rect 64558 11360 64682 11402
rect 64390 11320 64392 11360
rect 64392 11320 64434 11360
rect 64434 11320 64474 11360
rect 64474 11320 64514 11360
rect 64558 11320 64598 11360
rect 64598 11320 64638 11360
rect 64638 11320 64680 11360
rect 64680 11320 64682 11360
rect 64390 11278 64514 11320
rect 64558 11278 64682 11320
rect 76390 11360 76514 11402
rect 76558 11360 76682 11402
rect 76390 11320 76392 11360
rect 76392 11320 76434 11360
rect 76434 11320 76474 11360
rect 76474 11320 76514 11360
rect 76558 11320 76598 11360
rect 76598 11320 76638 11360
rect 76638 11320 76680 11360
rect 76680 11320 76682 11360
rect 76390 11278 76514 11320
rect 76558 11278 76682 11320
rect 3150 10604 3274 10646
rect 3318 10604 3442 10646
rect 3150 10564 3152 10604
rect 3152 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3274 10604
rect 3318 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3440 10604
rect 3440 10564 3442 10604
rect 3150 10522 3274 10564
rect 3318 10522 3442 10564
rect 15150 10604 15274 10646
rect 15318 10604 15442 10646
rect 15150 10564 15152 10604
rect 15152 10564 15194 10604
rect 15194 10564 15234 10604
rect 15234 10564 15274 10604
rect 15318 10564 15358 10604
rect 15358 10564 15398 10604
rect 15398 10564 15440 10604
rect 15440 10564 15442 10604
rect 15150 10522 15274 10564
rect 15318 10522 15442 10564
rect 27150 10604 27274 10646
rect 27318 10604 27442 10646
rect 27150 10564 27152 10604
rect 27152 10564 27194 10604
rect 27194 10564 27234 10604
rect 27234 10564 27274 10604
rect 27318 10564 27358 10604
rect 27358 10564 27398 10604
rect 27398 10564 27440 10604
rect 27440 10564 27442 10604
rect 27150 10522 27274 10564
rect 27318 10522 27442 10564
rect 39150 10604 39274 10646
rect 39318 10604 39442 10646
rect 39150 10564 39152 10604
rect 39152 10564 39194 10604
rect 39194 10564 39234 10604
rect 39234 10564 39274 10604
rect 39318 10564 39358 10604
rect 39358 10564 39398 10604
rect 39398 10564 39440 10604
rect 39440 10564 39442 10604
rect 39150 10522 39274 10564
rect 39318 10522 39442 10564
rect 51150 10604 51274 10646
rect 51318 10604 51442 10646
rect 51150 10564 51152 10604
rect 51152 10564 51194 10604
rect 51194 10564 51234 10604
rect 51234 10564 51274 10604
rect 51318 10564 51358 10604
rect 51358 10564 51398 10604
rect 51398 10564 51440 10604
rect 51440 10564 51442 10604
rect 51150 10522 51274 10564
rect 51318 10522 51442 10564
rect 63150 10604 63274 10646
rect 63318 10604 63442 10646
rect 63150 10564 63152 10604
rect 63152 10564 63194 10604
rect 63194 10564 63234 10604
rect 63234 10564 63274 10604
rect 63318 10564 63358 10604
rect 63358 10564 63398 10604
rect 63398 10564 63440 10604
rect 63440 10564 63442 10604
rect 63150 10522 63274 10564
rect 63318 10522 63442 10564
rect 75150 10604 75274 10646
rect 75318 10604 75442 10646
rect 75150 10564 75152 10604
rect 75152 10564 75194 10604
rect 75194 10564 75234 10604
rect 75234 10564 75274 10604
rect 75318 10564 75358 10604
rect 75358 10564 75398 10604
rect 75398 10564 75440 10604
rect 75440 10564 75442 10604
rect 75150 10522 75274 10564
rect 75318 10522 75442 10564
rect 4390 9848 4514 9890
rect 4558 9848 4682 9890
rect 4390 9808 4392 9848
rect 4392 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4514 9848
rect 4558 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4680 9848
rect 4680 9808 4682 9848
rect 4390 9766 4514 9808
rect 4558 9766 4682 9808
rect 16390 9848 16514 9890
rect 16558 9848 16682 9890
rect 16390 9808 16392 9848
rect 16392 9808 16434 9848
rect 16434 9808 16474 9848
rect 16474 9808 16514 9848
rect 16558 9808 16598 9848
rect 16598 9808 16638 9848
rect 16638 9808 16680 9848
rect 16680 9808 16682 9848
rect 16390 9766 16514 9808
rect 16558 9766 16682 9808
rect 28390 9848 28514 9890
rect 28558 9848 28682 9890
rect 28390 9808 28392 9848
rect 28392 9808 28434 9848
rect 28434 9808 28474 9848
rect 28474 9808 28514 9848
rect 28558 9808 28598 9848
rect 28598 9808 28638 9848
rect 28638 9808 28680 9848
rect 28680 9808 28682 9848
rect 28390 9766 28514 9808
rect 28558 9766 28682 9808
rect 40390 9848 40514 9890
rect 40558 9848 40682 9890
rect 40390 9808 40392 9848
rect 40392 9808 40434 9848
rect 40434 9808 40474 9848
rect 40474 9808 40514 9848
rect 40558 9808 40598 9848
rect 40598 9808 40638 9848
rect 40638 9808 40680 9848
rect 40680 9808 40682 9848
rect 40390 9766 40514 9808
rect 40558 9766 40682 9808
rect 52390 9848 52514 9890
rect 52558 9848 52682 9890
rect 52390 9808 52392 9848
rect 52392 9808 52434 9848
rect 52434 9808 52474 9848
rect 52474 9808 52514 9848
rect 52558 9808 52598 9848
rect 52598 9808 52638 9848
rect 52638 9808 52680 9848
rect 52680 9808 52682 9848
rect 52390 9766 52514 9808
rect 52558 9766 52682 9808
rect 64390 9848 64514 9890
rect 64558 9848 64682 9890
rect 64390 9808 64392 9848
rect 64392 9808 64434 9848
rect 64434 9808 64474 9848
rect 64474 9808 64514 9848
rect 64558 9808 64598 9848
rect 64598 9808 64638 9848
rect 64638 9808 64680 9848
rect 64680 9808 64682 9848
rect 64390 9766 64514 9808
rect 64558 9766 64682 9808
rect 76390 9848 76514 9890
rect 76558 9848 76682 9890
rect 76390 9808 76392 9848
rect 76392 9808 76434 9848
rect 76434 9808 76474 9848
rect 76474 9808 76514 9848
rect 76558 9808 76598 9848
rect 76598 9808 76638 9848
rect 76638 9808 76680 9848
rect 76680 9808 76682 9848
rect 76390 9766 76514 9808
rect 76558 9766 76682 9808
rect 3150 9092 3274 9134
rect 3318 9092 3442 9134
rect 3150 9052 3152 9092
rect 3152 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3274 9092
rect 3318 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3440 9092
rect 3440 9052 3442 9092
rect 3150 9010 3274 9052
rect 3318 9010 3442 9052
rect 15150 9092 15274 9134
rect 15318 9092 15442 9134
rect 15150 9052 15152 9092
rect 15152 9052 15194 9092
rect 15194 9052 15234 9092
rect 15234 9052 15274 9092
rect 15318 9052 15358 9092
rect 15358 9052 15398 9092
rect 15398 9052 15440 9092
rect 15440 9052 15442 9092
rect 15150 9010 15274 9052
rect 15318 9010 15442 9052
rect 27150 9092 27274 9134
rect 27318 9092 27442 9134
rect 27150 9052 27152 9092
rect 27152 9052 27194 9092
rect 27194 9052 27234 9092
rect 27234 9052 27274 9092
rect 27318 9052 27358 9092
rect 27358 9052 27398 9092
rect 27398 9052 27440 9092
rect 27440 9052 27442 9092
rect 27150 9010 27274 9052
rect 27318 9010 27442 9052
rect 39150 9092 39274 9134
rect 39318 9092 39442 9134
rect 39150 9052 39152 9092
rect 39152 9052 39194 9092
rect 39194 9052 39234 9092
rect 39234 9052 39274 9092
rect 39318 9052 39358 9092
rect 39358 9052 39398 9092
rect 39398 9052 39440 9092
rect 39440 9052 39442 9092
rect 39150 9010 39274 9052
rect 39318 9010 39442 9052
rect 51150 9092 51274 9134
rect 51318 9092 51442 9134
rect 51150 9052 51152 9092
rect 51152 9052 51194 9092
rect 51194 9052 51234 9092
rect 51234 9052 51274 9092
rect 51318 9052 51358 9092
rect 51358 9052 51398 9092
rect 51398 9052 51440 9092
rect 51440 9052 51442 9092
rect 51150 9010 51274 9052
rect 51318 9010 51442 9052
rect 63150 9092 63274 9134
rect 63318 9092 63442 9134
rect 63150 9052 63152 9092
rect 63152 9052 63194 9092
rect 63194 9052 63234 9092
rect 63234 9052 63274 9092
rect 63318 9052 63358 9092
rect 63358 9052 63398 9092
rect 63398 9052 63440 9092
rect 63440 9052 63442 9092
rect 63150 9010 63274 9052
rect 63318 9010 63442 9052
rect 75150 9092 75274 9134
rect 75318 9092 75442 9134
rect 75150 9052 75152 9092
rect 75152 9052 75194 9092
rect 75194 9052 75234 9092
rect 75234 9052 75274 9092
rect 75318 9052 75358 9092
rect 75358 9052 75398 9092
rect 75398 9052 75440 9092
rect 75440 9052 75442 9092
rect 75150 9010 75274 9052
rect 75318 9010 75442 9052
rect 4390 8336 4514 8378
rect 4558 8336 4682 8378
rect 4390 8296 4392 8336
rect 4392 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4514 8336
rect 4558 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4680 8336
rect 4680 8296 4682 8336
rect 4390 8254 4514 8296
rect 4558 8254 4682 8296
rect 16390 8336 16514 8378
rect 16558 8336 16682 8378
rect 16390 8296 16392 8336
rect 16392 8296 16434 8336
rect 16434 8296 16474 8336
rect 16474 8296 16514 8336
rect 16558 8296 16598 8336
rect 16598 8296 16638 8336
rect 16638 8296 16680 8336
rect 16680 8296 16682 8336
rect 16390 8254 16514 8296
rect 16558 8254 16682 8296
rect 28390 8336 28514 8378
rect 28558 8336 28682 8378
rect 28390 8296 28392 8336
rect 28392 8296 28434 8336
rect 28434 8296 28474 8336
rect 28474 8296 28514 8336
rect 28558 8296 28598 8336
rect 28598 8296 28638 8336
rect 28638 8296 28680 8336
rect 28680 8296 28682 8336
rect 28390 8254 28514 8296
rect 28558 8254 28682 8296
rect 40390 8336 40514 8378
rect 40558 8336 40682 8378
rect 40390 8296 40392 8336
rect 40392 8296 40434 8336
rect 40434 8296 40474 8336
rect 40474 8296 40514 8336
rect 40558 8296 40598 8336
rect 40598 8296 40638 8336
rect 40638 8296 40680 8336
rect 40680 8296 40682 8336
rect 40390 8254 40514 8296
rect 40558 8254 40682 8296
rect 52390 8336 52514 8378
rect 52558 8336 52682 8378
rect 52390 8296 52392 8336
rect 52392 8296 52434 8336
rect 52434 8296 52474 8336
rect 52474 8296 52514 8336
rect 52558 8296 52598 8336
rect 52598 8296 52638 8336
rect 52638 8296 52680 8336
rect 52680 8296 52682 8336
rect 52390 8254 52514 8296
rect 52558 8254 52682 8296
rect 64390 8336 64514 8378
rect 64558 8336 64682 8378
rect 64390 8296 64392 8336
rect 64392 8296 64434 8336
rect 64434 8296 64474 8336
rect 64474 8296 64514 8336
rect 64558 8296 64598 8336
rect 64598 8296 64638 8336
rect 64638 8296 64680 8336
rect 64680 8296 64682 8336
rect 64390 8254 64514 8296
rect 64558 8254 64682 8296
rect 76390 8336 76514 8378
rect 76558 8336 76682 8378
rect 76390 8296 76392 8336
rect 76392 8296 76434 8336
rect 76434 8296 76474 8336
rect 76474 8296 76514 8336
rect 76558 8296 76598 8336
rect 76598 8296 76638 8336
rect 76638 8296 76680 8336
rect 76680 8296 76682 8336
rect 76390 8254 76514 8296
rect 76558 8254 76682 8296
rect 3150 7580 3274 7622
rect 3318 7580 3442 7622
rect 3150 7540 3152 7580
rect 3152 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3274 7580
rect 3318 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3440 7580
rect 3440 7540 3442 7580
rect 3150 7498 3274 7540
rect 3318 7498 3442 7540
rect 15150 7580 15274 7622
rect 15318 7580 15442 7622
rect 15150 7540 15152 7580
rect 15152 7540 15194 7580
rect 15194 7540 15234 7580
rect 15234 7540 15274 7580
rect 15318 7540 15358 7580
rect 15358 7540 15398 7580
rect 15398 7540 15440 7580
rect 15440 7540 15442 7580
rect 15150 7498 15274 7540
rect 15318 7498 15442 7540
rect 27150 7580 27274 7622
rect 27318 7580 27442 7622
rect 27150 7540 27152 7580
rect 27152 7540 27194 7580
rect 27194 7540 27234 7580
rect 27234 7540 27274 7580
rect 27318 7540 27358 7580
rect 27358 7540 27398 7580
rect 27398 7540 27440 7580
rect 27440 7540 27442 7580
rect 27150 7498 27274 7540
rect 27318 7498 27442 7540
rect 39150 7580 39274 7622
rect 39318 7580 39442 7622
rect 39150 7540 39152 7580
rect 39152 7540 39194 7580
rect 39194 7540 39234 7580
rect 39234 7540 39274 7580
rect 39318 7540 39358 7580
rect 39358 7540 39398 7580
rect 39398 7540 39440 7580
rect 39440 7540 39442 7580
rect 39150 7498 39274 7540
rect 39318 7498 39442 7540
rect 51150 7580 51274 7622
rect 51318 7580 51442 7622
rect 51150 7540 51152 7580
rect 51152 7540 51194 7580
rect 51194 7540 51234 7580
rect 51234 7540 51274 7580
rect 51318 7540 51358 7580
rect 51358 7540 51398 7580
rect 51398 7540 51440 7580
rect 51440 7540 51442 7580
rect 51150 7498 51274 7540
rect 51318 7498 51442 7540
rect 63150 7580 63274 7622
rect 63318 7580 63442 7622
rect 63150 7540 63152 7580
rect 63152 7540 63194 7580
rect 63194 7540 63234 7580
rect 63234 7540 63274 7580
rect 63318 7540 63358 7580
rect 63358 7540 63398 7580
rect 63398 7540 63440 7580
rect 63440 7540 63442 7580
rect 63150 7498 63274 7540
rect 63318 7498 63442 7540
rect 75150 7580 75274 7622
rect 75318 7580 75442 7622
rect 75150 7540 75152 7580
rect 75152 7540 75194 7580
rect 75194 7540 75234 7580
rect 75234 7540 75274 7580
rect 75318 7540 75358 7580
rect 75358 7540 75398 7580
rect 75398 7540 75440 7580
rect 75440 7540 75442 7580
rect 75150 7498 75274 7540
rect 75318 7498 75442 7540
rect 4390 6824 4514 6866
rect 4558 6824 4682 6866
rect 4390 6784 4392 6824
rect 4392 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4514 6824
rect 4558 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4680 6824
rect 4680 6784 4682 6824
rect 4390 6742 4514 6784
rect 4558 6742 4682 6784
rect 16390 6824 16514 6866
rect 16558 6824 16682 6866
rect 16390 6784 16392 6824
rect 16392 6784 16434 6824
rect 16434 6784 16474 6824
rect 16474 6784 16514 6824
rect 16558 6784 16598 6824
rect 16598 6784 16638 6824
rect 16638 6784 16680 6824
rect 16680 6784 16682 6824
rect 16390 6742 16514 6784
rect 16558 6742 16682 6784
rect 28390 6824 28514 6866
rect 28558 6824 28682 6866
rect 28390 6784 28392 6824
rect 28392 6784 28434 6824
rect 28434 6784 28474 6824
rect 28474 6784 28514 6824
rect 28558 6784 28598 6824
rect 28598 6784 28638 6824
rect 28638 6784 28680 6824
rect 28680 6784 28682 6824
rect 28390 6742 28514 6784
rect 28558 6742 28682 6784
rect 40390 6824 40514 6866
rect 40558 6824 40682 6866
rect 40390 6784 40392 6824
rect 40392 6784 40434 6824
rect 40434 6784 40474 6824
rect 40474 6784 40514 6824
rect 40558 6784 40598 6824
rect 40598 6784 40638 6824
rect 40638 6784 40680 6824
rect 40680 6784 40682 6824
rect 40390 6742 40514 6784
rect 40558 6742 40682 6784
rect 52390 6824 52514 6866
rect 52558 6824 52682 6866
rect 52390 6784 52392 6824
rect 52392 6784 52434 6824
rect 52434 6784 52474 6824
rect 52474 6784 52514 6824
rect 52558 6784 52598 6824
rect 52598 6784 52638 6824
rect 52638 6784 52680 6824
rect 52680 6784 52682 6824
rect 52390 6742 52514 6784
rect 52558 6742 52682 6784
rect 64390 6824 64514 6866
rect 64558 6824 64682 6866
rect 64390 6784 64392 6824
rect 64392 6784 64434 6824
rect 64434 6784 64474 6824
rect 64474 6784 64514 6824
rect 64558 6784 64598 6824
rect 64598 6784 64638 6824
rect 64638 6784 64680 6824
rect 64680 6784 64682 6824
rect 64390 6742 64514 6784
rect 64558 6742 64682 6784
rect 76390 6824 76514 6866
rect 76558 6824 76682 6866
rect 76390 6784 76392 6824
rect 76392 6784 76434 6824
rect 76434 6784 76474 6824
rect 76474 6784 76514 6824
rect 76558 6784 76598 6824
rect 76598 6784 76638 6824
rect 76638 6784 76680 6824
rect 76680 6784 76682 6824
rect 76390 6742 76514 6784
rect 76558 6742 76682 6784
rect 3150 6068 3274 6110
rect 3318 6068 3442 6110
rect 3150 6028 3152 6068
rect 3152 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3274 6068
rect 3318 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3440 6068
rect 3440 6028 3442 6068
rect 3150 5986 3274 6028
rect 3318 5986 3442 6028
rect 15150 6068 15274 6110
rect 15318 6068 15442 6110
rect 15150 6028 15152 6068
rect 15152 6028 15194 6068
rect 15194 6028 15234 6068
rect 15234 6028 15274 6068
rect 15318 6028 15358 6068
rect 15358 6028 15398 6068
rect 15398 6028 15440 6068
rect 15440 6028 15442 6068
rect 15150 5986 15274 6028
rect 15318 5986 15442 6028
rect 27150 6068 27274 6110
rect 27318 6068 27442 6110
rect 27150 6028 27152 6068
rect 27152 6028 27194 6068
rect 27194 6028 27234 6068
rect 27234 6028 27274 6068
rect 27318 6028 27358 6068
rect 27358 6028 27398 6068
rect 27398 6028 27440 6068
rect 27440 6028 27442 6068
rect 27150 5986 27274 6028
rect 27318 5986 27442 6028
rect 39150 6068 39274 6110
rect 39318 6068 39442 6110
rect 39150 6028 39152 6068
rect 39152 6028 39194 6068
rect 39194 6028 39234 6068
rect 39234 6028 39274 6068
rect 39318 6028 39358 6068
rect 39358 6028 39398 6068
rect 39398 6028 39440 6068
rect 39440 6028 39442 6068
rect 39150 5986 39274 6028
rect 39318 5986 39442 6028
rect 51150 6068 51274 6110
rect 51318 6068 51442 6110
rect 51150 6028 51152 6068
rect 51152 6028 51194 6068
rect 51194 6028 51234 6068
rect 51234 6028 51274 6068
rect 51318 6028 51358 6068
rect 51358 6028 51398 6068
rect 51398 6028 51440 6068
rect 51440 6028 51442 6068
rect 51150 5986 51274 6028
rect 51318 5986 51442 6028
rect 63150 6068 63274 6110
rect 63318 6068 63442 6110
rect 63150 6028 63152 6068
rect 63152 6028 63194 6068
rect 63194 6028 63234 6068
rect 63234 6028 63274 6068
rect 63318 6028 63358 6068
rect 63358 6028 63398 6068
rect 63398 6028 63440 6068
rect 63440 6028 63442 6068
rect 63150 5986 63274 6028
rect 63318 5986 63442 6028
rect 75150 6068 75274 6110
rect 75318 6068 75442 6110
rect 75150 6028 75152 6068
rect 75152 6028 75194 6068
rect 75194 6028 75234 6068
rect 75234 6028 75274 6068
rect 75318 6028 75358 6068
rect 75358 6028 75398 6068
rect 75398 6028 75440 6068
rect 75440 6028 75442 6068
rect 75150 5986 75274 6028
rect 75318 5986 75442 6028
rect 4390 5312 4514 5354
rect 4558 5312 4682 5354
rect 4390 5272 4392 5312
rect 4392 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4514 5312
rect 4558 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4680 5312
rect 4680 5272 4682 5312
rect 4390 5230 4514 5272
rect 4558 5230 4682 5272
rect 16390 5312 16514 5354
rect 16558 5312 16682 5354
rect 16390 5272 16392 5312
rect 16392 5272 16434 5312
rect 16434 5272 16474 5312
rect 16474 5272 16514 5312
rect 16558 5272 16598 5312
rect 16598 5272 16638 5312
rect 16638 5272 16680 5312
rect 16680 5272 16682 5312
rect 16390 5230 16514 5272
rect 16558 5230 16682 5272
rect 28390 5312 28514 5354
rect 28558 5312 28682 5354
rect 28390 5272 28392 5312
rect 28392 5272 28434 5312
rect 28434 5272 28474 5312
rect 28474 5272 28514 5312
rect 28558 5272 28598 5312
rect 28598 5272 28638 5312
rect 28638 5272 28680 5312
rect 28680 5272 28682 5312
rect 28390 5230 28514 5272
rect 28558 5230 28682 5272
rect 40390 5312 40514 5354
rect 40558 5312 40682 5354
rect 40390 5272 40392 5312
rect 40392 5272 40434 5312
rect 40434 5272 40474 5312
rect 40474 5272 40514 5312
rect 40558 5272 40598 5312
rect 40598 5272 40638 5312
rect 40638 5272 40680 5312
rect 40680 5272 40682 5312
rect 40390 5230 40514 5272
rect 40558 5230 40682 5272
rect 52390 5312 52514 5354
rect 52558 5312 52682 5354
rect 52390 5272 52392 5312
rect 52392 5272 52434 5312
rect 52434 5272 52474 5312
rect 52474 5272 52514 5312
rect 52558 5272 52598 5312
rect 52598 5272 52638 5312
rect 52638 5272 52680 5312
rect 52680 5272 52682 5312
rect 52390 5230 52514 5272
rect 52558 5230 52682 5272
rect 64390 5312 64514 5354
rect 64558 5312 64682 5354
rect 64390 5272 64392 5312
rect 64392 5272 64434 5312
rect 64434 5272 64474 5312
rect 64474 5272 64514 5312
rect 64558 5272 64598 5312
rect 64598 5272 64638 5312
rect 64638 5272 64680 5312
rect 64680 5272 64682 5312
rect 64390 5230 64514 5272
rect 64558 5230 64682 5272
rect 76390 5312 76514 5354
rect 76558 5312 76682 5354
rect 76390 5272 76392 5312
rect 76392 5272 76434 5312
rect 76434 5272 76474 5312
rect 76474 5272 76514 5312
rect 76558 5272 76598 5312
rect 76598 5272 76638 5312
rect 76638 5272 76680 5312
rect 76680 5272 76682 5312
rect 76390 5230 76514 5272
rect 76558 5230 76682 5272
rect 3150 4556 3274 4598
rect 3318 4556 3442 4598
rect 3150 4516 3152 4556
rect 3152 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3274 4556
rect 3318 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3440 4556
rect 3440 4516 3442 4556
rect 3150 4474 3274 4516
rect 3318 4474 3442 4516
rect 15150 4556 15274 4598
rect 15318 4556 15442 4598
rect 15150 4516 15152 4556
rect 15152 4516 15194 4556
rect 15194 4516 15234 4556
rect 15234 4516 15274 4556
rect 15318 4516 15358 4556
rect 15358 4516 15398 4556
rect 15398 4516 15440 4556
rect 15440 4516 15442 4556
rect 15150 4474 15274 4516
rect 15318 4474 15442 4516
rect 27150 4556 27274 4598
rect 27318 4556 27442 4598
rect 27150 4516 27152 4556
rect 27152 4516 27194 4556
rect 27194 4516 27234 4556
rect 27234 4516 27274 4556
rect 27318 4516 27358 4556
rect 27358 4516 27398 4556
rect 27398 4516 27440 4556
rect 27440 4516 27442 4556
rect 27150 4474 27274 4516
rect 27318 4474 27442 4516
rect 39150 4556 39274 4598
rect 39318 4556 39442 4598
rect 39150 4516 39152 4556
rect 39152 4516 39194 4556
rect 39194 4516 39234 4556
rect 39234 4516 39274 4556
rect 39318 4516 39358 4556
rect 39358 4516 39398 4556
rect 39398 4516 39440 4556
rect 39440 4516 39442 4556
rect 39150 4474 39274 4516
rect 39318 4474 39442 4516
rect 51150 4556 51274 4598
rect 51318 4556 51442 4598
rect 51150 4516 51152 4556
rect 51152 4516 51194 4556
rect 51194 4516 51234 4556
rect 51234 4516 51274 4556
rect 51318 4516 51358 4556
rect 51358 4516 51398 4556
rect 51398 4516 51440 4556
rect 51440 4516 51442 4556
rect 51150 4474 51274 4516
rect 51318 4474 51442 4516
rect 63150 4556 63274 4598
rect 63318 4556 63442 4598
rect 63150 4516 63152 4556
rect 63152 4516 63194 4556
rect 63194 4516 63234 4556
rect 63234 4516 63274 4556
rect 63318 4516 63358 4556
rect 63358 4516 63398 4556
rect 63398 4516 63440 4556
rect 63440 4516 63442 4556
rect 63150 4474 63274 4516
rect 63318 4474 63442 4516
rect 75150 4556 75274 4598
rect 75318 4556 75442 4598
rect 75150 4516 75152 4556
rect 75152 4516 75194 4556
rect 75194 4516 75234 4556
rect 75234 4516 75274 4556
rect 75318 4516 75358 4556
rect 75358 4516 75398 4556
rect 75398 4516 75440 4556
rect 75440 4516 75442 4556
rect 75150 4474 75274 4516
rect 75318 4474 75442 4516
rect 4390 3800 4514 3842
rect 4558 3800 4682 3842
rect 4390 3760 4392 3800
rect 4392 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4514 3800
rect 4558 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4680 3800
rect 4680 3760 4682 3800
rect 4390 3718 4514 3760
rect 4558 3718 4682 3760
rect 16390 3800 16514 3842
rect 16558 3800 16682 3842
rect 16390 3760 16392 3800
rect 16392 3760 16434 3800
rect 16434 3760 16474 3800
rect 16474 3760 16514 3800
rect 16558 3760 16598 3800
rect 16598 3760 16638 3800
rect 16638 3760 16680 3800
rect 16680 3760 16682 3800
rect 16390 3718 16514 3760
rect 16558 3718 16682 3760
rect 28390 3800 28514 3842
rect 28558 3800 28682 3842
rect 28390 3760 28392 3800
rect 28392 3760 28434 3800
rect 28434 3760 28474 3800
rect 28474 3760 28514 3800
rect 28558 3760 28598 3800
rect 28598 3760 28638 3800
rect 28638 3760 28680 3800
rect 28680 3760 28682 3800
rect 28390 3718 28514 3760
rect 28558 3718 28682 3760
rect 40390 3800 40514 3842
rect 40558 3800 40682 3842
rect 40390 3760 40392 3800
rect 40392 3760 40434 3800
rect 40434 3760 40474 3800
rect 40474 3760 40514 3800
rect 40558 3760 40598 3800
rect 40598 3760 40638 3800
rect 40638 3760 40680 3800
rect 40680 3760 40682 3800
rect 40390 3718 40514 3760
rect 40558 3718 40682 3760
rect 52390 3800 52514 3842
rect 52558 3800 52682 3842
rect 52390 3760 52392 3800
rect 52392 3760 52434 3800
rect 52434 3760 52474 3800
rect 52474 3760 52514 3800
rect 52558 3760 52598 3800
rect 52598 3760 52638 3800
rect 52638 3760 52680 3800
rect 52680 3760 52682 3800
rect 52390 3718 52514 3760
rect 52558 3718 52682 3760
rect 64390 3800 64514 3842
rect 64558 3800 64682 3842
rect 64390 3760 64392 3800
rect 64392 3760 64434 3800
rect 64434 3760 64474 3800
rect 64474 3760 64514 3800
rect 64558 3760 64598 3800
rect 64598 3760 64638 3800
rect 64638 3760 64680 3800
rect 64680 3760 64682 3800
rect 64390 3718 64514 3760
rect 64558 3718 64682 3760
rect 76390 3800 76514 3842
rect 76558 3800 76682 3842
rect 76390 3760 76392 3800
rect 76392 3760 76434 3800
rect 76434 3760 76474 3800
rect 76474 3760 76514 3800
rect 76558 3760 76598 3800
rect 76598 3760 76638 3800
rect 76638 3760 76680 3800
rect 76680 3760 76682 3800
rect 76390 3718 76514 3760
rect 76558 3718 76682 3760
rect 3150 3044 3274 3086
rect 3318 3044 3442 3086
rect 3150 3004 3152 3044
rect 3152 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3274 3044
rect 3318 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3440 3044
rect 3440 3004 3442 3044
rect 3150 2962 3274 3004
rect 3318 2962 3442 3004
rect 15150 3044 15274 3086
rect 15318 3044 15442 3086
rect 15150 3004 15152 3044
rect 15152 3004 15194 3044
rect 15194 3004 15234 3044
rect 15234 3004 15274 3044
rect 15318 3004 15358 3044
rect 15358 3004 15398 3044
rect 15398 3004 15440 3044
rect 15440 3004 15442 3044
rect 15150 2962 15274 3004
rect 15318 2962 15442 3004
rect 27150 3044 27274 3086
rect 27318 3044 27442 3086
rect 27150 3004 27152 3044
rect 27152 3004 27194 3044
rect 27194 3004 27234 3044
rect 27234 3004 27274 3044
rect 27318 3004 27358 3044
rect 27358 3004 27398 3044
rect 27398 3004 27440 3044
rect 27440 3004 27442 3044
rect 27150 2962 27274 3004
rect 27318 2962 27442 3004
rect 39150 3044 39274 3086
rect 39318 3044 39442 3086
rect 39150 3004 39152 3044
rect 39152 3004 39194 3044
rect 39194 3004 39234 3044
rect 39234 3004 39274 3044
rect 39318 3004 39358 3044
rect 39358 3004 39398 3044
rect 39398 3004 39440 3044
rect 39440 3004 39442 3044
rect 39150 2962 39274 3004
rect 39318 2962 39442 3004
rect 51150 3044 51274 3086
rect 51318 3044 51442 3086
rect 51150 3004 51152 3044
rect 51152 3004 51194 3044
rect 51194 3004 51234 3044
rect 51234 3004 51274 3044
rect 51318 3004 51358 3044
rect 51358 3004 51398 3044
rect 51398 3004 51440 3044
rect 51440 3004 51442 3044
rect 51150 2962 51274 3004
rect 51318 2962 51442 3004
rect 63150 3044 63274 3086
rect 63318 3044 63442 3086
rect 63150 3004 63152 3044
rect 63152 3004 63194 3044
rect 63194 3004 63234 3044
rect 63234 3004 63274 3044
rect 63318 3004 63358 3044
rect 63358 3004 63398 3044
rect 63398 3004 63440 3044
rect 63440 3004 63442 3044
rect 63150 2962 63274 3004
rect 63318 2962 63442 3004
rect 75150 3044 75274 3086
rect 75318 3044 75442 3086
rect 75150 3004 75152 3044
rect 75152 3004 75194 3044
rect 75194 3004 75234 3044
rect 75234 3004 75274 3044
rect 75318 3004 75358 3044
rect 75358 3004 75398 3044
rect 75398 3004 75440 3044
rect 75440 3004 75442 3044
rect 75150 2962 75274 3004
rect 75318 2962 75442 3004
rect 4390 2288 4514 2330
rect 4558 2288 4682 2330
rect 4390 2248 4392 2288
rect 4392 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4514 2288
rect 4558 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4680 2288
rect 4680 2248 4682 2288
rect 4390 2206 4514 2248
rect 4558 2206 4682 2248
rect 16390 2288 16514 2330
rect 16558 2288 16682 2330
rect 16390 2248 16392 2288
rect 16392 2248 16434 2288
rect 16434 2248 16474 2288
rect 16474 2248 16514 2288
rect 16558 2248 16598 2288
rect 16598 2248 16638 2288
rect 16638 2248 16680 2288
rect 16680 2248 16682 2288
rect 16390 2206 16514 2248
rect 16558 2206 16682 2248
rect 28390 2288 28514 2330
rect 28558 2288 28682 2330
rect 28390 2248 28392 2288
rect 28392 2248 28434 2288
rect 28434 2248 28474 2288
rect 28474 2248 28514 2288
rect 28558 2248 28598 2288
rect 28598 2248 28638 2288
rect 28638 2248 28680 2288
rect 28680 2248 28682 2288
rect 28390 2206 28514 2248
rect 28558 2206 28682 2248
rect 40390 2288 40514 2330
rect 40558 2288 40682 2330
rect 40390 2248 40392 2288
rect 40392 2248 40434 2288
rect 40434 2248 40474 2288
rect 40474 2248 40514 2288
rect 40558 2248 40598 2288
rect 40598 2248 40638 2288
rect 40638 2248 40680 2288
rect 40680 2248 40682 2288
rect 40390 2206 40514 2248
rect 40558 2206 40682 2248
rect 52390 2288 52514 2330
rect 52558 2288 52682 2330
rect 52390 2248 52392 2288
rect 52392 2248 52434 2288
rect 52434 2248 52474 2288
rect 52474 2248 52514 2288
rect 52558 2248 52598 2288
rect 52598 2248 52638 2288
rect 52638 2248 52680 2288
rect 52680 2248 52682 2288
rect 52390 2206 52514 2248
rect 52558 2206 52682 2248
rect 64390 2288 64514 2330
rect 64558 2288 64682 2330
rect 64390 2248 64392 2288
rect 64392 2248 64434 2288
rect 64434 2248 64474 2288
rect 64474 2248 64514 2288
rect 64558 2248 64598 2288
rect 64598 2248 64638 2288
rect 64638 2248 64680 2288
rect 64680 2248 64682 2288
rect 64390 2206 64514 2248
rect 64558 2206 64682 2248
rect 76390 2288 76514 2330
rect 76558 2288 76682 2330
rect 76390 2248 76392 2288
rect 76392 2248 76434 2288
rect 76434 2248 76474 2288
rect 76474 2248 76514 2288
rect 76558 2248 76598 2288
rect 76598 2248 76638 2288
rect 76638 2248 76680 2288
rect 76680 2248 76682 2288
rect 76390 2206 76514 2248
rect 76558 2206 76682 2248
rect 3150 1532 3274 1574
rect 3318 1532 3442 1574
rect 3150 1492 3152 1532
rect 3152 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3274 1532
rect 3318 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3440 1532
rect 3440 1492 3442 1532
rect 3150 1450 3274 1492
rect 3318 1450 3442 1492
rect 15150 1532 15274 1574
rect 15318 1532 15442 1574
rect 15150 1492 15152 1532
rect 15152 1492 15194 1532
rect 15194 1492 15234 1532
rect 15234 1492 15274 1532
rect 15318 1492 15358 1532
rect 15358 1492 15398 1532
rect 15398 1492 15440 1532
rect 15440 1492 15442 1532
rect 15150 1450 15274 1492
rect 15318 1450 15442 1492
rect 27150 1532 27274 1574
rect 27318 1532 27442 1574
rect 27150 1492 27152 1532
rect 27152 1492 27194 1532
rect 27194 1492 27234 1532
rect 27234 1492 27274 1532
rect 27318 1492 27358 1532
rect 27358 1492 27398 1532
rect 27398 1492 27440 1532
rect 27440 1492 27442 1532
rect 27150 1450 27274 1492
rect 27318 1450 27442 1492
rect 39150 1532 39274 1574
rect 39318 1532 39442 1574
rect 39150 1492 39152 1532
rect 39152 1492 39194 1532
rect 39194 1492 39234 1532
rect 39234 1492 39274 1532
rect 39318 1492 39358 1532
rect 39358 1492 39398 1532
rect 39398 1492 39440 1532
rect 39440 1492 39442 1532
rect 39150 1450 39274 1492
rect 39318 1450 39442 1492
rect 51150 1532 51274 1574
rect 51318 1532 51442 1574
rect 51150 1492 51152 1532
rect 51152 1492 51194 1532
rect 51194 1492 51234 1532
rect 51234 1492 51274 1532
rect 51318 1492 51358 1532
rect 51358 1492 51398 1532
rect 51398 1492 51440 1532
rect 51440 1492 51442 1532
rect 51150 1450 51274 1492
rect 51318 1450 51442 1492
rect 63150 1532 63274 1574
rect 63318 1532 63442 1574
rect 63150 1492 63152 1532
rect 63152 1492 63194 1532
rect 63194 1492 63234 1532
rect 63234 1492 63274 1532
rect 63318 1492 63358 1532
rect 63358 1492 63398 1532
rect 63398 1492 63440 1532
rect 63440 1492 63442 1532
rect 63150 1450 63274 1492
rect 63318 1450 63442 1492
rect 75150 1532 75274 1574
rect 75318 1532 75442 1574
rect 75150 1492 75152 1532
rect 75152 1492 75194 1532
rect 75194 1492 75234 1532
rect 75234 1492 75274 1532
rect 75318 1492 75358 1532
rect 75358 1492 75398 1532
rect 75398 1492 75440 1532
rect 75440 1492 75442 1532
rect 75150 1450 75274 1492
rect 75318 1450 75442 1492
rect 4390 776 4514 818
rect 4558 776 4682 818
rect 4390 736 4392 776
rect 4392 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4514 776
rect 4558 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4680 776
rect 4680 736 4682 776
rect 4390 694 4514 736
rect 4558 694 4682 736
rect 16390 776 16514 818
rect 16558 776 16682 818
rect 16390 736 16392 776
rect 16392 736 16434 776
rect 16434 736 16474 776
rect 16474 736 16514 776
rect 16558 736 16598 776
rect 16598 736 16638 776
rect 16638 736 16680 776
rect 16680 736 16682 776
rect 16390 694 16514 736
rect 16558 694 16682 736
rect 28390 776 28514 818
rect 28558 776 28682 818
rect 28390 736 28392 776
rect 28392 736 28434 776
rect 28434 736 28474 776
rect 28474 736 28514 776
rect 28558 736 28598 776
rect 28598 736 28638 776
rect 28638 736 28680 776
rect 28680 736 28682 776
rect 28390 694 28514 736
rect 28558 694 28682 736
rect 40390 776 40514 818
rect 40558 776 40682 818
rect 40390 736 40392 776
rect 40392 736 40434 776
rect 40434 736 40474 776
rect 40474 736 40514 776
rect 40558 736 40598 776
rect 40598 736 40638 776
rect 40638 736 40680 776
rect 40680 736 40682 776
rect 40390 694 40514 736
rect 40558 694 40682 736
rect 52390 776 52514 818
rect 52558 776 52682 818
rect 52390 736 52392 776
rect 52392 736 52434 776
rect 52434 736 52474 776
rect 52474 736 52514 776
rect 52558 736 52598 776
rect 52598 736 52638 776
rect 52638 736 52680 776
rect 52680 736 52682 776
rect 52390 694 52514 736
rect 52558 694 52682 736
rect 64390 776 64514 818
rect 64558 776 64682 818
rect 64390 736 64392 776
rect 64392 736 64434 776
rect 64434 736 64474 776
rect 64474 736 64514 776
rect 64558 736 64598 776
rect 64598 736 64638 776
rect 64638 736 64680 776
rect 64680 736 64682 776
rect 64390 694 64514 736
rect 64558 694 64682 736
rect 76390 776 76514 818
rect 76558 776 76682 818
rect 76390 736 76392 776
rect 76392 736 76434 776
rect 76434 736 76474 776
rect 76474 736 76514 776
rect 76558 736 76598 776
rect 76598 736 76638 776
rect 76638 736 76680 776
rect 76680 736 76682 776
rect 76390 694 76514 736
rect 76558 694 76682 736
<< metal6 >>
rect 4316 38618 4756 38682
rect 3076 37862 3516 38600
rect 3076 37738 3150 37862
rect 3274 37738 3318 37862
rect 3442 37738 3516 37862
rect 3076 36350 3516 37738
rect 3076 36226 3150 36350
rect 3274 36226 3318 36350
rect 3442 36226 3516 36350
rect 3076 34838 3516 36226
rect 3076 34714 3150 34838
rect 3274 34714 3318 34838
rect 3442 34714 3516 34838
rect 3076 33326 3516 34714
rect 3076 33202 3150 33326
rect 3274 33202 3318 33326
rect 3442 33202 3516 33326
rect 3076 31814 3516 33202
rect 3076 31690 3150 31814
rect 3274 31690 3318 31814
rect 3442 31690 3516 31814
rect 3076 30302 3516 31690
rect 3076 30178 3150 30302
rect 3274 30178 3318 30302
rect 3442 30178 3516 30302
rect 3076 28790 3516 30178
rect 3076 28666 3150 28790
rect 3274 28666 3318 28790
rect 3442 28666 3516 28790
rect 3076 27278 3516 28666
rect 3076 27154 3150 27278
rect 3274 27154 3318 27278
rect 3442 27154 3516 27278
rect 3076 25766 3516 27154
rect 3076 25642 3150 25766
rect 3274 25642 3318 25766
rect 3442 25642 3516 25766
rect 3076 24254 3516 25642
rect 3076 24130 3150 24254
rect 3274 24130 3318 24254
rect 3442 24130 3516 24254
rect 3076 22742 3516 24130
rect 3076 22618 3150 22742
rect 3274 22618 3318 22742
rect 3442 22618 3516 22742
rect 3076 21230 3516 22618
rect 3076 21106 3150 21230
rect 3274 21106 3318 21230
rect 3442 21106 3516 21230
rect 3076 19718 3516 21106
rect 3076 19594 3150 19718
rect 3274 19594 3318 19718
rect 3442 19594 3516 19718
rect 3076 18206 3516 19594
rect 3076 18082 3150 18206
rect 3274 18082 3318 18206
rect 3442 18082 3516 18206
rect 3076 16694 3516 18082
rect 3076 16570 3150 16694
rect 3274 16570 3318 16694
rect 3442 16570 3516 16694
rect 3076 15182 3516 16570
rect 3076 15058 3150 15182
rect 3274 15058 3318 15182
rect 3442 15058 3516 15182
rect 3076 13670 3516 15058
rect 3076 13546 3150 13670
rect 3274 13546 3318 13670
rect 3442 13546 3516 13670
rect 3076 12158 3516 13546
rect 3076 12034 3150 12158
rect 3274 12034 3318 12158
rect 3442 12034 3516 12158
rect 3076 10646 3516 12034
rect 3076 10522 3150 10646
rect 3274 10522 3318 10646
rect 3442 10522 3516 10646
rect 3076 9134 3516 10522
rect 3076 9010 3150 9134
rect 3274 9010 3318 9134
rect 3442 9010 3516 9134
rect 3076 7622 3516 9010
rect 3076 7498 3150 7622
rect 3274 7498 3318 7622
rect 3442 7498 3516 7622
rect 3076 6110 3516 7498
rect 3076 5986 3150 6110
rect 3274 5986 3318 6110
rect 3442 5986 3516 6110
rect 3076 4598 3516 5986
rect 3076 4474 3150 4598
rect 3274 4474 3318 4598
rect 3442 4474 3516 4598
rect 3076 3086 3516 4474
rect 3076 2962 3150 3086
rect 3274 2962 3318 3086
rect 3442 2962 3516 3086
rect 3076 1574 3516 2962
rect 3076 1450 3150 1574
rect 3274 1450 3318 1574
rect 3442 1450 3516 1574
rect 3076 712 3516 1450
rect 4316 38494 4390 38618
rect 4514 38494 4558 38618
rect 4682 38494 4756 38618
rect 16316 38618 16756 38682
rect 4316 37106 4756 38494
rect 4316 36982 4390 37106
rect 4514 36982 4558 37106
rect 4682 36982 4756 37106
rect 4316 35594 4756 36982
rect 4316 35470 4390 35594
rect 4514 35470 4558 35594
rect 4682 35470 4756 35594
rect 4316 34082 4756 35470
rect 4316 33958 4390 34082
rect 4514 33958 4558 34082
rect 4682 33958 4756 34082
rect 4316 32570 4756 33958
rect 4316 32446 4390 32570
rect 4514 32446 4558 32570
rect 4682 32446 4756 32570
rect 4316 31058 4756 32446
rect 4316 30934 4390 31058
rect 4514 30934 4558 31058
rect 4682 30934 4756 31058
rect 4316 29546 4756 30934
rect 4316 29422 4390 29546
rect 4514 29422 4558 29546
rect 4682 29422 4756 29546
rect 4316 28034 4756 29422
rect 4316 27910 4390 28034
rect 4514 27910 4558 28034
rect 4682 27910 4756 28034
rect 4316 26522 4756 27910
rect 4316 26398 4390 26522
rect 4514 26398 4558 26522
rect 4682 26398 4756 26522
rect 4316 25010 4756 26398
rect 4316 24886 4390 25010
rect 4514 24886 4558 25010
rect 4682 24886 4756 25010
rect 4316 23498 4756 24886
rect 4316 23374 4390 23498
rect 4514 23374 4558 23498
rect 4682 23374 4756 23498
rect 4316 21986 4756 23374
rect 4316 21862 4390 21986
rect 4514 21862 4558 21986
rect 4682 21862 4756 21986
rect 4316 20474 4756 21862
rect 4316 20350 4390 20474
rect 4514 20350 4558 20474
rect 4682 20350 4756 20474
rect 4316 18962 4756 20350
rect 4316 18838 4390 18962
rect 4514 18838 4558 18962
rect 4682 18838 4756 18962
rect 4316 17450 4756 18838
rect 4316 17326 4390 17450
rect 4514 17326 4558 17450
rect 4682 17326 4756 17450
rect 4316 15938 4756 17326
rect 4316 15814 4390 15938
rect 4514 15814 4558 15938
rect 4682 15814 4756 15938
rect 4316 14426 4756 15814
rect 4316 14302 4390 14426
rect 4514 14302 4558 14426
rect 4682 14302 4756 14426
rect 4316 12914 4756 14302
rect 4316 12790 4390 12914
rect 4514 12790 4558 12914
rect 4682 12790 4756 12914
rect 4316 11402 4756 12790
rect 4316 11278 4390 11402
rect 4514 11278 4558 11402
rect 4682 11278 4756 11402
rect 4316 9890 4756 11278
rect 4316 9766 4390 9890
rect 4514 9766 4558 9890
rect 4682 9766 4756 9890
rect 4316 8378 4756 9766
rect 4316 8254 4390 8378
rect 4514 8254 4558 8378
rect 4682 8254 4756 8378
rect 4316 6866 4756 8254
rect 4316 6742 4390 6866
rect 4514 6742 4558 6866
rect 4682 6742 4756 6866
rect 4316 5354 4756 6742
rect 4316 5230 4390 5354
rect 4514 5230 4558 5354
rect 4682 5230 4756 5354
rect 4316 3842 4756 5230
rect 4316 3718 4390 3842
rect 4514 3718 4558 3842
rect 4682 3718 4756 3842
rect 4316 2330 4756 3718
rect 4316 2206 4390 2330
rect 4514 2206 4558 2330
rect 4682 2206 4756 2330
rect 4316 818 4756 2206
rect 4316 694 4390 818
rect 4514 694 4558 818
rect 4682 694 4756 818
rect 15076 37862 15516 38600
rect 15076 37738 15150 37862
rect 15274 37738 15318 37862
rect 15442 37738 15516 37862
rect 15076 36350 15516 37738
rect 15076 36226 15150 36350
rect 15274 36226 15318 36350
rect 15442 36226 15516 36350
rect 15076 34838 15516 36226
rect 15076 34714 15150 34838
rect 15274 34714 15318 34838
rect 15442 34714 15516 34838
rect 15076 33326 15516 34714
rect 15076 33202 15150 33326
rect 15274 33202 15318 33326
rect 15442 33202 15516 33326
rect 15076 31814 15516 33202
rect 15076 31690 15150 31814
rect 15274 31690 15318 31814
rect 15442 31690 15516 31814
rect 15076 30302 15516 31690
rect 15076 30178 15150 30302
rect 15274 30178 15318 30302
rect 15442 30178 15516 30302
rect 15076 28790 15516 30178
rect 15076 28666 15150 28790
rect 15274 28666 15318 28790
rect 15442 28666 15516 28790
rect 15076 27278 15516 28666
rect 15076 27154 15150 27278
rect 15274 27154 15318 27278
rect 15442 27154 15516 27278
rect 15076 25766 15516 27154
rect 15076 25642 15150 25766
rect 15274 25642 15318 25766
rect 15442 25642 15516 25766
rect 15076 24254 15516 25642
rect 15076 24130 15150 24254
rect 15274 24130 15318 24254
rect 15442 24130 15516 24254
rect 15076 22742 15516 24130
rect 15076 22618 15150 22742
rect 15274 22618 15318 22742
rect 15442 22618 15516 22742
rect 15076 21230 15516 22618
rect 15076 21106 15150 21230
rect 15274 21106 15318 21230
rect 15442 21106 15516 21230
rect 15076 19718 15516 21106
rect 15076 19594 15150 19718
rect 15274 19594 15318 19718
rect 15442 19594 15516 19718
rect 15076 18206 15516 19594
rect 15076 18082 15150 18206
rect 15274 18082 15318 18206
rect 15442 18082 15516 18206
rect 15076 16694 15516 18082
rect 15076 16570 15150 16694
rect 15274 16570 15318 16694
rect 15442 16570 15516 16694
rect 15076 15182 15516 16570
rect 15076 15058 15150 15182
rect 15274 15058 15318 15182
rect 15442 15058 15516 15182
rect 15076 13670 15516 15058
rect 15076 13546 15150 13670
rect 15274 13546 15318 13670
rect 15442 13546 15516 13670
rect 15076 12158 15516 13546
rect 15076 12034 15150 12158
rect 15274 12034 15318 12158
rect 15442 12034 15516 12158
rect 15076 10646 15516 12034
rect 15076 10522 15150 10646
rect 15274 10522 15318 10646
rect 15442 10522 15516 10646
rect 15076 9134 15516 10522
rect 15076 9010 15150 9134
rect 15274 9010 15318 9134
rect 15442 9010 15516 9134
rect 15076 7622 15516 9010
rect 15076 7498 15150 7622
rect 15274 7498 15318 7622
rect 15442 7498 15516 7622
rect 15076 6110 15516 7498
rect 15076 5986 15150 6110
rect 15274 5986 15318 6110
rect 15442 5986 15516 6110
rect 15076 4598 15516 5986
rect 15076 4474 15150 4598
rect 15274 4474 15318 4598
rect 15442 4474 15516 4598
rect 15076 3086 15516 4474
rect 15076 2962 15150 3086
rect 15274 2962 15318 3086
rect 15442 2962 15516 3086
rect 15076 1574 15516 2962
rect 15076 1450 15150 1574
rect 15274 1450 15318 1574
rect 15442 1450 15516 1574
rect 15076 712 15516 1450
rect 16316 38494 16390 38618
rect 16514 38494 16558 38618
rect 16682 38494 16756 38618
rect 28316 38618 28756 38682
rect 16316 37106 16756 38494
rect 16316 36982 16390 37106
rect 16514 36982 16558 37106
rect 16682 36982 16756 37106
rect 16316 35594 16756 36982
rect 16316 35470 16390 35594
rect 16514 35470 16558 35594
rect 16682 35470 16756 35594
rect 16316 34082 16756 35470
rect 16316 33958 16390 34082
rect 16514 33958 16558 34082
rect 16682 33958 16756 34082
rect 16316 32570 16756 33958
rect 16316 32446 16390 32570
rect 16514 32446 16558 32570
rect 16682 32446 16756 32570
rect 16316 31058 16756 32446
rect 16316 30934 16390 31058
rect 16514 30934 16558 31058
rect 16682 30934 16756 31058
rect 16316 29546 16756 30934
rect 16316 29422 16390 29546
rect 16514 29422 16558 29546
rect 16682 29422 16756 29546
rect 16316 28034 16756 29422
rect 16316 27910 16390 28034
rect 16514 27910 16558 28034
rect 16682 27910 16756 28034
rect 16316 26522 16756 27910
rect 16316 26398 16390 26522
rect 16514 26398 16558 26522
rect 16682 26398 16756 26522
rect 16316 25010 16756 26398
rect 16316 24886 16390 25010
rect 16514 24886 16558 25010
rect 16682 24886 16756 25010
rect 16316 23498 16756 24886
rect 16316 23374 16390 23498
rect 16514 23374 16558 23498
rect 16682 23374 16756 23498
rect 16316 21986 16756 23374
rect 16316 21862 16390 21986
rect 16514 21862 16558 21986
rect 16682 21862 16756 21986
rect 16316 20474 16756 21862
rect 16316 20350 16390 20474
rect 16514 20350 16558 20474
rect 16682 20350 16756 20474
rect 16316 18962 16756 20350
rect 16316 18838 16390 18962
rect 16514 18838 16558 18962
rect 16682 18838 16756 18962
rect 16316 17450 16756 18838
rect 16316 17326 16390 17450
rect 16514 17326 16558 17450
rect 16682 17326 16756 17450
rect 16316 15938 16756 17326
rect 16316 15814 16390 15938
rect 16514 15814 16558 15938
rect 16682 15814 16756 15938
rect 16316 14426 16756 15814
rect 16316 14302 16390 14426
rect 16514 14302 16558 14426
rect 16682 14302 16756 14426
rect 16316 12914 16756 14302
rect 16316 12790 16390 12914
rect 16514 12790 16558 12914
rect 16682 12790 16756 12914
rect 16316 11402 16756 12790
rect 16316 11278 16390 11402
rect 16514 11278 16558 11402
rect 16682 11278 16756 11402
rect 16316 9890 16756 11278
rect 16316 9766 16390 9890
rect 16514 9766 16558 9890
rect 16682 9766 16756 9890
rect 16316 8378 16756 9766
rect 16316 8254 16390 8378
rect 16514 8254 16558 8378
rect 16682 8254 16756 8378
rect 16316 6866 16756 8254
rect 16316 6742 16390 6866
rect 16514 6742 16558 6866
rect 16682 6742 16756 6866
rect 16316 5354 16756 6742
rect 16316 5230 16390 5354
rect 16514 5230 16558 5354
rect 16682 5230 16756 5354
rect 16316 3842 16756 5230
rect 16316 3718 16390 3842
rect 16514 3718 16558 3842
rect 16682 3718 16756 3842
rect 16316 2330 16756 3718
rect 16316 2206 16390 2330
rect 16514 2206 16558 2330
rect 16682 2206 16756 2330
rect 16316 818 16756 2206
rect 4316 630 4756 694
rect 16316 694 16390 818
rect 16514 694 16558 818
rect 16682 694 16756 818
rect 27076 37862 27516 38600
rect 27076 37738 27150 37862
rect 27274 37738 27318 37862
rect 27442 37738 27516 37862
rect 27076 36350 27516 37738
rect 27076 36226 27150 36350
rect 27274 36226 27318 36350
rect 27442 36226 27516 36350
rect 27076 34838 27516 36226
rect 27076 34714 27150 34838
rect 27274 34714 27318 34838
rect 27442 34714 27516 34838
rect 27076 33326 27516 34714
rect 27076 33202 27150 33326
rect 27274 33202 27318 33326
rect 27442 33202 27516 33326
rect 27076 31814 27516 33202
rect 27076 31690 27150 31814
rect 27274 31690 27318 31814
rect 27442 31690 27516 31814
rect 27076 30302 27516 31690
rect 27076 30178 27150 30302
rect 27274 30178 27318 30302
rect 27442 30178 27516 30302
rect 27076 28790 27516 30178
rect 27076 28666 27150 28790
rect 27274 28666 27318 28790
rect 27442 28666 27516 28790
rect 27076 27278 27516 28666
rect 27076 27154 27150 27278
rect 27274 27154 27318 27278
rect 27442 27154 27516 27278
rect 27076 25766 27516 27154
rect 27076 25642 27150 25766
rect 27274 25642 27318 25766
rect 27442 25642 27516 25766
rect 27076 24254 27516 25642
rect 27076 24130 27150 24254
rect 27274 24130 27318 24254
rect 27442 24130 27516 24254
rect 27076 22742 27516 24130
rect 27076 22618 27150 22742
rect 27274 22618 27318 22742
rect 27442 22618 27516 22742
rect 27076 21230 27516 22618
rect 27076 21106 27150 21230
rect 27274 21106 27318 21230
rect 27442 21106 27516 21230
rect 27076 19718 27516 21106
rect 27076 19594 27150 19718
rect 27274 19594 27318 19718
rect 27442 19594 27516 19718
rect 27076 18206 27516 19594
rect 27076 18082 27150 18206
rect 27274 18082 27318 18206
rect 27442 18082 27516 18206
rect 27076 16694 27516 18082
rect 27076 16570 27150 16694
rect 27274 16570 27318 16694
rect 27442 16570 27516 16694
rect 27076 15182 27516 16570
rect 27076 15058 27150 15182
rect 27274 15058 27318 15182
rect 27442 15058 27516 15182
rect 27076 13670 27516 15058
rect 27076 13546 27150 13670
rect 27274 13546 27318 13670
rect 27442 13546 27516 13670
rect 27076 12158 27516 13546
rect 27076 12034 27150 12158
rect 27274 12034 27318 12158
rect 27442 12034 27516 12158
rect 27076 10646 27516 12034
rect 27076 10522 27150 10646
rect 27274 10522 27318 10646
rect 27442 10522 27516 10646
rect 27076 9134 27516 10522
rect 27076 9010 27150 9134
rect 27274 9010 27318 9134
rect 27442 9010 27516 9134
rect 27076 7622 27516 9010
rect 27076 7498 27150 7622
rect 27274 7498 27318 7622
rect 27442 7498 27516 7622
rect 27076 6110 27516 7498
rect 27076 5986 27150 6110
rect 27274 5986 27318 6110
rect 27442 5986 27516 6110
rect 27076 4598 27516 5986
rect 27076 4474 27150 4598
rect 27274 4474 27318 4598
rect 27442 4474 27516 4598
rect 27076 3086 27516 4474
rect 27076 2962 27150 3086
rect 27274 2962 27318 3086
rect 27442 2962 27516 3086
rect 27076 1574 27516 2962
rect 27076 1450 27150 1574
rect 27274 1450 27318 1574
rect 27442 1450 27516 1574
rect 27076 712 27516 1450
rect 28316 38494 28390 38618
rect 28514 38494 28558 38618
rect 28682 38494 28756 38618
rect 40316 38618 40756 38682
rect 28316 37106 28756 38494
rect 28316 36982 28390 37106
rect 28514 36982 28558 37106
rect 28682 36982 28756 37106
rect 28316 35594 28756 36982
rect 28316 35470 28390 35594
rect 28514 35470 28558 35594
rect 28682 35470 28756 35594
rect 28316 34082 28756 35470
rect 28316 33958 28390 34082
rect 28514 33958 28558 34082
rect 28682 33958 28756 34082
rect 28316 32570 28756 33958
rect 28316 32446 28390 32570
rect 28514 32446 28558 32570
rect 28682 32446 28756 32570
rect 28316 31058 28756 32446
rect 28316 30934 28390 31058
rect 28514 30934 28558 31058
rect 28682 30934 28756 31058
rect 28316 29546 28756 30934
rect 28316 29422 28390 29546
rect 28514 29422 28558 29546
rect 28682 29422 28756 29546
rect 28316 28034 28756 29422
rect 28316 27910 28390 28034
rect 28514 27910 28558 28034
rect 28682 27910 28756 28034
rect 28316 26522 28756 27910
rect 28316 26398 28390 26522
rect 28514 26398 28558 26522
rect 28682 26398 28756 26522
rect 28316 25010 28756 26398
rect 28316 24886 28390 25010
rect 28514 24886 28558 25010
rect 28682 24886 28756 25010
rect 28316 23498 28756 24886
rect 28316 23374 28390 23498
rect 28514 23374 28558 23498
rect 28682 23374 28756 23498
rect 28316 21986 28756 23374
rect 28316 21862 28390 21986
rect 28514 21862 28558 21986
rect 28682 21862 28756 21986
rect 28316 20474 28756 21862
rect 28316 20350 28390 20474
rect 28514 20350 28558 20474
rect 28682 20350 28756 20474
rect 28316 18962 28756 20350
rect 28316 18838 28390 18962
rect 28514 18838 28558 18962
rect 28682 18838 28756 18962
rect 28316 17450 28756 18838
rect 28316 17326 28390 17450
rect 28514 17326 28558 17450
rect 28682 17326 28756 17450
rect 28316 15938 28756 17326
rect 28316 15814 28390 15938
rect 28514 15814 28558 15938
rect 28682 15814 28756 15938
rect 28316 14426 28756 15814
rect 28316 14302 28390 14426
rect 28514 14302 28558 14426
rect 28682 14302 28756 14426
rect 28316 12914 28756 14302
rect 28316 12790 28390 12914
rect 28514 12790 28558 12914
rect 28682 12790 28756 12914
rect 28316 11402 28756 12790
rect 28316 11278 28390 11402
rect 28514 11278 28558 11402
rect 28682 11278 28756 11402
rect 28316 9890 28756 11278
rect 28316 9766 28390 9890
rect 28514 9766 28558 9890
rect 28682 9766 28756 9890
rect 28316 8378 28756 9766
rect 28316 8254 28390 8378
rect 28514 8254 28558 8378
rect 28682 8254 28756 8378
rect 28316 6866 28756 8254
rect 28316 6742 28390 6866
rect 28514 6742 28558 6866
rect 28682 6742 28756 6866
rect 28316 5354 28756 6742
rect 28316 5230 28390 5354
rect 28514 5230 28558 5354
rect 28682 5230 28756 5354
rect 28316 3842 28756 5230
rect 28316 3718 28390 3842
rect 28514 3718 28558 3842
rect 28682 3718 28756 3842
rect 28316 2330 28756 3718
rect 28316 2206 28390 2330
rect 28514 2206 28558 2330
rect 28682 2206 28756 2330
rect 28316 818 28756 2206
rect 16316 630 16756 694
rect 28316 694 28390 818
rect 28514 694 28558 818
rect 28682 694 28756 818
rect 39076 37862 39516 38600
rect 39076 37738 39150 37862
rect 39274 37738 39318 37862
rect 39442 37738 39516 37862
rect 39076 36350 39516 37738
rect 39076 36226 39150 36350
rect 39274 36226 39318 36350
rect 39442 36226 39516 36350
rect 39076 34838 39516 36226
rect 39076 34714 39150 34838
rect 39274 34714 39318 34838
rect 39442 34714 39516 34838
rect 39076 33326 39516 34714
rect 39076 33202 39150 33326
rect 39274 33202 39318 33326
rect 39442 33202 39516 33326
rect 39076 31814 39516 33202
rect 39076 31690 39150 31814
rect 39274 31690 39318 31814
rect 39442 31690 39516 31814
rect 39076 30302 39516 31690
rect 39076 30178 39150 30302
rect 39274 30178 39318 30302
rect 39442 30178 39516 30302
rect 39076 28790 39516 30178
rect 39076 28666 39150 28790
rect 39274 28666 39318 28790
rect 39442 28666 39516 28790
rect 39076 27278 39516 28666
rect 39076 27154 39150 27278
rect 39274 27154 39318 27278
rect 39442 27154 39516 27278
rect 39076 25766 39516 27154
rect 39076 25642 39150 25766
rect 39274 25642 39318 25766
rect 39442 25642 39516 25766
rect 39076 24254 39516 25642
rect 39076 24130 39150 24254
rect 39274 24130 39318 24254
rect 39442 24130 39516 24254
rect 39076 22742 39516 24130
rect 39076 22618 39150 22742
rect 39274 22618 39318 22742
rect 39442 22618 39516 22742
rect 39076 21230 39516 22618
rect 39076 21106 39150 21230
rect 39274 21106 39318 21230
rect 39442 21106 39516 21230
rect 39076 19718 39516 21106
rect 39076 19594 39150 19718
rect 39274 19594 39318 19718
rect 39442 19594 39516 19718
rect 39076 18206 39516 19594
rect 39076 18082 39150 18206
rect 39274 18082 39318 18206
rect 39442 18082 39516 18206
rect 39076 16694 39516 18082
rect 39076 16570 39150 16694
rect 39274 16570 39318 16694
rect 39442 16570 39516 16694
rect 39076 15182 39516 16570
rect 39076 15058 39150 15182
rect 39274 15058 39318 15182
rect 39442 15058 39516 15182
rect 39076 13670 39516 15058
rect 39076 13546 39150 13670
rect 39274 13546 39318 13670
rect 39442 13546 39516 13670
rect 39076 12158 39516 13546
rect 39076 12034 39150 12158
rect 39274 12034 39318 12158
rect 39442 12034 39516 12158
rect 39076 10646 39516 12034
rect 39076 10522 39150 10646
rect 39274 10522 39318 10646
rect 39442 10522 39516 10646
rect 39076 9134 39516 10522
rect 39076 9010 39150 9134
rect 39274 9010 39318 9134
rect 39442 9010 39516 9134
rect 39076 7622 39516 9010
rect 39076 7498 39150 7622
rect 39274 7498 39318 7622
rect 39442 7498 39516 7622
rect 39076 6110 39516 7498
rect 39076 5986 39150 6110
rect 39274 5986 39318 6110
rect 39442 5986 39516 6110
rect 39076 4598 39516 5986
rect 39076 4474 39150 4598
rect 39274 4474 39318 4598
rect 39442 4474 39516 4598
rect 39076 3086 39516 4474
rect 39076 2962 39150 3086
rect 39274 2962 39318 3086
rect 39442 2962 39516 3086
rect 39076 1574 39516 2962
rect 39076 1450 39150 1574
rect 39274 1450 39318 1574
rect 39442 1450 39516 1574
rect 39076 712 39516 1450
rect 40316 38494 40390 38618
rect 40514 38494 40558 38618
rect 40682 38494 40756 38618
rect 52316 38618 52756 38682
rect 40316 37106 40756 38494
rect 40316 36982 40390 37106
rect 40514 36982 40558 37106
rect 40682 36982 40756 37106
rect 40316 35594 40756 36982
rect 40316 35470 40390 35594
rect 40514 35470 40558 35594
rect 40682 35470 40756 35594
rect 40316 34082 40756 35470
rect 40316 33958 40390 34082
rect 40514 33958 40558 34082
rect 40682 33958 40756 34082
rect 40316 32570 40756 33958
rect 40316 32446 40390 32570
rect 40514 32446 40558 32570
rect 40682 32446 40756 32570
rect 40316 31058 40756 32446
rect 40316 30934 40390 31058
rect 40514 30934 40558 31058
rect 40682 30934 40756 31058
rect 40316 29546 40756 30934
rect 40316 29422 40390 29546
rect 40514 29422 40558 29546
rect 40682 29422 40756 29546
rect 40316 28034 40756 29422
rect 40316 27910 40390 28034
rect 40514 27910 40558 28034
rect 40682 27910 40756 28034
rect 40316 26522 40756 27910
rect 40316 26398 40390 26522
rect 40514 26398 40558 26522
rect 40682 26398 40756 26522
rect 40316 25010 40756 26398
rect 40316 24886 40390 25010
rect 40514 24886 40558 25010
rect 40682 24886 40756 25010
rect 40316 23498 40756 24886
rect 40316 23374 40390 23498
rect 40514 23374 40558 23498
rect 40682 23374 40756 23498
rect 40316 21986 40756 23374
rect 40316 21862 40390 21986
rect 40514 21862 40558 21986
rect 40682 21862 40756 21986
rect 40316 20474 40756 21862
rect 40316 20350 40390 20474
rect 40514 20350 40558 20474
rect 40682 20350 40756 20474
rect 40316 18962 40756 20350
rect 40316 18838 40390 18962
rect 40514 18838 40558 18962
rect 40682 18838 40756 18962
rect 40316 17450 40756 18838
rect 40316 17326 40390 17450
rect 40514 17326 40558 17450
rect 40682 17326 40756 17450
rect 40316 15938 40756 17326
rect 40316 15814 40390 15938
rect 40514 15814 40558 15938
rect 40682 15814 40756 15938
rect 40316 14426 40756 15814
rect 40316 14302 40390 14426
rect 40514 14302 40558 14426
rect 40682 14302 40756 14426
rect 40316 12914 40756 14302
rect 40316 12790 40390 12914
rect 40514 12790 40558 12914
rect 40682 12790 40756 12914
rect 40316 11402 40756 12790
rect 40316 11278 40390 11402
rect 40514 11278 40558 11402
rect 40682 11278 40756 11402
rect 40316 9890 40756 11278
rect 40316 9766 40390 9890
rect 40514 9766 40558 9890
rect 40682 9766 40756 9890
rect 40316 8378 40756 9766
rect 40316 8254 40390 8378
rect 40514 8254 40558 8378
rect 40682 8254 40756 8378
rect 40316 6866 40756 8254
rect 40316 6742 40390 6866
rect 40514 6742 40558 6866
rect 40682 6742 40756 6866
rect 40316 5354 40756 6742
rect 40316 5230 40390 5354
rect 40514 5230 40558 5354
rect 40682 5230 40756 5354
rect 40316 3842 40756 5230
rect 40316 3718 40390 3842
rect 40514 3718 40558 3842
rect 40682 3718 40756 3842
rect 40316 2330 40756 3718
rect 40316 2206 40390 2330
rect 40514 2206 40558 2330
rect 40682 2206 40756 2330
rect 40316 818 40756 2206
rect 28316 630 28756 694
rect 40316 694 40390 818
rect 40514 694 40558 818
rect 40682 694 40756 818
rect 51076 37862 51516 38600
rect 51076 37738 51150 37862
rect 51274 37738 51318 37862
rect 51442 37738 51516 37862
rect 51076 36350 51516 37738
rect 51076 36226 51150 36350
rect 51274 36226 51318 36350
rect 51442 36226 51516 36350
rect 51076 34838 51516 36226
rect 51076 34714 51150 34838
rect 51274 34714 51318 34838
rect 51442 34714 51516 34838
rect 51076 33326 51516 34714
rect 51076 33202 51150 33326
rect 51274 33202 51318 33326
rect 51442 33202 51516 33326
rect 51076 31814 51516 33202
rect 51076 31690 51150 31814
rect 51274 31690 51318 31814
rect 51442 31690 51516 31814
rect 51076 30302 51516 31690
rect 51076 30178 51150 30302
rect 51274 30178 51318 30302
rect 51442 30178 51516 30302
rect 51076 28790 51516 30178
rect 51076 28666 51150 28790
rect 51274 28666 51318 28790
rect 51442 28666 51516 28790
rect 51076 27278 51516 28666
rect 51076 27154 51150 27278
rect 51274 27154 51318 27278
rect 51442 27154 51516 27278
rect 51076 25766 51516 27154
rect 51076 25642 51150 25766
rect 51274 25642 51318 25766
rect 51442 25642 51516 25766
rect 51076 15182 51516 25642
rect 51076 15058 51150 15182
rect 51274 15058 51318 15182
rect 51442 15058 51516 15182
rect 51076 13670 51516 15058
rect 51076 13546 51150 13670
rect 51274 13546 51318 13670
rect 51442 13546 51516 13670
rect 51076 12158 51516 13546
rect 51076 12034 51150 12158
rect 51274 12034 51318 12158
rect 51442 12034 51516 12158
rect 51076 10646 51516 12034
rect 51076 10522 51150 10646
rect 51274 10522 51318 10646
rect 51442 10522 51516 10646
rect 51076 9134 51516 10522
rect 51076 9010 51150 9134
rect 51274 9010 51318 9134
rect 51442 9010 51516 9134
rect 51076 7622 51516 9010
rect 51076 7498 51150 7622
rect 51274 7498 51318 7622
rect 51442 7498 51516 7622
rect 51076 6110 51516 7498
rect 51076 5986 51150 6110
rect 51274 5986 51318 6110
rect 51442 5986 51516 6110
rect 51076 4598 51516 5986
rect 51076 4474 51150 4598
rect 51274 4474 51318 4598
rect 51442 4474 51516 4598
rect 51076 3086 51516 4474
rect 51076 2962 51150 3086
rect 51274 2962 51318 3086
rect 51442 2962 51516 3086
rect 51076 1574 51516 2962
rect 51076 1450 51150 1574
rect 51274 1450 51318 1574
rect 51442 1450 51516 1574
rect 51076 712 51516 1450
rect 52316 38494 52390 38618
rect 52514 38494 52558 38618
rect 52682 38494 52756 38618
rect 64316 38618 64756 38682
rect 52316 37106 52756 38494
rect 52316 36982 52390 37106
rect 52514 36982 52558 37106
rect 52682 36982 52756 37106
rect 52316 35594 52756 36982
rect 52316 35470 52390 35594
rect 52514 35470 52558 35594
rect 52682 35470 52756 35594
rect 52316 34082 52756 35470
rect 52316 33958 52390 34082
rect 52514 33958 52558 34082
rect 52682 33958 52756 34082
rect 52316 32570 52756 33958
rect 52316 32446 52390 32570
rect 52514 32446 52558 32570
rect 52682 32446 52756 32570
rect 52316 31058 52756 32446
rect 52316 30934 52390 31058
rect 52514 30934 52558 31058
rect 52682 30934 52756 31058
rect 52316 29546 52756 30934
rect 52316 29422 52390 29546
rect 52514 29422 52558 29546
rect 52682 29422 52756 29546
rect 52316 28034 52756 29422
rect 52316 27910 52390 28034
rect 52514 27910 52558 28034
rect 52682 27910 52756 28034
rect 52316 26522 52756 27910
rect 52316 26398 52390 26522
rect 52514 26398 52558 26522
rect 52682 26398 52756 26522
rect 52316 25010 52756 26398
rect 52316 24886 52390 25010
rect 52514 24886 52558 25010
rect 52682 24886 52756 25010
rect 52316 14426 52756 24886
rect 52316 14302 52390 14426
rect 52514 14302 52558 14426
rect 52682 14302 52756 14426
rect 52316 12914 52756 14302
rect 52316 12790 52390 12914
rect 52514 12790 52558 12914
rect 52682 12790 52756 12914
rect 52316 11402 52756 12790
rect 52316 11278 52390 11402
rect 52514 11278 52558 11402
rect 52682 11278 52756 11402
rect 52316 9890 52756 11278
rect 52316 9766 52390 9890
rect 52514 9766 52558 9890
rect 52682 9766 52756 9890
rect 52316 8378 52756 9766
rect 52316 8254 52390 8378
rect 52514 8254 52558 8378
rect 52682 8254 52756 8378
rect 52316 6866 52756 8254
rect 52316 6742 52390 6866
rect 52514 6742 52558 6866
rect 52682 6742 52756 6866
rect 52316 5354 52756 6742
rect 52316 5230 52390 5354
rect 52514 5230 52558 5354
rect 52682 5230 52756 5354
rect 52316 3842 52756 5230
rect 52316 3718 52390 3842
rect 52514 3718 52558 3842
rect 52682 3718 52756 3842
rect 52316 2330 52756 3718
rect 52316 2206 52390 2330
rect 52514 2206 52558 2330
rect 52682 2206 52756 2330
rect 52316 818 52756 2206
rect 40316 630 40756 694
rect 52316 694 52390 818
rect 52514 694 52558 818
rect 52682 694 52756 818
rect 63076 37862 63516 38600
rect 63076 37738 63150 37862
rect 63274 37738 63318 37862
rect 63442 37738 63516 37862
rect 63076 36350 63516 37738
rect 63076 36226 63150 36350
rect 63274 36226 63318 36350
rect 63442 36226 63516 36350
rect 63076 34838 63516 36226
rect 63076 34714 63150 34838
rect 63274 34714 63318 34838
rect 63442 34714 63516 34838
rect 63076 33326 63516 34714
rect 63076 33202 63150 33326
rect 63274 33202 63318 33326
rect 63442 33202 63516 33326
rect 63076 31814 63516 33202
rect 63076 31690 63150 31814
rect 63274 31690 63318 31814
rect 63442 31690 63516 31814
rect 63076 30302 63516 31690
rect 63076 30178 63150 30302
rect 63274 30178 63318 30302
rect 63442 30178 63516 30302
rect 63076 28790 63516 30178
rect 63076 28666 63150 28790
rect 63274 28666 63318 28790
rect 63442 28666 63516 28790
rect 63076 27278 63516 28666
rect 63076 27154 63150 27278
rect 63274 27154 63318 27278
rect 63442 27154 63516 27278
rect 63076 25766 63516 27154
rect 63076 25642 63150 25766
rect 63274 25642 63318 25766
rect 63442 25642 63516 25766
rect 63076 19665 63516 25642
rect 63076 19541 63150 19665
rect 63274 19541 63318 19665
rect 63442 19541 63516 19665
rect 63076 19497 63516 19541
rect 63076 19373 63150 19497
rect 63274 19373 63318 19497
rect 63442 19373 63516 19497
rect 63076 19329 63516 19373
rect 63076 19205 63150 19329
rect 63274 19205 63318 19329
rect 63442 19205 63516 19329
rect 63076 19161 63516 19205
rect 63076 19037 63150 19161
rect 63274 19037 63318 19161
rect 63442 19037 63516 19161
rect 63076 18993 63516 19037
rect 63076 18869 63150 18993
rect 63274 18869 63318 18993
rect 63442 18869 63516 18993
rect 63076 18825 63516 18869
rect 63076 18701 63150 18825
rect 63274 18701 63318 18825
rect 63442 18701 63516 18825
rect 63076 18657 63516 18701
rect 63076 18533 63150 18657
rect 63274 18533 63318 18657
rect 63442 18533 63516 18657
rect 63076 18489 63516 18533
rect 63076 18365 63150 18489
rect 63274 18365 63318 18489
rect 63442 18365 63516 18489
rect 63076 18321 63516 18365
rect 63076 18197 63150 18321
rect 63274 18197 63318 18321
rect 63442 18197 63516 18321
rect 63076 18153 63516 18197
rect 63076 18029 63150 18153
rect 63274 18029 63318 18153
rect 63442 18029 63516 18153
rect 63076 17985 63516 18029
rect 63076 17861 63150 17985
rect 63274 17861 63318 17985
rect 63442 17861 63516 17985
rect 63076 17817 63516 17861
rect 63076 17693 63150 17817
rect 63274 17693 63318 17817
rect 63442 17693 63516 17817
rect 63076 17649 63516 17693
rect 63076 17525 63150 17649
rect 63274 17525 63318 17649
rect 63442 17525 63516 17649
rect 63076 15182 63516 17525
rect 63076 15058 63150 15182
rect 63274 15058 63318 15182
rect 63442 15058 63516 15182
rect 63076 13670 63516 15058
rect 63076 13546 63150 13670
rect 63274 13546 63318 13670
rect 63442 13546 63516 13670
rect 63076 12158 63516 13546
rect 63076 12034 63150 12158
rect 63274 12034 63318 12158
rect 63442 12034 63516 12158
rect 63076 10646 63516 12034
rect 63076 10522 63150 10646
rect 63274 10522 63318 10646
rect 63442 10522 63516 10646
rect 63076 9134 63516 10522
rect 63076 9010 63150 9134
rect 63274 9010 63318 9134
rect 63442 9010 63516 9134
rect 63076 7622 63516 9010
rect 63076 7498 63150 7622
rect 63274 7498 63318 7622
rect 63442 7498 63516 7622
rect 63076 6110 63516 7498
rect 63076 5986 63150 6110
rect 63274 5986 63318 6110
rect 63442 5986 63516 6110
rect 63076 4598 63516 5986
rect 63076 4474 63150 4598
rect 63274 4474 63318 4598
rect 63442 4474 63516 4598
rect 63076 3086 63516 4474
rect 63076 2962 63150 3086
rect 63274 2962 63318 3086
rect 63442 2962 63516 3086
rect 63076 1574 63516 2962
rect 63076 1450 63150 1574
rect 63274 1450 63318 1574
rect 63442 1450 63516 1574
rect 63076 712 63516 1450
rect 64316 38494 64390 38618
rect 64514 38494 64558 38618
rect 64682 38494 64756 38618
rect 76316 38618 76756 38682
rect 64316 37106 64756 38494
rect 64316 36982 64390 37106
rect 64514 36982 64558 37106
rect 64682 36982 64756 37106
rect 64316 35594 64756 36982
rect 64316 35470 64390 35594
rect 64514 35470 64558 35594
rect 64682 35470 64756 35594
rect 64316 34082 64756 35470
rect 64316 33958 64390 34082
rect 64514 33958 64558 34082
rect 64682 33958 64756 34082
rect 64316 32570 64756 33958
rect 64316 32446 64390 32570
rect 64514 32446 64558 32570
rect 64682 32446 64756 32570
rect 64316 31058 64756 32446
rect 64316 30934 64390 31058
rect 64514 30934 64558 31058
rect 64682 30934 64756 31058
rect 64316 29546 64756 30934
rect 64316 29422 64390 29546
rect 64514 29422 64558 29546
rect 64682 29422 64756 29546
rect 64316 28034 64756 29422
rect 64316 27910 64390 28034
rect 64514 27910 64558 28034
rect 64682 27910 64756 28034
rect 64316 26522 64756 27910
rect 64316 26398 64390 26522
rect 64514 26398 64558 26522
rect 64682 26398 64756 26522
rect 64316 25010 64756 26398
rect 64316 24886 64390 25010
rect 64514 24886 64558 25010
rect 64682 24886 64756 25010
rect 64316 22541 64756 24886
rect 75076 37862 75516 38600
rect 75076 37738 75150 37862
rect 75274 37738 75318 37862
rect 75442 37738 75516 37862
rect 75076 36350 75516 37738
rect 75076 36226 75150 36350
rect 75274 36226 75318 36350
rect 75442 36226 75516 36350
rect 75076 34838 75516 36226
rect 75076 34714 75150 34838
rect 75274 34714 75318 34838
rect 75442 34714 75516 34838
rect 75076 33326 75516 34714
rect 75076 33202 75150 33326
rect 75274 33202 75318 33326
rect 75442 33202 75516 33326
rect 75076 31814 75516 33202
rect 75076 31690 75150 31814
rect 75274 31690 75318 31814
rect 75442 31690 75516 31814
rect 75076 30302 75516 31690
rect 75076 30178 75150 30302
rect 75274 30178 75318 30302
rect 75442 30178 75516 30302
rect 75076 28790 75516 30178
rect 75076 28666 75150 28790
rect 75274 28666 75318 28790
rect 75442 28666 75516 28790
rect 75076 27278 75516 28666
rect 75076 27154 75150 27278
rect 75274 27154 75318 27278
rect 75442 27154 75516 27278
rect 75076 25766 75516 27154
rect 75076 25642 75150 25766
rect 75274 25642 75318 25766
rect 75442 25642 75516 25766
rect 74036 23162 74364 23264
rect 74036 23038 74138 23162
rect 74262 23038 74364 23162
rect 64316 22417 64390 22541
rect 64514 22417 64558 22541
rect 64682 22417 64756 22541
rect 64316 22373 64756 22417
rect 64316 22249 64390 22373
rect 64514 22249 64558 22373
rect 64682 22249 64756 22373
rect 64316 22205 64756 22249
rect 64316 22081 64390 22205
rect 64514 22081 64558 22205
rect 64682 22081 64756 22205
rect 64316 22037 64756 22081
rect 64316 21913 64390 22037
rect 64514 21913 64558 22037
rect 64682 21913 64756 22037
rect 64316 21869 64756 21913
rect 64316 21745 64390 21869
rect 64514 21745 64558 21869
rect 64682 21745 64756 21869
rect 64316 21701 64756 21745
rect 64316 21577 64390 21701
rect 64514 21577 64558 21701
rect 64682 21577 64756 21701
rect 64316 21533 64756 21577
rect 64316 21409 64390 21533
rect 64514 21409 64558 21533
rect 64682 21409 64756 21533
rect 64316 21365 64756 21409
rect 64316 21241 64390 21365
rect 64514 21241 64558 21365
rect 64682 21241 64756 21365
rect 64316 21197 64756 21241
rect 64316 21073 64390 21197
rect 64514 21073 64558 21197
rect 64682 21073 64756 21197
rect 64316 21029 64756 21073
rect 64316 20905 64390 21029
rect 64514 20905 64558 21029
rect 64682 20905 64756 21029
rect 64316 20861 64756 20905
rect 64316 20737 64390 20861
rect 64514 20737 64558 20861
rect 64682 20737 64756 20861
rect 64316 20693 64756 20737
rect 64316 20569 64390 20693
rect 64514 20569 64558 20693
rect 64682 20569 64756 20693
rect 64316 20525 64756 20569
rect 64316 20401 64390 20525
rect 64514 20401 64558 20525
rect 64682 20401 64756 20525
rect 64316 14426 64756 20401
rect 71756 22826 72084 22928
rect 71756 22702 71858 22826
rect 71982 22702 72084 22826
rect 71756 16442 72084 22702
rect 74036 17282 74364 23038
rect 74036 17158 74138 17282
rect 74262 17158 74364 17282
rect 74036 17056 74364 17158
rect 75076 19665 75516 25642
rect 75076 19541 75150 19665
rect 75274 19541 75318 19665
rect 75442 19541 75516 19665
rect 75076 19497 75516 19541
rect 75076 19373 75150 19497
rect 75274 19373 75318 19497
rect 75442 19373 75516 19497
rect 75076 19329 75516 19373
rect 75076 19205 75150 19329
rect 75274 19205 75318 19329
rect 75442 19205 75516 19329
rect 75076 19161 75516 19205
rect 75076 19037 75150 19161
rect 75274 19037 75318 19161
rect 75442 19037 75516 19161
rect 75076 18993 75516 19037
rect 75076 18869 75150 18993
rect 75274 18869 75318 18993
rect 75442 18869 75516 18993
rect 75076 18825 75516 18869
rect 75076 18701 75150 18825
rect 75274 18701 75318 18825
rect 75442 18701 75516 18825
rect 75076 18657 75516 18701
rect 75076 18533 75150 18657
rect 75274 18533 75318 18657
rect 75442 18533 75516 18657
rect 75076 18489 75516 18533
rect 75076 18365 75150 18489
rect 75274 18365 75318 18489
rect 75442 18365 75516 18489
rect 75076 18321 75516 18365
rect 75076 18197 75150 18321
rect 75274 18197 75318 18321
rect 75442 18197 75516 18321
rect 75076 18153 75516 18197
rect 75076 18029 75150 18153
rect 75274 18029 75318 18153
rect 75442 18029 75516 18153
rect 75076 17985 75516 18029
rect 75076 17861 75150 17985
rect 75274 17861 75318 17985
rect 75442 17861 75516 17985
rect 75076 17817 75516 17861
rect 75076 17693 75150 17817
rect 75274 17693 75318 17817
rect 75442 17693 75516 17817
rect 75076 17649 75516 17693
rect 75076 17525 75150 17649
rect 75274 17525 75318 17649
rect 75442 17525 75516 17649
rect 71756 16318 71858 16442
rect 71982 16318 72084 16442
rect 71756 16216 72084 16318
rect 64316 14302 64390 14426
rect 64514 14302 64558 14426
rect 64682 14302 64756 14426
rect 64316 12914 64756 14302
rect 64316 12790 64390 12914
rect 64514 12790 64558 12914
rect 64682 12790 64756 12914
rect 64316 11402 64756 12790
rect 64316 11278 64390 11402
rect 64514 11278 64558 11402
rect 64682 11278 64756 11402
rect 64316 9890 64756 11278
rect 64316 9766 64390 9890
rect 64514 9766 64558 9890
rect 64682 9766 64756 9890
rect 64316 8378 64756 9766
rect 64316 8254 64390 8378
rect 64514 8254 64558 8378
rect 64682 8254 64756 8378
rect 64316 6866 64756 8254
rect 64316 6742 64390 6866
rect 64514 6742 64558 6866
rect 64682 6742 64756 6866
rect 64316 5354 64756 6742
rect 64316 5230 64390 5354
rect 64514 5230 64558 5354
rect 64682 5230 64756 5354
rect 64316 3842 64756 5230
rect 64316 3718 64390 3842
rect 64514 3718 64558 3842
rect 64682 3718 64756 3842
rect 64316 2330 64756 3718
rect 64316 2206 64390 2330
rect 64514 2206 64558 2330
rect 64682 2206 64756 2330
rect 64316 818 64756 2206
rect 52316 630 52756 694
rect 64316 694 64390 818
rect 64514 694 64558 818
rect 64682 694 64756 818
rect 75076 15182 75516 17525
rect 75076 15058 75150 15182
rect 75274 15058 75318 15182
rect 75442 15058 75516 15182
rect 75076 13670 75516 15058
rect 75076 13546 75150 13670
rect 75274 13546 75318 13670
rect 75442 13546 75516 13670
rect 75076 12158 75516 13546
rect 75076 12034 75150 12158
rect 75274 12034 75318 12158
rect 75442 12034 75516 12158
rect 75076 10646 75516 12034
rect 75076 10522 75150 10646
rect 75274 10522 75318 10646
rect 75442 10522 75516 10646
rect 75076 9134 75516 10522
rect 75076 9010 75150 9134
rect 75274 9010 75318 9134
rect 75442 9010 75516 9134
rect 75076 7622 75516 9010
rect 75076 7498 75150 7622
rect 75274 7498 75318 7622
rect 75442 7498 75516 7622
rect 75076 6110 75516 7498
rect 75076 5986 75150 6110
rect 75274 5986 75318 6110
rect 75442 5986 75516 6110
rect 75076 4598 75516 5986
rect 75076 4474 75150 4598
rect 75274 4474 75318 4598
rect 75442 4474 75516 4598
rect 75076 3086 75516 4474
rect 75076 2962 75150 3086
rect 75274 2962 75318 3086
rect 75442 2962 75516 3086
rect 75076 1574 75516 2962
rect 75076 1450 75150 1574
rect 75274 1450 75318 1574
rect 75442 1450 75516 1574
rect 75076 712 75516 1450
rect 76316 38494 76390 38618
rect 76514 38494 76558 38618
rect 76682 38494 76756 38618
rect 76316 37106 76756 38494
rect 76316 36982 76390 37106
rect 76514 36982 76558 37106
rect 76682 36982 76756 37106
rect 76316 35594 76756 36982
rect 76316 35470 76390 35594
rect 76514 35470 76558 35594
rect 76682 35470 76756 35594
rect 76316 34082 76756 35470
rect 76316 33958 76390 34082
rect 76514 33958 76558 34082
rect 76682 33958 76756 34082
rect 76316 32570 76756 33958
rect 76316 32446 76390 32570
rect 76514 32446 76558 32570
rect 76682 32446 76756 32570
rect 76316 31058 76756 32446
rect 76316 30934 76390 31058
rect 76514 30934 76558 31058
rect 76682 30934 76756 31058
rect 76316 29546 76756 30934
rect 76316 29422 76390 29546
rect 76514 29422 76558 29546
rect 76682 29422 76756 29546
rect 76316 28034 76756 29422
rect 76316 27910 76390 28034
rect 76514 27910 76558 28034
rect 76682 27910 76756 28034
rect 76316 26522 76756 27910
rect 76316 26398 76390 26522
rect 76514 26398 76558 26522
rect 76682 26398 76756 26522
rect 76316 25010 76756 26398
rect 76316 24886 76390 25010
rect 76514 24886 76558 25010
rect 76682 24886 76756 25010
rect 76316 22541 76756 24886
rect 76316 22417 76390 22541
rect 76514 22417 76558 22541
rect 76682 22417 76756 22541
rect 76316 22373 76756 22417
rect 76316 22249 76390 22373
rect 76514 22249 76558 22373
rect 76682 22249 76756 22373
rect 76316 22205 76756 22249
rect 76316 22081 76390 22205
rect 76514 22081 76558 22205
rect 76682 22081 76756 22205
rect 76316 22037 76756 22081
rect 76316 21913 76390 22037
rect 76514 21913 76558 22037
rect 76682 21913 76756 22037
rect 76316 21869 76756 21913
rect 76316 21745 76390 21869
rect 76514 21745 76558 21869
rect 76682 21745 76756 21869
rect 76316 21701 76756 21745
rect 76316 21577 76390 21701
rect 76514 21577 76558 21701
rect 76682 21577 76756 21701
rect 76316 21533 76756 21577
rect 76316 21409 76390 21533
rect 76514 21409 76558 21533
rect 76682 21409 76756 21533
rect 76316 21365 76756 21409
rect 76316 21241 76390 21365
rect 76514 21241 76558 21365
rect 76682 21241 76756 21365
rect 76316 21197 76756 21241
rect 76316 21073 76390 21197
rect 76514 21073 76558 21197
rect 76682 21073 76756 21197
rect 76316 21029 76756 21073
rect 76316 20905 76390 21029
rect 76514 20905 76558 21029
rect 76682 20905 76756 21029
rect 76316 20861 76756 20905
rect 76316 20737 76390 20861
rect 76514 20737 76558 20861
rect 76682 20737 76756 20861
rect 76316 20693 76756 20737
rect 76316 20569 76390 20693
rect 76514 20569 76558 20693
rect 76682 20569 76756 20693
rect 76316 20525 76756 20569
rect 76316 20401 76390 20525
rect 76514 20401 76558 20525
rect 76682 20401 76756 20525
rect 76316 14426 76756 20401
rect 78596 23834 78924 23936
rect 78596 23710 78698 23834
rect 78822 23710 78924 23834
rect 78596 16274 78924 23710
rect 78596 16150 78698 16274
rect 78822 16150 78924 16274
rect 78596 16048 78924 16150
rect 76316 14302 76390 14426
rect 76514 14302 76558 14426
rect 76682 14302 76756 14426
rect 76316 12914 76756 14302
rect 76316 12790 76390 12914
rect 76514 12790 76558 12914
rect 76682 12790 76756 12914
rect 76316 11402 76756 12790
rect 76316 11278 76390 11402
rect 76514 11278 76558 11402
rect 76682 11278 76756 11402
rect 76316 9890 76756 11278
rect 76316 9766 76390 9890
rect 76514 9766 76558 9890
rect 76682 9766 76756 9890
rect 76316 8378 76756 9766
rect 76316 8254 76390 8378
rect 76514 8254 76558 8378
rect 76682 8254 76756 8378
rect 76316 6866 76756 8254
rect 76316 6742 76390 6866
rect 76514 6742 76558 6866
rect 76682 6742 76756 6866
rect 76316 5354 76756 6742
rect 76316 5230 76390 5354
rect 76514 5230 76558 5354
rect 76682 5230 76756 5354
rect 76316 3842 76756 5230
rect 76316 3718 76390 3842
rect 76514 3718 76558 3842
rect 76682 3718 76756 3842
rect 76316 2330 76756 3718
rect 76316 2206 76390 2330
rect 76514 2206 76558 2330
rect 76682 2206 76756 2330
rect 76316 818 76756 2206
rect 64316 630 64756 694
rect 76316 694 76390 818
rect 76514 694 76558 818
rect 76682 694 76756 818
rect 76316 630 76756 694
use sg13g2_inv_1  _0898_
timestamp 1676382929
transform -1 0 11136 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0899_
timestamp 1676382929
transform 1 0 4992 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _0900_
timestamp 1676382929
transform 1 0 51744 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0901_
timestamp 1676382929
transform 1 0 9696 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0902_
timestamp 1676382929
transform -1 0 13824 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0903_
timestamp 1676382929
transform 1 0 52416 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0904_
timestamp 1676382929
transform 1 0 6240 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0905_
timestamp 1676382929
transform -1 0 52704 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0906_
timestamp 1676382929
transform 1 0 2880 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0907_
timestamp 1676382929
transform 1 0 43392 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0908_
timestamp 1676382929
transform -1 0 47616 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0909_
timestamp 1676382929
transform 1 0 51744 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0910_
timestamp 1676382929
transform -1 0 51456 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0911_
timestamp 1676382929
transform -1 0 47520 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0912_
timestamp 1676382929
transform -1 0 45216 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0913_
timestamp 1676382929
transform -1 0 41088 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0914_
timestamp 1676382929
transform 1 0 38112 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0915_
timestamp 1676382929
transform 1 0 34560 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0916_
timestamp 1676382929
transform -1 0 33312 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0917_
timestamp 1676382929
transform -1 0 36960 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0918_
timestamp 1676382929
transform 1 0 38976 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0919_
timestamp 1676382929
transform 1 0 40992 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0920_
timestamp 1676382929
transform -1 0 43008 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0921_
timestamp 1676382929
transform 1 0 47712 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0922_
timestamp 1676382929
transform 1 0 47616 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0923_
timestamp 1676382929
transform -1 0 43680 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0924_
timestamp 1676382929
transform -1 0 47328 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0925_
timestamp 1676382929
transform 1 0 49248 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0926_
timestamp 1676382929
transform -1 0 52992 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0927_
timestamp 1676382929
transform 1 0 52128 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0928_
timestamp 1676382929
transform 1 0 50976 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0929_
timestamp 1676382929
transform -1 0 53664 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0930_
timestamp 1676382929
transform 1 0 56832 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0931_
timestamp 1676382929
transform 1 0 57120 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0932_
timestamp 1676382929
transform 1 0 56544 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0933_
timestamp 1676382929
transform 1 0 56160 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0934_
timestamp 1676382929
transform -1 0 53568 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0935_
timestamp 1676382929
transform 1 0 56544 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0936_
timestamp 1676382929
transform 1 0 57888 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0937_
timestamp 1676382929
transform 1 0 62112 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0938_
timestamp 1676382929
transform 1 0 63168 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _0939_
timestamp 1676382929
transform 1 0 62016 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0940_
timestamp 1676382929
transform -1 0 60672 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0941_
timestamp 1676382929
transform 1 0 60000 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0942_
timestamp 1676382929
transform 1 0 59424 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0943_
timestamp 1676382929
transform -1 0 67680 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0944_
timestamp 1676382929
transform 1 0 63744 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0945_
timestamp 1676382929
transform 1 0 63552 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0946_
timestamp 1676382929
transform 1 0 64800 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0947_
timestamp 1676382929
transform -1 0 66912 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0948_
timestamp 1676382929
transform 1 0 65568 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0949_
timestamp 1676382929
transform 1 0 66528 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0950_
timestamp 1676382929
transform 1 0 69792 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0951_
timestamp 1676382929
transform 1 0 69504 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0952_
timestamp 1676382929
transform 1 0 70176 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0953_
timestamp 1676382929
transform 1 0 68352 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0954_
timestamp 1676382929
transform 1 0 65952 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0955_
timestamp 1676382929
transform 1 0 72384 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0956_
timestamp 1676382929
transform 1 0 72096 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0957_
timestamp 1676382929
transform 1 0 73248 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0958_
timestamp 1676382929
transform 1 0 73824 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0959_
timestamp 1676382929
transform 1 0 74016 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0960_
timestamp 1676382929
transform 1 0 74400 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0961_
timestamp 1676382929
transform 1 0 74880 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0962_
timestamp 1676382929
transform 1 0 74208 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0963_
timestamp 1676382929
transform 1 0 74880 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _0964_
timestamp 1676382929
transform 1 0 76608 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _0965_
timestamp 1676382929
transform -1 0 77088 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0966_
timestamp 1676382929
transform 1 0 78624 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0967_
timestamp 1676382929
transform 1 0 77952 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0968_
timestamp 1676382929
transform -1 0 78336 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0969_
timestamp 1676382929
transform -1 0 78432 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0970_
timestamp 1676382929
transform 1 0 77664 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0971_
timestamp 1676382929
transform -1 0 77376 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0972_
timestamp 1676382929
transform -1 0 78336 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _0973_
timestamp 1676382929
transform -1 0 78720 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0974_
timestamp 1676382929
transform -1 0 78144 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0975_
timestamp 1676382929
transform -1 0 78240 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0976_
timestamp 1676382929
transform 1 0 76224 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0977_
timestamp 1676382929
transform -1 0 76992 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0978_
timestamp 1676382929
transform 1 0 75264 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0979_
timestamp 1676382929
transform 1 0 74688 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0980_
timestamp 1676382929
transform 1 0 72480 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0981_
timestamp 1676382929
transform -1 0 74592 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0982_
timestamp 1676382929
transform 1 0 73920 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0983_
timestamp 1676382929
transform -1 0 73824 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0984_
timestamp 1676382929
transform 1 0 73248 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0985_
timestamp 1676382929
transform -1 0 72960 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0986_
timestamp 1676382929
transform -1 0 72576 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0987_
timestamp 1676382929
transform -1 0 72192 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0988_
timestamp 1676382929
transform 1 0 64704 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0989_
timestamp 1676382929
transform 1 0 66432 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0990_
timestamp 1676382929
transform 1 0 67296 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0991_
timestamp 1676382929
transform 1 0 68928 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0992_
timestamp 1676382929
transform -1 0 69792 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0993_
timestamp 1676382929
transform 1 0 69216 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0994_
timestamp 1676382929
transform -1 0 65952 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0995_
timestamp 1676382929
transform 1 0 61632 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0996_
timestamp 1676382929
transform 1 0 57120 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0997_
timestamp 1676382929
transform 1 0 59808 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0998_
timestamp 1676382929
transform 1 0 65088 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0999_
timestamp 1676382929
transform 1 0 63840 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1000_
timestamp 1676382929
transform 1 0 62016 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1001_
timestamp 1676382929
transform -1 0 59328 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1002_
timestamp 1676382929
transform 1 0 56256 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1003_
timestamp 1676382929
transform -1 0 53280 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1004_
timestamp 1676382929
transform 1 0 51936 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1005_
timestamp 1676382929
transform 1 0 55008 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1006_
timestamp 1676382929
transform 1 0 57984 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1007_
timestamp 1676382929
transform -1 0 62976 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1008_
timestamp 1676382929
transform -1 0 62784 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1009_
timestamp 1676382929
transform -1 0 60480 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1010_
timestamp 1676382929
transform -1 0 57984 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1011_
timestamp 1676382929
transform -1 0 55200 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1012_
timestamp 1676382929
transform -1 0 53280 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1013_
timestamp 1676382929
transform 1 0 49152 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1014_
timestamp 1676382929
transform 1 0 48960 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1015_
timestamp 1676382929
transform -1 0 48960 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1016_
timestamp 1676382929
transform 1 0 52224 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1017_
timestamp 1676382929
transform -1 0 51360 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1018_
timestamp 1676382929
transform -1 0 47328 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1019_
timestamp 1676382929
transform 1 0 43296 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1020_
timestamp 1676382929
transform 1 0 44832 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1021_
timestamp 1676382929
transform -1 0 45792 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1022_
timestamp 1676382929
transform 1 0 43584 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1023_
timestamp 1676382929
transform 1 0 40896 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1024_
timestamp 1676382929
transform -1 0 39648 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1025_
timestamp 1676382929
transform -1 0 37632 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1026_
timestamp 1676382929
transform 1 0 37632 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1027_
timestamp 1676382929
transform -1 0 56160 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1028_
timestamp 1676382929
transform -1 0 55776 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1029_
timestamp 1676382929
transform 1 0 52128 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1030_
timestamp 1676382929
transform 1 0 51456 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1031_
timestamp 1676382929
transform 1 0 52128 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1032_
timestamp 1676382929
transform -1 0 43008 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1033_
timestamp 1676382929
transform -1 0 47328 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1034_
timestamp 1676382929
transform 1 0 50880 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1035_
timestamp 1676382929
transform 1 0 49536 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1036_
timestamp 1676382929
transform 1 0 45408 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1037_
timestamp 1676382929
transform 1 0 43008 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1038_
timestamp 1676382929
transform 1 0 41088 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1039_
timestamp 1676382929
transform 1 0 37440 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1040_
timestamp 1676382929
transform 1 0 33312 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1041_
timestamp 1676382929
transform -1 0 33600 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1042_
timestamp 1676382929
transform -1 0 36384 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1043_
timestamp 1676382929
transform -1 0 38592 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1044_
timestamp 1676382929
transform -1 0 41280 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1045_
timestamp 1676382929
transform -1 0 43392 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1046_
timestamp 1676382929
transform -1 0 45792 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1047_
timestamp 1676382929
transform 1 0 46176 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1048_
timestamp 1676382929
transform -1 0 44352 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1049_
timestamp 1676382929
transform -1 0 47040 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _1050_
timestamp 1676382929
transform -1 0 49440 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1051_
timestamp 1676382929
transform 1 0 52416 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1052_
timestamp 1676382929
transform 1 0 50496 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1053_
timestamp 1676382929
transform -1 0 50496 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1054_
timestamp 1676382929
transform 1 0 54336 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1055_
timestamp 1676382929
transform -1 0 55392 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1056_
timestamp 1676382929
transform 1 0 56352 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1057_
timestamp 1676382929
transform -1 0 55584 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1058_
timestamp 1676382929
transform 1 0 53760 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1059_
timestamp 1676382929
transform -1 0 53568 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1060_
timestamp 1676382929
transform -1 0 55968 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1061_
timestamp 1676382929
transform -1 0 58080 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1062_
timestamp 1676382929
transform -1 0 60384 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1063_
timestamp 1676382929
transform 1 0 62784 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1064_
timestamp 1676382929
transform 1 0 60384 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1065_
timestamp 1676382929
transform -1 0 58560 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1066_
timestamp 1676382929
transform -1 0 58368 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1067_
timestamp 1676382929
transform -1 0 59424 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1068_
timestamp 1676382929
transform 1 0 62496 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1069_
timestamp 1676382929
transform 1 0 62784 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1070_
timestamp 1676382929
transform 1 0 63168 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1071_
timestamp 1676382929
transform -1 0 64224 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _1072_
timestamp 1676382929
transform 1 0 64800 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _1073_
timestamp 1676382929
transform -1 0 65088 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1074_
timestamp 1676382929
transform -1 0 66336 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  _1075_
timestamp 1676382929
transform -1 0 69312 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1076_
timestamp 1676382929
transform -1 0 69504 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1077_
timestamp 1676382929
transform 1 0 67872 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _1078_
timestamp 1676382929
transform 1 0 66816 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1079_
timestamp 1676382929
transform -1 0 66624 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1080_
timestamp 1676382929
transform -1 0 68352 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1081_
timestamp 1676382929
transform -1 0 70752 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1082_
timestamp 1676382929
transform 1 0 72000 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1083_
timestamp 1676382929
transform -1 0 72288 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1084_
timestamp 1676382929
transform 1 0 72768 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1085_
timestamp 1676382929
transform 1 0 72576 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _1086_
timestamp 1676382929
transform 1 0 73056 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1087_
timestamp 1676382929
transform 1 0 72864 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1088_
timestamp 1676382929
transform -1 0 73632 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1089_
timestamp 1676382929
transform -1 0 78048 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1090_
timestamp 1676382929
transform -1 0 78240 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1091_
timestamp 1676382929
transform -1 0 78528 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1092_
timestamp 1676382929
transform -1 0 78240 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1093_
timestamp 1676382929
transform 1 0 77856 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1094_
timestamp 1676382929
transform 1 0 76128 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1095_
timestamp 1676382929
transform 1 0 75264 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1096_
timestamp 1676382929
transform -1 0 75744 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1097_
timestamp 1676382929
transform -1 0 76992 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1098_
timestamp 1676382929
transform 1 0 77664 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1099_
timestamp 1676382929
transform 1 0 77568 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1100_
timestamp 1676382929
transform -1 0 78336 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _1101_
timestamp 1676382929
transform -1 0 78144 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _1102_
timestamp 1676382929
transform -1 0 76704 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _1103_
timestamp 1676382929
transform 1 0 73152 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _1104_
timestamp 1676382929
transform 1 0 72000 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _1105_
timestamp 1676382929
transform 1 0 70848 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _1106_
timestamp 1676382929
transform 1 0 72480 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _1107_
timestamp 1676382929
transform 1 0 71712 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1108_
timestamp 1676382929
transform 1 0 70944 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _1109_
timestamp 1676382929
transform -1 0 71328 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1110_
timestamp 1676382929
transform 1 0 71040 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1111_
timestamp 1676382929
transform 1 0 68544 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1112_
timestamp 1676382929
transform 1 0 65376 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1113_
timestamp 1676382929
transform 1 0 64800 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1114_
timestamp 1676382929
transform 1 0 65568 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1115_
timestamp 1676382929
transform 1 0 67008 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1116_
timestamp 1676382929
transform 1 0 67968 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _1117_
timestamp 1676382929
transform -1 0 68352 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _1118_
timestamp 1676382929
transform 1 0 65664 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _1119_
timestamp 1676382929
transform 1 0 63744 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _1120_
timestamp 1676382929
transform 1 0 59808 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _1121_
timestamp 1676382929
transform -1 0 57792 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _1122_
timestamp 1676382929
transform -1 0 60384 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _1123_
timestamp 1676382929
transform -1 0 63744 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _1124_
timestamp 1676382929
transform 1 0 62688 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _1125_
timestamp 1676382929
transform 1 0 60288 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _1126_
timestamp 1676382929
transform 1 0 57024 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1127_
timestamp 1676382929
transform 1 0 55104 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _1128_
timestamp 1676382929
transform 1 0 51840 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _1129_
timestamp 1676382929
transform -1 0 52320 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _1130_
timestamp 1676382929
transform -1 0 55488 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _1131_
timestamp 1676382929
transform -1 0 58368 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _1132_
timestamp 1676382929
transform -1 0 60768 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1133_
timestamp 1676382929
transform 1 0 61728 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1134_
timestamp 1676382929
transform 1 0 58368 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1135_
timestamp 1676382929
transform 1 0 55776 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1136_
timestamp 1676382929
transform 1 0 53280 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1137_
timestamp 1676382929
transform 1 0 52128 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _1138_
timestamp 1676382929
transform 1 0 47904 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _1139_
timestamp 1676382929
transform -1 0 47520 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1140_
timestamp 1676382929
transform -1 0 49344 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1141_
timestamp 1676382929
transform -1 0 51168 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1142_
timestamp 1676382929
transform 1 0 49440 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1143_
timestamp 1676382929
transform 1 0 45792 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1144_
timestamp 1676382929
transform 1 0 43008 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1145_
timestamp 1676382929
transform -1 0 43584 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1146_
timestamp 1676382929
transform -1 0 44160 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1147_
timestamp 1676382929
transform 1 0 42048 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1148_
timestamp 1676382929
transform 1 0 39360 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1149_
timestamp 1676382929
transform 1 0 37632 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1150_
timestamp 1676382929
transform 1 0 36960 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1151_
timestamp 1676382929
transform 1 0 35136 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1152_
timestamp 1676382929
transform 1 0 31488 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1153_
timestamp 1676382929
transform 1 0 3648 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _1154_
timestamp 1676382929
transform -1 0 7104 0 1 15876
box -48 -56 336 834
use sg13g2_o21ai_1  _1155_
timestamp 1685175443
transform -1 0 43008 0 -1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1156_
timestamp 1677175127
transform 1 0 41856 0 -1 20412
box -48 -56 720 834
use sg13g2_nor2_1  _1157_
timestamp 1676627187
transform -1 0 1824 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1158_
timestamp 1683973020
transform -1 0 40416 0 -1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1159_
timestamp 1685173987
transform 1 0 40416 0 -1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1160_
timestamp 1685175443
transform -1 0 47232 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1161_
timestamp 1677175127
transform 1 0 46080 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1162_
timestamp 1683973020
transform -1 0 44448 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1163_
timestamp 1685173987
transform -1 0 45984 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1164_
timestamp 1685175443
transform -1 0 51360 0 -1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1165_
timestamp 1677175127
transform 1 0 49536 0 -1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1166_
timestamp 1683973020
transform -1 0 48192 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1167_
timestamp 1685173987
transform -1 0 48768 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1168_
timestamp 1685175443
transform -1 0 50880 0 1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1169_
timestamp 1677175127
transform -1 0 50496 0 1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1170_
timestamp 1683973020
transform 1 0 49056 0 -1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1171_
timestamp 1685173987
transform -1 0 50208 0 1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1172_
timestamp 1685175443
transform -1 0 47040 0 -1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1173_
timestamp 1677175127
transform -1 0 46464 0 1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1174_
timestamp 1683973020
transform 1 0 47232 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1175_
timestamp 1685173987
transform 1 0 46656 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1176_
timestamp 1685175443
transform 1 0 43968 0 1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1177_
timestamp 1677175127
transform -1 0 43968 0 1 17388
box -48 -56 720 834
use sg13g2_a21oi_1  _1178_
timestamp 1683973020
transform 1 0 44064 0 -1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1179_
timestamp 1685173987
transform 1 0 43200 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1180_
timestamp 1685175443
transform -1 0 41088 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1181_
timestamp 1677175127
transform 1 0 39936 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1182_
timestamp 1683973020
transform 1 0 41088 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1183_
timestamp 1685173987
transform -1 0 39936 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1184_
timestamp 1685175443
transform 1 0 37344 0 1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1185_
timestamp 1677175127
transform 1 0 36768 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1186_
timestamp 1683973020
transform 1 0 38016 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1187_
timestamp 1685173987
transform 1 0 36192 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1188_
timestamp 1685175443
transform -1 0 33792 0 1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1189_
timestamp 1677175127
transform 1 0 32736 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1190_
timestamp 1683973020
transform 1 0 33600 0 -1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1191_
timestamp 1685173987
transform 1 0 32736 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1192_
timestamp 1685175443
transform -1 0 33216 0 1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1193_
timestamp 1677175127
transform 1 0 32160 0 -1 17388
box -48 -56 720 834
use sg13g2_a21oi_1  _1194_
timestamp 1683973020
transform -1 0 32544 0 1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1195_
timestamp 1685173987
transform 1 0 31968 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1196_
timestamp 1685175443
transform -1 0 36480 0 1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1197_
timestamp 1677175127
transform 1 0 35424 0 -1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1198_
timestamp 1683973020
transform -1 0 34656 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1199_
timestamp 1685173987
transform -1 0 35232 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1200_
timestamp 1685175443
transform -1 0 38784 0 -1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1201_
timestamp 1677175127
transform 1 0 37632 0 -1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1202_
timestamp 1683973020
transform -1 0 37056 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1203_
timestamp 1685173987
transform -1 0 37536 0 1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1204_
timestamp 1685175443
transform -1 0 40992 0 -1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1205_
timestamp 1677175127
transform 1 0 39840 0 -1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1206_
timestamp 1683973020
transform -1 0 39072 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1207_
timestamp 1685173987
transform -1 0 39840 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1208_
timestamp 1685175443
transform -1 0 43392 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1209_
timestamp 1677175127
transform 1 0 42336 0 -1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1210_
timestamp 1683973020
transform -1 0 41664 0 -1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1211_
timestamp 1685173987
transform -1 0 42144 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1212_
timestamp 1685175443
transform -1 0 47136 0 -1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1213_
timestamp 1677175127
transform 1 0 44736 0 -1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1214_
timestamp 1683973020
transform -1 0 44160 0 -1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1215_
timestamp 1685173987
transform -1 0 44928 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1216_
timestamp 1685175443
transform 1 0 46272 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1217_
timestamp 1677175127
transform -1 0 47040 0 1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1218_
timestamp 1683973020
transform -1 0 46272 0 -1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1219_
timestamp 1685173987
transform 1 0 45600 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1220_
timestamp 1685175443
transform -1 0 44064 0 -1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1221_
timestamp 1677175127
transform 1 0 42912 0 -1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1222_
timestamp 1683973020
transform 1 0 44064 0 -1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1223_
timestamp 1685173987
transform 1 0 43008 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1224_
timestamp 1685175443
transform -1 0 46944 0 -1 9828
box -48 -56 538 834
use sg13g2_a21o_1  _1225_
timestamp 1677175127
transform 1 0 45792 0 -1 9828
box -48 -56 720 834
use sg13g2_a21oi_1  _1226_
timestamp 1683973020
transform -1 0 45216 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1227_
timestamp 1685173987
transform -1 0 45792 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1228_
timestamp 1685175443
transform -1 0 49440 0 1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1229_
timestamp 1677175127
transform 1 0 48288 0 1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1230_
timestamp 1683973020
transform -1 0 47904 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1231_
timestamp 1685173987
transform -1 0 48384 0 1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  _1232_
timestamp 1685175443
transform -1 0 52320 0 -1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1233_
timestamp 1677175127
transform 1 0 51168 0 1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1234_
timestamp 1683973020
transform -1 0 50496 0 1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1235_
timestamp 1685173987
transform -1 0 50976 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1236_
timestamp 1685175443
transform -1 0 51936 0 1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1237_
timestamp 1677175127
transform -1 0 51456 0 1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1238_
timestamp 1683973020
transform 1 0 51072 0 1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1239_
timestamp 1685173987
transform 1 0 50592 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1240_
timestamp 1685175443
transform -1 0 50112 0 -1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1241_
timestamp 1677175127
transform 1 0 49248 0 1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1242_
timestamp 1683973020
transform 1 0 49632 0 -1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1243_
timestamp 1685173987
transform -1 0 48576 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1244_
timestamp 1685175443
transform -1 0 53376 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1245_
timestamp 1677175127
transform 1 0 52224 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1246_
timestamp 1683973020
transform -1 0 51552 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1247_
timestamp 1685173987
transform -1 0 52224 0 1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1248_
timestamp 1685175443
transform -1 0 56160 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1249_
timestamp 1677175127
transform 1 0 55008 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1250_
timestamp 1683973020
transform -1 0 54336 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1251_
timestamp 1685173987
transform -1 0 54816 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1252_
timestamp 1685175443
transform -1 0 56832 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1253_
timestamp 1677175127
transform 1 0 55680 0 -1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1254_
timestamp 1683973020
transform 1 0 55392 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1255_
timestamp 1685173987
transform -1 0 55680 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1256_
timestamp 1685175443
transform -1 0 56352 0 1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1257_
timestamp 1677175127
transform -1 0 55968 0 1 9828
box -48 -56 720 834
use sg13g2_a21oi_1  _1258_
timestamp 1683973020
transform 1 0 55104 0 -1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1259_
timestamp 1685173987
transform -1 0 55296 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1260_
timestamp 1685175443
transform -1 0 56256 0 -1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1261_
timestamp 1677175127
transform -1 0 55296 0 -1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1262_
timestamp 1683973020
transform 1 0 54816 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1263_
timestamp 1685173987
transform 1 0 54048 0 -1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1264_
timestamp 1685175443
transform -1 0 53856 0 -1 6804
box -48 -56 538 834
use sg13g2_a21o_1  _1265_
timestamp 1677175127
transform 1 0 52224 0 -1 6804
box -48 -56 720 834
use sg13g2_a21oi_1  _1266_
timestamp 1683973020
transform 1 0 52896 0 -1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1267_
timestamp 1685173987
transform 1 0 52128 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _1268_
timestamp 1685175443
transform -1 0 56352 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1269_
timestamp 1677175127
transform 1 0 55104 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1270_
timestamp 1683973020
transform -1 0 54336 0 -1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _1271_
timestamp 1685173987
transform -1 0 54912 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _1272_
timestamp 1685175443
transform -1 0 58080 0 1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _1273_
timestamp 1677175127
transform 1 0 56928 0 1 3780
box -48 -56 720 834
use sg13g2_a21oi_1  _1274_
timestamp 1683973020
transform -1 0 56832 0 1 3780
box -48 -56 528 834
use sg13g2_a22oi_1  _1275_
timestamp 1685173987
transform -1 0 56832 0 1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1276_
timestamp 1685175443
transform -1 0 60960 0 -1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _1277_
timestamp 1677175127
transform 1 0 59712 0 -1 3780
box -48 -56 720 834
use sg13g2_a21oi_1  _1278_
timestamp 1683973020
transform -1 0 58848 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1279_
timestamp 1685173987
transform -1 0 59424 0 1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1280_
timestamp 1685175443
transform -1 0 62976 0 1 756
box -48 -56 538 834
use sg13g2_a21o_1  _1281_
timestamp 1677175127
transform 1 0 61632 0 1 2268
box -48 -56 720 834
use sg13g2_a21oi_1  _1282_
timestamp 1683973020
transform -1 0 60864 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1283_
timestamp 1685173987
transform -1 0 61440 0 1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1284_
timestamp 1685175443
transform -1 0 61920 0 1 6804
box -48 -56 538 834
use sg13g2_a21o_1  _1285_
timestamp 1677175127
transform 1 0 60864 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1286_
timestamp 1683973020
transform 1 0 61248 0 -1 3780
box -48 -56 528 834
use sg13g2_a22oi_1  _1287_
timestamp 1685173987
transform 1 0 60672 0 -1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _1288_
timestamp 1685175443
transform -1 0 60960 0 -1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1289_
timestamp 1677175127
transform -1 0 60000 0 -1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1290_
timestamp 1683973020
transform -1 0 60192 0 -1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1291_
timestamp 1685173987
transform 1 0 59616 0 1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  _1292_
timestamp 1685175443
transform -1 0 59904 0 1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1293_
timestamp 1677175127
transform 1 0 58848 0 1 9828
box -48 -56 720 834
use sg13g2_a21oi_1  _1294_
timestamp 1683973020
transform 1 0 59040 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1295_
timestamp 1685173987
transform -1 0 59040 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1296_
timestamp 1685175443
transform 1 0 58560 0 1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1297_
timestamp 1677175127
transform 1 0 58176 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1298_
timestamp 1683973020
transform 1 0 58368 0 1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1299_
timestamp 1685173987
transform 1 0 57984 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1300_
timestamp 1685175443
transform -1 0 62208 0 -1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1301_
timestamp 1677175127
transform 1 0 60960 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1302_
timestamp 1683973020
transform -1 0 59904 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1303_
timestamp 1685173987
transform -1 0 60864 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1304_
timestamp 1685175443
transform -1 0 63552 0 -1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1305_
timestamp 1677175127
transform 1 0 62496 0 1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1306_
timestamp 1683973020
transform 1 0 61440 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1307_
timestamp 1685173987
transform -1 0 62496 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1308_
timestamp 1685175443
transform -1 0 63840 0 -1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1309_
timestamp 1677175127
transform 1 0 62208 0 -1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1310_
timestamp 1683973020
transform 1 0 62112 0 1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1311_
timestamp 1685173987
transform -1 0 62208 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1312_
timestamp 1685175443
transform -1 0 64608 0 1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1313_
timestamp 1677175127
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1314_
timestamp 1683973020
transform 1 0 62592 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1315_
timestamp 1685173987
transform -1 0 63360 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1316_
timestamp 1685175443
transform -1 0 66624 0 -1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1317_
timestamp 1677175127
transform -1 0 65760 0 1 6804
box -48 -56 720 834
use sg13g2_a21oi_1  _1318_
timestamp 1683973020
transform -1 0 64704 0 1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1319_
timestamp 1685173987
transform -1 0 64992 0 1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _1320_
timestamp 1685175443
transform -1 0 65952 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1321_
timestamp 1677175127
transform 1 0 64512 0 -1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1322_
timestamp 1683973020
transform -1 0 64512 0 -1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _1323_
timestamp 1685173987
transform -1 0 64800 0 -1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _1324_
timestamp 1685175443
transform 1 0 65376 0 -1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _1325_
timestamp 1677175127
transform -1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_a21oi_1  _1326_
timestamp 1683973020
transform 1 0 64320 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1327_
timestamp 1685173987
transform -1 0 65376 0 1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1328_
timestamp 1685175443
transform -1 0 69888 0 1 756
box -48 -56 538 834
use sg13g2_a21o_1  _1329_
timestamp 1677175127
transform 1 0 68064 0 -1 2268
box -48 -56 720 834
use sg13g2_a21oi_1  _1330_
timestamp 1683973020
transform -1 0 67008 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1331_
timestamp 1685173987
transform -1 0 68064 0 -1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1332_
timestamp 1685175443
transform -1 0 69792 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1333_
timestamp 1677175127
transform 1 0 68544 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1334_
timestamp 1683973020
transform 1 0 68544 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1335_
timestamp 1685173987
transform 1 0 68256 0 1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _1336_
timestamp 1685175443
transform -1 0 69408 0 1 9828
box -48 -56 538 834
use sg13g2_a21o_1  _1337_
timestamp 1677175127
transform 1 0 68448 0 1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1338_
timestamp 1683973020
transform 1 0 68064 0 1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _1339_
timestamp 1685173987
transform 1 0 67872 0 -1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1340_
timestamp 1685175443
transform -1 0 68256 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1341_
timestamp 1677175127
transform 1 0 67296 0 -1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1342_
timestamp 1683973020
transform 1 0 67392 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1343_
timestamp 1685173987
transform -1 0 67488 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1344_
timestamp 1685175443
transform -1 0 66336 0 1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1345_
timestamp 1677175127
transform 1 0 65184 0 1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1346_
timestamp 1683973020
transform 1 0 65856 0 1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1347_
timestamp 1685173987
transform 1 0 65280 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1348_
timestamp 1685175443
transform -1 0 68352 0 -1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1349_
timestamp 1677175127
transform 1 0 67104 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1350_
timestamp 1683973020
transform 1 0 67200 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1351_
timestamp 1685173987
transform -1 0 67200 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1352_
timestamp 1685175443
transform -1 0 71520 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1353_
timestamp 1677175127
transform 1 0 69984 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1354_
timestamp 1683973020
transform -1 0 69216 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1355_
timestamp 1685173987
transform -1 0 70272 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1356_
timestamp 1685175443
transform -1 0 73056 0 1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1357_
timestamp 1677175127
transform 1 0 71616 0 1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1358_
timestamp 1683973020
transform -1 0 71616 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1359_
timestamp 1685173987
transform -1 0 71424 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1360_
timestamp 1685175443
transform -1 0 73920 0 1 11340
box -48 -56 538 834
use sg13g2_a21o_1  _1361_
timestamp 1677175127
transform -1 0 72960 0 1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1362_
timestamp 1683973020
transform 1 0 71520 0 1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1363_
timestamp 1685173987
transform -1 0 72192 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1364_
timestamp 1685175443
transform -1 0 74016 0 -1 9828
box -48 -56 538 834
use sg13g2_a21o_1  _1365_
timestamp 1677175127
transform 1 0 72480 0 -1 9828
box -48 -56 720 834
use sg13g2_a21oi_1  _1366_
timestamp 1683973020
transform 1 0 72192 0 1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1367_
timestamp 1685173987
transform -1 0 72480 0 -1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1368_
timestamp 1685175443
transform -1 0 74112 0 1 6804
box -48 -56 538 834
use sg13g2_a21o_1  _1369_
timestamp 1677175127
transform -1 0 72576 0 -1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1370_
timestamp 1683973020
transform 1 0 71424 0 -1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1371_
timestamp 1685173987
transform -1 0 72000 0 -1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  _1372_
timestamp 1685175443
transform -1 0 74688 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1373_
timestamp 1677175127
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1374_
timestamp 1683973020
transform 1 0 72192 0 -1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1375_
timestamp 1685173987
transform -1 0 72768 0 1 5292
box -48 -56 624 834
use sg13g2_o21ai_1  _1376_
timestamp 1685175443
transform -1 0 74400 0 -1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _1377_
timestamp 1677175127
transform -1 0 72672 0 1 3780
box -48 -56 720 834
use sg13g2_a21oi_1  _1378_
timestamp 1683973020
transform 1 0 70944 0 1 3780
box -48 -56 528 834
use sg13g2_a22oi_1  _1379_
timestamp 1685173987
transform -1 0 72000 0 1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _1380_
timestamp 1685175443
transform -1 0 74400 0 -1 2268
box -48 -56 538 834
use sg13g2_a21o_1  _1381_
timestamp 1677175127
transform 1 0 72288 0 1 2268
box -48 -56 720 834
use sg13g2_a21oi_1  _1382_
timestamp 1683973020
transform 1 0 71232 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1383_
timestamp 1685173987
transform -1 0 72288 0 1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1384_
timestamp 1685175443
transform 1 0 76416 0 1 756
box -48 -56 538 834
use sg13g2_a21o_1  _1385_
timestamp 1677175127
transform 1 0 76512 0 1 2268
box -48 -56 720 834
use sg13g2_a21oi_1  _1386_
timestamp 1683973020
transform -1 0 74880 0 -1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1387_
timestamp 1685173987
transform -1 0 75936 0 -1 2268
box -48 -56 624 834
use sg13g2_o21ai_1  _1388_
timestamp 1685175443
transform 1 0 77088 0 -1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1389_
timestamp 1677175127
transform 1 0 76224 0 1 3780
box -48 -56 720 834
use sg13g2_a21oi_1  _1390_
timestamp 1683973020
transform 1 0 77280 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _1391_
timestamp 1685173987
transform 1 0 76896 0 -1 3780
box -48 -56 624 834
use sg13g2_o21ai_1  _1392_
timestamp 1685175443
transform 1 0 77760 0 1 5292
box -48 -56 538 834
use sg13g2_a21o_1  _1393_
timestamp 1677175127
transform 1 0 77088 0 1 5292
box -48 -56 720 834
use sg13g2_a21oi_1  _1394_
timestamp 1683973020
transform 1 0 77568 0 -1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _1395_
timestamp 1685173987
transform 1 0 76416 0 -1 6804
box -48 -56 624 834
use sg13g2_o21ai_1  _1396_
timestamp 1685175443
transform -1 0 77952 0 1 9828
box -48 -56 538 834
use sg13g2_a21o_1  _1397_
timestamp 1677175127
transform 1 0 76896 0 -1 8316
box -48 -56 720 834
use sg13g2_a21oi_1  _1398_
timestamp 1683973020
transform 1 0 78144 0 1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _1399_
timestamp 1685173987
transform -1 0 76800 0 1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _1400_
timestamp 1685175443
transform -1 0 78048 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1401_
timestamp 1677175127
transform 1 0 77184 0 -1 11340
box -48 -56 720 834
use sg13g2_a21oi_1  _1402_
timestamp 1683973020
transform 1 0 77856 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1403_
timestamp 1685173987
transform -1 0 77472 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1404_
timestamp 1685175443
transform -1 0 77952 0 1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1405_
timestamp 1677175127
transform 1 0 76704 0 1 12852
box -48 -56 720 834
use sg13g2_a21oi_1  _1406_
timestamp 1683973020
transform 1 0 76416 0 1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1407_
timestamp 1685173987
transform -1 0 76896 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1408_
timestamp 1685175443
transform -1 0 77088 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1409_
timestamp 1677175127
transform -1 0 76128 0 -1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1410_
timestamp 1683973020
transform 1 0 75648 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1411_
timestamp 1685173987
transform -1 0 75744 0 1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1412_
timestamp 1685175443
transform 1 0 76512 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1413_
timestamp 1677175127
transform -1 0 76032 0 -1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1414_
timestamp 1683973020
transform 1 0 74784 0 1 23436
box -48 -56 528 834
use sg13g2_a22oi_1  _1415_
timestamp 1685173987
transform -1 0 75360 0 -1 24948
box -48 -56 624 834
use sg13g2_o21ai_1  _1416_
timestamp 1685175443
transform -1 0 77760 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1417_
timestamp 1677175127
transform 1 0 76128 0 -1 26460
box -48 -56 720 834
use sg13g2_a21oi_1  _1418_
timestamp 1683973020
transform -1 0 76224 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1419_
timestamp 1685173987
transform -1 0 76128 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1420_
timestamp 1685175443
transform -1 0 78048 0 1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1421_
timestamp 1677175127
transform 1 0 76992 0 1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1422_
timestamp 1683973020
transform 1 0 75648 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1423_
timestamp 1685173987
transform -1 0 76704 0 -1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1424_
timestamp 1685175443
transform -1 0 77856 0 -1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1425_
timestamp 1677175127
transform 1 0 76320 0 1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1426_
timestamp 1683973020
transform 1 0 76416 0 -1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1427_
timestamp 1685173987
transform -1 0 76320 0 1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _1428_
timestamp 1685175443
transform -1 0 77952 0 1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1429_
timestamp 1677175127
transform 1 0 76224 0 -1 32508
box -48 -56 720 834
use sg13g2_a21oi_1  _1430_
timestamp 1683973020
transform 1 0 76992 0 1 30996
box -48 -56 528 834
use sg13g2_a22oi_1  _1431_
timestamp 1685173987
transform 1 0 76416 0 1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _1432_
timestamp 1685175443
transform 1 0 78144 0 1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1433_
timestamp 1677175127
transform 1 0 77472 0 1 34020
box -48 -56 720 834
use sg13g2_a21oi_1  _1434_
timestamp 1683973020
transform 1 0 77568 0 -1 34020
box -48 -56 528 834
use sg13g2_a22oi_1  _1435_
timestamp 1685173987
transform 1 0 76992 0 -1 34020
box -48 -56 624 834
use sg13g2_o21ai_1  _1436_
timestamp 1685175443
transform 1 0 76224 0 1 35532
box -48 -56 538 834
use sg13g2_a21o_1  _1437_
timestamp 1677175127
transform -1 0 77376 0 1 35532
box -48 -56 720 834
use sg13g2_a21oi_1  _1438_
timestamp 1683973020
transform 1 0 77376 0 1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _1439_
timestamp 1685173987
transform 1 0 76032 0 -1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1440_
timestamp 1685175443
transform -1 0 74880 0 -1 38556
box -48 -56 538 834
use sg13g2_a21o_1  _1441_
timestamp 1677175127
transform 1 0 73056 0 1 37044
box -48 -56 720 834
use sg13g2_a21oi_1  _1442_
timestamp 1683973020
transform 1 0 73920 0 -1 38556
box -48 -56 528 834
use sg13g2_a22oi_1  _1443_
timestamp 1685173987
transform 1 0 73440 0 -1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1444_
timestamp 1685175443
transform -1 0 74208 0 1 35532
box -48 -56 538 834
use sg13g2_a21o_1  _1445_
timestamp 1677175127
transform -1 0 73056 0 1 35532
box -48 -56 720 834
use sg13g2_a21oi_1  _1446_
timestamp 1683973020
transform 1 0 72672 0 -1 37044
box -48 -56 528 834
use sg13g2_a22oi_1  _1447_
timestamp 1685173987
transform -1 0 72672 0 -1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1448_
timestamp 1685175443
transform -1 0 72192 0 -1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1449_
timestamp 1677175127
transform -1 0 71808 0 1 34020
box -48 -56 720 834
use sg13g2_a21oi_1  _1450_
timestamp 1683973020
transform -1 0 71712 0 1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _1451_
timestamp 1685173987
transform -1 0 72192 0 -1 35532
box -48 -56 624 834
use sg13g2_o21ai_1  _1452_
timestamp 1685175443
transform -1 0 74016 0 1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1453_
timestamp 1677175127
transform -1 0 72960 0 1 32508
box -48 -56 720 834
use sg13g2_a21oi_1  _1454_
timestamp 1683973020
transform -1 0 71712 0 -1 34020
box -48 -56 528 834
use sg13g2_a22oi_1  _1455_
timestamp 1685173987
transform -1 0 72000 0 -1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1456_
timestamp 1685175443
transform -1 0 73536 0 1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1457_
timestamp 1677175127
transform -1 0 72576 0 1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1458_
timestamp 1683973020
transform 1 0 72000 0 -1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _1459_
timestamp 1685173987
transform 1 0 71808 0 -1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _1460_
timestamp 1685175443
transform -1 0 73152 0 1 27972
box -48 -56 538 834
use sg13g2_a21o_1  _1461_
timestamp 1677175127
transform -1 0 71904 0 -1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1462_
timestamp 1683973020
transform 1 0 71040 0 1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1463_
timestamp 1685173987
transform 1 0 70848 0 1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1464_
timestamp 1685175443
transform -1 0 73056 0 -1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1465_
timestamp 1677175127
transform -1 0 72096 0 -1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1466_
timestamp 1683973020
transform -1 0 70848 0 1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1467_
timestamp 1685173987
transform -1 0 71328 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1468_
timestamp 1685175443
transform -1 0 72384 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1469_
timestamp 1677175127
transform -1 0 71616 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1470_
timestamp 1683973020
transform -1 0 71808 0 1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1471_
timestamp 1685173987
transform -1 0 71040 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1472_
timestamp 1685175443
transform -1 0 70368 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1473_
timestamp 1677175127
transform 1 0 68928 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1474_
timestamp 1683973020
transform 1 0 69408 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1475_
timestamp 1685173987
transform 1 0 68736 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1476_
timestamp 1685175443
transform -1 0 67392 0 -1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1477_
timestamp 1677175127
transform 1 0 66240 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1478_
timestamp 1683973020
transform 1 0 67104 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1479_
timestamp 1685173987
transform -1 0 66240 0 1 24948
box -48 -56 624 834
use sg13g2_o21ai_1  _1480_
timestamp 1685175443
transform -1 0 64608 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1481_
timestamp 1677175127
transform 1 0 63648 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1482_
timestamp 1683973020
transform 1 0 64512 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1483_
timestamp 1685173987
transform 1 0 63648 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1484_
timestamp 1685175443
transform 1 0 65760 0 -1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1485_
timestamp 1677175127
transform 1 0 64992 0 -1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1486_
timestamp 1683973020
transform 1 0 64320 0 1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1487_
timestamp 1685173987
transform -1 0 64992 0 -1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _1488_
timestamp 1685175443
transform -1 0 67008 0 -1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1489_
timestamp 1677175127
transform 1 0 65856 0 1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1490_
timestamp 1683973020
transform -1 0 65184 0 1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1491_
timestamp 1685173987
transform -1 0 65760 0 1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _1492_
timestamp 1685175443
transform 1 0 68064 0 -1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1493_
timestamp 1677175127
transform 1 0 67104 0 -1 32508
box -48 -56 720 834
use sg13g2_a21oi_1  _1494_
timestamp 1683973020
transform 1 0 66144 0 1 30996
box -48 -56 528 834
use sg13g2_a22oi_1  _1495_
timestamp 1685173987
transform -1 0 66912 0 -1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1496_
timestamp 1685175443
transform -1 0 69024 0 1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1497_
timestamp 1677175127
transform 1 0 67584 0 1 34020
box -48 -56 720 834
use sg13g2_a21oi_1  _1498_
timestamp 1683973020
transform 1 0 67200 0 -1 34020
box -48 -56 528 834
use sg13g2_a22oi_1  _1499_
timestamp 1685173987
transform -1 0 67584 0 1 34020
box -48 -56 624 834
use sg13g2_o21ai_1  _1500_
timestamp 1685175443
transform -1 0 69216 0 -1 37044
box -48 -56 538 834
use sg13g2_a21o_1  _1501_
timestamp 1677175127
transform -1 0 68256 0 -1 37044
box -48 -56 720 834
use sg13g2_a21oi_1  _1502_
timestamp 1683973020
transform 1 0 68256 0 -1 37044
box -48 -56 528 834
use sg13g2_a22oi_1  _1503_
timestamp 1685173987
transform -1 0 67584 0 -1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1504_
timestamp 1685175443
transform -1 0 65664 0 1 35532
box -48 -56 538 834
use sg13g2_a21o_1  _1505_
timestamp 1677175127
transform -1 0 64704 0 1 35532
box -48 -56 720 834
use sg13g2_a21oi_1  _1506_
timestamp 1683973020
transform 1 0 65184 0 -1 38556
box -48 -56 528 834
use sg13g2_a22oi_1  _1507_
timestamp 1685173987
transform 1 0 64032 0 1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1508_
timestamp 1685175443
transform -1 0 61632 0 1 35532
box -48 -56 538 834
use sg13g2_a21o_1  _1509_
timestamp 1677175127
transform -1 0 60768 0 -1 37044
box -48 -56 720 834
use sg13g2_a21oi_1  _1510_
timestamp 1683973020
transform 1 0 61152 0 -1 38556
box -48 -56 528 834
use sg13g2_a22oi_1  _1511_
timestamp 1685173987
transform -1 0 60096 0 -1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1512_
timestamp 1685175443
transform -1 0 57504 0 1 35532
box -48 -56 538 834
use sg13g2_a21o_1  _1513_
timestamp 1677175127
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_a21oi_1  _1514_
timestamp 1683973020
transform 1 0 57600 0 1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _1515_
timestamp 1685173987
transform 1 0 56448 0 1 37044
box -48 -56 624 834
use sg13g2_o21ai_1  _1516_
timestamp 1685175443
transform -1 0 59712 0 -1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1517_
timestamp 1677175127
transform 1 0 58848 0 -1 35532
box -48 -56 720 834
use sg13g2_a21oi_1  _1518_
timestamp 1683973020
transform -1 0 58560 0 1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _1519_
timestamp 1685173987
transform -1 0 58848 0 -1 35532
box -48 -56 624 834
use sg13g2_o21ai_1  _1520_
timestamp 1685175443
transform -1 0 64896 0 -1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1521_
timestamp 1677175127
transform -1 0 64128 0 1 34020
box -48 -56 720 834
use sg13g2_a21oi_1  _1522_
timestamp 1683973020
transform -1 0 61536 0 -1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _1523_
timestamp 1685173987
transform -1 0 62784 0 1 34020
box -48 -56 624 834
use sg13g2_o21ai_1  _1524_
timestamp 1685175443
transform -1 0 64128 0 1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1525_
timestamp 1677175127
transform -1 0 63648 0 1 32508
box -48 -56 720 834
use sg13g2_a21oi_1  _1526_
timestamp 1683973020
transform 1 0 62976 0 1 34020
box -48 -56 528 834
use sg13g2_a22oi_1  _1527_
timestamp 1685173987
transform -1 0 63264 0 -1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1528_
timestamp 1685175443
transform -1 0 61920 0 1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1529_
timestamp 1677175127
transform 1 0 60768 0 1 30996
box -48 -56 720 834
use sg13g2_a21oi_1  _1530_
timestamp 1683973020
transform 1 0 61440 0 -1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _1531_
timestamp 1685173987
transform 1 0 60672 0 -1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1532_
timestamp 1685175443
transform -1 0 58464 0 1 30996
box -48 -56 538 834
use sg13g2_a21o_1  _1533_
timestamp 1677175127
transform -1 0 57984 0 1 30996
box -48 -56 720 834
use sg13g2_a21oi_1  _1534_
timestamp 1683973020
transform 1 0 58560 0 1 30996
box -48 -56 528 834
use sg13g2_a22oi_1  _1535_
timestamp 1685173987
transform 1 0 57120 0 -1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1536_
timestamp 1685175443
transform -1 0 56256 0 1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _1537_
timestamp 1677175127
transform 1 0 54912 0 -1 34020
box -48 -56 720 834
use sg13g2_a21oi_1  _1538_
timestamp 1683973020
transform 1 0 55776 0 1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _1539_
timestamp 1685173987
transform 1 0 55008 0 1 32508
box -48 -56 624 834
use sg13g2_o21ai_1  _1540_
timestamp 1685175443
transform -1 0 53760 0 1 32508
box -48 -56 538 834
use sg13g2_a21o_1  _1541_
timestamp 1677175127
transform 1 0 50880 0 1 32508
box -48 -56 720 834
use sg13g2_a21oi_1  _1542_
timestamp 1683973020
transform 1 0 53760 0 1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _1543_
timestamp 1685173987
transform 1 0 51840 0 1 34020
box -48 -56 624 834
use sg13g2_o21ai_1  _1544_
timestamp 1685175443
transform -1 0 51840 0 1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1545_
timestamp 1677175127
transform 1 0 50880 0 1 30996
box -48 -56 720 834
use sg13g2_a21oi_1  _1546_
timestamp 1683973020
transform -1 0 50880 0 1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _1547_
timestamp 1685173987
transform 1 0 50304 0 1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _1548_
timestamp 1685175443
transform -1 0 55008 0 1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1549_
timestamp 1677175127
transform 1 0 53856 0 1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1550_
timestamp 1683973020
transform 1 0 51744 0 1 30996
box -48 -56 528 834
use sg13g2_a22oi_1  _1551_
timestamp 1685173987
transform -1 0 52800 0 1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _1552_
timestamp 1685175443
transform -1 0 57888 0 -1 27972
box -48 -56 538 834
use sg13g2_a21o_1  _1553_
timestamp 1677175127
transform 1 0 56928 0 -1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1554_
timestamp 1683973020
transform -1 0 56448 0 1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1555_
timestamp 1685173987
transform -1 0 56928 0 -1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _1556_
timestamp 1685175443
transform -1 0 62400 0 1 27972
box -48 -56 538 834
use sg13g2_a21o_1  _1557_
timestamp 1677175127
transform -1 0 61440 0 1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1558_
timestamp 1683973020
transform -1 0 59232 0 -1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1559_
timestamp 1685173987
transform -1 0 60288 0 1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1560_
timestamp 1685175443
transform -1 0 62112 0 -1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1561_
timestamp 1677175127
transform 1 0 60864 0 -1 26460
box -48 -56 720 834
use sg13g2_a21oi_1  _1562_
timestamp 1683973020
transform 1 0 61152 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1563_
timestamp 1685173987
transform -1 0 61152 0 -1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1564_
timestamp 1685175443
transform -1 0 60192 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1565_
timestamp 1677175127
transform 1 0 59040 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1566_
timestamp 1683973020
transform 1 0 59904 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1567_
timestamp 1685173987
transform 1 0 59232 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1568_
timestamp 1685175443
transform -1 0 57504 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1569_
timestamp 1677175127
transform -1 0 57120 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1570_
timestamp 1683973020
transform 1 0 57408 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1571_
timestamp 1685173987
transform 1 0 56064 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1572_
timestamp 1685175443
transform 1 0 54240 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1573_
timestamp 1677175127
transform -1 0 54240 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1574_
timestamp 1683973020
transform 1 0 54720 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1575_
timestamp 1685173987
transform 1 0 53568 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1576_
timestamp 1685175443
transform -1 0 53856 0 1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1577_
timestamp 1677175127
transform -1 0 52896 0 1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1578_
timestamp 1683973020
transform 1 0 52512 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1579_
timestamp 1685173987
transform -1 0 52512 0 -1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1580_
timestamp 1685175443
transform -1 0 49056 0 -1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1581_
timestamp 1677175127
transform -1 0 48576 0 -1 29484
box -48 -56 720 834
use sg13g2_a21oi_1  _1582_
timestamp 1683973020
transform 1 0 50880 0 -1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1583_
timestamp 1685173987
transform -1 0 48576 0 -1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _1584_
timestamp 1685175443
transform -1 0 48576 0 1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1585_
timestamp 1677175127
transform -1 0 48192 0 -1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1586_
timestamp 1683973020
transform 1 0 46560 0 -1 29484
box -48 -56 528 834
use sg13g2_a22oi_1  _1587_
timestamp 1685173987
transform -1 0 47616 0 -1 29484
box -48 -56 624 834
use sg13g2_o21ai_1  _1588_
timestamp 1685175443
transform -1 0 48576 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1589_
timestamp 1677175127
transform 1 0 47712 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1590_
timestamp 1683973020
transform 1 0 47040 0 1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1591_
timestamp 1685173987
transform -1 0 48096 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1592_
timestamp 1685175443
transform -1 0 52032 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1593_
timestamp 1677175127
transform -1 0 51456 0 1 23436
box -48 -56 720 834
use sg13g2_a21oi_1  _1594_
timestamp 1683973020
transform -1 0 50496 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1595_
timestamp 1685173987
transform -1 0 50784 0 1 23436
box -48 -56 624 834
use sg13g2_o21ai_1  _1596_
timestamp 1685175443
transform -1 0 50880 0 -1 21924
box -48 -56 538 834
use sg13g2_a21o_1  _1597_
timestamp 1677175127
transform 1 0 49248 0 1 21924
box -48 -56 720 834
use sg13g2_a21oi_1  _1598_
timestamp 1683973020
transform -1 0 50208 0 1 23436
box -48 -56 528 834
use sg13g2_a22oi_1  _1599_
timestamp 1685173987
transform 1 0 49632 0 -1 23436
box -48 -56 624 834
use sg13g2_o21ai_1  _1600_
timestamp 1685175443
transform -1 0 47136 0 -1 21924
box -48 -56 538 834
use sg13g2_a21o_1  _1601_
timestamp 1677175127
transform 1 0 46368 0 1 21924
box -48 -56 720 834
use sg13g2_a21oi_1  _1602_
timestamp 1683973020
transform 1 0 47328 0 1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1603_
timestamp 1685173987
transform 1 0 46080 0 -1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1604_
timestamp 1685175443
transform -1 0 43008 0 -1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1605_
timestamp 1677175127
transform 1 0 41952 0 1 21924
box -48 -56 720 834
use sg13g2_a21oi_1  _1606_
timestamp 1683973020
transform 1 0 42816 0 1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1607_
timestamp 1685173987
transform -1 0 41952 0 1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1608_
timestamp 1685175443
transform -1 0 44544 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1609_
timestamp 1677175127
transform -1 0 43968 0 1 23436
box -48 -56 720 834
use sg13g2_a21oi_1  _1610_
timestamp 1683973020
transform 1 0 40800 0 1 23436
box -48 -56 528 834
use sg13g2_a22oi_1  _1611_
timestamp 1685173987
transform -1 0 43104 0 1 23436
box -48 -56 624 834
use sg13g2_o21ai_1  _1612_
timestamp 1685175443
transform 1 0 44832 0 1 24948
box -48 -56 538 834
use sg13g2_a21o_1  _1613_
timestamp 1677175127
transform -1 0 44736 0 -1 26460
box -48 -56 720 834
use sg13g2_a21oi_1  _1614_
timestamp 1683973020
transform 1 0 42912 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1615_
timestamp 1685173987
transform -1 0 43968 0 -1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1616_
timestamp 1685175443
transform -1 0 43008 0 -1 29484
box -48 -56 538 834
use sg13g2_a21o_1  _1617_
timestamp 1677175127
transform -1 0 43104 0 -1 27972
box -48 -56 720 834
use sg13g2_a21oi_1  _1618_
timestamp 1683973020
transform 1 0 43104 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1619_
timestamp 1685173987
transform -1 0 42720 0 1 27972
box -48 -56 624 834
use sg13g2_o21ai_1  _1620_
timestamp 1685175443
transform 1 0 40224 0 1 26460
box -48 -56 538 834
use sg13g2_a21o_1  _1621_
timestamp 1677175127
transform 1 0 39648 0 1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1622_
timestamp 1683973020
transform 1 0 40512 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _1623_
timestamp 1685173987
transform 1 0 39648 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1624_
timestamp 1685175443
transform -1 0 39072 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1625_
timestamp 1677175127
transform -1 0 38400 0 -1 24948
box -48 -56 720 834
use sg13g2_a21oi_1  _1626_
timestamp 1683973020
transform 1 0 38304 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1627_
timestamp 1685173987
transform -1 0 38304 0 1 23436
box -48 -56 624 834
use sg13g2_o21ai_1  _1628_
timestamp 1685175443
transform -1 0 37056 0 1 23436
box -48 -56 538 834
use sg13g2_a21o_1  _1629_
timestamp 1677175127
transform 1 0 36288 0 -1 23436
box -48 -56 720 834
use sg13g2_a21oi_1  _1630_
timestamp 1683973020
transform 1 0 36096 0 1 23436
box -48 -56 528 834
use sg13g2_a22oi_1  _1631_
timestamp 1685173987
transform -1 0 36480 0 1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1632_
timestamp 1685175443
transform 1 0 36672 0 1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _1633_
timestamp 1677175127
transform -1 0 36672 0 -1 21924
box -48 -56 720 834
use sg13g2_a21oi_1  _1634_
timestamp 1683973020
transform 1 0 35424 0 1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1635_
timestamp 1685173987
transform -1 0 36000 0 1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1636_
timestamp 1685175443
transform -1 0 31104 0 -1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _1637_
timestamp 1677175127
transform 1 0 31104 0 -1 20412
box -48 -56 720 834
use sg13g2_a21oi_1  _1638_
timestamp 1683973020
transform 1 0 32928 0 1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  _1639_
timestamp 1685173987
transform 1 0 32352 0 1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1640_
timestamp 1685175443
transform -1 0 3840 0 -1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1641_
timestamp 1677175127
transform -1 0 4512 0 -1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1642_
timestamp 1683973020
transform -1 0 4704 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1643_
timestamp 1685173987
transform 1 0 4512 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1644_
timestamp 1685175443
transform 1 0 5952 0 -1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1645_
timestamp 1677175127
transform -1 0 7296 0 1 17388
box -48 -56 720 834
use sg13g2_a21oi_1  _1646_
timestamp 1683973020
transform -1 0 6720 0 1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1647_
timestamp 1685173987
transform -1 0 7008 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1648_
timestamp 1685175443
transform -1 0 11040 0 -1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1649_
timestamp 1677175127
transform -1 0 10464 0 1 17388
box -48 -56 720 834
use sg13g2_a21oi_1  _1650_
timestamp 1683973020
transform -1 0 10176 0 -1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1651_
timestamp 1685173987
transform -1 0 10848 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1652_
timestamp 1685175443
transform 1 0 12384 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1653_
timestamp 1677175127
transform -1 0 13536 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1654_
timestamp 1683973020
transform 1 0 13056 0 1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1655_
timestamp 1685173987
transform -1 0 12576 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1656_
timestamp 1685175443
transform 1 0 9696 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1657_
timestamp 1677175127
transform -1 0 10848 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1658_
timestamp 1683973020
transform 1 0 10848 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1659_
timestamp 1685173987
transform 1 0 9984 0 1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1660_
timestamp 1685175443
transform -1 0 8736 0 -1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _1661_
timestamp 1677175127
transform -1 0 7200 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1662_
timestamp 1683973020
transform 1 0 7200 0 1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1663_
timestamp 1685173987
transform 1 0 6528 0 1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1664_
timestamp 1685175443
transform 1 0 3072 0 1 20412
box -48 -56 538 834
use sg13g2_a21o_1  _1665_
timestamp 1677175127
transform -1 0 3936 0 -1 20412
box -48 -56 720 834
use sg13g2_a21oi_1  _1666_
timestamp 1683973020
transform 1 0 3936 0 -1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  _1667_
timestamp 1685173987
transform 1 0 3168 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1668_
timestamp 1685175443
transform 1 0 41376 0 -1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1669_
timestamp 1685175443
transform -1 0 46560 0 1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1670_
timestamp 1685175443
transform -1 0 50688 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1671_
timestamp 1685175443
transform -1 0 50976 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1672_
timestamp 1685175443
transform 1 0 46080 0 -1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1673_
timestamp 1685175443
transform -1 0 44928 0 1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1674_
timestamp 1685175443
transform 1 0 39456 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1675_
timestamp 1685175443
transform 1 0 36384 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1676_
timestamp 1685175443
transform -1 0 34560 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1677_
timestamp 1685175443
transform -1 0 33024 0 1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1678_
timestamp 1685175443
transform -1 0 35904 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1679_
timestamp 1685175443
transform -1 0 38016 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1680_
timestamp 1685175443
transform 1 0 39456 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1681_
timestamp 1685175443
transform -1 0 42816 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1682_
timestamp 1685175443
transform -1 0 45792 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1683_
timestamp 1685175443
transform -1 0 47040 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1684_
timestamp 1685175443
transform -1 0 42912 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1685_
timestamp 1685175443
transform 1 0 44832 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1686_
timestamp 1685175443
transform -1 0 48480 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1687_
timestamp 1685175443
transform -1 0 51840 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1688_
timestamp 1685175443
transform -1 0 51264 0 -1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1689_
timestamp 1685175443
transform 1 0 48960 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1690_
timestamp 1685175443
transform -1 0 52704 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1691_
timestamp 1685175443
transform -1 0 55488 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1692_
timestamp 1685175443
transform -1 0 56640 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1693_
timestamp 1685175443
transform -1 0 56160 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1694_
timestamp 1685175443
transform -1 0 55776 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1695_
timestamp 1685175443
transform 1 0 51648 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1696_
timestamp 1685175443
transform -1 0 55488 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1697_
timestamp 1685175443
transform 1 0 56832 0 -1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _1698_
timestamp 1685175443
transform -1 0 60576 0 1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _1699_
timestamp 1685175443
transform -1 0 62784 0 1 2268
box -48 -56 538 834
use sg13g2_o21ai_1  _1700_
timestamp 1685175443
transform 1 0 60576 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1701_
timestamp 1685175443
transform -1 0 60480 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1702_
timestamp 1685175443
transform -1 0 59328 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1703_
timestamp 1685175443
transform 1 0 57984 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1704_
timestamp 1685175443
transform -1 0 61344 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1705_
timestamp 1685175443
transform 1 0 62304 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1706_
timestamp 1685175443
transform -1 0 63360 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1707_
timestamp 1685175443
transform -1 0 63936 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1708_
timestamp 1685175443
transform -1 0 66144 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1709_
timestamp 1685175443
transform -1 0 65472 0 1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _1710_
timestamp 1685175443
transform -1 0 66336 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _1711_
timestamp 1685175443
transform -1 0 68544 0 1 2268
box -48 -56 538 834
use sg13g2_o21ai_1  _1712_
timestamp 1685175443
transform -1 0 68352 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1713_
timestamp 1685175443
transform 1 0 68160 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1714_
timestamp 1685175443
transform 1 0 67104 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1715_
timestamp 1685175443
transform -1 0 65856 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1716_
timestamp 1685175443
transform -1 0 67296 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1717_
timestamp 1685175443
transform -1 0 70272 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1718_
timestamp 1685175443
transform -1 0 72192 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1719_
timestamp 1685175443
transform -1 0 73440 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1720_
timestamp 1685175443
transform -1 0 73152 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1721_
timestamp 1685175443
transform -1 0 72768 0 1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1722_
timestamp 1685175443
transform -1 0 73152 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1723_
timestamp 1685175443
transform 1 0 72384 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _1724_
timestamp 1685175443
transform 1 0 71424 0 1 756
box -48 -56 538 834
use sg13g2_o21ai_1  _1725_
timestamp 1685175443
transform 1 0 76032 0 1 2268
box -48 -56 538 834
use sg13g2_o21ai_1  _1726_
timestamp 1685175443
transform -1 0 76224 0 1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _1727_
timestamp 1685175443
transform -1 0 76896 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1728_
timestamp 1685175443
transform -1 0 76896 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1729_
timestamp 1685175443
transform -1 0 77568 0 -1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1730_
timestamp 1685175443
transform 1 0 76416 0 -1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1731_
timestamp 1685175443
transform -1 0 76320 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1732_
timestamp 1685175443
transform -1 0 76512 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1733_
timestamp 1685175443
transform -1 0 77184 0 1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _1734_
timestamp 1685175443
transform -1 0 77568 0 1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _1735_
timestamp 1685175443
transform -1 0 77376 0 -1 29484
box -48 -56 538 834
use sg13g2_o21ai_1  _1736_
timestamp 1685175443
transform 1 0 75936 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1737_
timestamp 1685175443
transform 1 0 76512 0 -1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _1738_
timestamp 1685175443
transform 1 0 75552 0 -1 37044
box -48 -56 538 834
use sg13g2_o21ai_1  _1739_
timestamp 1685175443
transform -1 0 74496 0 -1 37044
box -48 -56 538 834
use sg13g2_o21ai_1  _1740_
timestamp 1685175443
transform -1 0 73248 0 -1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _1741_
timestamp 1685175443
transform -1 0 72288 0 1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _1742_
timestamp 1685175443
transform -1 0 73152 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1743_
timestamp 1685175443
transform -1 0 72672 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1744_
timestamp 1685175443
transform -1 0 72192 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1745_
timestamp 1685175443
transform -1 0 72192 0 -1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _1746_
timestamp 1685175443
transform -1 0 71616 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1747_
timestamp 1685175443
transform -1 0 69504 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1748_
timestamp 1685175443
transform 1 0 65856 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1749_
timestamp 1685175443
transform 1 0 62784 0 -1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _1750_
timestamp 1685175443
transform 1 0 65664 0 -1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1751_
timestamp 1685175443
transform -1 0 66720 0 -1 29484
box -48 -56 538 834
use sg13g2_o21ai_1  _1752_
timestamp 1685175443
transform -1 0 67488 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1753_
timestamp 1685175443
transform 1 0 66720 0 -1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _1754_
timestamp 1685175443
transform 1 0 69888 0 -1 38556
box -48 -56 538 834
use sg13g2_o21ai_1  _1755_
timestamp 1685175443
transform -1 0 65184 0 1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _1756_
timestamp 1685175443
transform -1 0 61248 0 -1 37044
box -48 -56 538 834
use sg13g2_o21ai_1  _1757_
timestamp 1685175443
transform -1 0 56352 0 1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _1758_
timestamp 1685175443
transform -1 0 58848 0 1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _1759_
timestamp 1685175443
transform -1 0 64416 0 -1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _1760_
timestamp 1685175443
transform -1 0 63648 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1761_
timestamp 1685175443
transform -1 0 61248 0 -1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1762_
timestamp 1685175443
transform 1 0 57312 0 -1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1763_
timestamp 1685175443
transform -1 0 55008 0 1 32508
box -48 -56 538 834
use sg13g2_o21ai_1  _1764_
timestamp 1685175443
transform -1 0 53280 0 1 32508
box -48 -56 538 834
use sg13g2_o21ai_1  _1765_
timestamp 1685175443
transform -1 0 50592 0 -1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _1766_
timestamp 1685175443
transform 1 0 53088 0 -1 29484
box -48 -56 538 834
use sg13g2_o21ai_1  _1767_
timestamp 1685175443
transform 1 0 56064 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1768_
timestamp 1685175443
transform -1 0 61920 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1769_
timestamp 1685175443
transform -1 0 61344 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1770_
timestamp 1685175443
transform -1 0 59712 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1771_
timestamp 1685175443
transform -1 0 57024 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1772_
timestamp 1685175443
transform -1 0 54240 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1773_
timestamp 1685175443
transform -1 0 53376 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1774_
timestamp 1685175443
transform -1 0 48576 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1775_
timestamp 1685175443
transform 1 0 48192 0 -1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _1776_
timestamp 1685175443
transform -1 0 47712 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1777_
timestamp 1685175443
transform -1 0 51936 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1778_
timestamp 1685175443
transform -1 0 50400 0 -1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1779_
timestamp 1685175443
transform 1 0 45888 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1780_
timestamp 1685175443
transform -1 0 42528 0 -1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1781_
timestamp 1685175443
transform -1 0 44256 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1782_
timestamp 1685175443
transform -1 0 44832 0 1 24948
box -48 -56 538 834
use sg13g2_o21ai_1  _1783_
timestamp 1685175443
transform -1 0 43488 0 -1 29484
box -48 -56 538 834
use sg13g2_o21ai_1  _1784_
timestamp 1685175443
transform 1 0 39456 0 -1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _1785_
timestamp 1685175443
transform -1 0 39552 0 1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1786_
timestamp 1685175443
transform 1 0 36864 0 1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1787_
timestamp 1685175443
transform 1 0 36864 0 -1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1788_
timestamp 1685175443
transform -1 0 31872 0 1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1789_
timestamp 1685175443
transform 1 0 4416 0 -1 21924
box -48 -56 538 834
use sg13g2_o21ai_1  _1790_
timestamp 1685175443
transform -1 0 7680 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1791_
timestamp 1685175443
transform 1 0 15168 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1792_
timestamp 1685175443
transform -1 0 13824 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1793_
timestamp 1685175443
transform 1 0 10752 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1794_
timestamp 1685175443
transform -1 0 8256 0 -1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1795_
timestamp 1685175443
transform -1 0 4128 0 -1 21924
box -48 -56 538 834
use sg13g2_dfrbpq_1  _1796_
timestamp 1746535128
transform 1 0 40128 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1797_
timestamp 1746535128
transform 1 0 45312 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1798_
timestamp 1746535128
transform 1 0 48288 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1799_
timestamp 1746535128
transform -1 0 50208 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1800_
timestamp 1746535128
transform 1 0 43008 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1801_
timestamp 1746535128
transform -1 0 43008 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1802_
timestamp 1746535128
transform -1 0 39936 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1803_
timestamp 1746535128
transform -1 0 37056 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1804_
timestamp 1746535128
transform -1 0 32736 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1805_
timestamp 1746535128
transform 1 0 31584 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1806_
timestamp 1746535128
transform 1 0 34368 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1807_
timestamp 1746535128
transform 1 0 36576 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1808_
timestamp 1746535128
transform 1 0 38688 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1809_
timestamp 1746535128
transform 1 0 41280 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1810_
timestamp 1746535128
transform 1 0 43968 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1811_
timestamp 1746535128
transform -1 0 46368 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1812_
timestamp 1746535128
transform 1 0 42528 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1813_
timestamp 1746535128
transform 1 0 45120 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1814_
timestamp 1746535128
transform 1 0 47808 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1815_
timestamp 1746535128
transform 1 0 49824 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1816_
timestamp 1746535128
transform 1 0 48192 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1817_
timestamp 1746535128
transform 1 0 48576 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1818_
timestamp 1746535128
transform 1 0 51456 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1819_
timestamp 1746535128
transform 1 0 54048 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1820_
timestamp 1746535128
transform -1 0 55872 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1821_
timestamp 1746535128
transform 1 0 53376 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1822_
timestamp 1746535128
transform 1 0 50592 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1823_
timestamp 1746535128
transform 1 0 51648 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1824_
timestamp 1746535128
transform 1 0 53760 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1825_
timestamp 1746535128
transform 1 0 55968 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1826_
timestamp 1746535128
transform 1 0 58272 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1827_
timestamp 1746535128
transform 1 0 59808 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1828_
timestamp 1746535128
transform -1 0 60768 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1829_
timestamp 1746535128
transform 1 0 57024 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1830_
timestamp 1746535128
transform 1 0 57024 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1831_
timestamp 1746535128
transform 1 0 57600 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1832_
timestamp 1746535128
transform 1 0 59904 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1833_
timestamp 1746535128
transform 1 0 60192 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1834_
timestamp 1746535128
transform 1 0 60576 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1835_
timestamp 1746535128
transform 1 0 62112 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1836_
timestamp 1746535128
transform -1 0 66240 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1837_
timestamp 1746535128
transform 1 0 63168 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1838_
timestamp 1746535128
transform 1 0 64896 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1839_
timestamp 1746535128
transform 1 0 66720 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1840_
timestamp 1746535128
transform 1 0 67872 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1841_
timestamp 1746535128
transform -1 0 68448 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1842_
timestamp 1746535128
transform -1 0 67296 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1843_
timestamp 1746535128
transform 1 0 64320 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1844_
timestamp 1746535128
transform 1 0 67104 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1845_
timestamp 1746535128
transform 1 0 68544 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1846_
timestamp 1746535128
transform 1 0 69408 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1847_
timestamp 1746535128
transform 1 0 69888 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1848_
timestamp 1746535128
transform -1 0 72192 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1849_
timestamp 1746535128
transform 1 0 69984 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1850_
timestamp 1746535128
transform 1 0 70464 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1851_
timestamp 1746535128
transform 1 0 69600 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1852_
timestamp 1746535128
transform 1 0 71328 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1853_
timestamp 1746535128
transform 1 0 75936 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1854_
timestamp 1746535128
transform 1 0 76896 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1855_
timestamp 1746535128
transform 1 0 76992 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1856_
timestamp 1746535128
transform 1 0 76800 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1857_
timestamp 1746535128
transform 1 0 74592 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1858_
timestamp 1746535128
transform 1 0 74112 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1859_
timestamp 1746535128
transform -1 0 75456 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1860_
timestamp 1746535128
transform 1 0 73152 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1861_
timestamp 1746535128
transform 1 0 74496 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1862_
timestamp 1746535128
transform 1 0 74400 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1863_
timestamp 1746535128
transform 1 0 74976 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1864_
timestamp 1746535128
transform 1 0 76320 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1865_
timestamp 1746535128
transform 1 0 76992 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1866_
timestamp 1746535128
transform 1 0 76704 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1867_
timestamp 1746535128
transform -1 0 72864 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1868_
timestamp 1746535128
transform -1 0 72096 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1869_
timestamp 1746535128
transform -1 0 71616 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1870_
timestamp 1746535128
transform 1 0 69696 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1871_
timestamp 1746535128
transform -1 0 71808 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1872_
timestamp 1746535128
transform -1 0 70944 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1873_
timestamp 1746535128
transform -1 0 70944 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1874_
timestamp 1746535128
transform -1 0 70560 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1875_
timestamp 1746535128
transform 1 0 66048 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1876_
timestamp 1746535128
transform -1 0 65760 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1877_
timestamp 1746535128
transform 1 0 62304 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1878_
timestamp 1746535128
transform 1 0 62976 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1879_
timestamp 1746535128
transform 1 0 63936 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1880_
timestamp 1746535128
transform 1 0 65376 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1881_
timestamp 1746535128
transform 1 0 66336 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1882_
timestamp 1746535128
transform -1 0 67296 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1883_
timestamp 1746535128
transform -1 0 64224 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1884_
timestamp 1746535128
transform -1 0 60000 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1885_
timestamp 1746535128
transform 1 0 56160 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1886_
timestamp 1746535128
transform 1 0 58560 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1887_
timestamp 1746535128
transform 1 0 61536 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1888_
timestamp 1746535128
transform -1 0 62688 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1889_
timestamp 1746535128
transform -1 0 60288 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1890_
timestamp 1746535128
transform -1 0 57024 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1891_
timestamp 1746535128
transform -1 0 54816 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1892_
timestamp 1746535128
transform -1 0 51840 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1893_
timestamp 1746535128
transform 1 0 50496 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1894_
timestamp 1746535128
transform 1 0 53568 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1895_
timestamp 1746535128
transform 1 0 56544 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1896_
timestamp 1746535128
transform 1 0 59232 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1897_
timestamp 1746535128
transform -1 0 61344 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1898_
timestamp 1746535128
transform -1 0 59232 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1899_
timestamp 1746535128
transform -1 0 56544 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1900_
timestamp 1746535128
transform -1 0 53376 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1901_
timestamp 1746535128
transform -1 0 52224 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1902_
timestamp 1746535128
transform -1 0 47904 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1903_
timestamp 1746535128
transform 1 0 45312 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1904_
timestamp 1746535128
transform 1 0 47712 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1905_
timestamp 1746535128
transform 1 0 48768 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1906_
timestamp 1746535128
transform -1 0 49920 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1907_
timestamp 1746535128
transform -1 0 46368 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1908_
timestamp 1746535128
transform 1 0 39936 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1909_
timestamp 1746535128
transform 1 0 40992 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1910_
timestamp 1746535128
transform 1 0 42048 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1911_
timestamp 1746535128
transform -1 0 42144 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1912_
timestamp 1746535128
transform -1 0 39456 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1913_
timestamp 1746535128
transform -1 0 37728 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1914_
timestamp 1746535128
transform -1 0 36288 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1915_
timestamp 1746535128
transform -1 0 36000 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1916_
timestamp 1746535128
transform -1 0 32352 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1917_
timestamp 1746535128
transform -1 0 6528 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1918_
timestamp 1746535128
transform 1 0 7008 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1919_
timestamp 1746535128
transform 1 0 10464 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1920_
timestamp 1746535128
transform 1 0 12576 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1921_
timestamp 1746535128
transform -1 0 11808 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1922_
timestamp 1746535128
transform -1 0 7776 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1923_
timestamp 1746535128
transform -1 0 3264 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1924_
timestamp 1746535128
transform 1 0 42720 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1925_
timestamp 1746535128
transform 1 0 46272 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1926_
timestamp 1746535128
transform 1 0 50208 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1927_
timestamp 1746535128
transform 1 0 50208 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1928_
timestamp 1746535128
transform 1 0 46464 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1929_
timestamp 1746535128
transform 1 0 43680 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1930_
timestamp 1746535128
transform 1 0 39936 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1931_
timestamp 1746535128
transform 1 0 36864 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1932_
timestamp 1746535128
transform 1 0 33504 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1933_
timestamp 1746535128
transform 1 0 32832 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1934_
timestamp 1746535128
transform 1 0 35520 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1935_
timestamp 1746535128
transform 1 0 38016 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1936_
timestamp 1746535128
transform 1 0 39936 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1937_
timestamp 1746535128
transform 1 0 42528 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1938_
timestamp 1746535128
transform 1 0 45792 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1939_
timestamp 1746535128
transform 1 0 46752 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1940_
timestamp 1746535128
transform 1 0 41184 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1941_
timestamp 1746535128
transform 1 0 45312 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1942_
timestamp 1746535128
transform 1 0 47904 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1943_
timestamp 1746535128
transform 1 0 51648 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1944_
timestamp 1746535128
transform 1 0 51264 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1945_
timestamp 1746535128
transform 1 0 48672 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1946_
timestamp 1746535128
transform 1 0 52416 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1947_
timestamp 1746535128
transform 1 0 55296 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1948_
timestamp 1746535128
transform 1 0 56640 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1949_
timestamp 1746535128
transform 1 0 56160 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1950_
timestamp 1746535128
transform 1 0 55584 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1951_
timestamp 1746535128
transform 1 0 52128 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1952_
timestamp 1746535128
transform 1 0 55488 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1953_
timestamp 1746535128
transform 1 0 57312 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1954_
timestamp 1746535128
transform 1 0 60576 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1955_
timestamp 1746535128
transform 1 0 62304 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1956_
timestamp 1746535128
transform 1 0 61056 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1957_
timestamp 1746535128
transform 1 0 59712 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1958_
timestamp 1746535128
transform 1 0 58848 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1959_
timestamp 1746535128
transform 1 0 57888 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1960_
timestamp 1746535128
transform 1 0 61056 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1961_
timestamp 1746535128
transform 1 0 62784 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1962_
timestamp 1746535128
transform 1 0 62688 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1963_
timestamp 1746535128
transform 1 0 63936 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1964_
timestamp 1746535128
transform 1 0 66048 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1965_
timestamp 1746535128
transform 1 0 65280 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1966_
timestamp 1746535128
transform 1 0 66336 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1967_
timestamp 1746535128
transform 1 0 68736 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1968_
timestamp 1746535128
transform 1 0 68352 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1969_
timestamp 1746535128
transform 1 0 68160 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1970_
timestamp 1746535128
transform 1 0 67584 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1971_
timestamp 1746535128
transform 1 0 64512 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1972_
timestamp 1746535128
transform 1 0 66816 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1973_
timestamp 1746535128
transform 1 0 70272 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1974_
timestamp 1746535128
transform 1 0 71808 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1975_
timestamp 1746535128
transform 1 0 72576 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1976_
timestamp 1746535128
transform 1 0 72768 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1977_
timestamp 1746535128
transform 1 0 72576 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1978_
timestamp 1746535128
transform 1 0 73152 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1979_
timestamp 1746535128
transform 1 0 72672 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1980_
timestamp 1746535128
transform 1 0 73152 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1981_
timestamp 1746535128
transform 1 0 76896 0 1 756
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1982_
timestamp 1746535128
transform 1 0 74496 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1983_
timestamp 1746535128
transform 1 0 75552 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1984_
timestamp 1746535128
transform 1 0 75264 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1985_
timestamp 1746535128
transform 1 0 76896 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1986_
timestamp 1746535128
transform 1 0 76896 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1987_
timestamp 1746535128
transform 1 0 76320 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1988_
timestamp 1746535128
transform 1 0 76512 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1989_
timestamp 1746535128
transform 1 0 76800 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1990_
timestamp 1746535128
transform 1 0 76992 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1991_
timestamp 1746535128
transform 1 0 76992 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1992_
timestamp 1746535128
transform 1 0 76896 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1993_
timestamp 1746535128
transform -1 0 77472 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1994_
timestamp 1746535128
transform 1 0 76608 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1995_
timestamp 1746535128
transform 1 0 73728 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1996_
timestamp 1746535128
transform 1 0 73248 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1997_
timestamp 1746535128
transform 1 0 72288 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1998_
timestamp 1746535128
transform 1 0 72768 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _1999_
timestamp 1746535128
transform 1 0 72384 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2000_
timestamp 1746535128
transform 1 0 72096 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2001_
timestamp 1746535128
transform 1 0 71904 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2002_
timestamp 1746535128
transform 1 0 71616 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2003_
timestamp 1746535128
transform 1 0 69024 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2004_
timestamp 1746535128
transform 1 0 66336 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2005_
timestamp 1746535128
transform 1 0 63264 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2006_
timestamp 1746535128
transform 1 0 65856 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2007_
timestamp 1746535128
transform 1 0 66624 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2008_
timestamp 1746535128
transform 1 0 67488 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2009_
timestamp 1746535128
transform 1 0 67680 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2010_
timestamp 1746535128
transform -1 0 70272 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2011_
timestamp 1746535128
transform 1 0 64224 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2012_
timestamp 1746535128
transform 1 0 60480 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2013_
timestamp 1746535128
transform 1 0 55008 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2014_
timestamp 1746535128
transform 1 0 58848 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2015_
timestamp 1746535128
transform 1 0 64224 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2016_
timestamp 1746535128
transform 1 0 63264 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2017_
timestamp 1746535128
transform 1 0 61248 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2018_
timestamp 1746535128
transform 1 0 57792 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2019_
timestamp 1746535128
transform 1 0 55584 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2020_
timestamp 1746535128
transform 1 0 52512 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2021_
timestamp 1746535128
transform 1 0 50592 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2022_
timestamp 1746535128
transform 1 0 53568 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2023_
timestamp 1746535128
transform 1 0 56544 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2024_
timestamp 1746535128
transform 1 0 61824 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2025_
timestamp 1746535128
transform 1 0 60864 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2026_
timestamp 1746535128
transform 1 0 59424 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2027_
timestamp 1746535128
transform 1 0 56544 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2028_
timestamp 1746535128
transform 1 0 53952 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2029_
timestamp 1746535128
transform 1 0 53088 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2030_
timestamp 1746535128
transform 1 0 48288 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2031_
timestamp 1746535128
transform 1 0 48672 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2032_
timestamp 1746535128
transform 1 0 46176 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2033_
timestamp 1746535128
transform 1 0 51360 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2034_
timestamp 1746535128
transform 1 0 49920 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2035_
timestamp 1746535128
transform 1 0 46368 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2036_
timestamp 1746535128
transform 1 0 42528 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2037_
timestamp 1746535128
transform 1 0 43584 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2038_
timestamp 1746535128
transform 1 0 44736 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2039_
timestamp 1746535128
transform 1 0 42720 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2040_
timestamp 1746535128
transform 1 0 39936 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2041_
timestamp 1746535128
transform 1 0 38400 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2042_
timestamp 1746535128
transform 1 0 37344 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2043_
timestamp 1746535128
transform 1 0 37344 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2044_
timestamp 1746535128
transform 1 0 30816 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2045_
timestamp 1746535128
transform 1 0 4896 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2046_
timestamp 1746535128
transform 1 0 7680 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2047_
timestamp 1746535128
transform 1 0 15648 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2048_
timestamp 1746535128
transform 1 0 13824 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2049_
timestamp 1746535128
transform 1 0 11136 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2050_
timestamp 1746535128
transform 1 0 7680 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _2051_
timestamp 1746535128
transform 1 0 3936 0 1 20412
box -48 -56 2640 834
use sg13g2_buf_1  _2060_
timestamp 1676381911
transform -1 0 29760 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _2061_
timestamp 1676381911
transform -1 0 1824 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _2062_
timestamp 1676381911
transform -1 0 1824 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _2063_
timestamp 1676381911
transform -1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2064_
timestamp 1676381911
transform -1 0 1824 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _2065_
timestamp 1676381911
transform -1 0 1824 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _2066_
timestamp 1676381911
transform -1 0 1920 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _2067_
timestamp 1676381911
transform -1 0 1824 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2068_
timestamp 1676381911
transform -1 0 1440 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _2069_
timestamp 1676381911
transform -1 0 2784 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _2070_
timestamp 1676381911
transform -1 0 1824 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2071_
timestamp 1676381911
transform -1 0 10656 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _2072_
timestamp 1676381911
transform -1 0 1824 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _2073_
timestamp 1676381911
transform -1 0 1440 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _2074_
timestamp 1676381911
transform -1 0 1824 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _2075_
timestamp 1676381911
transform -1 0 2304 0 1 18900
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 65376 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 63072 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 66240 0 1 15876
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 70368 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 76320 0 1 15876
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 71616 0 1 15876
box -48 -56 336 834
use sg13g2_buf_16  clkbuf_0_clk
timestamp 1676553496
transform -1 0 43968 0 1 18900
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_0__f_clk
timestamp 1676553496
transform -1 0 41472 0 1 14364
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_1__f_clk
timestamp 1676553496
transform 1 0 28992 0 -1 17388
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_2__f_clk
timestamp 1676553496
transform -1 0 55200 0 -1 15876
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_2_3__f_clk
timestamp 1676553496
transform -1 0 55200 0 1 30996
box -48 -56 2448 834
use sg13g2_buf_8  clkbuf_leaf_0_clk
timestamp 1676451365
transform 1 0 27456 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_1_clk
timestamp 1676451365
transform -1 0 8640 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_2_clk
timestamp 1676451365
transform 1 0 41280 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_3_clk
timestamp 1676451365
transform -1 0 50880 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_4_clk
timestamp 1676451365
transform -1 0 52800 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_5_clk
timestamp 1676451365
transform -1 0 67200 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_6_clk
timestamp 1676451365
transform 1 0 75744 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_7_clk
timestamp 1676451365
transform -1 0 69888 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_8_clk
timestamp 1676451365
transform -1 0 68640 0 -1 38556
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_9_clk
timestamp 1676451365
transform 1 0 48768 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_10_clk
timestamp 1676451365
transform 1 0 51552 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_11_clk
timestamp 1676451365
transform -1 0 73152 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_12_clk
timestamp 1676451365
transform -1 0 71424 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_13_clk
timestamp 1676451365
transform 1 0 72960 0 1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_14_clk
timestamp 1676451365
transform 1 0 61056 0 -1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_15_clk
timestamp 1676451365
transform 1 0 51840 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_16_clk
timestamp 1676451365
transform 1 0 45408 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_leaf_17_clk
timestamp 1676451365
transform -1 0 28512 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkload0
timestamp 1676451365
transform -1 0 30240 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkload1
timestamp 1676451365
transform 1 0 53088 0 -1 32508
box -48 -56 1296 834
use sg13g2_inv_4  clkload2
timestamp 1676383058
transform 1 0 48768 0 1 20412
box -48 -56 624 834
use sg13g2_inv_2  clkload3
timestamp 1676382947
transform 1 0 51264 0 1 14364
box -48 -56 432 834
use sg13g2_inv_2  clkload4
timestamp 1676382947
transform 1 0 53088 0 1 8316
box -48 -56 432 834
use sg13g2_buf_8  clkload5
timestamp 1676451365
transform 1 0 45408 0 -1 15876
box -48 -56 1296 834
use sg13g2_inv_4  clkload6
timestamp 1676383058
transform 1 0 26880 0 -1 20412
box -48 -56 624 834
use sg13g2_inv_8  clkload7
timestamp 1676383150
transform -1 0 8352 0 1 21924
box -48 -56 1008 834
use sg13g2_inv_8  clkload8
timestamp 1676383150
transform 1 0 27264 0 -1 15876
box -48 -56 1008 834
use sg13g2_inv_2  clkload9
timestamp 1676382947
transform -1 0 64800 0 -1 38556
box -48 -56 432 834
use sg13g2_inv_1  clkload10
timestamp 1676382929
transform -1 0 70176 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  clkload11
timestamp 1676382929
transform 1 0 59520 0 1 756
box -48 -56 336 834
use sg13g2_inv_1  clkload12
timestamp 1676382929
transform -1 0 75744 0 -1 38556
box -48 -56 336 834
use dac128module  dac
timestamp 0
transform 1 0 53240 0 1 17400
box 0 0 1 1
use sg13g2_inv_1  digitalen.g\[0\].u.inv1
timestamp 1676382929
transform -1 0 52800 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[0\].u.inv2
timestamp 1676382929
transform -1 0 52512 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv1
timestamp 1676382929
transform 1 0 78432 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[1\].u.inv2
timestamp 1676382929
transform 1 0 79296 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv1
timestamp 1676382929
transform 1 0 78912 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[2\].u.inv2
timestamp 1676382929
transform -1 0 78912 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv1
timestamp 1676382929
transform 1 0 52512 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  digitalen.g\[3\].u.inv2
timestamp 1676382929
transform -1 0 52800 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform -1 0 5472 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform -1 0 4800 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 34080 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform 1 0 37344 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 31872 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform -1 0 32352 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform 1 0 3552 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout30
timestamp 1676381911
transform 1 0 43008 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 45696 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 40992 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform -1 0 56352 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform 1 0 50208 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 48480 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform -1 0 49248 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform 1 0 40416 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 42432 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 42048 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform -1 0 50592 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform 1 0 56160 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform -1 0 51744 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 50496 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform -1 0 42912 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform 1 0 58560 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform -1 0 65088 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout47
timestamp 1676381911
transform -1 0 59328 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform 1 0 59904 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 60480 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout50
timestamp 1676381911
transform -1 0 69024 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform 1 0 69024 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout52
timestamp 1676381911
transform 1 0 77568 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform -1 0 69504 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 68352 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform 1 0 69216 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform 1 0 59520 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform -1 0 59520 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform 1 0 65184 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout59
timestamp 1676381911
transform -1 0 59904 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout60
timestamp 1676381911
transform 1 0 59136 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout61
timestamp 1676381911
transform -1 0 70272 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout62
timestamp 1676381911
transform 1 0 75168 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout63
timestamp 1676381911
transform 1 0 71520 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout64
timestamp 1676381911
transform 1 0 75360 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout65
timestamp 1676381911
transform 1 0 70656 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout66
timestamp 1676381911
transform 1 0 58368 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout67
timestamp 1676381911
transform 1 0 41664 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout68
timestamp 1676381911
transform 1 0 31680 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform 1 0 33216 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 6912 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform -1 0 44736 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform 1 0 49632 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform 1 0 50016 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform 1 0 44448 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform -1 0 43968 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform -1 0 52128 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform 1 0 50592 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform -1 0 45600 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 61344 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform -1 0 62112 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform -1 0 69216 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform 1 0 77568 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 69312 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform 1 0 61728 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 61728 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 71328 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 69984 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform 1 0 61728 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform 1 0 7296 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform -1 0 4224 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform 1 0 2688 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout92
timestamp 1676381911
transform 1 0 32352 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout93
timestamp 1676381911
transform -1 0 33696 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout94
timestamp 1676381911
transform -1 0 31392 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout95
timestamp 1676381911
transform 1 0 30048 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout96
timestamp 1676381911
transform 1 0 38592 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout97
timestamp 1676381911
transform -1 0 46944 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout98
timestamp 1676381911
transform -1 0 40128 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout99
timestamp 1676381911
transform 1 0 52320 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform -1 0 56352 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout101
timestamp 1676381911
transform -1 0 50496 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout102
timestamp 1676381911
transform 1 0 50880 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout103
timestamp 1676381911
transform 1 0 50496 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform 1 0 43776 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform 1 0 43392 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout106
timestamp 1676381911
transform 1 0 43008 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform -1 0 51648 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout108
timestamp 1676381911
transform 1 0 55008 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform 1 0 49920 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout110
timestamp 1676381911
transform 1 0 52032 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout111
timestamp 1676381911
transform -1 0 45024 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout112
timestamp 1676381911
transform -1 0 60384 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout113
timestamp 1676381911
transform -1 0 59904 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout114
timestamp 1676381911
transform -1 0 66144 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  fanout115
timestamp 1676381911
transform 1 0 61824 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout116
timestamp 1676381911
transform 1 0 62208 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout117
timestamp 1676381911
transform -1 0 73632 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout118
timestamp 1676381911
transform 1 0 73152 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout119
timestamp 1676381911
transform -1 0 69024 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout120
timestamp 1676381911
transform 1 0 69408 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout121
timestamp 1676381911
transform 1 0 75552 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout122
timestamp 1676381911
transform 1 0 70656 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout123
timestamp 1676381911
transform -1 0 60864 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout124
timestamp 1676381911
transform 1 0 60672 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout125
timestamp 1676381911
transform 1 0 63744 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout126
timestamp 1676381911
transform -1 0 62208 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout127
timestamp 1676381911
transform 1 0 60384 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout128
timestamp 1676381911
transform -1 0 69984 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout129
timestamp 1676381911
transform -1 0 78432 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout130
timestamp 1676381911
transform -1 0 72576 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout131
timestamp 1676381911
transform 1 0 73152 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  fanout132
timestamp 1676381911
transform 1 0 74208 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout133
timestamp 1676381911
transform -1 0 72960 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout134
timestamp 1676381911
transform 1 0 59904 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout135
timestamp 1676381911
transform 1 0 44160 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout136
timestamp 1676381911
transform 1 0 3264 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout137
timestamp 1676381911
transform -1 0 1920 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout138
timestamp 1676381911
transform -1 0 2304 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout139
timestamp 1676381911
transform -1 0 33312 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout140
timestamp 1676381911
transform 1 0 30432 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout141
timestamp 1676381911
transform 1 0 1728 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout142
timestamp 1676381911
transform 1 0 38976 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout143
timestamp 1676381911
transform 1 0 45024 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout144
timestamp 1676381911
transform -1 0 40032 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout145
timestamp 1676381911
transform -1 0 40416 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout146
timestamp 1676381911
transform 1 0 50688 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout147
timestamp 1676381911
transform 1 0 49248 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout148
timestamp 1676381911
transform -1 0 50112 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout149
timestamp 1676381911
transform 1 0 51264 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout150
timestamp 1676381911
transform 1 0 40512 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout151
timestamp 1676381911
transform -1 0 39648 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout152
timestamp 1676381911
transform 1 0 40704 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout153
timestamp 1676381911
transform 1 0 51168 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout154
timestamp 1676381911
transform -1 0 51264 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout155
timestamp 1676381911
transform -1 0 55776 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout156
timestamp 1676381911
transform 1 0 51936 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout157
timestamp 1676381911
transform -1 0 40512 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout158
timestamp 1676381911
transform -1 0 60288 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout159
timestamp 1676381911
transform 1 0 63072 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout160
timestamp 1676381911
transform 1 0 59904 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout161
timestamp 1676381911
transform -1 0 59232 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout162
timestamp 1676381911
transform 1 0 64992 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout163
timestamp 1676381911
transform 1 0 69792 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout164
timestamp 1676381911
transform 1 0 73824 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout165
timestamp 1676381911
transform 1 0 73920 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  fanout166
timestamp 1676381911
transform 1 0 69408 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout167
timestamp 1676381911
transform -1 0 70464 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout168
timestamp 1676381911
transform 1 0 75936 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout169
timestamp 1676381911
transform 1 0 59040 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout170
timestamp 1676381911
transform -1 0 60096 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout171
timestamp 1676381911
transform 1 0 61056 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout172
timestamp 1676381911
transform 1 0 66720 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout173
timestamp 1676381911
transform -1 0 61824 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout174
timestamp 1676381911
transform 1 0 60096 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout175
timestamp 1676381911
transform 1 0 68640 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout176
timestamp 1676381911
transform 1 0 76128 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout177
timestamp 1676381911
transform -1 0 68736 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout178
timestamp 1676381911
transform -1 0 73920 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout179
timestamp 1676381911
transform 1 0 74592 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout180
timestamp 1676381911
transform -1 0 69120 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout181
timestamp 1676381911
transform 1 0 58656 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout182
timestamp 1676381911
transform 1 0 2112 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout183
timestamp 1676381911
transform -1 0 6048 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout184
timestamp 1676381911
transform -1 0 1536 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout185
timestamp 1676381911
transform 1 0 30624 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout186
timestamp 1676381911
transform 1 0 30240 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout187
timestamp 1676381911
transform 1 0 29664 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout188
timestamp 1676381911
transform -1 0 47616 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout189
timestamp 1676381911
transform 1 0 40416 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout190
timestamp 1676381911
transform 1 0 40032 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout191
timestamp 1676381911
transform 1 0 49440 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout192
timestamp 1676381911
transform 1 0 56064 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout193
timestamp 1676381911
transform 1 0 51360 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout194
timestamp 1676381911
transform -1 0 56160 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout195
timestamp 1676381911
transform -1 0 52032 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout196
timestamp 1676381911
transform 1 0 40032 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout197
timestamp 1676381911
transform 1 0 45792 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout198
timestamp 1676381911
transform -1 0 40800 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout199
timestamp 1676381911
transform -1 0 49632 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout200
timestamp 1676381911
transform 1 0 54336 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout201
timestamp 1676381911
transform 1 0 57024 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout202
timestamp 1676381911
transform -1 0 50112 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout203
timestamp 1676381911
transform 1 0 39648 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout204
timestamp 1676381911
transform 1 0 61056 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout205
timestamp 1676381911
transform -1 0 64800 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout206
timestamp 1676381911
transform -1 0 61536 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout207
timestamp 1676381911
transform 1 0 61344 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout208
timestamp 1676381911
transform 1 0 60672 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout209
timestamp 1676381911
transform -1 0 78720 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  fanout210
timestamp 1676381911
transform -1 0 73632 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout211
timestamp 1676381911
transform -1 0 69024 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  fanout212
timestamp 1676381911
transform -1 0 70848 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout213
timestamp 1676381911
transform 1 0 73344 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  fanout214
timestamp 1676381911
transform 1 0 70848 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout215
timestamp 1676381911
transform 1 0 58752 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout216
timestamp 1676381911
transform 1 0 59136 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout217
timestamp 1676381911
transform 1 0 64800 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout218
timestamp 1676381911
transform 1 0 58752 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout219
timestamp 1676381911
transform -1 0 69216 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout220
timestamp 1676381911
transform -1 0 71136 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout221
timestamp 1676381911
transform 1 0 77184 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout222
timestamp 1676381911
transform 1 0 74496 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout223
timestamp 1676381911
transform 1 0 67296 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout224
timestamp 1676381911
transform 1 0 70368 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  fanout225
timestamp 1676381911
transform -1 0 60384 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  fanout226
timestamp 1676381911
transform 1 0 40320 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  fanout227
timestamp 1676381911
transform 1 0 1248 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_609
timestamp 1679577901
transform 1 0 59040 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_613
timestamp 1677579658
transform 1 0 59424 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_644
timestamp 1677579658
transform 1 0 62400 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_650
timestamp 1679581782
transform 1 0 62976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_657
timestamp 1679581782
transform 1 0 63648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_664
timestamp 1679581782
transform 1 0 64320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_671
timestamp 1679581782
transform 1 0 64992 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_678
timestamp 1679577901
transform 1 0 65664 0 1 756
box -48 -56 432 834
use sg13g2_decap_4  FILLER_0_685
timestamp 1679577901
transform 1 0 66336 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_716
timestamp 1677579658
transform 1 0 69312 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_783
timestamp 1679581782
transform 1 0 75744 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_822
timestamp 1677579658
transform 1 0 79488 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_595
timestamp 1679577901
transform 1 0 57696 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_599
timestamp 1677580104
transform 1 0 58080 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_628
timestamp 1677580104
transform 1 0 60864 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_774
timestamp 1679577901
transform 1 0 74880 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_778
timestamp 1677579658
transform 1 0 75264 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_819
timestamp 1679577901
transform 1 0 79200 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_578
timestamp 1677580104
transform 1 0 56064 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_586
timestamp 1679581782
transform 1 0 56832 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_593
timestamp 1677580104
transform 1 0 57504 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_595
timestamp 1677579658
transform 1 0 57696 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_599
timestamp 1677580104
transform 1 0 58080 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_601
timestamp 1677579658
transform 1 0 58272 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_634
timestamp 1677580104
transform 1 0 61440 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_651
timestamp 1677579658
transform 1 0 63072 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_662
timestamp 1677580104
transform 1 0 64128 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_675
timestamp 1677579658
transform 1 0 65376 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_683
timestamp 1679577901
transform 1 0 66144 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_692
timestamp 1679581782
transform 1 0 67008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_699
timestamp 1679577901
transform 1 0 67680 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_716
timestamp 1679581782
transform 1 0 69312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_723
timestamp 1679581782
transform 1 0 69984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_730
timestamp 1679577901
transform 1 0 70656 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_734
timestamp 1677580104
transform 1 0 71040 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_777
timestamp 1679581782
transform 1 0 75168 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_784
timestamp 1677580104
transform 1 0 75840 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_798
timestamp 1677579658
transform 1 0 77184 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_807
timestamp 1679581782
transform 1 0 78048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_814
timestamp 1679581782
transform 1 0 78720 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_821
timestamp 1677580104
transform 1 0 79392 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 6624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 7968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 8640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 9984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 10656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 12672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 18720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679581782
transform 1 0 19392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679581782
transform 1 0 20064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679581782
transform 1 0 20736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679581782
transform 1 0 21408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679581782
transform 1 0 22080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679581782
transform 1 0 22752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679581782
transform 1 0 23424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679581782
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 27456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 28128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679581782
transform 1 0 28800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679581782
transform 1 0 29472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679581782
transform 1 0 30144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679581782
transform 1 0 30816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679581782
transform 1 0 31488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_329
timestamp 1679581782
transform 1 0 32160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_336
timestamp 1679581782
transform 1 0 32832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_343
timestamp 1679581782
transform 1 0 33504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679581782
transform 1 0 34176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679581782
transform 1 0 34848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679581782
transform 1 0 35520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679581782
transform 1 0 36192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679581782
transform 1 0 36864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679581782
transform 1 0 37536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679581782
transform 1 0 38208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679581782
transform 1 0 38880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679581782
transform 1 0 39552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679581782
transform 1 0 40224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679581782
transform 1 0 40896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679581782
transform 1 0 41568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679581782
transform 1 0 42240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679581782
transform 1 0 42912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_448
timestamp 1679581782
transform 1 0 43584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_455
timestamp 1679581782
transform 1 0 44256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_462
timestamp 1679581782
transform 1 0 44928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_469
timestamp 1679581782
transform 1 0 45600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_476
timestamp 1679581782
transform 1 0 46272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679581782
transform 1 0 46944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679581782
transform 1 0 47616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_497
timestamp 1679581782
transform 1 0 48288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_504
timestamp 1679581782
transform 1 0 48960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_511
timestamp 1679581782
transform 1 0 49632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_518
timestamp 1679581782
transform 1 0 50304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_525
timestamp 1679581782
transform 1 0 50976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_532
timestamp 1679581782
transform 1 0 51648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_539
timestamp 1679581782
transform 1 0 52320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_546
timestamp 1679581782
transform 1 0 52992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_553
timestamp 1679581782
transform 1 0 53664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_560
timestamp 1679581782
transform 1 0 54336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_567
timestamp 1679581782
transform 1 0 55008 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_574
timestamp 1677580104
transform 1 0 55680 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_576
timestamp 1677579658
transform 1 0 55872 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_604
timestamp 1679581782
transform 1 0 58560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_611
timestamp 1679577901
transform 1 0 59232 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_615
timestamp 1677579658
transform 1 0 59616 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_623
timestamp 1677579658
transform 1 0 60384 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_629
timestamp 1677580104
transform 1 0 60960 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_631
timestamp 1677579658
transform 1 0 61152 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_662
timestamp 1677579658
transform 1 0 64128 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_672
timestamp 1677580104
transform 1 0 65088 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_674
timestamp 1677579658
transform 1 0 65280 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_716
timestamp 1677580104
transform 1 0 69312 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_718
timestamp 1677579658
transform 1 0 69504 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_746
timestamp 1677580104
transform 1 0 72192 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_756
timestamp 1677580104
transform 1 0 73152 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_761
timestamp 1677580104
transform 1 0 73632 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_763
timestamp 1677579658
transform 1 0 73824 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_769
timestamp 1679581782
transform 1 0 74400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_776
timestamp 1679581782
transform 1 0 75072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_783
timestamp 1679581782
transform 1 0 75744 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_790
timestamp 1677580104
transform 1 0 76416 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_801
timestamp 1677579658
transform 1 0 77472 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 17760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679581782
transform 1 0 18432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679581782
transform 1 0 19776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_207
timestamp 1679581782
transform 1 0 20448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_214
timestamp 1679581782
transform 1 0 21120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_221
timestamp 1679581782
transform 1 0 21792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_228
timestamp 1679581782
transform 1 0 22464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_235
timestamp 1679581782
transform 1 0 23136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_249
timestamp 1679581782
transform 1 0 24480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679581782
transform 1 0 25152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679581782
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_270
timestamp 1679581782
transform 1 0 26496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_277
timestamp 1679581782
transform 1 0 27168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_284
timestamp 1679581782
transform 1 0 27840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_291
timestamp 1679581782
transform 1 0 28512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_305
timestamp 1679581782
transform 1 0 29856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_312
timestamp 1679581782
transform 1 0 30528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_319
timestamp 1679581782
transform 1 0 31200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_326
timestamp 1679581782
transform 1 0 31872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_333
timestamp 1679581782
transform 1 0 32544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_340
timestamp 1679581782
transform 1 0 33216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_347
timestamp 1679581782
transform 1 0 33888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_354
timestamp 1679581782
transform 1 0 34560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_361
timestamp 1679581782
transform 1 0 35232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679581782
transform 1 0 35904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679581782
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679581782
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_389
timestamp 1679581782
transform 1 0 37920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_396
timestamp 1679581782
transform 1 0 38592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_403
timestamp 1679581782
transform 1 0 39264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_410
timestamp 1679581782
transform 1 0 39936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_417
timestamp 1679581782
transform 1 0 40608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_424
timestamp 1679581782
transform 1 0 41280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_431
timestamp 1679581782
transform 1 0 41952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_438
timestamp 1679581782
transform 1 0 42624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_445
timestamp 1679581782
transform 1 0 43296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_452
timestamp 1679581782
transform 1 0 43968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_459
timestamp 1679581782
transform 1 0 44640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_466
timestamp 1679581782
transform 1 0 45312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_473
timestamp 1679581782
transform 1 0 45984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_480
timestamp 1679581782
transform 1 0 46656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_487
timestamp 1679581782
transform 1 0 47328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_494
timestamp 1679581782
transform 1 0 48000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_501
timestamp 1679581782
transform 1 0 48672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_508
timestamp 1679581782
transform 1 0 49344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_515
timestamp 1679581782
transform 1 0 50016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_522
timestamp 1679581782
transform 1 0 50688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_529
timestamp 1679581782
transform 1 0 51360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_536
timestamp 1679581782
transform 1 0 52032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_543
timestamp 1679581782
transform 1 0 52704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_550
timestamp 1679577901
transform 1 0 53376 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_586
timestamp 1677579658
transform 1 0 56832 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_599
timestamp 1679581782
transform 1 0 58080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_606
timestamp 1679581782
transform 1 0 58752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_683
timestamp 1679581782
transform 1 0 66144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_690
timestamp 1679581782
transform 1 0 66816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_697
timestamp 1679581782
transform 1 0 67488 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_704
timestamp 1677579658
transform 1 0 68160 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_718
timestamp 1679581782
transform 1 0 69504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_725
timestamp 1679581782
transform 1 0 70176 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_732
timestamp 1677579658
transform 1 0 70848 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_778
timestamp 1679577901
transform 1 0 75264 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_782
timestamp 1677579658
transform 1 0 75648 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_822
timestamp 1677579658
transform 1 0 79488 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_536
timestamp 1677579658
transform 1 0 52032 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_543
timestamp 1679577901
transform 1 0 52704 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_547
timestamp 1677580104
transform 1 0 53088 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_552
timestamp 1677580104
transform 1 0 53568 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_554
timestamp 1677579658
transform 1 0 53760 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_566
timestamp 1679581782
transform 1 0 54912 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_573
timestamp 1677579658
transform 1 0 55584 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_577
timestamp 1679581782
transform 1 0 55968 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_584
timestamp 1677580104
transform 1 0 56640 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_618
timestamp 1679577901
transform 1 0 59904 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_622
timestamp 1677579658
transform 1 0 60288 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_632
timestamp 1677579658
transform 1 0 61248 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_644
timestamp 1679581782
transform 1 0 62400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_651
timestamp 1679581782
transform 1 0 63072 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_658
timestamp 1677580104
transform 1 0 63744 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_660
timestamp 1677579658
transform 1 0 63936 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_673
timestamp 1677579658
transform 1 0 65184 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_758
timestamp 1679581782
transform 1 0 73344 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_765
timestamp 1677580104
transform 1 0 74016 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_807
timestamp 1679581782
transform 1 0 78048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_814
timestamp 1679581782
transform 1 0 78720 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_821
timestamp 1677580104
transform 1 0 79392 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679581782
transform 1 0 5664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679581782
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679581782
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679581782
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679581782
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679581782
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679581782
transform 1 0 9696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679581782
transform 1 0 10368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679581782
transform 1 0 11040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 11712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 13728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 15744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_179
timestamp 1679581782
transform 1 0 17760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_186
timestamp 1679581782
transform 1 0 18432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_200
timestamp 1679581782
transform 1 0 19776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_207
timestamp 1679581782
transform 1 0 20448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_214
timestamp 1679581782
transform 1 0 21120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_221
timestamp 1679581782
transform 1 0 21792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_228
timestamp 1679581782
transform 1 0 22464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_235
timestamp 1679581782
transform 1 0 23136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_242
timestamp 1679581782
transform 1 0 23808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_249
timestamp 1679581782
transform 1 0 24480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_256
timestamp 1679581782
transform 1 0 25152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_263
timestamp 1679581782
transform 1 0 25824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_270
timestamp 1679581782
transform 1 0 26496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_277
timestamp 1679581782
transform 1 0 27168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_284
timestamp 1679581782
transform 1 0 27840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_291
timestamp 1679581782
transform 1 0 28512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_298
timestamp 1679581782
transform 1 0 29184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_305
timestamp 1679581782
transform 1 0 29856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_312
timestamp 1679581782
transform 1 0 30528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 31872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 32544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_340
timestamp 1679581782
transform 1 0 33216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_347
timestamp 1679581782
transform 1 0 33888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 34560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 35904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 36576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 37920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_396
timestamp 1679581782
transform 1 0 38592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_403
timestamp 1679581782
transform 1 0 39264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_410
timestamp 1679581782
transform 1 0 39936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_417
timestamp 1679581782
transform 1 0 40608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_424
timestamp 1679581782
transform 1 0 41280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_431
timestamp 1679581782
transform 1 0 41952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_438
timestamp 1679581782
transform 1 0 42624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_445
timestamp 1679581782
transform 1 0 43296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_452
timestamp 1679581782
transform 1 0 43968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_459
timestamp 1679581782
transform 1 0 44640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_466
timestamp 1679581782
transform 1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_473
timestamp 1679581782
transform 1 0 45984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_480
timestamp 1679581782
transform 1 0 46656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_487
timestamp 1679581782
transform 1 0 47328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_494
timestamp 1679581782
transform 1 0 48000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_501
timestamp 1679581782
transform 1 0 48672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_508
timestamp 1679581782
transform 1 0 49344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_515
timestamp 1679581782
transform 1 0 50016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_522
timestamp 1679581782
transform 1 0 50688 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_529
timestamp 1677580104
transform 1 0 51360 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_531
timestamp 1677579658
transform 1 0 51552 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_559
timestamp 1679581782
transform 1 0 54240 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_566
timestamp 1677580104
transform 1 0 54912 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_575
timestamp 1677579658
transform 1 0 55776 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_581
timestamp 1679581782
transform 1 0 56352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_588
timestamp 1679581782
transform 1 0 57024 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_595
timestamp 1677580104
transform 1 0 57696 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_627
timestamp 1677579658
transform 1 0 60768 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_635
timestamp 1679581782
transform 1 0 61536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_642
timestamp 1679581782
transform 1 0 62208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_649
timestamp 1679581782
transform 1 0 62880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_656
timestamp 1679581782
transform 1 0 63552 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_663
timestamp 1677580104
transform 1 0 64224 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_681
timestamp 1679581782
transform 1 0 65952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_688
timestamp 1679581782
transform 1 0 66624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_695
timestamp 1679581782
transform 1 0 67296 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_702
timestamp 1677579658
transform 1 0 67968 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_715
timestamp 1677579658
transform 1 0 69216 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_721
timestamp 1679581782
transform 1 0 69792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_728
timestamp 1679581782
transform 1 0 70464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_735
timestamp 1679581782
transform 1 0 71136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_742
timestamp 1679577901
transform 1 0 71808 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_752
timestamp 1677579658
transform 1 0 72768 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_760
timestamp 1679581782
transform 1 0 73536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_772
timestamp 1679581782
transform 1 0 74688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_779
timestamp 1679581782
transform 1 0 75360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_786
timestamp 1679581782
transform 1 0 76032 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_793
timestamp 1677579658
transform 1 0 76704 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_812
timestamp 1679581782
transform 1 0 78528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_819
timestamp 1679577901
transform 1 0 79200 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 9984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 10656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 12672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 20064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 22080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 22752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 23424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 24096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 24768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 25440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 26112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 26784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 27456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 28128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 28800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 29472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 30816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 31488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 32160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 32832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 33504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 34848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 35520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679581782
transform 1 0 36192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679581782
transform 1 0 36864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 37536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 38208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 38880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 39552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 40224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679581782
transform 1 0 40896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_427
timestamp 1679581782
transform 1 0 41568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_434
timestamp 1679581782
transform 1 0 42240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_441
timestamp 1679581782
transform 1 0 42912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_448
timestamp 1679581782
transform 1 0 43584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_455
timestamp 1679581782
transform 1 0 44256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_462
timestamp 1679581782
transform 1 0 44928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_469
timestamp 1679581782
transform 1 0 45600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_476
timestamp 1679581782
transform 1 0 46272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_483
timestamp 1679581782
transform 1 0 46944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_490
timestamp 1679581782
transform 1 0 47616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_497
timestamp 1679581782
transform 1 0 48288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_504
timestamp 1679581782
transform 1 0 48960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_511
timestamp 1679581782
transform 1 0 49632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_518
timestamp 1679581782
transform 1 0 50304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679581782
transform 1 0 50976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_532
timestamp 1679577901
transform 1 0 51648 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_536
timestamp 1677580104
transform 1 0 52032 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_555
timestamp 1679581782
transform 1 0 53856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_562
timestamp 1679577901
transform 1 0 54528 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_566
timestamp 1677579658
transform 1 0 54912 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_599
timestamp 1679581782
transform 1 0 58080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_606
timestamp 1679581782
transform 1 0 58752 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_613
timestamp 1677580104
transform 1 0 59424 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_615
timestamp 1677579658
transform 1 0 59616 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_621
timestamp 1679577901
transform 1 0 60192 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_684
timestamp 1679581782
transform 1 0 66240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_691
timestamp 1679581782
transform 1 0 66912 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_698
timestamp 1677580104
transform 1 0 67584 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_700
timestamp 1677579658
transform 1 0 67776 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_733
timestamp 1679577901
transform 1 0 70944 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_737
timestamp 1677579658
transform 1 0 71328 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_744
timestamp 1677580104
transform 1 0 72000 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_783
timestamp 1679581782
transform 1 0 75744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679581782
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679581782
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679581782
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679581782
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679581782
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679581782
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 11712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 13728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_144
timestamp 1679581782
transform 1 0 14400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_151
timestamp 1679581782
transform 1 0 15072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 15744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 17760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 18432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_200
timestamp 1679581782
transform 1 0 19776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_207
timestamp 1679581782
transform 1 0 20448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_214
timestamp 1679581782
transform 1 0 21120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_221
timestamp 1679581782
transform 1 0 21792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_228
timestamp 1679581782
transform 1 0 22464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_235
timestamp 1679581782
transform 1 0 23136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_242
timestamp 1679581782
transform 1 0 23808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_249
timestamp 1679581782
transform 1 0 24480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_256
timestamp 1679581782
transform 1 0 25152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_263
timestamp 1679581782
transform 1 0 25824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_270
timestamp 1679581782
transform 1 0 26496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_277
timestamp 1679581782
transform 1 0 27168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_284
timestamp 1679581782
transform 1 0 27840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_291
timestamp 1679581782
transform 1 0 28512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_298
timestamp 1679581782
transform 1 0 29184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_305
timestamp 1679581782
transform 1 0 29856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_312
timestamp 1679581782
transform 1 0 30528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_319
timestamp 1679581782
transform 1 0 31200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 31872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_333
timestamp 1679581782
transform 1 0 32544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_340
timestamp 1679581782
transform 1 0 33216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_347
timestamp 1679581782
transform 1 0 33888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 34560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_361
timestamp 1679581782
transform 1 0 35232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_368
timestamp 1679581782
transform 1 0 35904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_375
timestamp 1679581782
transform 1 0 36576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_382
timestamp 1679581782
transform 1 0 37248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_389
timestamp 1679581782
transform 1 0 37920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_396
timestamp 1679581782
transform 1 0 38592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_403
timestamp 1679581782
transform 1 0 39264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 39936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 40608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_424
timestamp 1679581782
transform 1 0 41280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_431
timestamp 1679581782
transform 1 0 41952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_438
timestamp 1679581782
transform 1 0 42624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_445
timestamp 1679581782
transform 1 0 43296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_452
timestamp 1679581782
transform 1 0 43968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_459
timestamp 1679581782
transform 1 0 44640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_466
timestamp 1679581782
transform 1 0 45312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_473
timestamp 1679581782
transform 1 0 45984 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_480
timestamp 1677579658
transform 1 0 46656 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_484
timestamp 1679581782
transform 1 0 47040 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_491
timestamp 1677579658
transform 1 0 47712 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_498
timestamp 1679581782
transform 1 0 48384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_505
timestamp 1679581782
transform 1 0 49056 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_512
timestamp 1677580104
transform 1 0 49728 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_514
timestamp 1677579658
transform 1 0 49920 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_520
timestamp 1679581782
transform 1 0 50496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_527
timestamp 1679577901
transform 1 0 51168 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_531
timestamp 1677579658
transform 1 0 51552 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_564
timestamp 1679581782
transform 1 0 54720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_571
timestamp 1679577901
transform 1 0 55392 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_575
timestamp 1677580104
transform 1 0 55776 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_581
timestamp 1677580104
transform 1 0 56352 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_586
timestamp 1677580104
transform 1 0 56832 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_621
timestamp 1679581782
transform 1 0 60192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_628
timestamp 1679577901
transform 1 0 60864 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_632
timestamp 1677580104
transform 1 0 61248 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_639
timestamp 1677579658
transform 1 0 61920 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_643
timestamp 1679581782
transform 1 0 62304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_650
timestamp 1679581782
transform 1 0 62976 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_657
timestamp 1677580104
transform 1 0 63648 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_659
timestamp 1677579658
transform 1 0 63840 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_668
timestamp 1677579658
transform 1 0 64704 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_679
timestamp 1677580104
transform 1 0 65760 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_681
timestamp 1677579658
transform 1 0 65952 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_713
timestamp 1679581782
transform 1 0 69024 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_720
timestamp 1677580104
transform 1 0 69696 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_722
timestamp 1677579658
transform 1 0 69888 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_753
timestamp 1679577901
transform 1 0 72864 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_766
timestamp 1679581782
transform 1 0 74112 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_773
timestamp 1677579658
transform 1 0 74784 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_777
timestamp 1679577901
transform 1 0 75168 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_816
timestamp 1679581782
transform 1 0 78912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679581782
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679581782
transform 1 0 3648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679581782
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 4992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679581782
transform 1 0 5664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679581782
transform 1 0 6336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679581782
transform 1 0 7008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679581782
transform 1 0 7680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679581782
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_123
timestamp 1679581782
transform 1 0 12384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679581782
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679581782
transform 1 0 13728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679581782
transform 1 0 14400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_151
timestamp 1679581782
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_158
timestamp 1679581782
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_165
timestamp 1679581782
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_172
timestamp 1679581782
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_179
timestamp 1679581782
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_186
timestamp 1679581782
transform 1 0 18432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_193
timestamp 1679581782
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_200
timestamp 1679581782
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1679581782
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_214
timestamp 1679581782
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_221
timestamp 1679581782
transform 1 0 21792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_228
timestamp 1679581782
transform 1 0 22464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_235
timestamp 1679581782
transform 1 0 23136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 23808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_249
timestamp 1679581782
transform 1 0 24480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_256
timestamp 1679581782
transform 1 0 25152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_263
timestamp 1679581782
transform 1 0 25824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_270
timestamp 1679581782
transform 1 0 26496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_277
timestamp 1679581782
transform 1 0 27168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_284
timestamp 1679581782
transform 1 0 27840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 28512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 29856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 30528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_319
timestamp 1679581782
transform 1 0 31200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 31872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_333
timestamp 1679581782
transform 1 0 32544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_340
timestamp 1679581782
transform 1 0 33216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_347
timestamp 1679581782
transform 1 0 33888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_354
timestamp 1679581782
transform 1 0 34560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679581782
transform 1 0 35232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679581782
transform 1 0 35904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679581782
transform 1 0 36576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_382
timestamp 1679581782
transform 1 0 37248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_389
timestamp 1679581782
transform 1 0 37920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_396
timestamp 1679581782
transform 1 0 38592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_403
timestamp 1679581782
transform 1 0 39264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679581782
transform 1 0 39936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679581782
transform 1 0 40608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679581782
transform 1 0 41280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679581782
transform 1 0 41952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_438
timestamp 1679581782
transform 1 0 42624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_445
timestamp 1679581782
transform 1 0 43296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_452
timestamp 1679581782
transform 1 0 43968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_459
timestamp 1679577901
transform 1 0 44640 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_463
timestamp 1677579658
transform 1 0 45024 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_491
timestamp 1677579658
transform 1 0 47712 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_519
timestamp 1677580104
transform 1 0 50400 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_548
timestamp 1677579658
transform 1 0 53184 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_552
timestamp 1677580104
transform 1 0 53568 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_580
timestamp 1679581782
transform 1 0 56256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_587
timestamp 1679581782
transform 1 0 56928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_594
timestamp 1679581782
transform 1 0 57600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_629
timestamp 1679581782
transform 1 0 60960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_636
timestamp 1679577901
transform 1 0 61632 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_640
timestamp 1677579658
transform 1 0 62016 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_672
timestamp 1679577901
transform 1 0 65088 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_676
timestamp 1677580104
transform 1 0 65472 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_691
timestamp 1679581782
transform 1 0 66912 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_698
timestamp 1677580104
transform 1 0 67584 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_700
timestamp 1677579658
transform 1 0 67776 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_707
timestamp 1677580104
transform 1 0 68448 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_717
timestamp 1679581782
transform 1 0 69408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_724
timestamp 1679581782
transform 1 0 70080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_731
timestamp 1679581782
transform 1 0 70752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_777
timestamp 1679581782
transform 1 0 75168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_784
timestamp 1679577901
transform 1 0 75840 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_788
timestamp 1677580104
transform 1 0 76224 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_809
timestamp 1679581782
transform 1 0 78240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_816
timestamp 1679581782
transform 1 0 78912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_53
timestamp 1679581782
transform 1 0 5664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_60
timestamp 1679581782
transform 1 0 6336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_67
timestamp 1679581782
transform 1 0 7008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_74
timestamp 1679581782
transform 1 0 7680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_81
timestamp 1679581782
transform 1 0 8352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_88
timestamp 1679581782
transform 1 0 9024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_95
timestamp 1679581782
transform 1 0 9696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_102
timestamp 1679581782
transform 1 0 10368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_109
timestamp 1679581782
transform 1 0 11040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 11712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_123
timestamp 1679581782
transform 1 0 12384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_130
timestamp 1679581782
transform 1 0 13056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_137
timestamp 1679581782
transform 1 0 13728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_144
timestamp 1679581782
transform 1 0 14400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_151
timestamp 1679581782
transform 1 0 15072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_158
timestamp 1679581782
transform 1 0 15744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_165
timestamp 1679581782
transform 1 0 16416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_172
timestamp 1679581782
transform 1 0 17088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_179
timestamp 1679581782
transform 1 0 17760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_186
timestamp 1679581782
transform 1 0 18432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_193
timestamp 1679581782
transform 1 0 19104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_200
timestamp 1679581782
transform 1 0 19776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_207
timestamp 1679581782
transform 1 0 20448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_214
timestamp 1679581782
transform 1 0 21120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_221
timestamp 1679581782
transform 1 0 21792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_228
timestamp 1679581782
transform 1 0 22464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_235
timestamp 1679581782
transform 1 0 23136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_242
timestamp 1679581782
transform 1 0 23808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_249
timestamp 1679581782
transform 1 0 24480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_256
timestamp 1679581782
transform 1 0 25152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_263
timestamp 1679581782
transform 1 0 25824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_270
timestamp 1679581782
transform 1 0 26496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_277
timestamp 1679581782
transform 1 0 27168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_284
timestamp 1679581782
transform 1 0 27840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_291
timestamp 1679581782
transform 1 0 28512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_298
timestamp 1679581782
transform 1 0 29184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1679581782
transform 1 0 29856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_312
timestamp 1679581782
transform 1 0 30528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_319
timestamp 1679581782
transform 1 0 31200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_326
timestamp 1679581782
transform 1 0 31872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_333
timestamp 1679581782
transform 1 0 32544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_340
timestamp 1679581782
transform 1 0 33216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_347
timestamp 1679581782
transform 1 0 33888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_354
timestamp 1679581782
transform 1 0 34560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_361
timestamp 1679581782
transform 1 0 35232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_368
timestamp 1679581782
transform 1 0 35904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_375
timestamp 1679581782
transform 1 0 36576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_382
timestamp 1679581782
transform 1 0 37248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_389
timestamp 1679581782
transform 1 0 37920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_396
timestamp 1679581782
transform 1 0 38592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_403
timestamp 1679581782
transform 1 0 39264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_410
timestamp 1679581782
transform 1 0 39936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_417
timestamp 1679581782
transform 1 0 40608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679581782
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679581782
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679581782
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679581782
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_452
timestamp 1679577901
transform 1 0 43968 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_471
timestamp 1679581782
transform 1 0 45792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_478
timestamp 1679581782
transform 1 0 46464 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_485
timestamp 1677580104
transform 1 0 47136 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_487
timestamp 1677579658
transform 1 0 47328 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_493
timestamp 1679577901
transform 1 0 47904 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_509
timestamp 1677580104
transform 1 0 49440 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_525
timestamp 1677580104
transform 1 0 50976 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_551
timestamp 1679581782
transform 1 0 53472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_558
timestamp 1679581782
transform 1 0 54144 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_600
timestamp 1677580104
transform 1 0 58176 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_602
timestamp 1677579658
transform 1 0 58368 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_614
timestamp 1677580104
transform 1 0 59520 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_643
timestamp 1679577901
transform 1 0 62304 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_647
timestamp 1677579658
transform 1 0 62688 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_654
timestamp 1677579658
transform 1 0 63360 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_667
timestamp 1679581782
transform 1 0 64608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_674
timestamp 1679577901
transform 1 0 65280 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_678
timestamp 1677580104
transform 1 0 65664 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_718
timestamp 1677579658
transform 1 0 69504 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_746
timestamp 1677579658
transform 1 0 72192 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_755
timestamp 1679581782
transform 1 0 73056 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_762
timestamp 1677580104
transform 1 0 73728 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_768
timestamp 1677579658
transform 1 0 74304 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_772
timestamp 1679581782
transform 1 0 74688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_779
timestamp 1679581782
transform 1 0 75360 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_786
timestamp 1677580104
transform 1 0 76032 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_821
timestamp 1677580104
transform 1 0 79392 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_32
timestamp 1679581782
transform 1 0 3648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679581782
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679581782
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679581782
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679581782
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679581782
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_95
timestamp 1679581782
transform 1 0 9696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_102
timestamp 1679581782
transform 1 0 10368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_109
timestamp 1679581782
transform 1 0 11040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_116
timestamp 1679581782
transform 1 0 11712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_137
timestamp 1679581782
transform 1 0 13728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679581782
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679581782
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_158
timestamp 1679581782
transform 1 0 15744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 17760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_186
timestamp 1679581782
transform 1 0 18432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_200
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_207
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679581782
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_221
timestamp 1679581782
transform 1 0 21792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_228
timestamp 1679581782
transform 1 0 22464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_235
timestamp 1679581782
transform 1 0 23136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_242
timestamp 1679581782
transform 1 0 23808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 24480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_263
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_270
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 27840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_291
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_298
timestamp 1679581782
transform 1 0 29184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1679581782
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1679581782
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_319
timestamp 1679581782
transform 1 0 31200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_326
timestamp 1679581782
transform 1 0 31872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_333
timestamp 1679581782
transform 1 0 32544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_340
timestamp 1679581782
transform 1 0 33216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 33888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 34560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_368
timestamp 1679581782
transform 1 0 35904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_375
timestamp 1679581782
transform 1 0 36576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_382
timestamp 1679581782
transform 1 0 37248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_389
timestamp 1679581782
transform 1 0 37920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_396
timestamp 1679581782
transform 1 0 38592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_410
timestamp 1679581782
transform 1 0 39936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_417
timestamp 1679581782
transform 1 0 40608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_424
timestamp 1679581782
transform 1 0 41280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_431
timestamp 1679577901
transform 1 0 41952 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_435
timestamp 1677580104
transform 1 0 42336 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_464
timestamp 1677579658
transform 1 0 45120 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_469
timestamp 1677580104
transform 1 0 45600 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_483
timestamp 1677579658
transform 1 0 46944 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_487
timestamp 1679581782
transform 1 0 47328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_499
timestamp 1679581782
transform 1 0 48480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_543
timestamp 1679581782
transform 1 0 52704 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_577
timestamp 1677579658
transform 1 0 55968 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_582
timestamp 1679577901
transform 1 0 56448 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_586
timestamp 1677580104
transform 1 0 56832 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_615
timestamp 1679577901
transform 1 0 59616 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679581782
transform 1 0 60384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679581782
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_641
timestamp 1679577901
transform 1 0 62112 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_645
timestamp 1677579658
transform 1 0 62496 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_687
timestamp 1679581782
transform 1 0 66528 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_694
timestamp 1677580104
transform 1 0 67200 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_731
timestamp 1679581782
transform 1 0 70752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_738
timestamp 1679577901
transform 1 0 71424 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_742
timestamp 1677579658
transform 1 0 71808 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_765
timestamp 1679581782
transform 1 0 74016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_772
timestamp 1679577901
transform 1 0 74688 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_776
timestamp 1677580104
transform 1 0 75072 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_814
timestamp 1679581782
transform 1 0 78720 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_821
timestamp 1677580104
transform 1 0 79392 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_4
timestamp 1679577901
transform 1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_8
timestamp 1677579658
transform 1 0 1344 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_13
timestamp 1679581782
transform 1 0 1824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_20
timestamp 1679581782
transform 1 0 2496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_27
timestamp 1679581782
transform 1 0 3168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_34
timestamp 1679581782
transform 1 0 3840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_41
timestamp 1679581782
transform 1 0 4512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_48
timestamp 1679581782
transform 1 0 5184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_55
timestamp 1679581782
transform 1 0 5856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_62
timestamp 1679581782
transform 1 0 6528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_69
timestamp 1679581782
transform 1 0 7200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_76
timestamp 1679581782
transform 1 0 7872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_83
timestamp 1679581782
transform 1 0 8544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_90
timestamp 1679581782
transform 1 0 9216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_97
timestamp 1679581782
transform 1 0 9888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_104
timestamp 1679581782
transform 1 0 10560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_111
timestamp 1679581782
transform 1 0 11232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_118
timestamp 1679581782
transform 1 0 11904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_125
timestamp 1679581782
transform 1 0 12576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_132
timestamp 1679581782
transform 1 0 13248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_139
timestamp 1679581782
transform 1 0 13920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_146
timestamp 1679581782
transform 1 0 14592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_153
timestamp 1679581782
transform 1 0 15264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_160
timestamp 1679581782
transform 1 0 15936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_167
timestamp 1679581782
transform 1 0 16608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_174
timestamp 1679581782
transform 1 0 17280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_181
timestamp 1679581782
transform 1 0 17952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_188
timestamp 1679581782
transform 1 0 18624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_195
timestamp 1679581782
transform 1 0 19296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_202
timestamp 1679581782
transform 1 0 19968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_209
timestamp 1679581782
transform 1 0 20640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_216
timestamp 1679581782
transform 1 0 21312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_223
timestamp 1679581782
transform 1 0 21984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_230
timestamp 1679581782
transform 1 0 22656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_237
timestamp 1679581782
transform 1 0 23328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_244
timestamp 1679581782
transform 1 0 24000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_251
timestamp 1679581782
transform 1 0 24672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_258
timestamp 1679581782
transform 1 0 25344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_265
timestamp 1679581782
transform 1 0 26016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_272
timestamp 1679581782
transform 1 0 26688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_279
timestamp 1679581782
transform 1 0 27360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_286
timestamp 1679581782
transform 1 0 28032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_293
timestamp 1679581782
transform 1 0 28704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_300
timestamp 1679581782
transform 1 0 29376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_307
timestamp 1679581782
transform 1 0 30048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_314
timestamp 1679581782
transform 1 0 30720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_321
timestamp 1679581782
transform 1 0 31392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_328
timestamp 1679581782
transform 1 0 32064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_335
timestamp 1679581782
transform 1 0 32736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_342
timestamp 1679581782
transform 1 0 33408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_349
timestamp 1679581782
transform 1 0 34080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_356
timestamp 1679581782
transform 1 0 34752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_363
timestamp 1679581782
transform 1 0 35424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_370
timestamp 1679581782
transform 1 0 36096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_377
timestamp 1679581782
transform 1 0 36768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_384
timestamp 1679581782
transform 1 0 37440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_391
timestamp 1679581782
transform 1 0 38112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_398
timestamp 1679581782
transform 1 0 38784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_405
timestamp 1679581782
transform 1 0 39456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_412
timestamp 1679581782
transform 1 0 40128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_419
timestamp 1679581782
transform 1 0 40800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_426
timestamp 1679581782
transform 1 0 41472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_433
timestamp 1679581782
transform 1 0 42144 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_440
timestamp 1677580104
transform 1 0 42816 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_448
timestamp 1679577901
transform 1 0 43584 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_452
timestamp 1677579658
transform 1 0 43968 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_456
timestamp 1677579658
transform 1 0 44352 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_520
timestamp 1677580104
transform 1 0 50496 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_531
timestamp 1677579658
transform 1 0 51552 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_559
timestamp 1679577901
transform 1 0 54240 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_563
timestamp 1677579658
transform 1 0 54624 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_581
timestamp 1679581782
transform 1 0 56352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_588
timestamp 1679581782
transform 1 0 57024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_595
timestamp 1679577901
transform 1 0 57696 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_622
timestamp 1677580104
transform 1 0 60288 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_624
timestamp 1677579658
transform 1 0 60480 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679581782
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_662
timestamp 1677580104
transform 1 0 64128 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_664
timestamp 1677579658
transform 1 0 64320 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_672
timestamp 1679581782
transform 1 0 65088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_679
timestamp 1679581782
transform 1 0 65760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_686
timestamp 1679577901
transform 1 0 66432 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_690
timestamp 1677579658
transform 1 0 66816 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_697
timestamp 1679581782
transform 1 0 67488 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_709
timestamp 1677580104
transform 1 0 68640 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_711
timestamp 1677579658
transform 1 0 68832 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_728
timestamp 1679581782
transform 1 0 70464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_735
timestamp 1679577901
transform 1 0 71136 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_739
timestamp 1677579658
transform 1 0 71520 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_751
timestamp 1677579658
transform 1 0 72672 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_779
timestamp 1679581782
transform 1 0 75360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_786
timestamp 1679577901
transform 1 0 76032 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_809
timestamp 1679581782
transform 1 0 78240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_816
timestamp 1679581782
transform 1 0 78912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679581782
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679581782
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679581782
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679581782
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679581782
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679581782
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679581782
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679581782
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679581782
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679581782
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_88
timestamp 1679581782
transform 1 0 9024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_95
timestamp 1679581782
transform 1 0 9696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_102
timestamp 1679581782
transform 1 0 10368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_109
timestamp 1679581782
transform 1 0 11040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_116
timestamp 1679581782
transform 1 0 11712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_123
timestamp 1679581782
transform 1 0 12384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_130
timestamp 1679581782
transform 1 0 13056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_137
timestamp 1679581782
transform 1 0 13728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_144
timestamp 1679581782
transform 1 0 14400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_151
timestamp 1679581782
transform 1 0 15072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_158
timestamp 1679581782
transform 1 0 15744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_165
timestamp 1679581782
transform 1 0 16416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_172
timestamp 1679581782
transform 1 0 17088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_179
timestamp 1679581782
transform 1 0 17760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_186
timestamp 1679581782
transform 1 0 18432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_193
timestamp 1679581782
transform 1 0 19104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_200
timestamp 1679581782
transform 1 0 19776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_207
timestamp 1679581782
transform 1 0 20448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_214
timestamp 1679581782
transform 1 0 21120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_221
timestamp 1679581782
transform 1 0 21792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_228
timestamp 1679581782
transform 1 0 22464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_235
timestamp 1679581782
transform 1 0 23136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_242
timestamp 1679581782
transform 1 0 23808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_249
timestamp 1679581782
transform 1 0 24480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_256
timestamp 1679581782
transform 1 0 25152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_263
timestamp 1679581782
transform 1 0 25824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_270
timestamp 1679581782
transform 1 0 26496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_277
timestamp 1679581782
transform 1 0 27168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_284
timestamp 1679581782
transform 1 0 27840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_291
timestamp 1679581782
transform 1 0 28512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_298
timestamp 1679581782
transform 1 0 29184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_305
timestamp 1679581782
transform 1 0 29856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_312
timestamp 1679581782
transform 1 0 30528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_319
timestamp 1679581782
transform 1 0 31200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_326
timestamp 1679581782
transform 1 0 31872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_333
timestamp 1679581782
transform 1 0 32544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_340
timestamp 1679581782
transform 1 0 33216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_347
timestamp 1679581782
transform 1 0 33888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_354
timestamp 1679581782
transform 1 0 34560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_361
timestamp 1679581782
transform 1 0 35232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_368
timestamp 1679581782
transform 1 0 35904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_375
timestamp 1679581782
transform 1 0 36576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_382
timestamp 1679581782
transform 1 0 37248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_389
timestamp 1679581782
transform 1 0 37920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_396
timestamp 1679581782
transform 1 0 38592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_403
timestamp 1679581782
transform 1 0 39264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_410
timestamp 1679581782
transform 1 0 39936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_417
timestamp 1679581782
transform 1 0 40608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_424
timestamp 1679581782
transform 1 0 41280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_431
timestamp 1679577901
transform 1 0 41952 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_435
timestamp 1677579658
transform 1 0 42336 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_458
timestamp 1679581782
transform 1 0 44544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_465
timestamp 1679577901
transform 1 0 45216 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_478
timestamp 1679581782
transform 1 0 46464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_485
timestamp 1679581782
transform 1 0 47136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_492
timestamp 1679581782
transform 1 0 47808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_499
timestamp 1679581782
transform 1 0 48480 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_506
timestamp 1677579658
transform 1 0 49152 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_510
timestamp 1679581782
transform 1 0 49536 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_527
timestamp 1677580104
transform 1 0 51168 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_546
timestamp 1679581782
transform 1 0 52992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_553
timestamp 1679581782
transform 1 0 53664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_560
timestamp 1679581782
transform 1 0 54336 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_567
timestamp 1677579658
transform 1 0 55008 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_573
timestamp 1677579658
transform 1 0 55584 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_606
timestamp 1677579658
transform 1 0 58752 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_634
timestamp 1677580104
transform 1 0 61440 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_659
timestamp 1679581782
transform 1 0 63840 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_666
timestamp 1677580104
transform 1 0 64512 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_702
timestamp 1679581782
transform 1 0 67968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_713
timestamp 1679581782
transform 1 0 69024 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_720
timestamp 1677580104
transform 1 0 69696 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_749
timestamp 1677580104
transform 1 0 72480 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_756
timestamp 1677579658
transform 1 0 73152 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_761
timestamp 1677580104
transform 1 0 73632 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_767
timestamp 1679577901
transform 1 0 74208 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_808
timestamp 1679581782
transform 1 0 78144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_815
timestamp 1679581782
transform 1 0 78816 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_822
timestamp 1677579658
transform 1 0 79488 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_4
timestamp 1679577901
transform 1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_8
timestamp 1677579658
transform 1 0 1344 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_13
timestamp 1679581782
transform 1 0 1824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_20
timestamp 1679581782
transform 1 0 2496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_27
timestamp 1679581782
transform 1 0 3168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_34
timestamp 1679581782
transform 1 0 3840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_41
timestamp 1679581782
transform 1 0 4512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_48
timestamp 1679581782
transform 1 0 5184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_55
timestamp 1679581782
transform 1 0 5856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_62
timestamp 1679581782
transform 1 0 6528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_69
timestamp 1679581782
transform 1 0 7200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_76
timestamp 1679581782
transform 1 0 7872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_83
timestamp 1679581782
transform 1 0 8544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_90
timestamp 1679581782
transform 1 0 9216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_97
timestamp 1679581782
transform 1 0 9888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_104
timestamp 1679581782
transform 1 0 10560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_111
timestamp 1679581782
transform 1 0 11232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_118
timestamp 1679581782
transform 1 0 11904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_125
timestamp 1679581782
transform 1 0 12576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_132
timestamp 1679581782
transform 1 0 13248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_139
timestamp 1679581782
transform 1 0 13920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_146
timestamp 1679581782
transform 1 0 14592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_153
timestamp 1679581782
transform 1 0 15264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_160
timestamp 1679581782
transform 1 0 15936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_167
timestamp 1679581782
transform 1 0 16608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_174
timestamp 1679581782
transform 1 0 17280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_181
timestamp 1679581782
transform 1 0 17952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_188
timestamp 1679581782
transform 1 0 18624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_195
timestamp 1679581782
transform 1 0 19296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_202
timestamp 1679581782
transform 1 0 19968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_209
timestamp 1679581782
transform 1 0 20640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_216
timestamp 1679581782
transform 1 0 21312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_223
timestamp 1679581782
transform 1 0 21984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_230
timestamp 1679581782
transform 1 0 22656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_237
timestamp 1679581782
transform 1 0 23328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_244
timestamp 1679581782
transform 1 0 24000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_251
timestamp 1679581782
transform 1 0 24672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_258
timestamp 1679581782
transform 1 0 25344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_265
timestamp 1679581782
transform 1 0 26016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_272
timestamp 1679581782
transform 1 0 26688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_279
timestamp 1679581782
transform 1 0 27360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_286
timestamp 1679581782
transform 1 0 28032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_293
timestamp 1679581782
transform 1 0 28704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_300
timestamp 1679581782
transform 1 0 29376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_307
timestamp 1679581782
transform 1 0 30048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_314
timestamp 1679581782
transform 1 0 30720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_321
timestamp 1679581782
transform 1 0 31392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_328
timestamp 1679581782
transform 1 0 32064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_335
timestamp 1679581782
transform 1 0 32736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_342
timestamp 1679581782
transform 1 0 33408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_349
timestamp 1679581782
transform 1 0 34080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_356
timestamp 1679581782
transform 1 0 34752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_363
timestamp 1679581782
transform 1 0 35424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_370
timestamp 1679581782
transform 1 0 36096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_377
timestamp 1679581782
transform 1 0 36768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_384
timestamp 1679581782
transform 1 0 37440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_391
timestamp 1679581782
transform 1 0 38112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_398
timestamp 1679581782
transform 1 0 38784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_405
timestamp 1679581782
transform 1 0 39456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_412
timestamp 1679581782
transform 1 0 40128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_419
timestamp 1679577901
transform 1 0 40800 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_484
timestamp 1679581782
transform 1 0 47040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_491
timestamp 1679577901
transform 1 0 47712 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_495
timestamp 1677579658
transform 1 0 48096 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_535
timestamp 1679581782
transform 1 0 51936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_542
timestamp 1679581782
transform 1 0 52608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_584
timestamp 1679581782
transform 1 0 56640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_591
timestamp 1679581782
transform 1 0 57312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_598
timestamp 1679581782
transform 1 0 57984 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_605
timestamp 1677580104
transform 1 0 58656 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_612
timestamp 1677579658
transform 1 0 59328 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_622
timestamp 1679581782
transform 1 0 60288 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_629
timestamp 1677580104
transform 1 0 60960 0 1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_14_635
timestamp 1679577901
transform 1 0 61536 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_639
timestamp 1677580104
transform 1 0 61920 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_646
timestamp 1677579658
transform 1 0 62592 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_685
timestamp 1679577901
transform 1 0 66336 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_689
timestamp 1677579658
transform 1 0 66720 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_725
timestamp 1679581782
transform 1 0 70176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_732
timestamp 1679581782
transform 1 0 70848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_764
timestamp 1679581782
transform 1 0 73920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_771
timestamp 1679581782
transform 1 0 74592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_778
timestamp 1679581782
transform 1 0 75264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_785
timestamp 1679577901
transform 1 0 75936 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_789
timestamp 1677579658
transform 1 0 76320 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_822
timestamp 1677579658
transform 1 0 79488 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_4
timestamp 1679577901
transform 1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_8
timestamp 1677579658
transform 1 0 1344 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_13
timestamp 1679581782
transform 1 0 1824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_20
timestamp 1679581782
transform 1 0 2496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_27
timestamp 1679581782
transform 1 0 3168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_34
timestamp 1679581782
transform 1 0 3840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_41
timestamp 1679581782
transform 1 0 4512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_48
timestamp 1679581782
transform 1 0 5184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_55
timestamp 1679581782
transform 1 0 5856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_62
timestamp 1679581782
transform 1 0 6528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_69
timestamp 1679581782
transform 1 0 7200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_76
timestamp 1679581782
transform 1 0 7872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_83
timestamp 1679581782
transform 1 0 8544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_90
timestamp 1679581782
transform 1 0 9216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_97
timestamp 1679581782
transform 1 0 9888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_104
timestamp 1679581782
transform 1 0 10560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_111
timestamp 1679581782
transform 1 0 11232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_118
timestamp 1679581782
transform 1 0 11904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_125
timestamp 1679581782
transform 1 0 12576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_132
timestamp 1679581782
transform 1 0 13248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_139
timestamp 1679581782
transform 1 0 13920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_146
timestamp 1679581782
transform 1 0 14592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_153
timestamp 1679581782
transform 1 0 15264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_160
timestamp 1679581782
transform 1 0 15936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_167
timestamp 1679581782
transform 1 0 16608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_174
timestamp 1679581782
transform 1 0 17280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_181
timestamp 1679581782
transform 1 0 17952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_188
timestamp 1679581782
transform 1 0 18624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_195
timestamp 1679581782
transform 1 0 19296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_202
timestamp 1679581782
transform 1 0 19968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_209
timestamp 1679581782
transform 1 0 20640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_216
timestamp 1679581782
transform 1 0 21312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_223
timestamp 1679581782
transform 1 0 21984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_230
timestamp 1679581782
transform 1 0 22656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_237
timestamp 1679581782
transform 1 0 23328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_244
timestamp 1679581782
transform 1 0 24000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_251
timestamp 1679581782
transform 1 0 24672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_258
timestamp 1679581782
transform 1 0 25344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_265
timestamp 1679581782
transform 1 0 26016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_272
timestamp 1679581782
transform 1 0 26688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_279
timestamp 1679581782
transform 1 0 27360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_286
timestamp 1679581782
transform 1 0 28032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_293
timestamp 1679581782
transform 1 0 28704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_300
timestamp 1679581782
transform 1 0 29376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_307
timestamp 1679581782
transform 1 0 30048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_314
timestamp 1679581782
transform 1 0 30720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_321
timestamp 1679581782
transform 1 0 31392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_328
timestamp 1679581782
transform 1 0 32064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_335
timestamp 1679581782
transform 1 0 32736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_342
timestamp 1679581782
transform 1 0 33408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_349
timestamp 1679581782
transform 1 0 34080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_356
timestamp 1679581782
transform 1 0 34752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_363
timestamp 1679581782
transform 1 0 35424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_370
timestamp 1679581782
transform 1 0 36096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_377
timestamp 1679581782
transform 1 0 36768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_384
timestamp 1679581782
transform 1 0 37440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_391
timestamp 1679581782
transform 1 0 38112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_398
timestamp 1679581782
transform 1 0 38784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_405
timestamp 1679581782
transform 1 0 39456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_412
timestamp 1679581782
transform 1 0 40128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_419
timestamp 1679577901
transform 1 0 40800 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_428
timestamp 1679581782
transform 1 0 41664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_435
timestamp 1679581782
transform 1 0 42336 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_442
timestamp 1677579658
transform 1 0 43008 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_454
timestamp 1677580104
transform 1 0 44160 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_462
timestamp 1679577901
transform 1 0 44928 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_466
timestamp 1677580104
transform 1 0 45312 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_508
timestamp 1677580104
transform 1 0 49344 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_510
timestamp 1677579658
transform 1 0 49536 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_516
timestamp 1679577901
transform 1 0 50112 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_555
timestamp 1679581782
transform 1 0 53856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_562
timestamp 1679577901
transform 1 0 54528 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_566
timestamp 1677580104
transform 1 0 54912 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_586
timestamp 1679581782
transform 1 0 56832 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_593
timestamp 1677579658
transform 1 0 57504 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_651
timestamp 1679577901
transform 1 0 63072 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_655
timestamp 1677579658
transform 1 0 63456 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_659
timestamp 1679577901
transform 1 0 63840 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_663
timestamp 1677579658
transform 1 0 64224 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_691
timestamp 1679581782
transform 1 0 66912 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_698
timestamp 1677580104
transform 1 0 67584 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_705
timestamp 1679581782
transform 1 0 68256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_712
timestamp 1679577901
transform 1 0 68928 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_716
timestamp 1677579658
transform 1 0 69312 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_747
timestamp 1677580104
transform 1 0 72288 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_749
timestamp 1677579658
transform 1 0 72480 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_777
timestamp 1679581782
transform 1 0 75168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_784
timestamp 1679577901
transform 1 0 75840 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_788
timestamp 1677579658
transform 1 0 76224 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_795
timestamp 1677580104
transform 1 0 76896 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_810
timestamp 1679581782
transform 1 0 78336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_817
timestamp 1679577901
transform 1 0 79008 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_821
timestamp 1677580104
transform 1 0 79392 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_4
timestamp 1679577901
transform 1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_8
timestamp 1677579658
transform 1 0 1344 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_13
timestamp 1679581782
transform 1 0 1824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_20
timestamp 1679581782
transform 1 0 2496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_27
timestamp 1679581782
transform 1 0 3168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_34
timestamp 1679581782
transform 1 0 3840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_41
timestamp 1679581782
transform 1 0 4512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_48
timestamp 1679581782
transform 1 0 5184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_55
timestamp 1679581782
transform 1 0 5856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_62
timestamp 1679581782
transform 1 0 6528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_69
timestamp 1679581782
transform 1 0 7200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_76
timestamp 1679581782
transform 1 0 7872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_83
timestamp 1679581782
transform 1 0 8544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_90
timestamp 1679581782
transform 1 0 9216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_97
timestamp 1679581782
transform 1 0 9888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_104
timestamp 1679581782
transform 1 0 10560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_111
timestamp 1679581782
transform 1 0 11232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_118
timestamp 1679581782
transform 1 0 11904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_125
timestamp 1679581782
transform 1 0 12576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_132
timestamp 1679581782
transform 1 0 13248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_139
timestamp 1679581782
transform 1 0 13920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_146
timestamp 1679581782
transform 1 0 14592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_153
timestamp 1679581782
transform 1 0 15264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_160
timestamp 1679581782
transform 1 0 15936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_167
timestamp 1679581782
transform 1 0 16608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_174
timestamp 1679581782
transform 1 0 17280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_181
timestamp 1679581782
transform 1 0 17952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_188
timestamp 1679581782
transform 1 0 18624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_195
timestamp 1679581782
transform 1 0 19296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_202
timestamp 1679581782
transform 1 0 19968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_209
timestamp 1679581782
transform 1 0 20640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_216
timestamp 1679581782
transform 1 0 21312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_223
timestamp 1679581782
transform 1 0 21984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_230
timestamp 1679581782
transform 1 0 22656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_237
timestamp 1679581782
transform 1 0 23328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_244
timestamp 1679581782
transform 1 0 24000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_251
timestamp 1679581782
transform 1 0 24672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_258
timestamp 1679581782
transform 1 0 25344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_265
timestamp 1679581782
transform 1 0 26016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_272
timestamp 1679581782
transform 1 0 26688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_279
timestamp 1679581782
transform 1 0 27360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_286
timestamp 1679581782
transform 1 0 28032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_293
timestamp 1679581782
transform 1 0 28704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_300
timestamp 1679581782
transform 1 0 29376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_307
timestamp 1679581782
transform 1 0 30048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_314
timestamp 1679581782
transform 1 0 30720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_321
timestamp 1679581782
transform 1 0 31392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_328
timestamp 1679581782
transform 1 0 32064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_335
timestamp 1679581782
transform 1 0 32736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_342
timestamp 1679581782
transform 1 0 33408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_349
timestamp 1679581782
transform 1 0 34080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_356
timestamp 1679581782
transform 1 0 34752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_363
timestamp 1679581782
transform 1 0 35424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_370
timestamp 1679581782
transform 1 0 36096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_377
timestamp 1679581782
transform 1 0 36768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_384
timestamp 1679581782
transform 1 0 37440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_391
timestamp 1679577901
transform 1 0 38112 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_395
timestamp 1677580104
transform 1 0 38496 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_451
timestamp 1677579658
transform 1 0 43872 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_484
timestamp 1679577901
transform 1 0 47040 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_488
timestamp 1677580104
transform 1 0 47424 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_493
timestamp 1679581782
transform 1 0 47904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_500
timestamp 1679581782
transform 1 0 48576 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_514
timestamp 1677580104
transform 1 0 49920 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_516
timestamp 1677579658
transform 1 0 50112 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_520
timestamp 1679577901
transform 1 0 50496 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_524
timestamp 1677580104
transform 1 0 50880 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_544
timestamp 1679581782
transform 1 0 52800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_551
timestamp 1679581782
transform 1 0 53472 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_558
timestamp 1677579658
transform 1 0 54144 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_565
timestamp 1677580104
transform 1 0 54816 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_567
timestamp 1677579658
transform 1 0 55008 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_576
timestamp 1677580104
transform 1 0 55872 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_578
timestamp 1677579658
transform 1 0 56064 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_611
timestamp 1679581782
transform 1 0 59232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_628
timestamp 1679577901
transform 1 0 60864 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_632
timestamp 1677580104
transform 1 0 61248 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_652
timestamp 1679581782
transform 1 0 63168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_659
timestamp 1679581782
transform 1 0 63840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_666
timestamp 1679581782
transform 1 0 64512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_699
timestamp 1679577901
transform 1 0 67680 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_706
timestamp 1677580104
transform 1 0 68352 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_747
timestamp 1677580104
transform 1 0 72288 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_749
timestamp 1677579658
transform 1 0 72480 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_755
timestamp 1679581782
transform 1 0 73056 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_762
timestamp 1677579658
transform 1 0 73728 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_800
timestamp 1677579658
transform 1 0 77376 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_806
timestamp 1677580104
transform 1 0 77952 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679581782
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_818
timestamp 1679577901
transform 1 0 79104 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_822
timestamp 1677579658
transform 1 0 79488 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_7
timestamp 1677580104
transform 1 0 1248 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_13
timestamp 1679581782
transform 1 0 1824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_20
timestamp 1679581782
transform 1 0 2496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_27
timestamp 1679581782
transform 1 0 3168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_34
timestamp 1679581782
transform 1 0 3840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_41
timestamp 1679581782
transform 1 0 4512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_48
timestamp 1679581782
transform 1 0 5184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_55
timestamp 1679581782
transform 1 0 5856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_62
timestamp 1679581782
transform 1 0 6528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_69
timestamp 1679581782
transform 1 0 7200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_76
timestamp 1679581782
transform 1 0 7872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_83
timestamp 1679581782
transform 1 0 8544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_90
timestamp 1679581782
transform 1 0 9216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_97
timestamp 1679581782
transform 1 0 9888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_104
timestamp 1679581782
transform 1 0 10560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_111
timestamp 1679581782
transform 1 0 11232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_118
timestamp 1679581782
transform 1 0 11904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_125
timestamp 1679581782
transform 1 0 12576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_132
timestamp 1679581782
transform 1 0 13248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_139
timestamp 1679581782
transform 1 0 13920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_146
timestamp 1679581782
transform 1 0 14592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_153
timestamp 1679581782
transform 1 0 15264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_160
timestamp 1679581782
transform 1 0 15936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_167
timestamp 1679581782
transform 1 0 16608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_174
timestamp 1679581782
transform 1 0 17280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_181
timestamp 1679581782
transform 1 0 17952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_188
timestamp 1679581782
transform 1 0 18624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_195
timestamp 1679581782
transform 1 0 19296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_202
timestamp 1679581782
transform 1 0 19968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_209
timestamp 1679581782
transform 1 0 20640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_216
timestamp 1679581782
transform 1 0 21312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_223
timestamp 1679581782
transform 1 0 21984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_230
timestamp 1679581782
transform 1 0 22656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_237
timestamp 1679581782
transform 1 0 23328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_244
timestamp 1679581782
transform 1 0 24000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_251
timestamp 1679581782
transform 1 0 24672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_258
timestamp 1679581782
transform 1 0 25344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_265
timestamp 1679581782
transform 1 0 26016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_272
timestamp 1679581782
transform 1 0 26688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_279
timestamp 1679581782
transform 1 0 27360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_286
timestamp 1679581782
transform 1 0 28032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_293
timestamp 1679581782
transform 1 0 28704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_300
timestamp 1679581782
transform 1 0 29376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_307
timestamp 1679581782
transform 1 0 30048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_314
timestamp 1679581782
transform 1 0 30720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_321
timestamp 1679581782
transform 1 0 31392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_328
timestamp 1679581782
transform 1 0 32064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_335
timestamp 1679581782
transform 1 0 32736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_342
timestamp 1679581782
transform 1 0 33408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_349
timestamp 1679581782
transform 1 0 34080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_356
timestamp 1679581782
transform 1 0 34752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_363
timestamp 1679581782
transform 1 0 35424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_370
timestamp 1679577901
transform 1 0 36096 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_374
timestamp 1677579658
transform 1 0 36480 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_402
timestamp 1677579658
transform 1 0 39168 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_424
timestamp 1677580104
transform 1 0 41280 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_426
timestamp 1677579658
transform 1 0 41472 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_433
timestamp 1677580104
transform 1 0 42144 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_442
timestamp 1679581782
transform 1 0 43008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_449
timestamp 1679581782
transform 1 0 43680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_456
timestamp 1679577901
transform 1 0 44352 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_485
timestamp 1679581782
transform 1 0 47136 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_492
timestamp 1677580104
transform 1 0 47808 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_527
timestamp 1677580104
transform 1 0 51168 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_529
timestamp 1677579658
transform 1 0 51360 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_584
timestamp 1679581782
transform 1 0 56640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_591
timestamp 1679581782
transform 1 0 57312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_604
timestamp 1679577901
transform 1 0 58560 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_608
timestamp 1677580104
transform 1 0 58944 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_648
timestamp 1677580104
transform 1 0 62784 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_650
timestamp 1677579658
transform 1 0 62976 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_656
timestamp 1679581782
transform 1 0 63552 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_663
timestamp 1677580104
transform 1 0 64224 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_665
timestamp 1677579658
transform 1 0 64416 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_726
timestamp 1677580104
transform 1 0 70272 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_731
timestamp 1677579658
transform 1 0 70752 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_738
timestamp 1679577901
transform 1 0 71424 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_769
timestamp 1679581782
transform 1 0 74400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_776
timestamp 1679577901
transform 1 0 75072 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_780
timestamp 1677580104
transform 1 0 75456 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_822
timestamp 1677579658
transform 1 0 79488 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679581782
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679581782
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679581782
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679581782
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_32
timestamp 1679581782
transform 1 0 3648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_39
timestamp 1679581782
transform 1 0 4320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_46
timestamp 1679581782
transform 1 0 4992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_53
timestamp 1679581782
transform 1 0 5664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_60
timestamp 1679581782
transform 1 0 6336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679581782
transform 1 0 7008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_74
timestamp 1679581782
transform 1 0 7680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_81
timestamp 1679581782
transform 1 0 8352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_88
timestamp 1679581782
transform 1 0 9024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_95
timestamp 1679581782
transform 1 0 9696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_102
timestamp 1679581782
transform 1 0 10368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_109
timestamp 1679581782
transform 1 0 11040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_116
timestamp 1679581782
transform 1 0 11712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_123
timestamp 1679581782
transform 1 0 12384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_130
timestamp 1679581782
transform 1 0 13056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_137
timestamp 1679581782
transform 1 0 13728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_144
timestamp 1679581782
transform 1 0 14400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_151
timestamp 1679581782
transform 1 0 15072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_158
timestamp 1679581782
transform 1 0 15744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_165
timestamp 1679581782
transform 1 0 16416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_172
timestamp 1679581782
transform 1 0 17088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_179
timestamp 1679581782
transform 1 0 17760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_186
timestamp 1679581782
transform 1 0 18432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_193
timestamp 1679581782
transform 1 0 19104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_200
timestamp 1679581782
transform 1 0 19776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_207
timestamp 1679581782
transform 1 0 20448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_214
timestamp 1679581782
transform 1 0 21120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_221
timestamp 1679581782
transform 1 0 21792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_228
timestamp 1679581782
transform 1 0 22464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_235
timestamp 1679581782
transform 1 0 23136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_242
timestamp 1679581782
transform 1 0 23808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_249
timestamp 1679581782
transform 1 0 24480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_256
timestamp 1679581782
transform 1 0 25152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_263
timestamp 1679581782
transform 1 0 25824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_270
timestamp 1679581782
transform 1 0 26496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_277
timestamp 1679581782
transform 1 0 27168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_284
timestamp 1679581782
transform 1 0 27840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_291
timestamp 1679581782
transform 1 0 28512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_298
timestamp 1679581782
transform 1 0 29184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_305
timestamp 1679581782
transform 1 0 29856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_312
timestamp 1679581782
transform 1 0 30528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_319
timestamp 1679581782
transform 1 0 31200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_326
timestamp 1679581782
transform 1 0 31872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_333
timestamp 1679581782
transform 1 0 32544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_340
timestamp 1679581782
transform 1 0 33216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_347
timestamp 1679577901
transform 1 0 33888 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_351
timestamp 1677579658
transform 1 0 34272 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_385
timestamp 1679581782
transform 1 0 37536 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_392
timestamp 1677579658
transform 1 0 38208 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_426
timestamp 1679581782
transform 1 0 41472 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_433
timestamp 1677580104
transform 1 0 42144 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_440
timestamp 1677579658
transform 1 0 42816 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_446
timestamp 1679581782
transform 1 0 43392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_453
timestamp 1679581782
transform 1 0 44064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_460
timestamp 1679577901
transform 1 0 44736 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_464
timestamp 1677580104
transform 1 0 45120 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_498
timestamp 1677580104
transform 1 0 48384 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_500
timestamp 1677579658
transform 1 0 48576 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_553
timestamp 1677580104
transform 1 0 53664 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_563
timestamp 1679577901
transform 1 0 54624 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_579
timestamp 1679581782
transform 1 0 56160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_586
timestamp 1679581782
transform 1 0 56832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_593
timestamp 1679581782
transform 1 0 57504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_611
timestamp 1679581782
transform 1 0 59232 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_618
timestamp 1677580104
transform 1 0 59904 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_624
timestamp 1679577901
transform 1 0 60480 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_628
timestamp 1677579658
transform 1 0 60864 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_636
timestamp 1677580104
transform 1 0 61632 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_642
timestamp 1677579658
transform 1 0 62208 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_680
timestamp 1679581782
transform 1 0 65856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_687
timestamp 1679577901
transform 1 0 66528 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_691
timestamp 1677580104
transform 1 0 66912 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_700
timestamp 1679577901
transform 1 0 67776 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_704
timestamp 1677580104
transform 1 0 68160 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_719
timestamp 1679577901
transform 1 0 69600 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_739
timestamp 1677580104
transform 1 0 71520 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_746
timestamp 1679581782
transform 1 0 72192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_753
timestamp 1679577901
transform 1 0 72864 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_757
timestamp 1677579658
transform 1 0 73248 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_762
timestamp 1679581782
transform 1 0 73728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_769
timestamp 1679581782
transform 1 0 74400 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_776
timestamp 1677579658
transform 1 0 75072 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_783
timestamp 1677579658
transform 1 0 75744 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_789
timestamp 1677580104
transform 1 0 76320 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_791
timestamp 1677579658
transform 1 0 76512 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_797
timestamp 1679581782
transform 1 0 77088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_804
timestamp 1679581782
transform 1 0 77760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_811
timestamp 1679581782
transform 1 0 78432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_818
timestamp 1679577901
transform 1 0 79104 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_822
timestamp 1677579658
transform 1 0 79488 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_4
timestamp 1679577901
transform 1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_8
timestamp 1677579658
transform 1 0 1344 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_13
timestamp 1679581782
transform 1 0 1824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_20
timestamp 1679581782
transform 1 0 2496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_27
timestamp 1679581782
transform 1 0 3168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_34
timestamp 1679581782
transform 1 0 3840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_41
timestamp 1679581782
transform 1 0 4512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_48
timestamp 1679581782
transform 1 0 5184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_55
timestamp 1679581782
transform 1 0 5856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_62
timestamp 1679581782
transform 1 0 6528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_69
timestamp 1679581782
transform 1 0 7200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_76
timestamp 1679581782
transform 1 0 7872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_83
timestamp 1679581782
transform 1 0 8544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_90
timestamp 1679581782
transform 1 0 9216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_97
timestamp 1679581782
transform 1 0 9888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_104
timestamp 1679581782
transform 1 0 10560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_111
timestamp 1679581782
transform 1 0 11232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_118
timestamp 1679581782
transform 1 0 11904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_125
timestamp 1679581782
transform 1 0 12576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_132
timestamp 1679581782
transform 1 0 13248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_139
timestamp 1679581782
transform 1 0 13920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_146
timestamp 1679581782
transform 1 0 14592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_153
timestamp 1679581782
transform 1 0 15264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_160
timestamp 1679581782
transform 1 0 15936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_167
timestamp 1679581782
transform 1 0 16608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_174
timestamp 1679581782
transform 1 0 17280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_181
timestamp 1679581782
transform 1 0 17952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_188
timestamp 1679581782
transform 1 0 18624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_195
timestamp 1679581782
transform 1 0 19296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_202
timestamp 1679581782
transform 1 0 19968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_209
timestamp 1679581782
transform 1 0 20640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_216
timestamp 1679581782
transform 1 0 21312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_223
timestamp 1679581782
transform 1 0 21984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_230
timestamp 1679581782
transform 1 0 22656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_237
timestamp 1679581782
transform 1 0 23328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_244
timestamp 1679581782
transform 1 0 24000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_251
timestamp 1679581782
transform 1 0 24672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_258
timestamp 1679581782
transform 1 0 25344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_265
timestamp 1679581782
transform 1 0 26016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_272
timestamp 1679577901
transform 1 0 26688 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_276
timestamp 1677580104
transform 1 0 27072 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_288
timestamp 1679581782
transform 1 0 28224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_295
timestamp 1679581782
transform 1 0 28896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_302
timestamp 1679581782
transform 1 0 29568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_309
timestamp 1679581782
transform 1 0 30240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_316
timestamp 1679581782
transform 1 0 30912 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_361
timestamp 1677580104
transform 1 0 35232 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_373
timestamp 1677580104
transform 1 0 36384 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_380
timestamp 1679577901
transform 1 0 37056 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_384
timestamp 1677580104
transform 1 0 37440 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_398
timestamp 1679581782
transform 1 0 38784 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_464
timestamp 1677580104
transform 1 0 45120 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_466
timestamp 1677579658
transform 1 0 45312 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_494
timestamp 1679581782
transform 1 0 48000 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_501
timestamp 1677580104
transform 1 0 48672 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_503
timestamp 1677579658
transform 1 0 48864 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_509
timestamp 1677580104
transform 1 0 49440 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_516
timestamp 1679581782
transform 1 0 50112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_523
timestamp 1679581782
transform 1 0 50784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_530
timestamp 1679581782
transform 1 0 51456 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_537
timestamp 1677579658
transform 1 0 52128 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_543
timestamp 1677579658
transform 1 0 52704 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_569
timestamp 1677579658
transform 1 0 55200 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_624
timestamp 1679577901
transform 1 0 60480 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_646
timestamp 1679581782
transform 1 0 62592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_653
timestamp 1679581782
transform 1 0 63264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_660
timestamp 1679581782
transform 1 0 63936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_667
timestamp 1679577901
transform 1 0 64608 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_675
timestamp 1679581782
transform 1 0 65376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_682
timestamp 1679581782
transform 1 0 66048 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_689
timestamp 1677579658
transform 1 0 66720 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_695
timestamp 1677579658
transform 1 0 67296 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_699
timestamp 1677580104
transform 1 0 67680 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_709
timestamp 1679581782
transform 1 0 68640 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_716
timestamp 1677579658
transform 1 0 69312 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_787
timestamp 1677580104
transform 1 0 76128 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_816
timestamp 1679581782
transform 1 0 78912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_4
timestamp 1679577901
transform 1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_8
timestamp 1677579658
transform 1 0 1344 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_13
timestamp 1679581782
transform 1 0 1824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_20
timestamp 1679581782
transform 1 0 2496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_27
timestamp 1679581782
transform 1 0 3168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_34
timestamp 1679581782
transform 1 0 3840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_41
timestamp 1679581782
transform 1 0 4512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_48
timestamp 1679581782
transform 1 0 5184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_55
timestamp 1679577901
transform 1 0 5856 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_64
timestamp 1677579658
transform 1 0 6720 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_68
timestamp 1679581782
transform 1 0 7104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_75
timestamp 1679581782
transform 1 0 7776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_82
timestamp 1679581782
transform 1 0 8448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_89
timestamp 1679581782
transform 1 0 9120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_96
timestamp 1679577901
transform 1 0 9792 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_100
timestamp 1677579658
transform 1 0 10176 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_105
timestamp 1679581782
transform 1 0 10656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_112
timestamp 1679581782
transform 1 0 11328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_119
timestamp 1679581782
transform 1 0 12000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_126
timestamp 1679581782
transform 1 0 12672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_133
timestamp 1679581782
transform 1 0 13344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_140
timestamp 1679581782
transform 1 0 14016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_147
timestamp 1679581782
transform 1 0 14688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_154
timestamp 1679581782
transform 1 0 15360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_161
timestamp 1679581782
transform 1 0 16032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_168
timestamp 1679581782
transform 1 0 16704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_175
timestamp 1679581782
transform 1 0 17376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_182
timestamp 1679581782
transform 1 0 18048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_189
timestamp 1679581782
transform 1 0 18720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_196
timestamp 1679581782
transform 1 0 19392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_203
timestamp 1679581782
transform 1 0 20064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_210
timestamp 1679581782
transform 1 0 20736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_217
timestamp 1679581782
transform 1 0 21408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_224
timestamp 1679581782
transform 1 0 22080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_231
timestamp 1679581782
transform 1 0 22752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_238
timestamp 1679581782
transform 1 0 23424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_245
timestamp 1679581782
transform 1 0 24096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1679581782
transform 1 0 24768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_259
timestamp 1679581782
transform 1 0 25440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679581782
transform 1 0 26112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_273
timestamp 1679577901
transform 1 0 26784 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_277
timestamp 1677579658
transform 1 0 27168 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_291
timestamp 1679577901
transform 1 0 28512 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_295
timestamp 1677579658
transform 1 0 28896 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_309
timestamp 1679581782
transform 1 0 30240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_316
timestamp 1679581782
transform 1 0 30912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_323
timestamp 1679577901
transform 1 0 31584 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_333
timestamp 1677580104
transform 1 0 32544 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_340
timestamp 1677579658
transform 1 0 33216 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_344
timestamp 1679581782
transform 1 0 33600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_351
timestamp 1679581782
transform 1 0 34272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_358
timestamp 1679577901
transform 1 0 34944 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_362
timestamp 1677579658
transform 1 0 35328 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_368
timestamp 1677579658
transform 1 0 35904 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_374
timestamp 1677580104
transform 1 0 36480 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_379
timestamp 1679577901
transform 1 0 36960 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_383
timestamp 1677580104
transform 1 0 37344 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_417
timestamp 1679577901
transform 1 0 40608 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_424
timestamp 1679581782
transform 1 0 41280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_431
timestamp 1679581782
transform 1 0 41952 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_438
timestamp 1677579658
transform 1 0 42624 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_469
timestamp 1677580104
transform 1 0 45600 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_505
timestamp 1679577901
transform 1 0 49056 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_509
timestamp 1677579658
transform 1 0 49440 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_528
timestamp 1679581782
transform 1 0 51264 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_535
timestamp 1677580104
transform 1 0 51936 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_572
timestamp 1677580104
transform 1 0 55488 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_574
timestamp 1677579658
transform 1 0 55680 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_582
timestamp 1677579658
transform 1 0 56448 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_592
timestamp 1679577901
transform 1 0 57408 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_596
timestamp 1677580104
transform 1 0 57792 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_603
timestamp 1677579658
transform 1 0 58464 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_616
timestamp 1677580104
transform 1 0 59712 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_618
timestamp 1677579658
transform 1 0 59904 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_622
timestamp 1677579658
transform 1 0 60288 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_657
timestamp 1677579658
transform 1 0 63648 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_661
timestamp 1679581782
transform 1 0 64032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_668
timestamp 1679581782
transform 1 0 64704 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_675
timestamp 1677580104
transform 1 0 65376 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_680
timestamp 1677579658
transform 1 0 65856 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_717
timestamp 1677579658
transform 1 0 69408 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_736
timestamp 1679577901
transform 1 0 71232 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_743
timestamp 1677580104
transform 1 0 71904 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_751
timestamp 1679577901
transform 1 0 72672 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_755
timestamp 1677580104
transform 1 0 73056 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_760
timestamp 1679577901
transform 1 0 73536 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_764
timestamp 1677579658
transform 1 0 73920 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_768
timestamp 1679581782
transform 1 0 74304 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_775
timestamp 1677580104
transform 1 0 74976 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_777
timestamp 1677579658
transform 1 0 75168 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_792
timestamp 1679581782
transform 1 0 76608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_799
timestamp 1679577901
transform 1 0 77280 0 1 15876
box -48 -56 432 834
use sg13g2_decap_4  FILLER_20_806
timestamp 1679577901
transform 1 0 77952 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_810
timestamp 1677579658
transform 1 0 78336 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_814
timestamp 1679577901
transform 1 0 78720 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_818
timestamp 1677580104
transform 1 0 79104 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_8
timestamp 1679581782
transform 1 0 1344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_15
timestamp 1679577901
transform 1 0 2016 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_23
timestamp 1679581782
transform 1 0 2784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_30
timestamp 1679581782
transform 1 0 3456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_37
timestamp 1679581782
transform 1 0 4128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_44
timestamp 1679581782
transform 1 0 4800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_51
timestamp 1679577901
transform 1 0 5472 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_55
timestamp 1677579658
transform 1 0 5856 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_94
timestamp 1677579658
transform 1 0 9600 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_100
timestamp 1677579658
transform 1 0 10176 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_110
timestamp 1679581782
transform 1 0 11136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_117
timestamp 1679581782
transform 1 0 11808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_124
timestamp 1679581782
transform 1 0 12480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_131
timestamp 1679581782
transform 1 0 13152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_138
timestamp 1679581782
transform 1 0 13824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_145
timestamp 1679581782
transform 1 0 14496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_152
timestamp 1679581782
transform 1 0 15168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_159
timestamp 1679581782
transform 1 0 15840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_166
timestamp 1679581782
transform 1 0 16512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_173
timestamp 1679581782
transform 1 0 17184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_180
timestamp 1679581782
transform 1 0 17856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_187
timestamp 1679581782
transform 1 0 18528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_194
timestamp 1679581782
transform 1 0 19200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_201
timestamp 1679581782
transform 1 0 19872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_208
timestamp 1679581782
transform 1 0 20544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_215
timestamp 1679581782
transform 1 0 21216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_222
timestamp 1679581782
transform 1 0 21888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_229
timestamp 1679581782
transform 1 0 22560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_236
timestamp 1679581782
transform 1 0 23232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_243
timestamp 1679581782
transform 1 0 23904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_250
timestamp 1679581782
transform 1 0 24576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_257
timestamp 1679581782
transform 1 0 25248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_264
timestamp 1679581782
transform 1 0 25920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_271
timestamp 1679581782
transform 1 0 26592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_278
timestamp 1679581782
transform 1 0 27264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_285
timestamp 1679581782
transform 1 0 27936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_292
timestamp 1679577901
transform 1 0 28608 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_321
timestamp 1679581782
transform 1 0 31392 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_328
timestamp 1677579658
transform 1 0 32064 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_363
timestamp 1677579658
transform 1 0 35424 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_391
timestamp 1679581782
transform 1 0 38112 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_398
timestamp 1677580104
transform 1 0 38784 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_403
timestamp 1679581782
transform 1 0 39264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_410
timestamp 1679577901
transform 1 0 39936 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_414
timestamp 1677579658
transform 1 0 40320 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_425
timestamp 1679581782
transform 1 0 41376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_432
timestamp 1679581782
transform 1 0 42048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_439
timestamp 1679577901
transform 1 0 42720 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_443
timestamp 1677579658
transform 1 0 43104 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_450
timestamp 1677580104
transform 1 0 43776 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_452
timestamp 1677579658
transform 1 0 43968 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_458
timestamp 1679581782
transform 1 0 44544 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_465
timestamp 1677580104
transform 1 0 45216 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_484
timestamp 1677580104
transform 1 0 47040 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_489
timestamp 1677579658
transform 1 0 47520 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_4
timestamp 1677579658
transform 1 0 960 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_13
timestamp 1679581782
transform 1 0 1824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_20
timestamp 1679581782
transform 1 0 2496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_27
timestamp 1679577901
transform 1 0 3168 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_31
timestamp 1677579658
transform 1 0 3552 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_62
timestamp 1677579658
transform 1 0 6528 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_95
timestamp 1677579658
transform 1 0 9696 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_138
timestamp 1679581782
transform 1 0 13824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_145
timestamp 1679581782
transform 1 0 14496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_152
timestamp 1679581782
transform 1 0 15168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_159
timestamp 1679581782
transform 1 0 15840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_166
timestamp 1679581782
transform 1 0 16512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_173
timestamp 1679581782
transform 1 0 17184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_180
timestamp 1679581782
transform 1 0 17856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_187
timestamp 1679581782
transform 1 0 18528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_194
timestamp 1679581782
transform 1 0 19200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_201
timestamp 1679581782
transform 1 0 19872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_208
timestamp 1679581782
transform 1 0 20544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_215
timestamp 1679581782
transform 1 0 21216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_222
timestamp 1679581782
transform 1 0 21888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_229
timestamp 1679581782
transform 1 0 22560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_236
timestamp 1679581782
transform 1 0 23232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_243
timestamp 1679581782
transform 1 0 23904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_250
timestamp 1679581782
transform 1 0 24576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_257
timestamp 1679581782
transform 1 0 25248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_264
timestamp 1679581782
transform 1 0 25920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_271
timestamp 1679581782
transform 1 0 26592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_278
timestamp 1679581782
transform 1 0 27264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_285
timestamp 1679581782
transform 1 0 27936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_292
timestamp 1679581782
transform 1 0 28608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_299
timestamp 1679581782
transform 1 0 29280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_306
timestamp 1679581782
transform 1 0 29952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_313
timestamp 1679581782
transform 1 0 30624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_320
timestamp 1679577901
transform 1 0 31296 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_346
timestamp 1679581782
transform 1 0 33792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_353
timestamp 1679581782
transform 1 0 34464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_360
timestamp 1679581782
transform 1 0 35136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_367
timestamp 1679581782
transform 1 0 35808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_374
timestamp 1679581782
transform 1 0 36480 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_381
timestamp 1677580104
transform 1 0 37152 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_388
timestamp 1677580104
transform 1 0 37824 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_390
timestamp 1677579658
transform 1 0 38016 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_394
timestamp 1679581782
transform 1 0 38400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_401
timestamp 1679577901
transform 1 0 39072 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_405
timestamp 1677580104
transform 1 0 39456 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_465
timestamp 1679581782
transform 1 0 45216 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_472
timestamp 1677580104
transform 1 0 45888 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_479
timestamp 1679581782
transform 1 0 46560 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_486
timestamp 1677579658
transform 1 0 47232 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_490
timestamp 1679581782
transform 1 0 47616 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_497
timestamp 1677580104
transform 1 0 48288 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_517
timestamp 1677580104
transform 1 0 50208 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_530
timestamp 1679581782
transform 1 0 51456 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_537
timestamp 1677579658
transform 1 0 52128 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_4
timestamp 1677579658
transform 1 0 960 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_13
timestamp 1679581782
transform 1 0 1824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_20
timestamp 1679581782
transform 1 0 2496 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_27
timestamp 1677580104
transform 1 0 3168 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_51
timestamp 1679581782
transform 1 0 5472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_58
timestamp 1679577901
transform 1 0 6144 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_66
timestamp 1677580104
transform 1 0 6912 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_68
timestamp 1677579658
transform 1 0 7104 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_101
timestamp 1677580104
transform 1 0 10272 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_103
timestamp 1677579658
transform 1 0 10464 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679581782
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_116
timestamp 1677580104
transform 1 0 11712 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_118
timestamp 1677579658
transform 1 0 11904 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_184
timestamp 1679581782
transform 1 0 18240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_191
timestamp 1679581782
transform 1 0 18912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_198
timestamp 1679581782
transform 1 0 19584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_205
timestamp 1679581782
transform 1 0 20256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_212
timestamp 1679581782
transform 1 0 20928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_219
timestamp 1679581782
transform 1 0 21600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_226
timestamp 1679581782
transform 1 0 22272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_233
timestamp 1679581782
transform 1 0 22944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_240
timestamp 1679581782
transform 1 0 23616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_247
timestamp 1679581782
transform 1 0 24288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_254
timestamp 1679581782
transform 1 0 24960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_261
timestamp 1679581782
transform 1 0 25632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_268
timestamp 1679581782
transform 1 0 26304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_275
timestamp 1679581782
transform 1 0 26976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_282
timestamp 1679581782
transform 1 0 27648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_289
timestamp 1679581782
transform 1 0 28320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_296
timestamp 1679581782
transform 1 0 28992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_303
timestamp 1679577901
transform 1 0 29664 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_307
timestamp 1677579658
transform 1 0 30048 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_357
timestamp 1679581782
transform 1 0 34848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_364
timestamp 1679581782
transform 1 0 35520 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_371
timestamp 1677580104
transform 1 0 36192 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_503
timestamp 1677580104
transform 1 0 48864 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_522
timestamp 1677580104
transform 1 0 50688 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679581782
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_543
timestamp 1677579658
transform 1 0 52704 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_4
timestamp 1677580104
transform 1 0 960 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_18
timestamp 1679577901
transform 1 0 2304 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_22
timestamp 1677580104
transform 1 0 2688 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_33
timestamp 1677579658
transform 1 0 3744 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_43
timestamp 1679581782
transform 1 0 4704 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_50
timestamp 1677580104
transform 1 0 5376 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_52
timestamp 1677579658
transform 1 0 5568 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_57
timestamp 1677580104
transform 1 0 6048 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679581782
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_112
timestamp 1679581782
transform 1 0 11328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_119
timestamp 1679577901
transform 1 0 12000 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_135
timestamp 1679581782
transform 1 0 13536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_142
timestamp 1679581782
transform 1 0 14208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_149
timestamp 1679581782
transform 1 0 14880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_156
timestamp 1679581782
transform 1 0 15552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_163
timestamp 1679581782
transform 1 0 16224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_170
timestamp 1679581782
transform 1 0 16896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_177
timestamp 1679581782
transform 1 0 17568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_184
timestamp 1679581782
transform 1 0 18240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_191
timestamp 1679581782
transform 1 0 18912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_198
timestamp 1679581782
transform 1 0 19584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_205
timestamp 1679581782
transform 1 0 20256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_212
timestamp 1679581782
transform 1 0 20928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_219
timestamp 1679581782
transform 1 0 21600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_226
timestamp 1679581782
transform 1 0 22272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_233
timestamp 1679581782
transform 1 0 22944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_240
timestamp 1679581782
transform 1 0 23616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_247
timestamp 1679581782
transform 1 0 24288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_254
timestamp 1679581782
transform 1 0 24960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_261
timestamp 1679581782
transform 1 0 25632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_268
timestamp 1679581782
transform 1 0 26304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_275
timestamp 1679581782
transform 1 0 26976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_282
timestamp 1679581782
transform 1 0 27648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_289
timestamp 1679581782
transform 1 0 28320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_296
timestamp 1679581782
transform 1 0 28992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_303
timestamp 1679581782
transform 1 0 29664 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_310
timestamp 1677580104
transform 1 0 30336 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_312
timestamp 1677579658
transform 1 0 30528 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_317
timestamp 1679577901
transform 1 0 31008 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_321
timestamp 1677579658
transform 1 0 31392 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_325
timestamp 1679577901
transform 1 0 31776 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_329
timestamp 1677580104
transform 1 0 32160 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_342
timestamp 1677579658
transform 1 0 33408 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_370
timestamp 1677579658
transform 1 0 36096 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_387
timestamp 1677580104
transform 1 0 37728 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_389
timestamp 1677579658
transform 1 0 37920 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_395
timestamp 1677579658
transform 1 0 38496 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_457
timestamp 1679577901
transform 1 0 44448 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_461
timestamp 1677580104
transform 1 0 44832 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_473
timestamp 1677579658
transform 1 0 45984 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_490
timestamp 1677579658
transform 1 0 47616 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_515
timestamp 1677580104
transform 1 0 50016 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_0
timestamp 1677579658
transform 1 0 576 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_44
timestamp 1679577901
transform 1 0 4800 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_85
timestamp 1679577901
transform 1 0 8736 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_89
timestamp 1677579658
transform 1 0 9120 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_117
timestamp 1679581782
transform 1 0 11808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_124
timestamp 1679581782
transform 1 0 12480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_131
timestamp 1679581782
transform 1 0 13152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_138
timestamp 1679581782
transform 1 0 13824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_145
timestamp 1679581782
transform 1 0 14496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_152
timestamp 1679581782
transform 1 0 15168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_159
timestamp 1679581782
transform 1 0 15840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_166
timestamp 1679581782
transform 1 0 16512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_173
timestamp 1679581782
transform 1 0 17184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_180
timestamp 1679581782
transform 1 0 17856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_187
timestamp 1679581782
transform 1 0 18528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_194
timestamp 1679581782
transform 1 0 19200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_201
timestamp 1679581782
transform 1 0 19872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_208
timestamp 1679581782
transform 1 0 20544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_215
timestamp 1679581782
transform 1 0 21216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_222
timestamp 1679581782
transform 1 0 21888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_229
timestamp 1679581782
transform 1 0 22560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_236
timestamp 1679581782
transform 1 0 23232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_243
timestamp 1679581782
transform 1 0 23904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_250
timestamp 1679581782
transform 1 0 24576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_257
timestamp 1679581782
transform 1 0 25248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_264
timestamp 1679581782
transform 1 0 25920 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_271
timestamp 1677580104
transform 1 0 26592 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_273
timestamp 1677579658
transform 1 0 26784 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_293
timestamp 1679581782
transform 1 0 28704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_300
timestamp 1679581782
transform 1 0 29376 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_307
timestamp 1677580104
transform 1 0 30048 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_325
timestamp 1677579658
transform 1 0 31776 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_330
timestamp 1679581782
transform 1 0 32256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_349
timestamp 1679577901
transform 1 0 34080 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_380
timestamp 1677580104
transform 1 0 37056 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_382
timestamp 1677579658
transform 1 0 37248 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_410
timestamp 1677579658
transform 1 0 39936 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_437
timestamp 1677580104
transform 1 0 42528 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_25_493
timestamp 1679577901
transform 1 0 47904 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_536
timestamp 1679581782
transform 1 0 52032 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_543
timestamp 1677579658
transform 1 0 52704 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_4
timestamp 1677580104
transform 1 0 960 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_6
timestamp 1677579658
transform 1 0 1152 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_18
timestamp 1679577901
transform 1 0 2304 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_68
timestamp 1677580104
transform 1 0 7104 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_70
timestamp 1677579658
transform 1 0 7296 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_84
timestamp 1679581782
transform 1 0 8640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_91
timestamp 1679577901
transform 1 0 9312 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_104
timestamp 1677580104
transform 1 0 10560 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_111
timestamp 1679581782
transform 1 0 11232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_118
timestamp 1679581782
transform 1 0 11904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_125
timestamp 1679581782
transform 1 0 12576 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_132
timestamp 1677579658
transform 1 0 13248 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679581782
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679581782
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679581782
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679581782
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679581782
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_256
timestamp 1679581782
transform 1 0 25152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_263
timestamp 1679581782
transform 1 0 25824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_270
timestamp 1679581782
transform 1 0 26496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679581782
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679581782
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679581782
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_298
timestamp 1677580104
transform 1 0 29184 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_342
timestamp 1679581782
transform 1 0 33408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_349
timestamp 1679581782
transform 1 0 34080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_356
timestamp 1679577901
transform 1 0 34752 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_369
timestamp 1679581782
transform 1 0 36000 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_381
timestamp 1677580104
transform 1 0 37152 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_387
timestamp 1679581782
transform 1 0 37728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_394
timestamp 1679581782
transform 1 0 38400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_401
timestamp 1679581782
transform 1 0 39072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_442
timestamp 1679577901
transform 1 0 43008 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_446
timestamp 1677580104
transform 1 0 43392 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679581782
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679581782
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679581782
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_473
timestamp 1679577901
transform 1 0 45984 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_477
timestamp 1677580104
transform 1 0 46368 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_483
timestamp 1677579658
transform 1 0 46944 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679581782
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679581782
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_501
timestamp 1677579658
transform 1 0 48672 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_508
timestamp 1677579658
transform 1 0 49344 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_524
timestamp 1679581782
transform 1 0 50880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_531
timestamp 1679577901
transform 1 0 51552 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_535
timestamp 1677580104
transform 1 0 51936 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_543
timestamp 1677579658
transform 1 0 52704 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_37
timestamp 1677580104
transform 1 0 4128 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_39
timestamp 1677579658
transform 1 0 4320 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_72
timestamp 1677580104
transform 1 0 7488 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_101
timestamp 1679581782
transform 1 0 10272 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_108
timestamp 1677580104
transform 1 0 10944 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_137
timestamp 1679581782
transform 1 0 13728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_144
timestamp 1679581782
transform 1 0 14400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_151
timestamp 1679581782
transform 1 0 15072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_158
timestamp 1679581782
transform 1 0 15744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_165
timestamp 1679581782
transform 1 0 16416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_172
timestamp 1679581782
transform 1 0 17088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_179
timestamp 1679581782
transform 1 0 17760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_186
timestamp 1679581782
transform 1 0 18432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_193
timestamp 1679581782
transform 1 0 19104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_200
timestamp 1679581782
transform 1 0 19776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_207
timestamp 1679581782
transform 1 0 20448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_214
timestamp 1679581782
transform 1 0 21120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_221
timestamp 1679581782
transform 1 0 21792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_228
timestamp 1679581782
transform 1 0 22464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_235
timestamp 1679581782
transform 1 0 23136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_242
timestamp 1679581782
transform 1 0 23808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_249
timestamp 1679581782
transform 1 0 24480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_256
timestamp 1679581782
transform 1 0 25152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_263
timestamp 1679581782
transform 1 0 25824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_270
timestamp 1679581782
transform 1 0 26496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_277
timestamp 1679581782
transform 1 0 27168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_284
timestamp 1679581782
transform 1 0 27840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_291
timestamp 1679581782
transform 1 0 28512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_298
timestamp 1679577901
transform 1 0 29184 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_302
timestamp 1677579658
transform 1 0 29568 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_376
timestamp 1677580104
transform 1 0 36672 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_415
timestamp 1679581782
transform 1 0 40416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_422
timestamp 1679581782
transform 1 0 41088 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_429
timestamp 1677580104
transform 1 0 41760 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_431
timestamp 1677579658
transform 1 0 41952 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_464
timestamp 1679581782
transform 1 0 45120 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_485
timestamp 1677580104
transform 1 0 47136 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_524
timestamp 1677580104
transform 1 0 50880 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_529
timestamp 1677579658
transform 1 0 51360 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_536
timestamp 1677579658
transform 1 0 52032 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_543
timestamp 1677579658
transform 1 0 52704 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_67
timestamp 1679577901
transform 1 0 7008 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679581782
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679581782
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679581782
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679581782
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679581782
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679581782
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_144
timestamp 1679581782
transform 1 0 14400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_151
timestamp 1679581782
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_158
timestamp 1679581782
transform 1 0 15744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_165
timestamp 1679581782
transform 1 0 16416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_172
timestamp 1679581782
transform 1 0 17088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_179
timestamp 1679581782
transform 1 0 17760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_186
timestamp 1679581782
transform 1 0 18432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_193
timestamp 1679581782
transform 1 0 19104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_200
timestamp 1679581782
transform 1 0 19776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_207
timestamp 1679581782
transform 1 0 20448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_214
timestamp 1679581782
transform 1 0 21120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_221
timestamp 1679581782
transform 1 0 21792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_228
timestamp 1679581782
transform 1 0 22464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_235
timestamp 1679581782
transform 1 0 23136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_242
timestamp 1679581782
transform 1 0 23808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_249
timestamp 1679581782
transform 1 0 24480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_256
timestamp 1679581782
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_263
timestamp 1679581782
transform 1 0 25824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_270
timestamp 1679581782
transform 1 0 26496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_277
timestamp 1679581782
transform 1 0 27168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_284
timestamp 1679581782
transform 1 0 27840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_291
timestamp 1679581782
transform 1 0 28512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_298
timestamp 1679581782
transform 1 0 29184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_305
timestamp 1679581782
transform 1 0 29856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_312
timestamp 1679577901
transform 1 0 30528 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_316
timestamp 1677579658
transform 1 0 30912 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_326
timestamp 1677579658
transform 1 0 31872 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_331
timestamp 1679581782
transform 1 0 32352 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_338
timestamp 1677580104
transform 1 0 33024 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_344
timestamp 1679581782
transform 1 0 33600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_351
timestamp 1679581782
transform 1 0 34272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_358
timestamp 1679577901
transform 1 0 34944 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_362
timestamp 1677579658
transform 1 0 35328 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_374
timestamp 1679577901
transform 1 0 36480 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_389
timestamp 1679581782
transform 1 0 37920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_396
timestamp 1679581782
transform 1 0 38592 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_403
timestamp 1677579658
transform 1 0 39264 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_407
timestamp 1679581782
transform 1 0 39648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_414
timestamp 1679581782
transform 1 0 40320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_421
timestamp 1679577901
transform 1 0 40992 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_438
timestamp 1677580104
transform 1 0 42624 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_448
timestamp 1677580104
transform 1 0 43584 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_492
timestamp 1679581782
transform 1 0 47808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_499
timestamp 1679581782
transform 1 0 48480 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_506
timestamp 1677579658
transform 1 0 49152 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_4
timestamp 1679577901
transform 1 0 960 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_8
timestamp 1677579658
transform 1 0 1344 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_13
timestamp 1679581782
transform 1 0 1824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_20
timestamp 1679581782
transform 1 0 2496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_27
timestamp 1679581782
transform 1 0 3168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_34
timestamp 1679581782
transform 1 0 3840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_41
timestamp 1679581782
transform 1 0 4512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_48
timestamp 1679581782
transform 1 0 5184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_55
timestamp 1679581782
transform 1 0 5856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_62
timestamp 1679581782
transform 1 0 6528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_69
timestamp 1679581782
transform 1 0 7200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_76
timestamp 1679581782
transform 1 0 7872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_83
timestamp 1679581782
transform 1 0 8544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_90
timestamp 1679581782
transform 1 0 9216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_97
timestamp 1679581782
transform 1 0 9888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_104
timestamp 1679581782
transform 1 0 10560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_111
timestamp 1679581782
transform 1 0 11232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_118
timestamp 1679581782
transform 1 0 11904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_125
timestamp 1679581782
transform 1 0 12576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_132
timestamp 1679581782
transform 1 0 13248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_139
timestamp 1679581782
transform 1 0 13920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_146
timestamp 1679581782
transform 1 0 14592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_153
timestamp 1679581782
transform 1 0 15264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_160
timestamp 1679581782
transform 1 0 15936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_167
timestamp 1679581782
transform 1 0 16608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_174
timestamp 1679581782
transform 1 0 17280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_181
timestamp 1679581782
transform 1 0 17952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_188
timestamp 1679581782
transform 1 0 18624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_195
timestamp 1679581782
transform 1 0 19296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_202
timestamp 1679581782
transform 1 0 19968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_209
timestamp 1679581782
transform 1 0 20640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_216
timestamp 1679581782
transform 1 0 21312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_223
timestamp 1679581782
transform 1 0 21984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_230
timestamp 1679581782
transform 1 0 22656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_237
timestamp 1679581782
transform 1 0 23328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_244
timestamp 1679581782
transform 1 0 24000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_251
timestamp 1679581782
transform 1 0 24672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_258
timestamp 1679581782
transform 1 0 25344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_265
timestamp 1679581782
transform 1 0 26016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_272
timestamp 1679581782
transform 1 0 26688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_279
timestamp 1679581782
transform 1 0 27360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_286
timestamp 1679581782
transform 1 0 28032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_293
timestamp 1679581782
transform 1 0 28704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_300
timestamp 1679581782
transform 1 0 29376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_307
timestamp 1679581782
transform 1 0 30048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_314
timestamp 1679581782
transform 1 0 30720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_321
timestamp 1679581782
transform 1 0 31392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_328
timestamp 1679581782
transform 1 0 32064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_335
timestamp 1679581782
transform 1 0 32736 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_342
timestamp 1677580104
transform 1 0 33408 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_344
timestamp 1677579658
transform 1 0 33600 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_382
timestamp 1677579658
transform 1 0 37248 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_448
timestamp 1677580104
transform 1 0 43584 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_455
timestamp 1679577901
transform 1 0 44256 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_459
timestamp 1677580104
transform 1 0 44640 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_464
timestamp 1679581782
transform 1 0 45120 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_471
timestamp 1677579658
transform 1 0 45792 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_504
timestamp 1677580104
transform 1 0 48960 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_509
timestamp 1677580104
transform 1 0 49440 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_525
timestamp 1677580104
transform 1 0 50976 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_527
timestamp 1677579658
transform 1 0 51168 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_532
timestamp 1677580104
transform 1 0 51648 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_534
timestamp 1677579658
transform 1 0 51840 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_4
timestamp 1679577901
transform 1 0 960 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_8
timestamp 1677580104
transform 1 0 1344 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_18
timestamp 1679581782
transform 1 0 2304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_25
timestamp 1679581782
transform 1 0 2976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_32
timestamp 1679581782
transform 1 0 3648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_39
timestamp 1679581782
transform 1 0 4320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_46
timestamp 1679581782
transform 1 0 4992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_53
timestamp 1679581782
transform 1 0 5664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_60
timestamp 1679581782
transform 1 0 6336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_67
timestamp 1679581782
transform 1 0 7008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_74
timestamp 1679581782
transform 1 0 7680 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_81
timestamp 1679581782
transform 1 0 8352 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_88
timestamp 1679581782
transform 1 0 9024 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_95
timestamp 1679581782
transform 1 0 9696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_102
timestamp 1679581782
transform 1 0 10368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_109
timestamp 1679581782
transform 1 0 11040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_116
timestamp 1679581782
transform 1 0 11712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_123
timestamp 1679581782
transform 1 0 12384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_130
timestamp 1679581782
transform 1 0 13056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_137
timestamp 1679581782
transform 1 0 13728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_144
timestamp 1679581782
transform 1 0 14400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_151
timestamp 1679581782
transform 1 0 15072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_158
timestamp 1679581782
transform 1 0 15744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_165
timestamp 1679581782
transform 1 0 16416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_172
timestamp 1679581782
transform 1 0 17088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_179
timestamp 1679581782
transform 1 0 17760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_186
timestamp 1679581782
transform 1 0 18432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_193
timestamp 1679581782
transform 1 0 19104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_200
timestamp 1679581782
transform 1 0 19776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_207
timestamp 1679581782
transform 1 0 20448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_214
timestamp 1679581782
transform 1 0 21120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_221
timestamp 1679581782
transform 1 0 21792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_228
timestamp 1679581782
transform 1 0 22464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_235
timestamp 1679581782
transform 1 0 23136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_242
timestamp 1679581782
transform 1 0 23808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_249
timestamp 1679581782
transform 1 0 24480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_256
timestamp 1679581782
transform 1 0 25152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_263
timestamp 1679581782
transform 1 0 25824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_270
timestamp 1679581782
transform 1 0 26496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_277
timestamp 1679581782
transform 1 0 27168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_284
timestamp 1679581782
transform 1 0 27840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_291
timestamp 1679581782
transform 1 0 28512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_298
timestamp 1679581782
transform 1 0 29184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_305
timestamp 1679581782
transform 1 0 29856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_312
timestamp 1679581782
transform 1 0 30528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_319
timestamp 1679581782
transform 1 0 31200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_326
timestamp 1679581782
transform 1 0 31872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_333
timestamp 1679581782
transform 1 0 32544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_340
timestamp 1679581782
transform 1 0 33216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_347
timestamp 1679581782
transform 1 0 33888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_354
timestamp 1679581782
transform 1 0 34560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_361
timestamp 1679581782
transform 1 0 35232 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_368
timestamp 1677580104
transform 1 0 35904 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_380
timestamp 1679581782
transform 1 0 37056 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_393
timestamp 1677580104
transform 1 0 38304 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_395
timestamp 1677579658
transform 1 0 38496 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_406
timestamp 1679581782
transform 1 0 39552 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_413
timestamp 1677580104
transform 1 0 40224 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_443
timestamp 1677580104
transform 1 0 43104 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_452
timestamp 1677579658
transform 1 0 43968 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_458
timestamp 1679581782
transform 1 0 44544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_465
timestamp 1679581782
transform 1 0 45216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_472
timestamp 1679581782
transform 1 0 45888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_479
timestamp 1679581782
transform 1 0 46560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_491
timestamp 1679577901
transform 1 0 47712 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_500
timestamp 1677579658
transform 1 0 48576 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_504
timestamp 1679581782
transform 1 0 48960 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_511
timestamp 1677579658
transform 1 0 49632 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679581782
transform 1 0 52320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_549
timestamp 1679577901
transform 1 0 53280 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_553
timestamp 1677579658
transform 1 0 53664 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_559
timestamp 1679581782
transform 1 0 54240 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_569
timestamp 1677580104
transform 1 0 55200 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_571
timestamp 1677579658
transform 1 0 55392 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_575
timestamp 1677579658
transform 1 0 55776 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_579
timestamp 1677579658
transform 1 0 56160 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_593
timestamp 1677580104
transform 1 0 57504 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_598
timestamp 1679581782
transform 1 0 57984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_605
timestamp 1679577901
transform 1 0 58656 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_609
timestamp 1677580104
transform 1 0 59040 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_624
timestamp 1679577901
transform 1 0 60480 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_633
timestamp 1679581782
transform 1 0 61344 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_643
timestamp 1677580104
transform 1 0 62304 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_648
timestamp 1677580104
transform 1 0 62784 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_650
timestamp 1677579658
transform 1 0 62976 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_654
timestamp 1679577901
transform 1 0 63360 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_658
timestamp 1677579658
transform 1 0 63744 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_667
timestamp 1677579658
transform 1 0 64608 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_671
timestamp 1677579658
transform 1 0 64992 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_678
timestamp 1677580104
transform 1 0 65664 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_712
timestamp 1677579658
transform 1 0 68928 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_718
timestamp 1679577901
transform 1 0 69504 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_727
timestamp 1679581782
transform 1 0 70368 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_734
timestamp 1677579658
transform 1 0 71040 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_740
timestamp 1677580104
transform 1 0 71616 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_742
timestamp 1677579658
transform 1 0 71808 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_746
timestamp 1677579658
transform 1 0 72192 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_750
timestamp 1677579658
transform 1 0 72576 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_754
timestamp 1679581782
transform 1 0 72960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_761
timestamp 1679581782
transform 1 0 73632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_768
timestamp 1679577901
transform 1 0 74304 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_772
timestamp 1677579658
transform 1 0 74688 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_778
timestamp 1677580104
transform 1 0 75264 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_783
timestamp 1677580104
transform 1 0 75744 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_785
timestamp 1677579658
transform 1 0 75936 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_796
timestamp 1677579658
transform 1 0 76992 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679581782
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_807
timestamp 1679577901
transform 1 0 78048 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_811
timestamp 1677580104
transform 1 0 78432 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_819
timestamp 1679577901
transform 1 0 79200 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_4
timestamp 1679581782
transform 1 0 960 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_11
timestamp 1677579658
transform 1 0 1632 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_20
timestamp 1679581782
transform 1 0 2496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_27
timestamp 1679581782
transform 1 0 3168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_34
timestamp 1679581782
transform 1 0 3840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_41
timestamp 1679581782
transform 1 0 4512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_48
timestamp 1679581782
transform 1 0 5184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_55
timestamp 1679581782
transform 1 0 5856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_62
timestamp 1679581782
transform 1 0 6528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_69
timestamp 1679581782
transform 1 0 7200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_76
timestamp 1679581782
transform 1 0 7872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_83
timestamp 1679581782
transform 1 0 8544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_90
timestamp 1679581782
transform 1 0 9216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_97
timestamp 1679581782
transform 1 0 9888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_104
timestamp 1679581782
transform 1 0 10560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_111
timestamp 1679581782
transform 1 0 11232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_118
timestamp 1679581782
transform 1 0 11904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_125
timestamp 1679581782
transform 1 0 12576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_132
timestamp 1679581782
transform 1 0 13248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_139
timestamp 1679581782
transform 1 0 13920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_146
timestamp 1679581782
transform 1 0 14592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_153
timestamp 1679581782
transform 1 0 15264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_160
timestamp 1679581782
transform 1 0 15936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_167
timestamp 1679581782
transform 1 0 16608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_174
timestamp 1679581782
transform 1 0 17280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_181
timestamp 1679581782
transform 1 0 17952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_188
timestamp 1679581782
transform 1 0 18624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_195
timestamp 1679581782
transform 1 0 19296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_202
timestamp 1679581782
transform 1 0 19968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_209
timestamp 1679581782
transform 1 0 20640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_216
timestamp 1679581782
transform 1 0 21312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_223
timestamp 1679581782
transform 1 0 21984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_230
timestamp 1679581782
transform 1 0 22656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_237
timestamp 1679581782
transform 1 0 23328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_244
timestamp 1679581782
transform 1 0 24000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_251
timestamp 1679581782
transform 1 0 24672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_258
timestamp 1679581782
transform 1 0 25344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_265
timestamp 1679581782
transform 1 0 26016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_272
timestamp 1679581782
transform 1 0 26688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_279
timestamp 1679581782
transform 1 0 27360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_286
timestamp 1679581782
transform 1 0 28032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_293
timestamp 1679581782
transform 1 0 28704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_300
timestamp 1679581782
transform 1 0 29376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_307
timestamp 1679581782
transform 1 0 30048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_314
timestamp 1679581782
transform 1 0 30720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_321
timestamp 1679581782
transform 1 0 31392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_328
timestamp 1679581782
transform 1 0 32064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_335
timestamp 1679581782
transform 1 0 32736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_342
timestamp 1679581782
transform 1 0 33408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_349
timestamp 1679581782
transform 1 0 34080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_356
timestamp 1679577901
transform 1 0 34752 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_610
timestamp 1677580104
transform 1 0 59136 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_612
timestamp 1677579658
transform 1 0 59328 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_640
timestamp 1679581782
transform 1 0 62016 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_647
timestamp 1677579658
transform 1 0 62688 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_680
timestamp 1679581782
transform 1 0 65856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_687
timestamp 1679577901
transform 1 0 66528 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_696
timestamp 1679581782
transform 1 0 67392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_703
timestamp 1679577901
transform 1 0 68064 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_707
timestamp 1677580104
transform 1 0 68448 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_767
timestamp 1679577901
transform 1 0 74208 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_771
timestamp 1677580104
transform 1 0 74592 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_786
timestamp 1677579658
transform 1 0 76032 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_818
timestamp 1679577901
transform 1 0 79104 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_822
timestamp 1677579658
transform 1 0 79488 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_4
timestamp 1679581782
transform 1 0 960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_11
timestamp 1679581782
transform 1 0 1632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_18
timestamp 1679581782
transform 1 0 2304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_25
timestamp 1679581782
transform 1 0 2976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1679581782
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_39
timestamp 1679581782
transform 1 0 4320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_46
timestamp 1679581782
transform 1 0 4992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_53
timestamp 1679581782
transform 1 0 5664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_60
timestamp 1679581782
transform 1 0 6336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679581782
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679581782
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679581782
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679581782
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_109
timestamp 1679581782
transform 1 0 11040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_116
timestamp 1679581782
transform 1 0 11712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_123
timestamp 1679581782
transform 1 0 12384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_130
timestamp 1679581782
transform 1 0 13056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_137
timestamp 1679581782
transform 1 0 13728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_144
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_151
timestamp 1679581782
transform 1 0 15072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_158
timestamp 1679581782
transform 1 0 15744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_165
timestamp 1679581782
transform 1 0 16416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679581782
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679581782
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679581782
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679581782
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679581782
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679581782
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679581782
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_221
timestamp 1679581782
transform 1 0 21792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679581782
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679581782
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_242
timestamp 1679581782
transform 1 0 23808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_249
timestamp 1679581782
transform 1 0 24480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_256
timestamp 1679581782
transform 1 0 25152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_263
timestamp 1679581782
transform 1 0 25824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_270
timestamp 1679581782
transform 1 0 26496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_277
timestamp 1679581782
transform 1 0 27168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_284
timestamp 1679581782
transform 1 0 27840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_291
timestamp 1679581782
transform 1 0 28512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_298
timestamp 1679581782
transform 1 0 29184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_305
timestamp 1679581782
transform 1 0 29856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_312
timestamp 1679581782
transform 1 0 30528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_319
timestamp 1679581782
transform 1 0 31200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_326
timestamp 1679581782
transform 1 0 31872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_333
timestamp 1679581782
transform 1 0 32544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_340
timestamp 1679581782
transform 1 0 33216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_347
timestamp 1679581782
transform 1 0 33888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_354
timestamp 1679581782
transform 1 0 34560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_361
timestamp 1679581782
transform 1 0 35232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_368
timestamp 1679581782
transform 1 0 35904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_375
timestamp 1679581782
transform 1 0 36576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_382
timestamp 1679577901
transform 1 0 37248 0 1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_32_389
timestamp 1679577901
transform 1 0 37920 0 1 24948
box -48 -56 432 834
use sg13g2_decap_4  FILLER_32_398
timestamp 1679577901
transform 1 0 38784 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_402
timestamp 1677579658
transform 1 0 39168 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_414
timestamp 1677580104
transform 1 0 40320 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_423
timestamp 1679577901
transform 1 0 41184 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_427
timestamp 1677579658
transform 1 0 41568 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_440
timestamp 1677580104
transform 1 0 42816 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_454
timestamp 1677580104
transform 1 0 44160 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_466
timestamp 1677580104
transform 1 0 45312 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_471
timestamp 1679581782
transform 1 0 45792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_478
timestamp 1679581782
transform 1 0 46464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_485
timestamp 1679577901
transform 1 0 47136 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_489
timestamp 1677580104
transform 1 0 47520 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_498
timestamp 1679581782
transform 1 0 48384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_508
timestamp 1679581782
transform 1 0 49344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_540
timestamp 1679581782
transform 1 0 52416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_547
timestamp 1679577901
transform 1 0 53088 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_551
timestamp 1677579658
transform 1 0 53472 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_564
timestamp 1679581782
transform 1 0 54720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_571
timestamp 1679581782
transform 1 0 55392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_578
timestamp 1679577901
transform 1 0 56064 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_589
timestamp 1677580104
transform 1 0 57120 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_591
timestamp 1677579658
transform 1 0 57312 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_597
timestamp 1679577901
transform 1 0 57888 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_601
timestamp 1677579658
transform 1 0 58272 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_655
timestamp 1677580104
transform 1 0 63456 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_664
timestamp 1677580104
transform 1 0 64320 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_671
timestamp 1679577901
transform 1 0 64992 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_691
timestamp 1677580104
transform 1 0 66912 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_698
timestamp 1679581782
transform 1 0 67584 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_705
timestamp 1677580104
transform 1 0 68256 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_707
timestamp 1677579658
transform 1 0 68448 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_711
timestamp 1677579658
transform 1 0 68832 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_727
timestamp 1679577901
transform 1 0 70368 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_731
timestamp 1677580104
transform 1 0 70752 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_740
timestamp 1677580104
transform 1 0 71616 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_742
timestamp 1677579658
transform 1 0 71808 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_748
timestamp 1679581782
transform 1 0 72384 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_755
timestamp 1677579658
transform 1 0 73056 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_788
timestamp 1679577901
transform 1 0 76224 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_792
timestamp 1677579658
transform 1 0 76608 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_798
timestamp 1677579658
transform 1 0 77184 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_804
timestamp 1677580104
transform 1 0 77760 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_806
timestamp 1677579658
transform 1 0 77952 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_810
timestamp 1679581782
transform 1 0 78336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_817
timestamp 1679577901
transform 1 0 79008 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_821
timestamp 1677580104
transform 1 0 79392 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_4
timestamp 1679581782
transform 1 0 960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_11
timestamp 1679581782
transform 1 0 1632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_18
timestamp 1679581782
transform 1 0 2304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_25
timestamp 1679581782
transform 1 0 2976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_32
timestamp 1679581782
transform 1 0 3648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_39
timestamp 1679581782
transform 1 0 4320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679581782
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_53
timestamp 1679581782
transform 1 0 5664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_60
timestamp 1679581782
transform 1 0 6336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_67
timestamp 1679581782
transform 1 0 7008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_74
timestamp 1679581782
transform 1 0 7680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_81
timestamp 1679581782
transform 1 0 8352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_88
timestamp 1679581782
transform 1 0 9024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_95
timestamp 1679581782
transform 1 0 9696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_102
timestamp 1679581782
transform 1 0 10368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_109
timestamp 1679581782
transform 1 0 11040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_116
timestamp 1679581782
transform 1 0 11712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_123
timestamp 1679581782
transform 1 0 12384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_130
timestamp 1679581782
transform 1 0 13056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_137
timestamp 1679581782
transform 1 0 13728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_144
timestamp 1679581782
transform 1 0 14400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_151
timestamp 1679581782
transform 1 0 15072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_158
timestamp 1679581782
transform 1 0 15744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_165
timestamp 1679581782
transform 1 0 16416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_172
timestamp 1679581782
transform 1 0 17088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_179
timestamp 1679581782
transform 1 0 17760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_186
timestamp 1679581782
transform 1 0 18432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_193
timestamp 1679581782
transform 1 0 19104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_200
timestamp 1679581782
transform 1 0 19776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_207
timestamp 1679581782
transform 1 0 20448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_214
timestamp 1679581782
transform 1 0 21120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_221
timestamp 1679581782
transform 1 0 21792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_228
timestamp 1679581782
transform 1 0 22464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_235
timestamp 1679581782
transform 1 0 23136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_242
timestamp 1679581782
transform 1 0 23808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_249
timestamp 1679581782
transform 1 0 24480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_256
timestamp 1679581782
transform 1 0 25152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_263
timestamp 1679581782
transform 1 0 25824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_270
timestamp 1679581782
transform 1 0 26496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_277
timestamp 1679581782
transform 1 0 27168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_284
timestamp 1679581782
transform 1 0 27840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_291
timestamp 1679581782
transform 1 0 28512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_298
timestamp 1679581782
transform 1 0 29184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_305
timestamp 1679581782
transform 1 0 29856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_312
timestamp 1679581782
transform 1 0 30528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_319
timestamp 1679581782
transform 1 0 31200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_326
timestamp 1679581782
transform 1 0 31872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_333
timestamp 1679581782
transform 1 0 32544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_340
timestamp 1679581782
transform 1 0 33216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_347
timestamp 1679581782
transform 1 0 33888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_354
timestamp 1679581782
transform 1 0 34560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_361
timestamp 1679581782
transform 1 0 35232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_368
timestamp 1679581782
transform 1 0 35904 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_375
timestamp 1677580104
transform 1 0 36576 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_377
timestamp 1677579658
transform 1 0 36768 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_452
timestamp 1677579658
transform 1 0 43968 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_487
timestamp 1679577901
transform 1 0 47328 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679581782
transform 1 0 50304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679581782
transform 1 0 50976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679581782
transform 1 0 51648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679581782
transform 1 0 52320 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_558
timestamp 1677580104
transform 1 0 54144 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_569
timestamp 1679577901
transform 1 0 55200 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_573
timestamp 1677580104
transform 1 0 55584 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_617
timestamp 1677579658
transform 1 0 59808 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_627
timestamp 1677579658
transform 1 0 60768 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_635
timestamp 1677579658
transform 1 0 61536 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_641
timestamp 1679581782
transform 1 0 62112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_648
timestamp 1679577901
transform 1 0 62784 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_679
timestamp 1677580104
transform 1 0 65760 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_681
timestamp 1677579658
transform 1 0 65952 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_709
timestamp 1677579658
transform 1 0 68640 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_716
timestamp 1677579658
transform 1 0 69312 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_726
timestamp 1677580104
transform 1 0 70272 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_737
timestamp 1679577901
transform 1 0 71328 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_746
timestamp 1679577901
transform 1 0 72192 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_755
timestamp 1677580104
transform 1 0 73056 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_760
timestamp 1679581782
transform 1 0 73536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_767
timestamp 1679581782
transform 1 0 74208 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_774
timestamp 1677580104
transform 1 0 74880 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_776
timestamp 1677579658
transform 1 0 75072 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_821
timestamp 1677580104
transform 1 0 79392 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679581782
transform 1 0 10656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679581782
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679581782
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679581782
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679581782
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679581782
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679581782
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679581782
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679581782
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679581782
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679581782
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679581782
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679581782
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679581782
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679581782
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679581782
transform 1 0 28800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679581782
transform 1 0 29472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679581782
transform 1 0 30144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679581782
transform 1 0 30816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679581782
transform 1 0 31488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679581782
transform 1 0 32160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679581782
transform 1 0 32832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679581782
transform 1 0 33504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679581782
transform 1 0 34176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679581782
transform 1 0 34848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679581782
transform 1 0 35520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679581782
transform 1 0 36192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679581782
transform 1 0 36864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679581782
transform 1 0 37536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679581782
transform 1 0 38208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_399
timestamp 1679577901
transform 1 0 38880 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_403
timestamp 1677579658
transform 1 0 39264 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_422
timestamp 1679581782
transform 1 0 41088 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_429
timestamp 1677580104
transform 1 0 41760 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_431
timestamp 1677579658
transform 1 0 41952 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_463
timestamp 1679581782
transform 1 0 45024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_470
timestamp 1679581782
transform 1 0 45696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_477
timestamp 1679581782
transform 1 0 46368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_500
timestamp 1679577901
transform 1 0 48576 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_507
timestamp 1679581782
transform 1 0 49248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_514
timestamp 1679581782
transform 1 0 49920 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_521
timestamp 1677580104
transform 1 0 50592 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_555
timestamp 1677579658
transform 1 0 53856 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_583
timestamp 1679581782
transform 1 0 56544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_590
timestamp 1679581782
transform 1 0 57216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_597
timestamp 1679577901
transform 1 0 57888 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_601
timestamp 1677579658
transform 1 0 58272 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_640
timestamp 1679581782
transform 1 0 62016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_647
timestamp 1679581782
transform 1 0 62688 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_654
timestamp 1677580104
transform 1 0 63360 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_656
timestamp 1677579658
transform 1 0 63552 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_663
timestamp 1677579658
transform 1 0 64224 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679581782
transform 1 0 65088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679581782
transform 1 0 65760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679581782
transform 1 0 66432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_693
timestamp 1679581782
transform 1 0 67104 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_700
timestamp 1677580104
transform 1 0 67776 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_729
timestamp 1677580104
transform 1 0 70560 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_742
timestamp 1677579658
transform 1 0 71808 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_814
timestamp 1679581782
transform 1 0 78720 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_821
timestamp 1677580104
transform 1 0 79392 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679581782
transform 1 0 37536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679581782
transform 1 0 38208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679581782
transform 1 0 38880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_406
timestamp 1679577901
transform 1 0 39552 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_410
timestamp 1677580104
transform 1 0 39936 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_421
timestamp 1679581782
transform 1 0 40992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_428
timestamp 1679577901
transform 1 0 41664 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_435
timestamp 1677579658
transform 1 0 42336 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_458
timestamp 1679581782
transform 1 0 44544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_465
timestamp 1679577901
transform 1 0 45216 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_469
timestamp 1677580104
transform 1 0 45600 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_475
timestamp 1679581782
transform 1 0 46176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_482
timestamp 1679577901
transform 1 0 46848 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_35_528
timestamp 1679581782
transform 1 0 51264 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_546
timestamp 1677579658
transform 1 0 52992 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679581782
transform 1 0 55680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679581782
transform 1 0 56352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_588
timestamp 1679577901
transform 1 0 57024 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_597
timestamp 1677579658
transform 1 0 57888 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_601
timestamp 1679577901
transform 1 0 58272 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_605
timestamp 1677579658
transform 1 0 58656 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_622
timestamp 1677580104
transform 1 0 60288 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_624
timestamp 1677579658
transform 1 0 60480 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_636
timestamp 1679581782
transform 1 0 61632 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_670
timestamp 1677579658
transform 1 0 64896 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_683
timestamp 1677580104
transform 1 0 66144 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_685
timestamp 1677579658
transform 1 0 66336 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_689
timestamp 1679581782
transform 1 0 66720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_696
timestamp 1679581782
transform 1 0 67392 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_703
timestamp 1677580104
transform 1 0 68064 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_705
timestamp 1677579658
transform 1 0 68256 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_733
timestamp 1677579658
transform 1 0 70944 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_737
timestamp 1677579658
transform 1 0 71328 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_745
timestamp 1679581782
transform 1 0 72096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_752
timestamp 1679581782
transform 1 0 72768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_759
timestamp 1679581782
transform 1 0 73440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_766
timestamp 1679581782
transform 1 0 74112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_773
timestamp 1679581782
transform 1 0 74784 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_780
timestamp 1677580104
transform 1 0 75456 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679581782
transform 1 0 38880 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_493
timestamp 1677580104
transform 1 0 47904 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_500
timestamp 1679581782
transform 1 0 48576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_507
timestamp 1679577901
transform 1 0 49248 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_550
timestamp 1679581782
transform 1 0 53376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_557
timestamp 1679581782
transform 1 0 54048 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_564
timestamp 1677580104
transform 1 0 54720 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_566
timestamp 1677579658
transform 1 0 54912 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_570
timestamp 1679581782
transform 1 0 55296 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_577
timestamp 1677579658
transform 1 0 55968 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_610
timestamp 1679577901
transform 1 0 59136 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_614
timestamp 1677580104
transform 1 0 59520 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_622
timestamp 1677580104
transform 1 0 60288 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_644
timestamp 1677580104
transform 1 0 62400 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_646
timestamp 1677579658
transform 1 0 62592 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_707
timestamp 1679577901
transform 1 0 68448 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_715
timestamp 1679581782
transform 1 0 69216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_722
timestamp 1679577901
transform 1 0 69888 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_726
timestamp 1677579658
transform 1 0 70272 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_738
timestamp 1677580104
transform 1 0 71424 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_740
timestamp 1677579658
transform 1 0 71616 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_750
timestamp 1677579658
transform 1 0 72576 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_756
timestamp 1679577901
transform 1 0 73152 0 1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_36_763
timestamp 1679577901
transform 1 0 73824 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_767
timestamp 1677580104
transform 1 0 74208 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_806
timestamp 1679581782
transform 1 0 77952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_813
timestamp 1679581782
transform 1 0 78624 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_820
timestamp 1677580104
transform 1 0 79296 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_822
timestamp 1677579658
transform 1 0 79488 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679581782
transform 1 0 38880 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_406
timestamp 1677579658
transform 1 0 39552 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_419
timestamp 1679581782
transform 1 0 40800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_426
timestamp 1679581782
transform 1 0 41472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_433
timestamp 1679577901
transform 1 0 42144 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_447
timestamp 1679581782
transform 1 0 43488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_454
timestamp 1679581782
transform 1 0 44160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_461
timestamp 1679581782
transform 1 0 44832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_468
timestamp 1679581782
transform 1 0 45504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_475
timestamp 1679577901
transform 1 0 46176 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_490
timestamp 1677580104
transform 1 0 47616 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_492
timestamp 1677579658
transform 1 0 47808 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_505
timestamp 1677580104
transform 1 0 49056 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_540
timestamp 1679581782
transform 1 0 52416 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_579
timestamp 1677580104
transform 1 0 56160 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_594
timestamp 1679577901
transform 1 0 57600 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_598
timestamp 1677579658
transform 1 0 57984 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_602
timestamp 1679577901
transform 1 0 58368 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_671
timestamp 1677580104
transform 1 0 64992 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_677
timestamp 1677580104
transform 1 0 65568 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_693
timestamp 1677580104
transform 1 0 67104 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_698
timestamp 1679581782
transform 1 0 67584 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_705
timestamp 1677579658
transform 1 0 68256 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_743
timestamp 1677580104
transform 1 0 71904 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_772
timestamp 1679581782
transform 1 0 74688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_779
timestamp 1679581782
transform 1 0 75360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_786
timestamp 1679577901
transform 1 0 76032 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_808
timestamp 1679581782
transform 1 0 78144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_815
timestamp 1679581782
transform 1 0 78816 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_822
timestamp 1677579658
transform 1 0 79488 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679581782
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679581782
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_413
timestamp 1677579658
transform 1 0 40224 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_418
timestamp 1679581782
transform 1 0 40704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_425
timestamp 1679581782
transform 1 0 41376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_432
timestamp 1679581782
transform 1 0 42048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_439
timestamp 1679581782
transform 1 0 42720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_446
timestamp 1679581782
transform 1 0 43392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_453
timestamp 1679581782
transform 1 0 44064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_460
timestamp 1679577901
transform 1 0 44736 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_464
timestamp 1677580104
transform 1 0 45120 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_496
timestamp 1677579658
transform 1 0 48192 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_528
timestamp 1677579658
transform 1 0 51264 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_534
timestamp 1677580104
transform 1 0 51840 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679581782
transform 1 0 52320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679581782
transform 1 0 52992 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_553
timestamp 1677580104
transform 1 0 53664 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_575
timestamp 1677580104
transform 1 0 55776 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_582
timestamp 1677579658
transform 1 0 56448 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_618
timestamp 1679581782
transform 1 0 59904 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_625
timestamp 1677579658
transform 1 0 60576 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_642
timestamp 1679581782
transform 1 0 62208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_649
timestamp 1679581782
transform 1 0 62880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_656
timestamp 1679581782
transform 1 0 63552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_663
timestamp 1679577901
transform 1 0 64224 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_667
timestamp 1677579658
transform 1 0 64608 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_679
timestamp 1677579658
transform 1 0 65760 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_687
timestamp 1677579658
transform 1 0 66528 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_715
timestamp 1679581782
transform 1 0 69216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_722
timestamp 1679581782
transform 1 0 69888 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_729
timestamp 1677579658
transform 1 0 70560 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_754
timestamp 1677579658
transform 1 0 72960 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_767
timestamp 1679581782
transform 1 0 74208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_774
timestamp 1679577901
transform 1 0 74880 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_778
timestamp 1677579658
transform 1 0 75264 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679581782
transform 1 0 40896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679581782
transform 1 0 41568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679581782
transform 1 0 42240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679581782
transform 1 0 42912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679581782
transform 1 0 43584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679581782
transform 1 0 44256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679581782
transform 1 0 44928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679581782
transform 1 0 46272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679581782
transform 1 0 46944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_490
timestamp 1679577901
transform 1 0 47616 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_500
timestamp 1679581782
transform 1 0 48576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_507
timestamp 1679581782
transform 1 0 49248 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_514
timestamp 1677580104
transform 1 0 49920 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_548
timestamp 1679577901
transform 1 0 53184 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_583
timestamp 1679581782
transform 1 0 56544 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_590
timestamp 1677579658
transform 1 0 57216 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_623
timestamp 1679577901
transform 1 0 60384 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_659
timestamp 1677579658
transform 1 0 63840 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_695
timestamp 1679581782
transform 1 0 67296 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_702
timestamp 1677579658
transform 1 0 67968 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_708
timestamp 1679577901
transform 1 0 68544 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_805
timestamp 1679581782
transform 1 0 77856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_812
timestamp 1679581782
transform 1 0 78528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_819
timestamp 1679577901
transform 1 0 79200 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679581782
transform 1 0 39552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679581782
transform 1 0 40224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679581782
transform 1 0 41568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679581782
transform 1 0 42912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679581782
transform 1 0 43584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679581782
transform 1 0 44256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679581782
transform 1 0 44928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679581782
transform 1 0 45600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679581782
transform 1 0 46272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679581782
transform 1 0 48288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679581782
transform 1 0 48960 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_511
timestamp 1677580104
transform 1 0 49632 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_513
timestamp 1677579658
transform 1 0 49824 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_531
timestamp 1677580104
transform 1 0 51552 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_572
timestamp 1679581782
transform 1 0 55488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_579
timestamp 1679581782
transform 1 0 56160 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_586
timestamp 1677580104
transform 1 0 56832 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_603
timestamp 1677579658
transform 1 0 58464 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_612
timestamp 1679581782
transform 1 0 59328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_619
timestamp 1679581782
transform 1 0 60000 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_626
timestamp 1677579658
transform 1 0 60672 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_639
timestamp 1679581782
transform 1 0 61920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_646
timestamp 1679577901
transform 1 0 62592 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_650
timestamp 1677580104
transform 1 0 62976 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_662
timestamp 1679581782
transform 1 0 64128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_669
timestamp 1679581782
transform 1 0 64800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_676
timestamp 1679581782
transform 1 0 65472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_688
timestamp 1679577901
transform 1 0 66624 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_724
timestamp 1677580104
transform 1 0 70080 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_726
timestamp 1677579658
transform 1 0 70272 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_730
timestamp 1679581782
transform 1 0 70656 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_744
timestamp 1677580104
transform 1 0 72000 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_765
timestamp 1677580104
transform 1 0 74016 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_767
timestamp 1677579658
transform 1 0 74208 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_771
timestamp 1679581782
transform 1 0 74592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_778
timestamp 1679581782
transform 1 0 75264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_809
timestamp 1679581782
transform 1 0 78240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_816
timestamp 1679581782
transform 1 0 78912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679581782
transform 1 0 40224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679581782
transform 1 0 42240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679581782
transform 1 0 42912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679581782
transform 1 0 43584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679581782
transform 1 0 44256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679581782
transform 1 0 44928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679581782
transform 1 0 45600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679581782
transform 1 0 46272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679581782
transform 1 0 46944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679581782
transform 1 0 47616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679581782
transform 1 0 48288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679581782
transform 1 0 48960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679581782
transform 1 0 49632 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_518
timestamp 1677580104
transform 1 0 50304 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_560
timestamp 1677579658
transform 1 0 54336 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_588
timestamp 1677579658
transform 1 0 57024 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_625
timestamp 1677579658
transform 1 0 60576 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_632
timestamp 1677580104
transform 1 0 61248 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_639
timestamp 1679581782
transform 1 0 61920 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_646
timestamp 1677579658
transform 1 0 62592 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_680
timestamp 1679577901
transform 1 0 65856 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_684
timestamp 1677579658
transform 1 0 66240 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_691
timestamp 1677580104
transform 1 0 66912 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_700
timestamp 1679577901
transform 1 0 67776 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_704
timestamp 1677580104
transform 1 0 68160 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679581782
transform 1 0 69120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679581782
transform 1 0 69792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_728
timestamp 1679581782
transform 1 0 70464 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_735
timestamp 1677580104
transform 1 0 71136 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_737
timestamp 1677579658
transform 1 0 71328 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679581782
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_786
timestamp 1677580104
transform 1 0 76032 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_822
timestamp 1677579658
transform 1 0 79488 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679581782
transform 1 0 42240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679581782
transform 1 0 42912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679581782
transform 1 0 43584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679581782
transform 1 0 44256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679581782
transform 1 0 44928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679581782
transform 1 0 45600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679581782
transform 1 0 46272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679581782
transform 1 0 46944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679581782
transform 1 0 47616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679581782
transform 1 0 48288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679581782
transform 1 0 48960 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_511
timestamp 1677579658
transform 1 0 49632 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_516
timestamp 1677580104
transform 1 0 50112 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_518
timestamp 1677579658
transform 1 0 50304 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_559
timestamp 1677580104
transform 1 0 54240 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_561
timestamp 1677579658
transform 1 0 54432 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_573
timestamp 1677580104
transform 1 0 55584 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_580
timestamp 1679581782
transform 1 0 56256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_587
timestamp 1679581782
transform 1 0 56928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_594
timestamp 1679581782
transform 1 0 57600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_601
timestamp 1679581782
transform 1 0 58272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_608
timestamp 1679581782
transform 1 0 58944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_615
timestamp 1679577901
transform 1 0 59616 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_619
timestamp 1677579658
transform 1 0 60000 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_657
timestamp 1677579658
transform 1 0 63648 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_662
timestamp 1679581782
transform 1 0 64128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_669
timestamp 1679577901
transform 1 0 64800 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_673
timestamp 1677580104
transform 1 0 65184 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_705
timestamp 1679581782
transform 1 0 68256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_712
timestamp 1679581782
transform 1 0 68928 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_719
timestamp 1677579658
transform 1 0 69600 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_754
timestamp 1679581782
transform 1 0 72960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_761
timestamp 1679581782
transform 1 0 73632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_768
timestamp 1679581782
transform 1 0 74304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_775
timestamp 1679581782
transform 1 0 74976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_782
timestamp 1679581782
transform 1 0 75648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_816
timestamp 1679581782
transform 1 0 78912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679581782
transform 1 0 46272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679581782
transform 1 0 46944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679581782
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679581782
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_504
timestamp 1677580104
transform 1 0 48960 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_506
timestamp 1677579658
transform 1 0 49152 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_537
timestamp 1677579658
transform 1 0 52128 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_565
timestamp 1677579658
transform 1 0 54816 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_600
timestamp 1679581782
transform 1 0 58176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_607
timestamp 1679577901
transform 1 0 58848 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_616
timestamp 1677579658
transform 1 0 59712 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_620
timestamp 1679581782
transform 1 0 60096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_627
timestamp 1679581782
transform 1 0 60768 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_634
timestamp 1677580104
transform 1 0 61440 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_636
timestamp 1677579658
transform 1 0 61632 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_641
timestamp 1679581782
transform 1 0 62112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_648
timestamp 1679581782
transform 1 0 62784 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_658
timestamp 1677580104
transform 1 0 63744 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_670
timestamp 1679581782
transform 1 0 64896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_677
timestamp 1679581782
transform 1 0 65568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_684
timestamp 1679577901
transform 1 0 66240 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_688
timestamp 1677579658
transform 1 0 66624 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_726
timestamp 1679581782
transform 1 0 70272 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_733
timestamp 1677580104
transform 1 0 70944 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_735
timestamp 1677579658
transform 1 0 71136 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_746
timestamp 1677580104
transform 1 0 72192 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_748
timestamp 1677579658
transform 1 0 72384 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_752
timestamp 1679581782
transform 1 0 72768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_759
timestamp 1679581782
transform 1 0 73440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_766
timestamp 1679577901
transform 1 0 74112 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_770
timestamp 1677580104
transform 1 0 74496 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_775
timestamp 1679581782
transform 1 0 74976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_782
timestamp 1679577901
transform 1 0 75648 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_786
timestamp 1677580104
transform 1 0 76032 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_810
timestamp 1679581782
transform 1 0 78336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_817
timestamp 1679577901
transform 1 0 79008 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_821
timestamp 1677580104
transform 1 0 79392 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679581782
transform 1 0 45600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679581782
transform 1 0 46272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679581782
transform 1 0 46944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679581782
transform 1 0 47616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679581782
transform 1 0 48288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679581782
transform 1 0 48960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679581782
transform 1 0 50304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679581782
transform 1 0 50976 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_532
timestamp 1677580104
transform 1 0 51648 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_540
timestamp 1677579658
transform 1 0 52416 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_571
timestamp 1679577901
transform 1 0 55392 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_580
timestamp 1679581782
transform 1 0 56256 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_587
timestamp 1677580104
transform 1 0 56928 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_592
timestamp 1679581782
transform 1 0 57408 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_599
timestamp 1677580104
transform 1 0 58080 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_601
timestamp 1677579658
transform 1 0 58272 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_634
timestamp 1679581782
transform 1 0 61440 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_641
timestamp 1677579658
transform 1 0 62112 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_648
timestamp 1677580104
transform 1 0 62784 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_662
timestamp 1677579658
transform 1 0 64128 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_690
timestamp 1677580104
transform 1 0 66816 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_705
timestamp 1677580104
transform 1 0 68256 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_707
timestamp 1677579658
transform 1 0 68448 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_713
timestamp 1679577901
transform 1 0 69024 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_717
timestamp 1677579658
transform 1 0 69408 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679581782
transform 1 0 69792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_728
timestamp 1679577901
transform 1 0 70464 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_813
timestamp 1679581782
transform 1 0 78624 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_820
timestamp 1677580104
transform 1 0 79296 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_822
timestamp 1677579658
transform 1 0 79488 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679581782
transform 1 0 48288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679581782
transform 1 0 48960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679581782
transform 1 0 49632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679581782
transform 1 0 50304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679581782
transform 1 0 50976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679581782
transform 1 0 51648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679581782
transform 1 0 52320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679581782
transform 1 0 52992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679581782
transform 1 0 53664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679581782
transform 1 0 54336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_594
timestamp 1679581782
transform 1 0 57600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_614
timestamp 1679577901
transform 1 0 59520 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_618
timestamp 1677580104
transform 1 0 59904 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_662
timestamp 1679581782
transform 1 0 64128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_669
timestamp 1679581782
transform 1 0 64800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_676
timestamp 1679581782
transform 1 0 65472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_683
timestamp 1679581782
transform 1 0 66144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_690
timestamp 1679581782
transform 1 0 66816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_697
timestamp 1679577901
transform 1 0 67488 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_701
timestamp 1677580104
transform 1 0 67872 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_706
timestamp 1679581782
transform 1 0 68352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_746
timestamp 1679577901
transform 1 0 72192 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_750
timestamp 1677580104
transform 1 0 72576 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679581782
transform 1 0 75840 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_791
timestamp 1677580104
transform 1 0 76512 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_574
timestamp 1677580104
transform 1 0 55680 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_593
timestamp 1677579658
transform 1 0 57504 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_639
timestamp 1679581782
transform 1 0 61920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_646
timestamp 1679581782
transform 1 0 62592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_653
timestamp 1679577901
transform 1 0 63264 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_657
timestamp 1677579658
transform 1 0 63648 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_681
timestamp 1679577901
transform 1 0 65952 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_712
timestamp 1679581782
transform 1 0 68928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_719
timestamp 1679581782
transform 1 0 69600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_726
timestamp 1679581782
transform 1 0 70272 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_733
timestamp 1677580104
transform 1 0 70944 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_735
timestamp 1677579658
transform 1 0 71136 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_741
timestamp 1677580104
transform 1 0 71712 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_743
timestamp 1677579658
transform 1 0 71904 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_747
timestamp 1677579658
transform 1 0 72288 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_755
timestamp 1679581782
transform 1 0 73056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_775
timestamp 1679581782
transform 1 0 74976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_782
timestamp 1679577901
transform 1 0 75648 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_786
timestamp 1677580104
transform 1 0 76032 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_808
timestamp 1679581782
transform 1 0 78144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_815
timestamp 1679581782
transform 1 0 78816 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_822
timestamp 1677579658
transform 1 0 79488 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_574
timestamp 1679577901
transform 1 0 55680 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_578
timestamp 1677579658
transform 1 0 56064 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_632
timestamp 1679577901
transform 1 0 61248 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_690
timestamp 1677580104
transform 1 0 66816 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_47_774
timestamp 1679577901
transform 1 0 74880 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_4  FILLER_47_819
timestamp 1679577901
transform 1 0 79200 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_581
timestamp 1677579658
transform 1 0 56352 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_623
timestamp 1677579658
transform 1 0 60384 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_658
timestamp 1677580104
transform 1 0 63744 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_660
timestamp 1677579658
transform 1 0 63936 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_667
timestamp 1677579658
transform 1 0 64608 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_753
timestamp 1677580104
transform 1 0 72864 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_789
timestamp 1677579658
transform 1 0 76320 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_820
timestamp 1677580104
transform 1 0 79296 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_822
timestamp 1677579658
transform 1 0 79488 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 1632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_25
timestamp 1679581782
transform 1 0 2976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_32
timestamp 1679581782
transform 1 0 3648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_39
timestamp 1679581782
transform 1 0 4320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_46
timestamp 1679581782
transform 1 0 4992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_53
timestamp 1679581782
transform 1 0 5664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_60
timestamp 1679581782
transform 1 0 6336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_67
timestamp 1679581782
transform 1 0 7008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_74
timestamp 1679581782
transform 1 0 7680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_81
timestamp 1679581782
transform 1 0 8352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_88
timestamp 1679581782
transform 1 0 9024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_95
timestamp 1679581782
transform 1 0 9696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_102
timestamp 1679581782
transform 1 0 10368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_109
timestamp 1679581782
transform 1 0 11040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_116
timestamp 1679581782
transform 1 0 11712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_123
timestamp 1679581782
transform 1 0 12384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_130
timestamp 1679581782
transform 1 0 13056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_137
timestamp 1679581782
transform 1 0 13728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_144
timestamp 1679581782
transform 1 0 14400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_151
timestamp 1679581782
transform 1 0 15072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_158
timestamp 1679581782
transform 1 0 15744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_165
timestamp 1679581782
transform 1 0 16416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_172
timestamp 1679581782
transform 1 0 17088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_179
timestamp 1679581782
transform 1 0 17760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_186
timestamp 1679581782
transform 1 0 18432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_193
timestamp 1679581782
transform 1 0 19104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_200
timestamp 1679581782
transform 1 0 19776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_207
timestamp 1679581782
transform 1 0 20448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_214
timestamp 1679581782
transform 1 0 21120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_221
timestamp 1679581782
transform 1 0 21792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_228
timestamp 1679581782
transform 1 0 22464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_235
timestamp 1679581782
transform 1 0 23136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_242
timestamp 1679581782
transform 1 0 23808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_249
timestamp 1679581782
transform 1 0 24480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_256
timestamp 1679581782
transform 1 0 25152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_263
timestamp 1679581782
transform 1 0 25824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_270
timestamp 1679581782
transform 1 0 26496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_277
timestamp 1679581782
transform 1 0 27168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_284
timestamp 1679581782
transform 1 0 27840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_291
timestamp 1679581782
transform 1 0 28512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_298
timestamp 1679581782
transform 1 0 29184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_305
timestamp 1679581782
transform 1 0 29856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_312
timestamp 1679581782
transform 1 0 30528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_319
timestamp 1679581782
transform 1 0 31200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_326
timestamp 1679581782
transform 1 0 31872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_333
timestamp 1679581782
transform 1 0 32544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_340
timestamp 1679581782
transform 1 0 33216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_347
timestamp 1679581782
transform 1 0 33888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_354
timestamp 1679581782
transform 1 0 34560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_361
timestamp 1679581782
transform 1 0 35232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_368
timestamp 1679581782
transform 1 0 35904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_375
timestamp 1679581782
transform 1 0 36576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_382
timestamp 1679581782
transform 1 0 37248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_389
timestamp 1679581782
transform 1 0 37920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_396
timestamp 1679581782
transform 1 0 38592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_403
timestamp 1679581782
transform 1 0 39264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_410
timestamp 1679581782
transform 1 0 39936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_417
timestamp 1679581782
transform 1 0 40608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_424
timestamp 1679581782
transform 1 0 41280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_431
timestamp 1679581782
transform 1 0 41952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_438
timestamp 1679581782
transform 1 0 42624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_445
timestamp 1679581782
transform 1 0 43296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_452
timestamp 1679581782
transform 1 0 43968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_459
timestamp 1679581782
transform 1 0 44640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_466
timestamp 1679581782
transform 1 0 45312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_473
timestamp 1679581782
transform 1 0 45984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_480
timestamp 1679581782
transform 1 0 46656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_487
timestamp 1679581782
transform 1 0 47328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_494
timestamp 1679581782
transform 1 0 48000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_501
timestamp 1679581782
transform 1 0 48672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_508
timestamp 1679581782
transform 1 0 49344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_515
timestamp 1679581782
transform 1 0 50016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_522
timestamp 1679581782
transform 1 0 50688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_529
timestamp 1679581782
transform 1 0 51360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_536
timestamp 1679581782
transform 1 0 52032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_543
timestamp 1679581782
transform 1 0 52704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_550
timestamp 1679581782
transform 1 0 53376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_557
timestamp 1679581782
transform 1 0 54048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_564
timestamp 1679581782
transform 1 0 54720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_571
timestamp 1679581782
transform 1 0 55392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_578
timestamp 1679581782
transform 1 0 56064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_585
timestamp 1679581782
transform 1 0 56736 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_592
timestamp 1677579658
transform 1 0 57408 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_596
timestamp 1679581782
transform 1 0 57792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_603
timestamp 1679581782
transform 1 0 58464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_610
timestamp 1679581782
transform 1 0 59136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_620
timestamp 1679581782
transform 1 0 60096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_627
timestamp 1679577901
transform 1 0 60768 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_636
timestamp 1679581782
transform 1 0 61632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_643
timestamp 1679581782
transform 1 0 62304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_650
timestamp 1679581782
transform 1 0 62976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_657
timestamp 1679581782
transform 1 0 63648 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_664
timestamp 1677579658
transform 1 0 64320 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_694
timestamp 1677580104
transform 1 0 67200 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_763
timestamp 1677579658
transform 1 0 73824 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_774
timestamp 1679577901
transform 1 0 74880 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_778
timestamp 1677580104
transform 1 0 75264 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_796
timestamp 1677580104
transform 1 0 76992 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_802
timestamp 1679581782
transform 1 0 77568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_809
timestamp 1679581782
transform 1 0 78240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_816
timestamp 1679581782
transform 1 0 78912 0 -1 38556
box -48 -56 720 834
use sg13g2_tiehi  heichips25_pudding_228
timestamp 1680000651
transform -1 0 1344 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_229
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_230
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_231
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_232
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_233
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_234
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 576 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 576 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 576 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 576 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 576 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
use analog_wires  wires
timestamp 0
transform 1 0 80000 0 1 800
box 0 0 1 1
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 16316 630 16756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 28316 630 28756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 40316 630 40756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 52316 630 52756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64316 630 64756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 76316 630 76756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 15076 712 15516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 27076 712 27516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 39076 712 39516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 51076 712 51516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63076 712 63516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 75076 712 75516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 99920 21586 100000 21726 0 FreeSans 640 0 0 0 i_in
port 4 nsew signal bidirectional
flabel metal3 s 99920 19949 100000 20089 0 FreeSans 640 0 0 0 i_out
port 5 nsew signal bidirectional
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 6 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 7 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 8 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 9 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 10 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 11 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 12 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 13 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 14 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 15 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 16 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 17 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 18 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 19 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 20 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 21 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 22 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 23 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 24 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 25 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 26 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 27 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 28 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 29 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 30 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 31 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 32 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 33 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 34 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 35 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 36 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 37 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 38 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 39 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 40 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 41 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 42 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 43 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 44 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 45 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 46 nsew signal output
rlabel via5 76620 22479 76620 22479 0 VGND
rlabel via5 75380 19603 75380 19603 0 VPWR
rlabel metal2 54048 16926 54048 16926 0 _0000_
rlabel metal2 62832 28140 62832 28140 0 _0001_
rlabel metal3 61872 23772 61872 23772 0 _0002_
rlabel metal3 59952 23604 59952 23604 0 _0003_
rlabel metal2 56832 23856 56832 23856 0 _0004_
rlabel metal2 63165 22828 63165 22828 0 _0005_
rlabel metal2 62765 22828 62765 22828 0 _0006_
rlabel metal2 62365 22828 62365 22828 0 _0007_
rlabel metal3 61942 22764 61942 22764 0 _0008_
rlabel metal3 61022 22764 61022 22764 0 _0009_
rlabel metal2 61165 22828 61165 22828 0 _0010_
rlabel metal4 36768 15498 36768 15498 0 _0011_
rlabel metal2 60765 22732 60765 22732 0 _0012_
rlabel metal2 60278 22764 60278 22764 0 _0013_
rlabel metal3 42336 21462 42336 21462 0 _0014_
rlabel metal2 59565 22828 59565 22828 0 _0015_
rlabel via3 59150 22764 59150 22764 0 _0016_
rlabel metal2 58765 22828 58765 22828 0 _0017_
rlabel metal3 58174 22932 58174 22932 0 _0018_
rlabel metal2 39456 22050 39456 22050 0 _0019_
rlabel metal3 38160 22092 38160 22092 0 _0020_
rlabel metal2 37776 22092 37776 22092 0 _0021_
rlabel metal3 39984 16968 39984 16968 0 _0022_
rlabel metal3 55968 22974 55968 22974 0 _0023_
rlabel metal5 5800 21546 5800 21546 0 _0024_
rlabel metal2 7680 18480 7680 18480 0 _0025_
rlabel metal3 15360 18690 15360 18690 0 _0026_
rlabel metal2 13632 20874 13632 20874 0 _0027_
rlabel metal4 10944 20664 10944 20664 0 _0028_
rlabel metal2 8064 19530 8064 19530 0 _0029_
rlabel metal4 5952 21504 5952 21504 0 _0030_
rlabel metal2 39648 15582 39648 15582 0 _0031_
rlabel metal2 42624 14952 42624 14952 0 _0032_
rlabel metal4 59712 16296 59712 16296 0 _0033_
rlabel metal2 57600 14028 57600 14028 0 _0034_
rlabel metal2 42720 11172 42720 11172 0 _0035_
rlabel metal2 57408 14028 57408 14028 0 _0036_
rlabel metal3 58944 13650 58944 13650 0 _0037_
rlabel metal3 61536 14196 61536 14196 0 _0038_
rlabel metal2 54475 17336 54475 17336 0 _0039_
rlabel metal4 61920 16590 61920 16590 0 _0040_
rlabel metal4 62016 16590 62016 16590 0 _0041_
rlabel metal3 58176 14952 58176 14952 0 _0042_
rlabel metal3 60144 16464 60144 16464 0 _0043_
rlabel metal2 57312 16632 57312 16632 0 _0044_
rlabel metal4 60576 15666 60576 15666 0 _0045_
rlabel metal4 56352 16800 56352 16800 0 _0046_
rlabel metal2 64875 17366 64875 17366 0 _0047_
rlabel metal2 58512 14196 58512 14196 0 _0048_
rlabel metal2 58128 5712 58128 5712 0 _0049_
rlabel metal2 54816 16422 54816 16422 0 _0050_
rlabel metal2 62304 6426 62304 6426 0 _0051_
rlabel metal4 66336 15750 66336 15750 0 _0052_
rlabel metal2 62208 7224 62208 7224 0 _0053_
rlabel metal4 60480 16548 60480 16548 0 _0054_
rlabel metal2 67680 16338 67680 16338 0 _0055_
rlabel metal2 59616 16758 59616 16758 0 _0056_
rlabel metal3 62256 15540 62256 15540 0 _0057_
rlabel metal2 62592 15792 62592 15792 0 _0058_
rlabel metal2 63264 11550 63264 11550 0 _0059_
rlabel metal2 69696 12810 69696 12810 0 _0060_
rlabel metal2 55200 16842 55200 16842 0 _0061_
rlabel metal4 70176 15456 70176 15456 0 _0062_
rlabel metal2 65760 16506 65760 16506 0 _0063_
rlabel metal2 66720 16002 66720 16002 0 _0064_
rlabel metal2 69984 15960 69984 15960 0 _0065_
rlabel metal3 68736 16212 68736 16212 0 _0066_
rlabel metal4 72576 15750 72576 15750 0 _0067_
rlabel metal3 70704 15456 70704 15456 0 _0068_
rlabel metal2 66144 16506 66144 16506 0 _0069_
rlabel metal2 72576 16002 72576 16002 0 _0070_
rlabel metal2 73728 16422 73728 16422 0 _0071_
rlabel metal2 55680 16674 55680 16674 0 _0072_
rlabel metal2 74016 16758 74016 16758 0 _0073_
rlabel metal3 74256 13440 74256 13440 0 _0074_
rlabel metal3 73920 16044 73920 16044 0 _0075_
rlabel metal3 74981 17136 74981 17136 0 _0076_
rlabel metal3 75456 7056 75456 7056 0 _0077_
rlabel metal3 75264 15960 75264 15960 0 _0078_
rlabel metal3 75312 2856 75312 2856 0 _0079_
rlabel metal3 76800 17262 76800 17262 0 _0080_
rlabel metal3 77088 14364 77088 14364 0 _0081_
rlabel metal3 78384 15876 78384 15876 0 _0082_
rlabel metal3 56064 16422 56064 16422 0 _0083_
rlabel metal2 78061 17052 78061 17052 0 _0084_
rlabel metal3 78288 12264 78288 12264 0 _0085_
rlabel metal3 76608 14070 76608 14070 0 _0086_
rlabel metal2 77856 16800 77856 16800 0 _0087_
rlabel metal2 79165 22828 79165 22828 0 _0088_
rlabel metal2 78765 22732 78765 22732 0 _0089_
rlabel metal2 78365 22828 78365 22828 0 _0090_
rlabel via3 77958 22764 77958 22764 0 _0091_
rlabel metal2 76128 31374 76128 31374 0 _0092_
rlabel metal2 77165 22690 77165 22690 0 _0093_
rlabel metal4 40896 16296 40896 16296 0 _0094_
rlabel metal2 75744 36414 75744 36414 0 _0095_
rlabel metal2 76342 22764 76342 22764 0 _0096_
rlabel metal3 75312 33432 75312 33432 0 _0097_
rlabel metal2 75510 22764 75510 22764 0 _0098_
rlabel metal2 75165 22828 75165 22828 0 _0099_
rlabel metal3 74486 22764 74486 22764 0 _0100_
rlabel metal3 74238 23016 74238 23016 0 _0101_
rlabel metal2 73942 22932 73942 22932 0 _0102_
rlabel metal2 73565 22828 73565 22828 0 _0103_
rlabel metal2 73165 22828 73165 22828 0 _0104_
rlabel metal4 38304 17010 38304 17010 0 _0105_
rlabel metal2 72765 22828 72765 22828 0 _0106_
rlabel metal2 62976 23982 62976 23982 0 _0107_
rlabel metal2 71965 22828 71965 22828 0 _0108_
rlabel metal3 71302 22848 71302 22848 0 _0109_
rlabel metal2 71150 22764 71150 22764 0 _0110_
rlabel metal2 66912 33642 66912 33642 0 _0111_
rlabel metal2 70224 25872 70224 25872 0 _0112_
rlabel metal2 65760 35364 65760 35364 0 _0113_
rlabel metal2 61824 35196 61824 35196 0 _0114_
rlabel metal2 69165 22828 69165 22828 0 _0115_
rlabel metal4 34752 17640 34752 17640 0 _0116_
rlabel metal2 60000 34020 60000 34020 0 _0117_
rlabel metal2 65280 24360 65280 24360 0 _0118_
rlabel metal2 67965 22828 67965 22828 0 _0119_
rlabel metal2 62208 24192 62208 24192 0 _0120_
rlabel metal2 57504 30912 57504 30912 0 _0121_
rlabel metal2 56448 24108 56448 24108 0 _0122_
rlabel metal2 66365 22690 66365 22690 0 _0123_
rlabel metal3 65382 22932 65382 22932 0 _0124_
rlabel metal2 55200 28056 55200 28056 0 _0125_
rlabel metal2 56256 27846 56256 27846 0 _0126_
rlabel metal4 33216 16548 33216 16548 0 _0127_
rlabel metal2 40704 20076 40704 20076 0 _0128_
rlabel metal2 45408 19908 45408 19908 0 _0129_
rlabel metal2 48432 20076 48432 20076 0 _0130_
rlabel metal2 49920 17514 49920 17514 0 _0131_
rlabel metal2 43104 15750 43104 15750 0 _0132_
rlabel metal2 42912 17262 42912 17262 0 _0133_
rlabel metal2 39744 20076 39744 20076 0 _0134_
rlabel metal2 36960 19908 36960 19908 0 _0135_
rlabel metal2 32640 18396 32640 18396 0 _0136_
rlabel metal3 31968 16380 31968 16380 0 _0137_
rlabel metal3 34704 14700 34704 14700 0 _0138_
rlabel metal2 37248 14658 37248 14658 0 _0139_
rlabel metal3 39168 13188 39168 13188 0 _0140_
rlabel metal3 41616 13188 41616 13188 0 _0141_
rlabel metal3 44352 12684 44352 12684 0 _0142_
rlabel metal2 45888 11172 45888 11172 0 _0143_
rlabel metal2 42624 9954 42624 9954 0 _0144_
rlabel metal2 45504 8442 45504 8442 0 _0145_
rlabel metal2 47904 7812 47904 7812 0 _0146_
rlabel metal2 49920 9156 49920 9156 0 _0147_
rlabel metal3 49584 10836 49584 10836 0 _0148_
rlabel metal2 48672 13902 48672 13902 0 _0149_
rlabel metal3 51744 14868 51744 14868 0 _0150_
rlabel metal2 54144 13860 54144 13860 0 _0151_
rlabel metal2 55776 11865 55776 11865 0 _0152_
rlabel metal3 54240 10332 54240 10332 0 _0153_
rlabel metal2 54336 7896 54336 7896 0 _0154_
rlabel metal3 52080 4788 52080 4788 0 _0155_
rlabel metal2 53856 4158 53856 4158 0 _0156_
rlabel metal3 56304 2772 56304 2772 0 _0157_
rlabel metal2 59136 2394 59136 2394 0 _0158_
rlabel metal3 60480 1092 60480 1092 0 _0159_
rlabel metal2 60960 4746 60960 4746 0 _0160_
rlabel metal3 58512 7140 58512 7140 0 _0161_
rlabel metal3 57936 9492 57936 9492 0 _0162_
rlabel metal3 57984 13860 57984 13860 0 _0163_
rlabel metal2 60000 13986 60000 13986 0 _0164_
rlabel metal3 61248 13356 61248 13356 0 _0165_
rlabel metal2 60672 10500 60672 10500 0 _0166_
rlabel metal2 63072 8442 63072 8442 0 _0167_
rlabel metal2 66144 6132 66144 6132 0 _0168_
rlabel metal2 63264 3654 63264 3654 0 _0169_
rlabel metal2 65088 2394 65088 2394 0 _0170_
rlabel metal2 67776 1428 67776 1428 0 _0171_
rlabel metal2 67968 4788 67968 4788 0 _0172_
rlabel metal2 68160 8190 68160 8190 0 _0173_
rlabel metal2 67200 10668 67200 10668 0 _0174_
rlabel metal2 64416 12180 64416 12180 0 _0175_
rlabel metal2 67056 14028 67056 14028 0 _0176_
rlabel metal2 68640 13524 68640 13524 0 _0177_
rlabel metal3 70896 13356 70896 13356 0 _0178_
rlabel metal3 70944 11004 70944 11004 0 _0179_
rlabel metal2 72144 8652 72144 8652 0 _0180_
rlabel metal3 70896 6300 70896 6300 0 _0181_
rlabel metal2 72480 5418 72480 5418 0 _0182_
rlabel metal3 70704 4284 70704 4284 0 _0183_
rlabel metal2 72000 2562 72000 2562 0 _0184_
rlabel metal2 76032 1806 76032 1806 0 _0185_
rlabel metal2 77184 3654 77184 3654 0 _0186_
rlabel metal2 77088 6342 77088 6342 0 _0187_
rlabel metal2 76896 8736 76896 8736 0 _0188_
rlabel metal3 75936 11004 75936 11004 0 _0189_
rlabel metal3 75552 13356 75552 13356 0 _0190_
rlabel metal2 75360 15414 75360 15414 0 _0191_
rlabel metal2 75072 24822 75072 24822 0 _0192_
rlabel metal2 75840 26082 75840 26082 0 _0193_
rlabel metal3 75456 27468 75456 27468 0 _0194_
rlabel metal2 75072 30576 75072 30576 0 _0195_
rlabel metal2 76416 32718 76416 32718 0 _0196_
rlabel metal2 77280 34356 77280 34356 0 _0197_
rlabel metal2 76320 36708 76320 36708 0 _0198_
rlabel metal2 73728 36708 73728 36708 0 _0199_
rlabel metal2 72000 36582 72000 36582 0 _0200_
rlabel metal2 71520 35112 71520 35112 0 _0201_
rlabel metal2 71712 32382 71712 32382 0 _0202_
rlabel metal3 71904 30660 71904 30660 0 _0203_
rlabel metal2 70848 29022 70848 29022 0 _0204_
rlabel metal2 70944 27636 70944 27636 0 _0205_
rlabel metal2 70752 26334 70752 26334 0 _0206_
rlabel metal3 67584 26124 67584 26124 0 _0207_
rlabel metal3 65808 26124 65808 26124 0 _0208_
rlabel metal2 62400 27300 62400 27300 0 _0209_
rlabel metal2 63072 28434 63072 28434 0 _0210_
rlabel metal2 64032 30450 64032 30450 0 _0211_
rlabel metal3 66048 32004 66048 32004 0 _0212_
rlabel metal3 66864 35784 66864 35784 0 _0213_
rlabel metal2 67296 36918 67296 36918 0 _0214_
rlabel metal2 64320 37204 64320 37204 0 _0215_
rlabel metal2 59808 36918 59808 36918 0 _0216_
rlabel metal2 56736 37023 56736 37023 0 _0217_
rlabel metal2 58560 35406 58560 35406 0 _0218_
rlabel metal2 61632 35154 61632 35154 0 _0219_
rlabel metal2 62976 31962 62976 31962 0 _0220_
rlabel metal3 60576 32172 60576 32172 0 _0221_
rlabel metal2 56928 32298 56928 32298 0 _0222_
rlabel metal3 55056 33432 55056 33432 0 _0223_
rlabel metal3 51936 34524 51936 34524 0 _0224_
rlabel metal2 50592 31836 50592 31836 0 _0225_
rlabel metal2 53664 31122 53664 31122 0 _0226_
rlabel metal2 56640 29358 56640 29358 0 _0227_
rlabel metal2 59328 29064 59328 29064 0 _0228_
rlabel metal2 61296 26796 61296 26796 0 _0229_
rlabel metal3 59328 26208 59328 26208 0 _0230_
rlabel metal2 56352 26082 56352 26082 0 _0231_
rlabel metal2 53856 26166 53856 26166 0 _0232_
rlabel metal2 52224 27594 52224 27594 0 _0233_
rlabel metal2 47808 29946 47808 29946 0 _0234_
rlabel metal2 45408 28644 45408 28644 0 _0235_
rlabel metal2 47808 26586 47808 26586 0 _0236_
rlabel metal2 48864 24528 48864 24528 0 _0237_
rlabel metal2 49920 22302 49920 22302 0 _0238_
rlabel metal2 46368 21798 46368 21798 0 _0239_
rlabel metal3 40848 23100 40848 23100 0 _0240_
rlabel metal3 41952 24696 41952 24696 0 _0241_
rlabel metal2 42144 26334 42144 26334 0 _0242_
rlabel metal2 42048 28434 42048 28434 0 _0243_
rlabel metal2 39936 27006 39936 27006 0 _0244_
rlabel metal2 37632 24276 37632 24276 0 _0245_
rlabel metal2 36192 22764 36192 22764 0 _0246_
rlabel metal2 35808 21588 35808 21588 0 _0247_
rlabel metal2 32256 20874 32256 20874 0 _0248_
rlabel metal2 6432 18060 6432 18060 0 _0249_
rlabel metal3 6912 17052 6912 17052 0 _0250_
rlabel metal2 10560 17262 10560 17262 0 _0251_
rlabel metal2 12672 18438 12672 18438 0 _0252_
rlabel metal3 10992 20916 10992 20916 0 _0253_
rlabel metal2 7680 20538 7680 20538 0 _0254_
rlabel metal2 3168 19950 3168 19950 0 _0255_
rlabel metal3 42288 20412 42288 20412 0 _0256_
rlabel metal2 46176 17892 46176 17892 0 _0257_
rlabel metal2 50304 18942 50304 18942 0 _0258_
rlabel metal2 50592 16464 50592 16464 0 _0259_
rlabel metal2 46512 16212 46512 16212 0 _0260_
rlabel metal2 44544 17892 44544 17892 0 _0261_
rlabel metal2 39936 18564 39936 18564 0 _0262_
rlabel metal2 36864 18564 36864 18564 0 _0263_
rlabel metal2 34224 18732 34224 18732 0 _0264_
rlabel metal2 32928 17346 32928 17346 0 _0265_
rlabel metal2 35520 16632 35520 16632 0 _0266_
rlabel metal3 37872 16128 37872 16128 0 _0267_
rlabel metal2 40032 15666 40032 15666 0 _0268_
rlabel metal2 42432 14868 42432 14868 0 _0269_
rlabel metal3 45648 14616 45648 14616 0 _0270_
rlabel metal2 46656 12990 46656 12990 0 _0271_
rlabel metal2 42480 11172 42480 11172 0 _0272_
rlabel metal2 45312 10080 45312 10080 0 _0273_
rlabel metal2 48048 9660 48048 9660 0 _0274_
rlabel metal2 51744 10458 51744 10458 0 _0275_
rlabel metal2 51360 12642 51360 12642 0 _0276_
rlabel metal3 49056 14700 49056 14700 0 _0277_
rlabel metal2 52416 15708 52416 15708 0 _0278_
rlabel metal2 55392 15834 55392 15834 0 _0279_
rlabel metal2 56256 13272 56256 13272 0 _0280_
rlabel metal3 56016 11004 56016 11004 0 _0281_
rlabel metal2 55488 8148 55488 8148 0 _0282_
rlabel metal2 52128 7140 52128 7140 0 _0283_
rlabel metal3 55344 6552 55344 6552 0 _0284_
rlabel metal2 57312 4956 57312 4956 0 _0285_
rlabel metal3 60432 4032 60432 4032 0 _0286_
rlabel metal2 62400 2226 62400 2226 0 _0287_
rlabel metal3 61056 6468 61056 6468 0 _0288_
rlabel metal2 60096 8358 60096 8358 0 _0289_
rlabel metal2 58944 11298 58944 11298 0 _0290_
rlabel metal2 57984 15708 57984 15708 0 _0291_
rlabel metal2 61056 15708 61056 15708 0 _0292_
rlabel metal2 62784 14616 62784 14616 0 _0293_
rlabel metal2 62976 11382 62976 11382 0 _0294_
rlabel metal2 64032 9618 64032 9618 0 _0295_
rlabel metal2 66144 7266 66144 7266 0 _0296_
rlabel metal2 65376 5250 65376 5250 0 _0297_
rlabel metal3 66192 3444 66192 3444 0 _0298_
rlabel metal2 68832 2226 68832 2226 0 _0299_
rlabel metal3 68208 6468 68208 6468 0 _0300_
rlabel metal2 68256 9786 68256 9786 0 _0301_
rlabel metal2 67584 11592 67584 11592 0 _0302_
rlabel metal2 64608 14154 64608 14154 0 _0303_
rlabel metal2 66912 15918 66912 15918 0 _0304_
rlabel metal2 70368 15666 70368 15666 0 _0305_
rlabel metal2 71856 14112 71856 14112 0 _0306_
rlabel metal2 73008 11676 73008 11676 0 _0307_
rlabel metal2 72816 10164 72816 10164 0 _0308_
rlabel metal2 72672 8274 72672 8274 0 _0309_
rlabel metal2 73248 6594 73248 6594 0 _0310_
rlabel metal2 72768 3822 72768 3822 0 _0311_
rlabel metal3 72528 1008 72528 1008 0 _0312_
rlabel metal2 76992 1764 76992 1764 0 _0313_
rlabel metal2 75840 4284 75840 4284 0 _0314_
rlabel metal3 76080 7140 76080 7140 0 _0315_
rlabel metal2 75360 9786 75360 9786 0 _0316_
rlabel metal2 76992 12096 76992 12096 0 _0317_
rlabel metal2 76896 14028 76896 14028 0 _0318_
rlabel metal3 76176 14700 76176 14700 0 _0319_
rlabel metal3 76320 23604 76320 23604 0 _0320_
rlabel metal2 76800 25704 76800 25704 0 _0321_
rlabel metal2 77136 26796 77136 26796 0 _0322_
rlabel metal3 76992 29274 76992 29274 0 _0323_
rlabel metal2 76128 31164 76128 31164 0 _0324_
rlabel metal2 76896 33894 76896 33894 0 _0325_
rlabel metal3 76320 36708 76320 36708 0 _0326_
rlabel metal2 74112 37086 74112 37086 0 _0327_
rlabel metal3 73104 35280 73104 35280 0 _0328_
rlabel metal3 72144 34272 72144 34272 0 _0329_
rlabel metal2 72768 31710 72768 31710 0 _0330_
rlabel metal2 72480 30954 72480 30954 0 _0331_
rlabel metal3 72000 28308 72000 28308 0 _0332_
rlabel metal2 71808 26502 71808 26502 0 _0333_
rlabel metal2 71232 23940 71232 23940 0 _0334_
rlabel metal2 69120 24192 69120 24192 0 _0335_
rlabel metal2 66336 23688 66336 23688 0 _0336_
rlabel metal2 63264 24612 63264 24612 0 _0337_
rlabel metal2 66000 27804 66000 27804 0 _0338_
rlabel metal2 66336 29358 66336 29358 0 _0339_
rlabel metal3 67296 31164 67296 31164 0 _0340_
rlabel metal3 67440 33684 67440 33684 0 _0341_
rlabel metal2 70224 37380 70224 37380 0 _0342_
rlabel metal2 64800 36288 64800 36288 0 _0343_
rlabel metal2 60864 37086 60864 37086 0 _0344_
rlabel metal3 55536 35280 55536 35280 0 _0345_
rlabel metal2 58704 34188 58704 34188 0 _0346_
rlabel metal2 64032 34062 64032 34062 0 _0347_
rlabel metal2 63264 31374 63264 31374 0 _0348_
rlabel metal2 61344 30786 61344 30786 0 _0349_
rlabel metal2 57888 30786 57888 30786 0 _0350_
rlabel metal3 55152 33348 55152 33348 0 _0351_
rlabel metal2 52752 34272 52752 34272 0 _0352_
rlabel metal3 50448 30660 50448 30660 0 _0353_
rlabel metal2 53568 29148 53568 29148 0 _0354_
rlabel metal2 56544 28224 56544 28224 0 _0355_
rlabel metal2 61536 28728 61536 28728 0 _0356_
rlabel metal2 60960 24486 60960 24486 0 _0357_
rlabel metal2 59328 24192 59328 24192 0 _0358_
rlabel metal2 56640 24192 56640 24192 0 _0359_
rlabel metal2 53856 23982 53856 23982 0 _0360_
rlabel metal2 53184 27888 53184 27888 0 _0361_
rlabel metal2 48192 28602 48192 28602 0 _0362_
rlabel metal3 48672 27636 48672 27636 0 _0363_
rlabel metal3 46800 23772 46800 23772 0 _0364_
rlabel metal2 51504 23772 51504 23772 0 _0365_
rlabel metal2 50016 21966 50016 21966 0 _0366_
rlabel metal2 46368 23100 46368 23100 0 _0367_
rlabel metal2 42624 21714 42624 21714 0 _0368_
rlabel metal2 43776 23268 43776 23268 0 _0369_
rlabel metal2 44448 25704 44448 25704 0 _0370_
rlabel metal2 42816 28434 42816 28434 0 _0371_
rlabel metal2 39936 26124 39936 26124 0 _0372_
rlabel metal2 39168 23898 39168 23898 0 _0373_
rlabel metal2 37248 22302 37248 22302 0 _0374_
rlabel metal3 37344 21672 37344 21672 0 _0375_
rlabel metal3 31200 21672 31200 21672 0 _0376_
rlabel metal2 4896 21588 4896 21588 0 _0377_
rlabel metal2 7776 18438 7776 18438 0 _0378_
rlabel metal2 15648 18564 15648 18564 0 _0379_
rlabel metal2 13680 20580 13680 20580 0 _0380_
rlabel metal2 11184 20748 11184 20748 0 _0381_
rlabel metal2 7872 20874 7872 20874 0 _0382_
rlabel metal2 4032 20580 4032 20580 0 _0383_
rlabel metal3 56064 13020 56064 13020 0 _0384_
rlabel metal2 55584 12990 55584 12990 0 _0385_
rlabel metal2 55584 10752 55584 10752 0 _0386_
rlabel metal2 55872 10290 55872 10290 0 _0387_
rlabel metal2 54912 10500 54912 10500 0 _0388_
rlabel metal3 55392 7980 55392 7980 0 _0389_
rlabel metal3 54720 7728 54720 7728 0 _0390_
rlabel metal3 54720 7896 54720 7896 0 _0391_
rlabel metal3 53040 6468 53040 6468 0 _0392_
rlabel metal3 52128 6300 52128 6300 0 _0393_
rlabel metal2 52512 4998 52512 4998 0 _0394_
rlabel metal2 55968 5712 55968 5712 0 _0395_
rlabel metal2 55200 5334 55200 5334 0 _0396_
rlabel metal2 54528 4788 54528 4788 0 _0397_
rlabel metal3 57504 4116 57504 4116 0 _0398_
rlabel metal2 56832 2856 56832 2856 0 _0399_
rlabel metal2 56448 2784 56448 2784 0 _0400_
rlabel metal3 60336 3444 60336 3444 0 _0401_
rlabel metal2 59808 3528 59808 3528 0 _0402_
rlabel metal2 59040 2730 59040 2730 0 _0403_
rlabel metal2 62592 1134 62592 1134 0 _0404_
rlabel metal3 62112 2772 62112 2772 0 _0405_
rlabel metal2 61056 2730 61056 2730 0 _0406_
rlabel metal2 61248 5964 61248 5964 0 _0407_
rlabel metal2 60912 5796 60912 5796 0 _0408_
rlabel metal2 61440 3990 61440 3990 0 _0409_
rlabel metal3 60096 7980 60096 7980 0 _0410_
rlabel metal2 59856 7728 59856 7728 0 _0411_
rlabel metal2 60000 6930 60000 6930 0 _0412_
rlabel metal2 59232 10500 59232 10500 0 _0413_
rlabel metal2 58896 10332 58896 10332 0 _0414_
rlabel metal2 58656 8778 58656 8778 0 _0415_
rlabel metal2 58560 15246 58560 15246 0 _0416_
rlabel metal2 58272 15582 58272 15582 0 _0417_
rlabel metal2 58416 10416 58416 10416 0 _0418_
rlabel metal2 61344 14784 61344 14784 0 _0419_
rlabel metal3 60864 14868 60864 14868 0 _0420_
rlabel metal2 60480 13524 60480 13524 0 _0421_
rlabel metal2 62880 13608 62880 13608 0 _0422_
rlabel metal2 62544 13440 62544 13440 0 _0423_
rlabel metal3 61872 13272 61872 13272 0 _0424_
rlabel metal3 63024 11004 63024 11004 0 _0425_
rlabel metal3 62688 10752 62688 10752 0 _0426_
rlabel metal2 61824 11277 61824 11277 0 _0427_
rlabel metal2 64224 8694 64224 8694 0 _0428_
rlabel metal2 63552 8778 63552 8778 0 _0429_
rlabel metal3 62832 8736 62832 8736 0 _0430_
rlabel metal2 65376 7728 65376 7728 0 _0431_
rlabel metal2 65616 7308 65616 7308 0 _0432_
rlabel metal2 64608 5796 64608 5796 0 _0433_
rlabel metal3 65232 4956 65232 4956 0 _0434_
rlabel metal2 64608 4956 64608 4956 0 _0435_
rlabel metal2 64416 3486 64416 3486 0 _0436_
rlabel metal2 65760 3024 65760 3024 0 _0437_
rlabel metal2 66048 2730 66048 2730 0 _0438_
rlabel metal3 64752 2688 64752 2688 0 _0439_
rlabel metal3 68976 1092 68976 1092 0 _0440_
rlabel metal2 68208 1764 68208 1764 0 _0441_
rlabel metal2 66816 2226 66816 2226 0 _0442_
rlabel metal2 69408 5712 69408 5712 0 _0443_
rlabel metal2 68640 5124 68640 5124 0 _0444_
rlabel metal2 68640 3528 68640 3528 0 _0445_
rlabel metal2 68832 8820 68832 8820 0 _0446_
rlabel metal2 68544 9324 68544 9324 0 _0447_
rlabel metal2 68256 5712 68256 5712 0 _0448_
rlabel metal2 67680 11214 67680 11214 0 _0449_
rlabel metal2 67392 11256 67392 11256 0 _0450_
rlabel metal2 67584 9702 67584 9702 0 _0451_
rlabel metal3 65760 12936 65760 12936 0 _0452_
rlabel metal2 65328 13440 65328 13440 0 _0453_
rlabel metal2 65664 11802 65664 11802 0 _0454_
rlabel metal3 67728 14700 67728 14700 0 _0455_
rlabel metal2 67248 14868 67248 14868 0 _0456_
rlabel metal2 66816 13314 66816 13314 0 _0457_
rlabel metal3 70752 14700 70752 14700 0 _0458_
rlabel metal2 70080 14406 70080 14406 0 _0459_
rlabel metal3 69456 13944 69456 13944 0 _0460_
rlabel metal3 72336 13188 72336 13188 0 _0461_
rlabel metal3 71472 13944 71472 13944 0 _0462_
rlabel metal2 71520 13818 71520 13818 0 _0463_
rlabel via2 73532 11676 73532 11676 0 _0464_
rlabel metal3 72432 11844 72432 11844 0 _0465_
rlabel metal2 71808 10878 71808 10878 0 _0466_
rlabel metal3 73248 9492 73248 9492 0 _0467_
rlabel metal2 72672 10395 72672 10395 0 _0468_
rlabel metal2 72096 9702 72096 9702 0 _0469_
rlabel metal2 73728 7560 73728 7560 0 _0470_
rlabel metal3 72144 7728 72144 7728 0 _0471_
rlabel metal2 71616 7056 71616 7056 0 _0472_
rlabel metal2 74304 5712 74304 5712 0 _0473_
rlabel metal2 72576 5754 72576 5754 0 _0474_
rlabel metal2 72384 5964 72384 5964 0 _0475_
rlabel metal2 74016 3696 74016 3696 0 _0476_
rlabel metal2 72624 4284 72624 4284 0 _0477_
rlabel metal2 71616 4074 71616 4074 0 _0478_
rlabel metal3 73344 2100 73344 2100 0 _0479_
rlabel metal2 72096 2058 72096 2058 0 _0480_
rlabel metal2 71904 2562 71904 2562 0 _0481_
rlabel metal2 76848 1092 76848 1092 0 _0482_
rlabel metal3 76032 2604 76032 2604 0 _0483_
rlabel metal2 75552 1806 75552 1806 0 _0484_
rlabel metal3 77040 4116 77040 4116 0 _0485_
rlabel metal2 76320 4116 76320 4116 0 _0486_
rlabel metal2 77328 2856 77328 2856 0 _0487_
rlabel metal3 77808 5628 77808 5628 0 _0488_
rlabel metal2 76608 6132 76608 6132 0 _0489_
rlabel metal2 77760 5754 77760 5754 0 _0490_
rlabel metal2 77280 8232 77280 8232 0 _0491_
rlabel metal2 76608 8862 76608 8862 0 _0492_
rlabel metal2 78336 7938 78336 7938 0 _0493_
rlabel metal2 77568 11760 77568 11760 0 _0494_
rlabel metal2 77280 11676 77280 11676 0 _0495_
rlabel metal2 78000 9660 78000 9660 0 _0496_
rlabel metal2 77568 13272 77568 13272 0 _0497_
rlabel metal2 76752 13440 76752 13440 0 _0498_
rlabel metal2 76512 12180 76512 12180 0 _0499_
rlabel metal2 76704 15120 76704 15120 0 _0500_
rlabel metal2 76032 14994 76032 14994 0 _0501_
rlabel metal3 75600 14196 75600 14196 0 _0502_
rlabel metal3 76992 23604 76992 23604 0 _0503_
rlabel metal2 75936 24486 75936 24486 0 _0504_
rlabel metal2 74928 24024 74928 24024 0 _0505_
rlabel metal3 76944 25284 76944 25284 0 _0506_
rlabel metal3 76560 25956 76560 25956 0 _0507_
rlabel metal2 75936 25536 75936 25536 0 _0508_
rlabel metal2 77664 27132 77664 27132 0 _0509_
rlabel metal2 77088 28434 77088 28434 0 _0510_
rlabel metal2 76320 27468 76320 27468 0 _0511_
rlabel metal2 77424 29316 77424 29316 0 _0512_
rlabel metal2 76128 29526 76128 29526 0 _0513_
rlabel metal3 76272 29316 76272 29316 0 _0514_
rlabel metal2 77568 31500 77568 31500 0 _0515_
rlabel metal2 76272 31332 76272 31332 0 _0516_
rlabel metal2 76800 31458 76800 31458 0 _0517_
rlabel metal3 78192 34356 78192 34356 0 _0518_
rlabel metal2 77184 33726 77184 33726 0 _0519_
rlabel metal2 77376 33558 77376 33558 0 _0520_
rlabel metal2 76608 35952 76608 35952 0 _0521_
rlabel metal3 76752 36624 76752 36624 0 _0522_
rlabel metal3 76944 36120 76944 36120 0 _0523_
rlabel metal2 74496 37800 74496 37800 0 _0524_
rlabel metal2 74208 36666 74208 36666 0 _0525_
rlabel metal2 73824 36876 73824 36876 0 _0526_
rlabel metal2 73824 35952 73824 35952 0 _0527_
rlabel metal2 72960 36246 72960 36246 0 _0528_
rlabel metal2 72288 36750 72288 36750 0 _0529_
rlabel metal2 71808 34104 71808 34104 0 _0530_
rlabel metal2 72000 34440 72000 34440 0 _0531_
rlabel metal2 71808 35406 71808 35406 0 _0532_
rlabel metal4 73632 31920 73632 31920 0 _0533_
rlabel metal2 72864 31500 72864 31500 0 _0534_
rlabel metal2 71616 32760 71616 32760 0 _0535_
rlabel metal3 72672 29820 72672 29820 0 _0536_
rlabel metal3 72240 30576 72240 30576 0 _0537_
rlabel metal2 72192 30702 72192 30702 0 _0538_
rlabel metal2 72768 28392 72768 28392 0 _0539_
rlabel metal2 71904 28602 71904 28602 0 _0540_
rlabel metal2 71232 29022 71232 29022 0 _0541_
rlabel metal2 72672 26838 72672 26838 0 _0542_
rlabel metal2 71904 26334 71904 26334 0 _0543_
rlabel metal4 70944 27678 70944 27678 0 _0544_
rlabel metal3 71616 25284 71616 25284 0 _0545_
rlabel metal2 71424 25452 71424 25452 0 _0546_
rlabel metal3 71136 26040 71136 26040 0 _0547_
rlabel metal2 69984 24108 69984 24108 0 _0548_
rlabel metal2 69120 25452 69120 25452 0 _0549_
rlabel metal2 69120 25998 69120 25998 0 _0550_
rlabel metal2 67008 24528 67008 24528 0 _0551_
rlabel metal2 66048 25242 66048 25242 0 _0552_
rlabel metal2 65856 25410 65856 25410 0 _0553_
rlabel metal2 64224 24108 64224 24108 0 _0554_
rlabel metal3 63408 25452 63408 25452 0 _0555_
rlabel metal2 64608 25746 64608 25746 0 _0556_
rlabel metal2 65376 27888 65376 27888 0 _0557_
rlabel metal2 65088 27846 65088 27846 0 _0558_
rlabel metal2 64416 27426 64416 27426 0 _0559_
rlabel metal3 66432 29820 66432 29820 0 _0560_
rlabel metal2 65952 29778 65952 29778 0 _0561_
rlabel metal2 65376 29946 65376 29946 0 _0562_
rlabel metal2 68448 31290 68448 31290 0 _0563_
rlabel metal2 67200 31626 67200 31626 0 _0564_
rlabel metal2 66240 31626 66240 31626 0 _0565_
rlabel metal3 68304 34356 68304 34356 0 _0566_
rlabel metal3 67200 34440 67200 34440 0 _0567_
rlabel via1 67401 33852 67401 33852 0 _0568_
rlabel metal3 68352 36708 68352 36708 0 _0569_
rlabel metal2 68160 36708 68160 36708 0 _0570_
rlabel metal2 67200 36582 67200 36582 0 _0571_
rlabel metal2 65280 35952 65280 35952 0 _0572_
rlabel metal2 64608 35952 64608 35952 0 _0573_
rlabel metal3 64848 37464 64848 37464 0 _0574_
rlabel metal2 61248 36288 61248 36288 0 _0575_
rlabel metal2 60672 36582 60672 36582 0 _0576_
rlabel metal2 59712 36750 59712 36750 0 _0577_
rlabel metal3 56928 35868 56928 35868 0 _0578_
rlabel metal2 56448 36498 56448 36498 0 _0579_
rlabel metal3 57216 35784 57216 35784 0 _0580_
rlabel metal2 59280 33852 59280 33852 0 _0581_
rlabel metal2 58656 35070 58656 35070 0 _0582_
rlabel metal2 58464 35406 58464 35406 0 _0583_
rlabel metal3 64128 33852 64128 33852 0 _0584_
rlabel metal3 62592 34482 62592 34482 0 _0585_
rlabel metal2 62400 34692 62400 34692 0 _0586_
rlabel metal2 63744 31626 63744 31626 0 _0587_
rlabel metal2 63552 32550 63552 32550 0 _0588_
rlabel metal2 63072 34188 63072 34188 0 _0589_
rlabel metal2 61536 31416 61536 31416 0 _0590_
rlabel metal2 60816 31500 60816 31500 0 _0591_
rlabel metal2 61056 32046 61056 32046 0 _0592_
rlabel metal3 57888 31332 57888 31332 0 _0593_
rlabel metal2 57888 31794 57888 31794 0 _0594_
rlabel metal2 58656 31836 58656 31836 0 _0595_
rlabel metal2 55296 33810 55296 33810 0 _0596_
rlabel metal2 55200 32886 55200 32886 0 _0597_
rlabel metal2 55392 32970 55392 32970 0 _0598_
rlabel metal3 52320 32844 52320 32844 0 _0599_
rlabel metal2 52032 34230 52032 34230 0 _0600_
rlabel metal3 52656 34440 52656 34440 0 _0601_
rlabel metal2 51456 29946 51456 29946 0 _0602_
rlabel metal2 50496 31290 50496 31290 0 _0603_
rlabel metal2 50688 32046 50688 32046 0 _0604_
rlabel metal2 54624 29988 54624 29988 0 _0605_
rlabel metal2 53952 30744 53952 30744 0 _0606_
rlabel metal2 52416 31500 52416 31500 0 _0607_
rlabel metal2 57504 28098 57504 28098 0 _0608_
rlabel metal2 56736 29022 56736 29022 0 _0609_
rlabel metal2 56544 29022 56544 29022 0 _0610_
rlabel metal3 61536 28308 61536 28308 0 _0611_
rlabel metal2 61344 28434 61344 28434 0 _0612_
rlabel metal2 59904 28644 59904 28644 0 _0613_
rlabel metal2 61248 26040 61248 26040 0 _0614_
rlabel metal2 61008 25956 61008 25956 0 _0615_
rlabel metal2 60768 27342 60768 27342 0 _0616_
rlabel metal2 59808 24318 59808 24318 0 _0617_
rlabel metal2 59136 24612 59136 24612 0 _0618_
rlabel metal2 59616 25998 59616 25998 0 _0619_
rlabel metal2 57120 24108 57120 24108 0 _0620_
rlabel metal2 57024 25788 57024 25788 0 _0621_
rlabel metal3 56976 25536 56976 25536 0 _0622_
rlabel metal2 54624 25368 54624 25368 0 _0623_
rlabel metal2 54144 24591 54144 24591 0 _0624_
rlabel metal2 53952 25998 53952 25998 0 _0625_
rlabel metal2 53472 27552 53472 27552 0 _0626_
rlabel metal3 52512 28476 52512 28476 0 _0627_
rlabel metal2 52128 27510 52128 27510 0 _0628_
rlabel metal2 48192 29190 48192 29190 0 _0629_
rlabel metal2 48528 28980 48528 28980 0 _0630_
rlabel metal2 51072 29568 51072 29568 0 _0631_
rlabel metal2 48192 27216 48192 27216 0 _0632_
rlabel metal2 48000 28413 48000 28413 0 _0633_
rlabel metal2 47232 29190 47232 29190 0 _0634_
rlabel metal2 48144 23772 48144 23772 0 _0635_
rlabel metal3 47616 25452 47616 25452 0 _0636_
rlabel metal3 47472 26880 47472 26880 0 _0637_
rlabel metal2 51072 24276 51072 24276 0 _0638_
rlabel metal3 50976 24024 50976 24024 0 _0639_
rlabel metal2 50400 24486 50400 24486 0 _0640_
rlabel metal2 50496 21924 50496 21924 0 _0641_
rlabel metal3 49728 22428 49728 22428 0 _0642_
rlabel metal2 50016 23310 50016 23310 0 _0643_
rlabel metal2 46752 22008 46752 22008 0 _0644_
rlabel metal2 46320 22512 46320 22512 0 _0645_
rlabel metal3 46992 21504 46992 21504 0 _0646_
rlabel metal3 42480 22092 42480 22092 0 _0647_
rlabel metal2 41760 22008 41760 22008 0 _0648_
rlabel metal2 41568 22386 41568 22386 0 _0649_
rlabel metal3 43872 23772 43872 23772 0 _0650_
rlabel metal2 42912 23730 42912 23730 0 _0651_
rlabel metal3 41856 23856 41856 23856 0 _0652_
rlabel metal2 45216 25620 45216 25620 0 _0653_
rlabel metal2 44592 25872 44592 25872 0 _0654_
rlabel metal2 43104 26124 43104 26124 0 _0655_
rlabel metal2 42720 28056 42720 28056 0 _0656_
rlabel metal2 42528 28560 42528 28560 0 _0657_
rlabel metal2 43104 27930 43104 27930 0 _0658_
rlabel metal2 40032 25620 40032 25620 0 _0659_
rlabel metal2 39744 25830 39744 25830 0 _0660_
rlabel metal3 40320 26880 40320 26880 0 _0661_
rlabel metal2 38688 23898 38688 23898 0 _0662_
rlabel metal3 38208 23856 38208 23856 0 _0663_
rlabel metal2 37920 23751 37920 23751 0 _0664_
rlabel metal2 36672 23352 36672 23352 0 _0665_
rlabel metal2 36288 22302 36288 22302 0 _0666_
rlabel metal2 36192 23604 36192 23604 0 _0667_
rlabel metal3 36672 20748 36672 20748 0 _0668_
rlabel metal3 36192 21336 36192 21336 0 _0669_
rlabel metal2 35616 21462 35616 21462 0 _0670_
rlabel metal3 31104 20076 31104 20076 0 _0671_
rlabel metal2 32544 20538 32544 20538 0 _0672_
rlabel metal2 32736 20937 32736 20937 0 _0673_
rlabel metal3 3792 18564 3792 18564 0 _0674_
rlabel metal2 4704 18522 4704 18522 0 _0675_
rlabel metal2 4896 18942 4896 18942 0 _0676_
rlabel metal2 6960 17724 6960 17724 0 _0677_
rlabel metal2 7104 18312 7104 18312 0 _0678_
rlabel metal2 6624 16716 6624 16716 0 _0679_
rlabel metal2 10080 18144 10080 18144 0 _0680_
rlabel metal2 10368 18144 10368 18144 0 _0681_
rlabel metal2 10464 16926 10464 16926 0 _0682_
rlabel metal3 12960 19236 12960 19236 0 _0683_
rlabel metal3 12912 19404 12912 19404 0 _0684_
rlabel metal3 12672 17976 12672 17976 0 _0685_
rlabel metal3 10272 19236 10272 19236 0 _0686_
rlabel metal2 11040 20118 11040 20118 0 _0687_
rlabel metal2 11040 19278 11040 19278 0 _0688_
rlabel metal2 8352 19656 8352 19656 0 _0689_
rlabel metal2 6912 19782 6912 19782 0 _0690_
rlabel metal2 7344 19488 7344 19488 0 _0691_
rlabel metal2 3552 20328 3552 20328 0 _0692_
rlabel metal2 3840 19950 3840 19950 0 _0693_
rlabel metal2 3552 19362 3552 19362 0 _0694_
rlabel metal3 10368 17724 10368 17724 0 _0695_
rlabel metal3 6288 3612 6288 3612 0 _0696_
rlabel metal2 10080 20454 10080 20454 0 _0697_
rlabel metal2 12480 18606 12480 18606 0 _0698_
rlabel metal2 6480 19488 6480 19488 0 _0699_
rlabel metal2 3024 19488 3024 19488 0 _0700_
rlabel via2 42432 20246 42432 20246 0 _0701_
rlabel via1 46656 18997 46656 18997 0 _0702_
rlabel via2 50112 18803 50112 18803 0 _0703_
rlabel via1 49920 16042 49920 16042 0 _0704_
rlabel via2 45888 16042 45888 16042 0 _0705_
rlabel via2 43392 17554 43392 17554 0 _0706_
rlabel via2 40512 19066 40512 19066 0 _0707_
rlabel metal3 36960 19236 36960 19236 0 _0708_
rlabel metal2 33312 18871 33312 18871 0 _0709_
rlabel metal2 32736 17180 32736 17180 0 _0710_
rlabel metal3 35664 15708 35664 15708 0 _0711_
rlabel metal2 38352 14952 38352 14952 0 _0712_
rlabel via2 40416 14198 40416 14198 0 _0713_
rlabel metal2 42048 14070 42048 14070 0 _0714_
rlabel metal2 45408 14200 45408 14200 0 _0715_
rlabel metal2 46416 11172 46416 11172 0 _0716_
rlabel metal2 44112 10164 44112 10164 0 _0717_
rlabel metal2 45696 8022 45696 8022 0 _0718_
rlabel metal2 48864 8524 48864 8524 0 _0719_
rlabel via2 51744 8413 51744 8413 0 _0720_
rlabel metal2 50880 11884 50880 11884 0 _0721_
rlabel metal2 49824 13522 49824 13522 0 _0722_
rlabel via2 52800 14530 52800 14530 0 _0723_
rlabel metal3 55392 13440 55392 13440 0 _0724_
rlabel metal2 56256 12308 56256 12308 0 _0725_
rlabel metal2 55392 9421 55392 9421 0 _0726_
rlabel metal2 54144 8064 54144 8064 0 _0727_
rlabel metal2 52224 4914 52224 4914 0 _0728_
rlabel metal3 55296 5124 55296 5124 0 _0729_
rlabel metal3 56736 2730 56736 2730 0 _0730_
rlabel metal2 60240 2856 60240 2856 0 _0731_
rlabel via2 62208 2434 62208 2434 0 _0732_
rlabel metal2 60768 4998 60768 4998 0 _0733_
rlabel via2 59424 8150 59424 8150 0 _0734_
rlabel via2 59424 9994 59424 9994 0 _0735_
rlabel metal2 58752 14167 58752 14167 0 _0736_
rlabel metal3 61728 13860 61728 13860 0 _0737_
rlabel via1 63072 12961 63072 12961 0 _0738_
rlabel metal2 62112 10962 62112 10962 0 _0739_
rlabel metal2 63264 8568 63264 8568 0 _0740_
rlabel metal2 64992 6594 64992 6594 0 _0741_
rlabel metal2 64992 3612 64992 3612 0 _0742_
rlabel metal2 65568 1861 65568 1861 0 _0743_
rlabel via2 68640 2171 68640 2171 0 _0744_
rlabel metal2 69216 4368 69216 4368 0 _0745_
rlabel metal2 67968 8148 67968 8148 0 _0746_
rlabel via2 67872 11243 67872 11243 0 _0747_
rlabel metal2 65760 13060 65760 13060 0 _0748_
rlabel metal3 67632 13188 67632 13188 0 _0749_
rlabel metal2 70560 14335 70560 14335 0 _0750_
rlabel metal3 71760 13356 71760 13356 0 _0751_
rlabel metal2 72096 10857 72096 10857 0 _0752_
rlabel metal2 73056 9284 73056 9284 0 _0753_
rlabel metal3 72528 7140 72528 7140 0 _0754_
rlabel metal2 73440 5542 73440 5542 0 _0755_
rlabel metal2 71904 3864 71904 3864 0 _0756_
rlabel via2 72864 2602 72864 2602 0 _0757_
rlabel metal2 77088 2155 77088 2155 0 _0758_
rlabel metal3 77520 3444 77520 3444 0 _0759_
rlabel via2 77664 5458 77664 5458 0 _0760_
rlabel metal2 77472 8345 77472 8345 0 _0761_
rlabel metal3 77712 10752 77712 10752 0 _0762_
rlabel metal2 76320 13368 76320 13368 0 _0763_
rlabel metal2 75504 15766 75504 15766 0 _0764_
rlabel metal2 75264 24486 75264 24486 0 _0765_
rlabel via1 76704 26294 76704 26294 0 _0766_
rlabel metal3 77232 27636 77232 27636 0 _0767_
rlabel metal2 76224 29778 76224 29778 0 _0768_
rlabel via2 76800 32411 76800 32411 0 _0769_
rlabel metal2 78048 34228 78048 34228 0 _0770_
rlabel metal2 76128 36372 76128 36372 0 _0771_
rlabel metal2 73536 36792 73536 36792 0 _0772_
rlabel metal2 72192 36162 72192 36162 0 _0773_
rlabel metal2 71040 34902 71040 34902 0 _0774_
rlabel via2 72384 32605 72384 32605 0 _0775_
rlabel metal2 71904 30912 71904 30912 0 _0776_
rlabel metal2 71088 28896 71088 28896 0 _0777_
rlabel metal3 71328 27804 71328 27804 0 _0778_
rlabel metal2 70944 26208 70944 26208 0 _0779_
rlabel metal2 68784 25536 68784 25536 0 _0780_
rlabel metal3 65856 25284 65856 25284 0 _0781_
rlabel metal3 64368 26796 64368 26796 0 _0782_
rlabel metal2 65664 28560 65664 28560 0 _0783_
rlabel via2 66432 29650 66432 29650 0 _0784_
rlabel metal2 67680 32537 67680 32537 0 _0785_
rlabel metal2 68160 34564 68160 34564 0 _0786_
rlabel metal2 67488 37338 67488 37338 0 _0787_
rlabel metal2 63936 36750 63936 36750 0 _0788_
rlabel metal2 60000 37338 60000 37338 0 _0789_
rlabel metal3 57072 37380 57072 37380 0 _0790_
rlabel via2 59424 35366 59424 35366 0 _0791_
rlabel metal2 63552 34104 63552 34104 0 _0792_
rlabel via2 63072 32674 63072 32674 0 _0793_
rlabel metal2 60768 32004 60768 32004 0 _0794_
rlabel metal2 57216 31878 57216 31878 0 _0795_
rlabel metal2 55200 34188 55200 34188 0 _0796_
rlabel metal3 51792 33432 51792 33432 0 _0797_
rlabel metal2 51456 31051 51456 31051 0 _0798_
rlabel via1 54432 29650 54432 29650 0 _0799_
rlabel via2 57504 29318 57504 29318 0 _0800_
rlabel metal3 60384 28308 60384 28308 0 _0801_
rlabel metal2 61920 27342 61920 27342 0 _0802_
rlabel via2 59616 25114 59616 25114 0 _0803_
rlabel metal3 56256 25956 56256 25956 0 _0804_
rlabel metal2 53568 26124 53568 26124 0 _0805_
rlabel metal2 52320 28516 52320 28516 0 _0806_
rlabel metal2 48096 29946 48096 29946 0 _0807_
rlabel metal2 47424 27804 47424 27804 0 _0808_
rlabel metal2 48288 25156 48288 25156 0 _0809_
rlabel metal2 50880 24358 50880 24358 0 _0810_
rlabel metal2 49824 21979 49824 21979 0 _0811_
rlabel metal2 45984 21672 45984 21672 0 _0812_
rlabel metal2 42528 22468 42528 22468 0 _0813_
rlabel metal2 43344 23268 43344 23268 0 _0814_
rlabel metal2 43920 26124 43920 26124 0 _0815_
rlabel metal2 42624 28056 42624 28056 0 _0816_
rlabel metal3 39984 26796 39984 26796 0 _0817_
rlabel metal3 38016 25116 38016 25116 0 _0818_
rlabel metal2 36624 22260 36624 22260 0 _0819_
rlabel metal2 35952 20748 35952 20748 0 _0820_
rlabel metal2 31680 20525 31680 20525 0 _0821_
rlabel metal2 3936 18356 3936 18356 0 _0822_
rlabel metal2 6816 17472 6816 17472 0 _0823_
rlabel metal2 42624 18942 42624 18942 0 _0824_
rlabel metal2 41760 20097 41760 20097 0 _0825_
rlabel metal3 4368 23016 4368 23016 0 _0826_
rlabel metal2 40608 20076 40608 20076 0 _0827_
rlabel metal2 46848 18984 46848 18984 0 _0828_
rlabel metal2 46128 19404 46128 19404 0 _0829_
rlabel metal2 45600 19362 45600 19362 0 _0830_
rlabel metal3 50448 18564 50448 18564 0 _0831_
rlabel metal2 49632 18858 49632 18858 0 _0832_
rlabel metal2 48384 19404 48384 19404 0 _0833_
rlabel metal2 50160 16212 50160 16212 0 _0834_
rlabel metal2 50688 16380 50688 16380 0 _0835_
rlabel metal2 49824 17934 49824 17934 0 _0836_
rlabel metal2 46080 16254 46080 16254 0 _0837_
rlabel metal2 46368 15918 46368 15918 0 _0838_
rlabel metal2 47040 15372 47040 15372 0 _0839_
rlabel metal2 44160 17556 44160 17556 0 _0840_
rlabel metal2 43776 17577 43776 17577 0 _0841_
rlabel metal2 43584 16905 43584 16905 0 _0842_
rlabel metal3 40512 19236 40512 19236 0 _0843_
rlabel metal2 39744 18942 39744 18942 0 _0844_
rlabel metal2 39552 19362 39552 19362 0 _0845_
rlabel metal2 37728 18228 37728 18228 0 _0846_
rlabel metal2 36384 19194 36384 19194 0 _0847_
rlabel metal2 36576 19362 36576 19362 0 _0848_
rlabel metal2 33408 17766 33408 17766 0 _0849_
rlabel metal3 34272 18522 34272 18522 0 _0850_
rlabel metal2 33696 18186 33696 18186 0 _0851_
rlabel metal2 32688 16212 32688 16212 0 _0852_
rlabel metal2 32256 17094 32256 17094 0 _0853_
rlabel metal2 32352 16926 32352 16926 0 _0854_
rlabel metal2 35808 15792 35808 15792 0 _0855_
rlabel metal2 35568 15372 35568 15372 0 _0856_
rlabel metal2 34848 15414 34848 15414 0 _0857_
rlabel metal2 38016 15582 38016 15582 0 _0858_
rlabel metal2 37728 15036 37728 15036 0 _0859_
rlabel metal2 37152 15036 37152 15036 0 _0860_
rlabel metal3 40416 14028 40416 14028 0 _0861_
rlabel metal2 39648 14196 39648 14196 0 _0862_
rlabel metal2 39456 14238 39456 14238 0 _0863_
rlabel metal2 42720 14271 42720 14271 0 _0864_
rlabel metal2 42480 13860 42480 13860 0 _0865_
rlabel metal2 41616 12348 41616 12348 0 _0866_
rlabel metal2 45120 14070 45120 14070 0 _0867_
rlabel metal2 44832 14154 44832 14154 0 _0868_
rlabel metal2 44544 12390 44544 12390 0 _0869_
rlabel metal2 46656 12096 46656 12096 0 _0870_
rlabel metal3 46896 13356 46896 13356 0 _0871_
rlabel metal2 45984 11592 45984 11592 0 _0872_
rlabel metal2 43296 11046 43296 11046 0 _0873_
rlabel metal2 43008 10710 43008 10710 0 _0874_
rlabel metal2 43392 10500 43392 10500 0 _0875_
rlabel metal3 46368 9492 46368 9492 0 _0876_
rlabel metal2 45888 9492 45888 9492 0 _0877_
rlabel metal2 45408 8820 45408 8820 0 _0878_
rlabel metal3 48864 8484 48864 8484 0 _0879_
rlabel metal2 48384 8778 48384 8778 0 _0880_
rlabel metal2 48000 7350 48000 7350 0 _0881_
rlabel metal2 51552 9366 51552 9366 0 _0882_
rlabel metal3 51456 8904 51456 8904 0 _0883_
rlabel metal3 50496 7392 50496 7392 0 _0884_
rlabel metal3 51312 11592 51312 11592 0 _0885_
rlabel metal2 51264 11403 51264 11403 0 _0886_
rlabel metal2 51072 10416 51072 10416 0 _0887_
rlabel metal2 49632 14364 49632 14364 0 _0888_
rlabel metal2 48384 14028 48384 14028 0 _0889_
rlabel metal2 49824 12726 49824 12726 0 _0890_
rlabel metal2 52992 14784 52992 14784 0 _0891_
rlabel metal2 52368 14952 52368 14952 0 _0892_
rlabel metal3 51648 13440 51648 13440 0 _0893_
rlabel metal2 55776 14784 55776 14784 0 _0894_
rlabel metal3 54864 14868 54864 14868 0 _0895_
rlabel metal2 54432 13440 54432 13440 0 _0896_
rlabel metal2 56064 12558 56064 12558 0 _0897_
rlabel metal3 18366 36708 18366 36708 0 clk
rlabel metal2 39264 14826 39264 14826 0 clknet_0_clk
rlabel metal2 41280 14280 41280 14280 0 clknet_2_0__leaf_clk
rlabel metal3 35136 23772 35136 23772 0 clknet_2_1__leaf_clk
rlabel metal2 61344 1890 61344 1890 0 clknet_2_2__leaf_clk
rlabel metal2 75936 38304 75936 38304 0 clknet_2_3__leaf_clk
rlabel metal3 12864 18564 12864 18564 0 clknet_leaf_0_clk
rlabel metal2 53760 15120 53760 15120 0 clknet_leaf_10_clk
rlabel metal2 78192 14028 78192 14028 0 clknet_leaf_11_clk
rlabel metal2 70176 1092 70176 1092 0 clknet_leaf_12_clk
rlabel metal2 78240 1512 78240 1512 0 clknet_leaf_13_clk
rlabel metal3 60768 1932 60768 1932 0 clknet_leaf_14_clk
rlabel metal3 57984 3444 57984 3444 0 clknet_leaf_15_clk
rlabel metal2 42528 12318 42528 12318 0 clknet_leaf_16_clk
rlabel metal2 9024 18522 9024 18522 0 clknet_leaf_17_clk
rlabel metal3 3600 20748 3600 20748 0 clknet_leaf_1_clk
rlabel metal2 38592 20832 38592 20832 0 clknet_leaf_2_clk
rlabel metal2 54912 28728 54912 28728 0 clknet_leaf_3_clk
rlabel metal3 51312 33684 51312 33684 0 clknet_leaf_4_clk
rlabel metal2 59904 35112 59904 35112 0 clknet_leaf_5_clk
rlabel metal3 73872 34356 73872 34356 0 clknet_leaf_6_clk
rlabel metal2 62976 28728 62976 28728 0 clknet_leaf_7_clk
rlabel metal3 56592 24612 56592 24612 0 clknet_leaf_8_clk
rlabel metal2 51264 22638 51264 22638 0 clknet_leaf_9_clk
rlabel metal3 43488 19236 43488 19236 0 daisychain\[0\]
rlabel metal2 61536 27720 61536 27720 0 daisychain\[100\]
rlabel metal3 59568 26124 59568 26124 0 daisychain\[101\]
rlabel metal2 57792 25368 57792 25368 0 daisychain\[102\]
rlabel metal2 55104 26376 55104 26376 0 daisychain\[103\]
rlabel metal2 53376 26292 53376 26292 0 daisychain\[104\]
rlabel metal2 51264 29064 51264 29064 0 daisychain\[105\]
rlabel metal3 46176 29148 46176 29148 0 daisychain\[106\]
rlabel metal3 47616 27636 47616 27636 0 daisychain\[107\]
rlabel metal2 50112 25578 50112 25578 0 daisychain\[108\]
rlabel metal3 50544 24528 50544 24528 0 daisychain\[109\]
rlabel metal2 36672 15246 36672 15246 0 daisychain\[10\]
rlabel metal3 48480 21336 48480 21336 0 daisychain\[110\]
rlabel metal3 44880 22092 44880 22092 0 daisychain\[111\]
rlabel metal3 41808 23268 41808 23268 0 daisychain\[112\]
rlabel metal2 43440 24780 43440 24780 0 daisychain\[113\]
rlabel metal2 44064 27342 44064 27342 0 daisychain\[114\]
rlabel metal3 40272 27636 40272 27636 0 daisychain\[115\]
rlabel metal2 38688 26040 38688 26040 0 daisychain\[116\]
rlabel via2 36480 24528 36480 24528 0 daisychain\[117\]
rlabel metal2 35760 22680 35760 22680 0 daisychain\[118\]
rlabel metal3 34272 20748 34272 20748 0 daisychain\[119\]
rlabel metal2 38688 14574 38688 14574 0 daisychain\[11\]
rlabel metal2 4310 19186 4310 19186 0 daisychain\[120\]
rlabel metal2 3744 17766 3744 17766 0 daisychain\[121\]
rlabel metal2 7008 16254 7008 16254 0 daisychain\[122\]
rlabel metal2 11040 16674 11040 16674 0 daisychain\[123\]
rlabel metal2 1728 17892 1728 17892 0 daisychain\[124\]
rlabel metal2 1344 18732 1344 18732 0 daisychain\[125\]
rlabel metal3 3024 20076 3024 20076 0 daisychain\[126\]
rlabel metal3 1488 19320 1488 19320 0 daisychain\[127\]
rlabel metal2 41280 12738 41280 12738 0 daisychain\[12\]
rlabel metal3 43536 12516 43536 12516 0 daisychain\[13\]
rlabel metal3 46176 13020 46176 13020 0 daisychain\[14\]
rlabel metal2 44448 11256 44448 11256 0 daisychain\[15\]
rlabel metal2 45024 9702 45024 9702 0 daisychain\[16\]
rlabel metal3 47280 7728 47280 7728 0 daisychain\[17\]
rlabel metal3 49968 8148 49968 8148 0 daisychain\[18\]
rlabel metal2 52272 9660 52272 9660 0 daisychain\[19\]
rlabel metal2 47808 20370 47808 20370 0 daisychain\[1\]
rlabel metal2 50592 12222 50592 12222 0 daisychain\[20\]
rlabel metal2 51072 13188 51072 13188 0 daisychain\[21\]
rlabel metal2 53952 14448 53952 14448 0 daisychain\[22\]
rlabel metal2 55776 13482 55776 13482 0 daisychain\[23\]
rlabel metal2 55488 11382 55488 11382 0 daisychain\[24\]
rlabel metal2 55488 8946 55488 8946 0 daisychain\[25\]
rlabel metal2 53856 7812 53856 7812 0 daisychain\[26\]
rlabel metal2 53952 5208 53952 5208 0 daisychain\[27\]
rlabel metal2 56256 4620 56256 4620 0 daisychain\[28\]
rlabel metal2 58224 2604 58224 2604 0 daisychain\[29\]
rlabel metal2 50928 17724 50928 17724 0 daisychain\[2\]
rlabel metal2 60480 2352 60480 2352 0 daisychain\[30\]
rlabel metal3 62256 2604 62256 2604 0 daisychain\[31\]
rlabel metal2 59808 5712 59808 5712 0 daisychain\[32\]
rlabel metal2 59424 8526 59424 8526 0 daisychain\[33\]
rlabel metal3 59136 10164 59136 10164 0 daisychain\[34\]
rlabel metal2 59520 13356 59520 13356 0 daisychain\[35\]
rlabel metal3 62112 13776 62112 13776 0 daisychain\[36\]
rlabel metal2 62688 11970 62688 11970 0 daisychain\[37\]
rlabel metal2 63264 10206 63264 10206 0 daisychain\[38\]
rlabel metal2 64320 7434 64320 7434 0 daisychain\[39\]
rlabel metal2 47616 16170 47616 16170 0 daisychain\[3\]
rlabel metal3 64320 6636 64320 6636 0 daisychain\[40\]
rlabel metal2 64752 2604 64752 2604 0 daisychain\[41\]
rlabel metal3 66816 1680 66816 1680 0 daisychain\[42\]
rlabel metal2 69264 2604 69264 2604 0 daisychain\[43\]
rlabel metal2 70368 5376 70368 5376 0 daisychain\[44\]
rlabel metal2 67776 9198 67776 9198 0 daisychain\[45\]
rlabel metal2 66240 11424 66240 11424 0 daisychain\[46\]
rlabel metal3 67295 13104 67295 13104 0 daisychain\[47\]
rlabel metal3 68928 13776 68928 13776 0 daisychain\[48\]
rlabel metal2 71040 13524 71040 13524 0 daisychain\[49\]
rlabel metal3 44976 17052 44976 17052 0 daisychain\[4\]
rlabel metal2 72096 12474 72096 12474 0 daisychain\[50\]
rlabel metal2 72288 11172 72288 11172 0 daisychain\[51\]
rlabel metal2 71808 8358 71808 8358 0 daisychain\[52\]
rlabel metal2 72672 7056 72672 7056 0 daisychain\[53\]
rlabel metal3 72144 4704 72144 4704 0 daisychain\[54\]
rlabel metal3 71856 3192 71856 3192 0 daisychain\[55\]
rlabel metal2 73824 2226 73824 2226 0 daisychain\[56\]
rlabel metal3 78192 2604 78192 2604 0 daisychain\[57\]
rlabel via2 78144 4200 78144 4200 0 daisychain\[58\]
rlabel metal3 79008 6636 79008 6636 0 daisychain\[59\]
rlabel metal2 40512 17766 40512 17766 0 daisychain\[5\]
rlabel metal2 78192 7980 78192 7980 0 daisychain\[60\]
rlabel metal2 76992 11172 76992 11172 0 daisychain\[61\]
rlabel metal2 76224 13734 76224 13734 0 daisychain\[62\]
rlabel metal5 74684 23100 74684 23100 0 daisychain\[63\]
rlabel metal2 75696 25116 75696 25116 0 daisychain\[64\]
rlabel metal2 76896 27342 76896 27342 0 daisychain\[65\]
rlabel metal2 76848 28560 76848 28560 0 daisychain\[66\]
rlabel metal2 77424 30828 77424 30828 0 daisychain\[67\]
rlabel metal3 78528 33684 78528 33684 0 daisychain\[68\]
rlabel metal3 78768 35868 78768 35868 0 daisychain\[69\]
rlabel metal2 38400 19110 38400 19110 0 daisychain\[6\]
rlabel metal2 76608 37338 76608 37338 0 daisychain\[70\]
rlabel metal2 73056 36960 73056 36960 0 daisychain\[71\]
rlabel metal3 70464 35868 70464 35868 0 daisychain\[72\]
rlabel metal2 70944 34650 70944 34650 0 daisychain\[73\]
rlabel metal2 72384 32256 72384 32256 0 daisychain\[74\]
rlabel metal2 71424 30114 71424 30114 0 daisychain\[75\]
rlabel metal2 70464 28602 70464 28602 0 daisychain\[76\]
rlabel metal2 71232 27594 71232 27594 0 daisychain\[77\]
rlabel metal2 69792 26376 69792 26376 0 daisychain\[78\]
rlabel metal2 68592 25284 68592 25284 0 daisychain\[79\]
rlabel metal3 36048 19824 36048 19824 0 daisychain\[7\]
rlabel metal2 64896 25620 64896 25620 0 daisychain\[80\]
rlabel metal2 64752 26796 64752 26796 0 daisychain\[81\]
rlabel metal2 65424 28560 65424 28560 0 daisychain\[82\]
rlabel metal2 66432 30912 66432 30912 0 daisychain\[83\]
rlabel metal2 67584 33402 67584 33402 0 daisychain\[84\]
rlabel metal3 68544 35700 68544 35700 0 daisychain\[85\]
rlabel metal2 65568 38052 65568 38052 0 daisychain\[86\]
rlabel metal2 61728 36372 61728 36372 0 daisychain\[87\]
rlabel metal3 58608 37212 58608 37212 0 daisychain\[88\]
rlabel metal2 58608 36540 58608 36540 0 daisychain\[89\]
rlabel metal2 33408 18270 33408 18270 0 daisychain\[8\]
rlabel metal2 60288 35238 60288 35238 0 daisychain\[90\]
rlabel metal2 63370 34491 63370 34491 0 daisychain\[91\]
rlabel metal2 61824 32424 61824 32424 0 daisychain\[92\]
rlabel metal2 58944 31626 58944 31626 0 daisychain\[93\]
rlabel metal2 56160 32298 56160 32298 0 daisychain\[94\]
rlabel metal3 54672 34356 54672 34356 0 daisychain\[95\]
rlabel metal3 49920 33432 49920 33432 0 daisychain\[96\]
rlabel metal2 52128 31626 52128 31626 0 daisychain\[97\]
rlabel metal3 55728 30828 55728 30828 0 daisychain\[98\]
rlabel metal2 58848 29400 58848 29400 0 daisychain\[99\]
rlabel metal2 34080 15960 34080 15960 0 daisychain\[9\]
rlabel metal2 53616 16968 53616 16968 0 digitalen.g\[0\].u.OUTN
rlabel metal2 53472 17010 53472 17010 0 digitalen.g\[0\].u.OUTP
rlabel metal2 79392 16254 79392 16254 0 digitalen.g\[1\].u.OUTN
rlabel metal2 79488 16758 79488 16758 0 digitalen.g\[1\].u.OUTP
rlabel metal2 79565 22828 79565 22828 0 digitalen.g\[2\].u.OUTN
rlabel metal3 79197 23016 79197 23016 0 digitalen.g\[2\].u.OUTP
rlabel metal2 52704 22638 52704 22638 0 digitalen.g\[3\].u.OUTN
rlabel metal2 53675 22828 53675 22828 0 digitalen.g\[3\].u.OUTP
rlabel metal3 99924 21672 99924 21672 0 i_in
rlabel metal3 99924 19992 99924 19992 0 i_out
rlabel metal3 366 15708 366 15708 0 net
rlabel metal2 864 37704 864 37704 0 net1
rlabel metal3 1200 11760 1200 11760 0 net10
rlabel metal2 56256 6300 56256 6300 0 net100
rlabel metal2 50112 18564 50112 18564 0 net101
rlabel metal2 56064 15162 56064 15162 0 net102
rlabel metal3 57792 14700 57792 14700 0 net103
rlabel metal2 42912 18642 42912 18642 0 net104
rlabel metal3 42768 27636 42768 27636 0 net105
rlabel metal2 46896 22260 46896 22260 0 net106
rlabel metal3 54048 25284 54048 25284 0 net107
rlabel metal2 56160 34314 56160 34314 0 net108
rlabel metal2 55392 33474 55392 33474 0 net109
rlabel metal2 864 12726 864 12726 0 net11
rlabel metal2 49920 27300 49920 27300 0 net110
rlabel metal2 39888 20832 39888 20832 0 net111
rlabel metal2 62832 2352 62832 2352 0 net112
rlabel metal2 62688 10962 62688 10962 0 net113
rlabel metal2 65664 2742 65664 2742 0 net114
rlabel metal2 62112 14322 62112 14322 0 net115
rlabel metal2 61920 15036 61920 15036 0 net116
rlabel metal2 72768 2646 72768 2646 0 net117
rlabel metal2 77856 6300 77856 6300 0 net118
rlabel metal2 72096 7182 72096 7182 0 net119
rlabel metal3 1200 13272 1200 13272 0 net12
rlabel metal2 77664 11340 77664 11340 0 net120
rlabel metal2 77856 13272 77856 13272 0 net121
rlabel metal2 77376 8106 77376 8106 0 net122
rlabel metal2 62016 25620 62016 25620 0 net123
rlabel metal2 61536 35826 61536 35826 0 net124
rlabel metal2 68064 33936 68064 33936 0 net125
rlabel metal3 60048 33936 60048 33936 0 net126
rlabel metal2 62112 29400 62112 29400 0 net127
rlabel metal2 69696 25158 69696 25158 0 net128
rlabel via2 77952 27048 77952 27048 0 net129
rlabel metal2 1104 18144 1104 18144 0 net13
rlabel metal2 71328 34440 71328 34440 0 net130
rlabel metal2 76800 29862 76800 29862 0 net131
rlabel metal2 76320 35784 76320 35784 0 net132
rlabel metal2 73536 34524 73536 34524 0 net133
rlabel metal2 60480 26292 60480 26292 0 net134
rlabel metal4 61920 15078 61920 15078 0 net135
rlabel metal2 2784 21084 2784 21084 0 net136
rlabel metal2 4512 21546 4512 21546 0 net137
rlabel metal2 1920 23604 1920 23604 0 net138
rlabel metal2 36192 16758 36192 16758 0 net139
rlabel metal2 864 15414 864 15414 0 net14
rlabel metal2 36960 20664 36960 20664 0 net140
rlabel metal2 2016 24108 2016 24108 0 net141
rlabel metal2 42816 11046 42816 11046 0 net142
rlabel metal2 46944 19068 46944 19068 0 net143
rlabel metal2 39552 18858 39552 18858 0 net144
rlabel metal2 40128 17514 40128 17514 0 net145
rlabel metal2 56064 5208 56064 5208 0 net146
rlabel metal2 53088 14574 53088 14574 0 net147
rlabel metal2 55440 16212 55440 16212 0 net148
rlabel metal2 55680 8190 55680 8190 0 net149
rlabel metal2 720 2688 720 2688 0 net15
rlabel metal3 42624 21588 42624 21588 0 net150
rlabel metal2 40608 25242 40608 25242 0 net151
rlabel metal2 42720 28896 42720 28896 0 net152
rlabel via1 51844 23780 51844 23780 0 net153
rlabel metal2 55968 34440 55968 34440 0 net154
rlabel metal3 56544 30072 56544 30072 0 net155
rlabel metal3 54672 25284 54672 25284 0 net156
rlabel metal3 40272 17808 40272 17808 0 net157
rlabel metal2 62688 1848 62688 1848 0 net158
rlabel metal2 63840 9408 63840 9408 0 net159
rlabel metal3 1680 3360 1680 3360 0 net16
rlabel metal2 60144 10248 60144 10248 0 net160
rlabel metal2 58896 14952 58896 14952 0 net161
rlabel metal3 67632 15540 67632 15540 0 net162
rlabel metal3 68976 2604 68976 2604 0 net163
rlabel metal2 74112 2184 74112 2184 0 net164
rlabel metal2 76800 7560 76800 7560 0 net165
rlabel metal2 73536 8904 73536 8904 0 net166
rlabel metal2 77664 13074 77664 13074 0 net167
rlabel metal2 76512 13986 76512 13986 0 net168
rlabel metal2 65088 15624 65088 15624 0 net169
rlabel metal3 1152 4200 1152 4200 0 net17
rlabel metal2 61248 24108 61248 24108 0 net170
rlabel metal2 59424 33600 59424 33600 0 net171
rlabel metal2 65376 35070 65376 35070 0 net172
rlabel metal2 59040 34020 59040 34020 0 net173
rlabel metal3 60576 25536 60576 25536 0 net174
rlabel metal2 76800 23898 76800 23898 0 net175
rlabel metal2 76416 24066 76416 24066 0 net176
rlabel metal2 71904 33474 71904 33474 0 net177
rlabel metal2 77424 29148 77424 29148 0 net178
rlabel metal2 74880 35658 74880 35658 0 net179
rlabel metal2 912 4872 912 4872 0 net18
rlabel metal2 68640 32214 68640 32214 0 net180
rlabel metal2 58944 25410 58944 25410 0 net181
rlabel metal2 2400 24990 2400 24990 0 net182
rlabel metal2 6048 17892 6048 17892 0 net183
rlabel metal2 2784 19782 2784 19782 0 net184
rlabel metal2 34848 14364 34848 14364 0 net185
rlabel metal2 39600 21588 39600 21588 0 net186
rlabel metal2 36000 16842 36000 16842 0 net187
rlabel metal2 46272 14490 46272 14490 0 net188
rlabel metal2 39216 13272 39216 13272 0 net189
rlabel metal3 1248 5712 1248 5712 0 net19
rlabel metal2 43008 9744 43008 9744 0 net190
rlabel metal2 50304 9534 50304 9534 0 net191
rlabel metal2 57552 7140 57552 7140 0 net192
rlabel metal2 54528 13944 54528 13944 0 net193
rlabel metal2 55776 15792 55776 15792 0 net194
rlabel metal2 56112 16296 56112 16296 0 net195
rlabel metal2 43008 21042 43008 21042 0 net196
rlabel metal2 45792 21168 45792 21168 0 net197
rlabel metal2 40416 26166 40416 26166 0 net198
rlabel metal2 53568 27468 53568 27468 0 net199
rlabel metal2 912 22932 912 22932 0 net2
rlabel metal2 960 18312 960 18312 0 net20
rlabel metal3 56544 26796 56544 26796 0 net200
rlabel metal2 56640 36498 56640 36498 0 net201
rlabel metal2 52992 34104 52992 34104 0 net202
rlabel metal2 40704 29190 40704 29190 0 net203
rlabel metal2 60288 1302 60288 1302 0 net204
rlabel metal2 64416 9576 64416 9576 0 net205
rlabel metal2 61152 9912 61152 9912 0 net206
rlabel metal2 61632 15162 61632 15162 0 net207
rlabel metal2 64992 14994 64992 14994 0 net208
rlabel metal2 76416 2016 76416 2016 0 net209
rlabel metal2 1488 18312 1488 18312 0 net21
rlabel metal2 76032 7182 76032 7182 0 net210
rlabel metal3 71808 1974 71808 1974 0 net211
rlabel metal2 69024 13230 69024 13230 0 net212
rlabel metal4 77376 13104 77376 13104 0 net213
rlabel metal2 73459 14739 73459 14739 0 net214
rlabel metal2 59040 27132 59040 27132 0 net215
rlabel metal2 62112 35196 62112 35196 0 net216
rlabel metal2 66816 35952 66816 35952 0 net217
rlabel metal2 59328 34398 59328 34398 0 net218
rlabel metal2 74976 26754 74976 26754 0 net219
rlabel metal3 1584 17304 1584 17304 0 net22
rlabel metal2 71136 35280 71136 35280 0 net220
rlabel metal2 77472 35028 77472 35028 0 net221
rlabel metal2 77136 36708 77136 36708 0 net222
rlabel metal2 74592 36750 74592 36750 0 net223
rlabel metal2 77472 27846 77472 27846 0 net224
rlabel metal2 60096 37170 60096 37170 0 net225
rlabel metal5 40032 19992 40032 19992 0 net226
rlabel metal2 5952 20370 5952 20370 0 net227
rlabel metal3 558 16548 558 16548 0 net228
rlabel metal3 366 17388 366 17388 0 net229
rlabel metal2 5232 18312 5232 18312 0 net23
rlabel metal3 366 18228 366 18228 0 net230
rlabel metal3 366 19068 366 19068 0 net231
rlabel metal3 366 19908 366 19908 0 net232
rlabel metal3 366 20748 366 20748 0 net233
rlabel metal3 366 21588 366 21588 0 net234
rlabel metal2 6816 19908 6816 19908 0 net24
rlabel metal3 38784 19236 38784 19236 0 net25
rlabel metal2 36672 19362 36672 19362 0 net26
rlabel metal2 40560 27636 40560 27636 0 net27
rlabel metal2 35952 22260 35952 22260 0 net28
rlabel metal2 4704 19950 4704 19950 0 net29
rlabel metal3 1200 23100 1200 23100 0 net3
rlabel metal3 42240 18396 42240 18396 0 net30
rlabel metal2 47136 16170 47136 16170 0 net31
rlabel metal2 41280 19404 41280 19404 0 net32
rlabel metal3 58176 2604 58176 2604 0 net33
rlabel metal2 54144 4872 54144 4872 0 net34
rlabel metal3 54240 14742 54240 14742 0 net35
rlabel metal3 58368 11172 58368 11172 0 net36
rlabel metal3 41184 22260 41184 22260 0 net37
rlabel metal2 42720 25158 42720 25158 0 net38
rlabel metal2 42528 25452 42528 25452 0 net39
rlabel metal3 1536 24528 1536 24528 0 net4
rlabel metal2 54048 25998 54048 25998 0 net40
rlabel metal3 58080 35868 58080 35868 0 net41
rlabel metal2 51456 29064 51456 29064 0 net42
rlabel metal3 56928 33600 56928 33600 0 net43
rlabel metal3 41760 25368 41760 25368 0 net44
rlabel metal3 60192 2604 60192 2604 0 net45
rlabel metal3 67248 2604 67248 2604 0 net46
rlabel metal2 59040 8358 59040 8358 0 net47
rlabel metal3 59952 13440 59952 13440 0 net48
rlabel metal2 60000 13398 60000 13398 0 net49
rlabel metal3 2208 21504 2208 21504 0 net5
rlabel metal2 68688 2604 68688 2604 0 net50
rlabel metal2 72000 9786 72000 9786 0 net51
rlabel metal3 75120 1932 75120 1932 0 net52
rlabel metal2 77664 7854 77664 7854 0 net53
rlabel metal2 76512 11592 76512 11592 0 net54
rlabel metal2 69504 13734 69504 13734 0 net55
rlabel metal2 65760 25242 65760 25242 0 net56
rlabel metal2 61440 35154 61440 35154 0 net57
rlabel metal2 67104 36750 67104 36750 0 net58
rlabel metal2 62928 34356 62928 34356 0 net59
rlabel metal2 864 26418 864 26418 0 net6
rlabel metal2 59808 29652 59808 29652 0 net60
rlabel metal2 69984 26250 69984 26250 0 net61
rlabel metal2 75648 25788 75648 25788 0 net62
rlabel metal2 71616 35910 71616 35910 0 net63
rlabel metal2 77520 35868 77520 35868 0 net64
rlabel metal2 73920 36540 73920 36540 0 net65
rlabel metal2 58656 26544 58656 26544 0 net66
rlabel metal3 42384 26040 42384 26040 0 net67
rlabel metal2 40128 21504 40128 21504 0 net68
rlabel metal2 33504 22050 33504 22050 0 net69
rlabel metal3 15168 9408 15168 9408 0 net7
rlabel metal2 4416 19320 4416 19320 0 net70
rlabel metal2 44928 8736 44928 8736 0 net71
rlabel metal2 58560 2688 58560 2688 0 net72
rlabel metal3 53664 13062 53664 13062 0 net73
rlabel metal2 49920 11676 49920 11676 0 net74
rlabel metal2 43104 22596 43104 22596 0 net75
rlabel metal2 51168 29232 51168 29232 0 net76
rlabel metal2 56160 29694 56160 29694 0 net77
rlabel metal3 44208 20832 44208 20832 0 net78
rlabel metal2 64608 2520 64608 2520 0 net79
rlabel metal2 864 10290 864 10290 0 net8
rlabel metal3 60672 13188 60672 13188 0 net80
rlabel metal2 74592 2478 74592 2478 0 net81
rlabel metal2 77568 2742 77568 2742 0 net82
rlabel metal2 75936 13650 75936 13650 0 net83
rlabel metal2 61248 35364 61248 35364 0 net84
rlabel metal2 61440 27804 61440 27804 0 net85
rlabel metal2 77280 31458 77280 31458 0 net86
rlabel metal2 74448 35868 74448 35868 0 net87
rlabel metal2 76320 35112 76320 35112 0 net88
rlabel metal2 6816 18354 6816 18354 0 net89
rlabel metal2 864 11214 864 11214 0 net9
rlabel metal2 6816 17766 6816 17766 0 net90
rlabel metal2 6720 19446 6720 19446 0 net91
rlabel metal2 37440 18228 37440 18228 0 net92
rlabel metal2 33408 19572 33408 19572 0 net93
rlabel metal2 31056 20076 31056 20076 0 net94
rlabel metal2 33648 19992 33648 19992 0 net95
rlabel metal2 42816 13986 42816 13986 0 net96
rlabel metal2 46560 19908 46560 19908 0 net97
rlabel metal2 39888 20580 39888 20580 0 net98
rlabel metal3 55920 10164 55920 10164 0 net99
rlabel metal3 366 37548 366 37548 0 rst_n
rlabel metal3 42912 18501 42912 18501 0 state\[0\]
rlabel metal2 62880 28350 62880 28350 0 state\[100\]
rlabel metal2 62688 23814 62688 23814 0 state\[101\]
rlabel metal2 61920 23982 61920 23982 0 state\[102\]
rlabel metal2 59040 24276 59040 24276 0 state\[103\]
rlabel metal2 63275 22828 63275 22828 0 state\[104\]
rlabel metal2 62875 22690 62875 22690 0 state\[105\]
rlabel metal2 62475 22690 62475 22690 0 state\[106\]
rlabel metal2 62075 22828 62075 22828 0 state\[107\]
rlabel metal2 61675 22828 61675 22828 0 state\[108\]
rlabel metal2 61275 22828 61275 22828 0 state\[109\]
rlabel metal4 38016 16926 38016 16926 0 state\[10\]
rlabel metal4 57120 22932 57120 22932 0 state\[110\]
rlabel metal3 48048 22260 48048 22260 0 state\[111\]
rlabel metal3 42816 23226 42816 23226 0 state\[112\]
rlabel metal2 59675 22828 59675 22828 0 state\[113\]
rlabel metal2 59275 22828 59275 22828 0 state\[114\]
rlabel metal2 58875 22828 58875 22828 0 state\[115\]
rlabel metal2 40944 25284 40944 25284 0 state\[116\]
rlabel metal2 39216 22260 39216 22260 0 state\[117\]
rlabel metal2 57675 22690 57675 22690 0 state\[118\]
rlabel metal2 37680 22260 37680 22260 0 state\[119\]
rlabel metal2 40512 16506 40512 16506 0 state\[11\]
rlabel metal2 33360 21336 33360 21336 0 state\[120\]
rlabel metal2 3648 18438 3648 18438 0 state\[121\]
rlabel metal2 6144 14406 6144 14406 0 state\[122\]
rlabel metal2 18144 18228 18144 18228 0 state\[123\]
rlabel metal3 12288 19236 12288 19236 0 state\[124\]
rlabel metal2 13632 21294 13632 21294 0 state\[125\]
rlabel metal2 1824 19656 1824 19656 0 state\[126\]
rlabel metal2 3264 20790 3264 20790 0 state\[127\]
rlabel metal2 42432 16380 42432 16380 0 state\[12\]
rlabel metal3 54432 15330 54432 15330 0 state\[13\]
rlabel metal4 59424 16464 59424 16464 0 state\[14\]
rlabel metal2 59808 15624 59808 15624 0 state\[15\]
rlabel metal3 57552 14280 57552 14280 0 state\[16\]
rlabel metal3 48384 10416 48384 10416 0 state\[17\]
rlabel metal4 60960 15960 60960 15960 0 state\[18\]
rlabel metal3 61248 14112 61248 14112 0 state\[19\]
rlabel metal2 54336 15666 54336 15666 0 state\[1\]
rlabel metal2 53424 16212 53424 16212 0 state\[20\]
rlabel metal3 61152 16086 61152 16086 0 state\[21\]
rlabel metal2 54912 16674 54912 16674 0 state\[22\]
rlabel metal2 57792 15834 57792 15834 0 state\[23\]
rlabel metal2 63648 14658 63648 14658 0 state\[24\]
rlabel metal2 63936 16884 63936 16884 0 state\[25\]
rlabel metal3 57216 13692 57216 13692 0 state\[26\]
rlabel metal2 54624 7434 54624 7434 0 state\[27\]
rlabel metal2 57984 6762 57984 6762 0 state\[28\]
rlabel metal2 59856 4788 59856 4788 0 state\[29\]
rlabel metal2 54765 17378 54765 17378 0 state\[2\]
rlabel metal3 62400 13020 62400 13020 0 state\[30\]
rlabel metal3 65520 2100 65520 2100 0 state\[31\]
rlabel metal2 62112 6930 62112 6930 0 state\[32\]
rlabel metal2 60576 16170 60576 16170 0 state\[33\]
rlabel metal2 60096 16590 60096 16590 0 state\[34\]
rlabel metal2 60384 16002 60384 16002 0 state\[35\]
rlabel metal2 62016 15802 62016 15802 0 state\[36\]
rlabel metal2 65280 15036 65280 15036 0 state\[37\]
rlabel metal2 65184 13440 65184 13440 0 state\[38\]
rlabel metal2 69486 17052 69486 17052 0 state\[39\]
rlabel metal2 55104 16926 55104 16926 0 state\[3\]
rlabel metal2 68496 7392 68496 7392 0 state\[40\]
rlabel metal2 65760 5796 65760 5796 0 state\[41\]
rlabel metal2 66624 16464 66624 16464 0 state\[42\]
rlabel metal2 71232 2394 71232 2394 0 state\[43\]
rlabel metal2 69600 16170 69600 16170 0 state\[44\]
rlabel metal3 70704 13860 70704 13860 0 state\[45\]
rlabel metal3 68448 15582 68448 15582 0 state\[46\]
rlabel metal3 66528 14196 66528 14196 0 state\[47\]
rlabel metal2 73165 17366 73165 17366 0 state\[48\]
rlabel metal2 73536 16716 73536 16716 0 state\[49\]
rlabel metal2 55584 16506 55584 16506 0 state\[4\]
rlabel metal2 73920 16716 73920 16716 0 state\[50\]
rlabel metal2 74112 15708 74112 15708 0 state\[51\]
rlabel metal3 74448 16212 74448 16212 0 state\[52\]
rlabel metal2 75022 17052 75022 17052 0 state\[53\]
rlabel metal2 75024 15288 75024 15288 0 state\[54\]
rlabel metal2 75504 14532 75504 14532 0 state\[55\]
rlabel metal2 74976 2688 74976 2688 0 state\[56\]
rlabel metal2 76608 1596 76608 1596 0 state\[57\]
rlabel via3 77174 17304 77174 17304 0 state\[58\]
rlabel metal3 78240 14280 78240 14280 0 state\[59\]
rlabel metal2 55968 16590 55968 16590 0 state\[5\]
rlabel metal3 78384 15120 78384 15120 0 state\[60\]
rlabel metal3 78240 13398 78240 13398 0 state\[61\]
rlabel metal3 79056 14196 79056 14196 0 state\[62\]
rlabel metal3 79008 15708 79008 15708 0 state\[63\]
rlabel metal2 79275 22828 79275 22828 0 state\[64\]
rlabel metal3 78576 22932 78576 22932 0 state\[65\]
rlabel metal2 78475 22828 78475 22828 0 state\[66\]
rlabel metal2 78075 22690 78075 22690 0 state\[67\]
rlabel metal2 77675 22828 77675 22828 0 state\[68\]
rlabel metal2 76320 33768 76320 33768 0 state\[69\]
rlabel metal3 41664 18480 41664 18480 0 state\[6\]
rlabel metal2 76875 22690 76875 22690 0 state\[70\]
rlabel metal2 76445 22848 76445 22848 0 state\[71\]
rlabel metal3 75957 22764 75957 22764 0 state\[72\]
rlabel metal2 74688 34188 74688 34188 0 state\[73\]
rlabel metal2 75120 31920 75120 31920 0 state\[74\]
rlabel metal2 74875 22732 74875 22732 0 state\[75\]
rlabel metal2 74475 22828 74475 22828 0 state\[76\]
rlabel metal2 73776 22932 73776 22932 0 state\[77\]
rlabel metal2 73675 22690 73675 22690 0 state\[78\]
rlabel metal2 73275 22828 73275 22828 0 state\[79\]
rlabel metal3 39360 18270 39360 18270 0 state\[7\]
rlabel metal2 72875 22828 72875 22828 0 state\[80\]
rlabel metal2 72475 22828 72475 22828 0 state\[81\]
rlabel metal2 72075 22828 72075 22828 0 state\[82\]
rlabel metal2 67392 29316 67392 29316 0 state\[83\]
rlabel metal2 71275 22828 71275 22828 0 state\[84\]
rlabel metal3 70717 22764 70717 22764 0 state\[85\]
rlabel metal3 69168 36708 69168 36708 0 state\[86\]
rlabel metal2 66672 36456 66672 36456 0 state\[87\]
rlabel metal2 69675 22828 69675 22828 0 state\[88\]
rlabel metal2 57216 34188 57216 34188 0 state\[89\]
rlabel metal2 36000 18480 36000 18480 0 state\[8\]
rlabel metal3 61728 34188 61728 34188 0 state\[90\]
rlabel metal2 67296 24360 67296 24360 0 state\[91\]
rlabel metal2 68075 22828 68075 22828 0 state\[92\]
rlabel metal4 62688 30954 62688 30954 0 state\[93\]
rlabel metal2 60288 30366 60288 30366 0 state\[94\]
rlabel metal2 58080 34104 58080 34104 0 state\[95\]
rlabel metal3 54624 33180 54624 33180 0 state\[96\]
rlabel metal2 58272 23562 58272 23562 0 state\[97\]
rlabel metal2 56064 28812 56064 28812 0 state\[98\]
rlabel metal2 59040 27930 59040 27930 0 state\[99\]
rlabel metal4 35328 16884 35328 16884 0 state\[9\]
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 25788 366 25788 0 ui_in[4]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal2 672 6720 672 6720 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
