* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

.subckt heichips25_template VGND VPWR analog_pin0 analog_pin1 analog_pin2 analog_pin3
+ clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_28_907 VPWR VGND sg13g2_decap_8
XFILLER_39_266 VPWR VGND sg13g2_decap_8
XFILLER_27_406 VPWR VGND sg13g2_decap_8
XFILLER_36_973 VPWR VGND sg13g2_decap_8
XFILLER_35_483 VPWR VGND sg13g2_decap_8
XFILLER_23_634 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_19_907 VPWR VGND sg13g2_decap_8
XFILLER_18_417 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_42_910 VPWR VGND sg13g2_decap_8
XFILLER_26_74 VPWR VGND sg13g2_decap_8
XFILLER_14_634 VPWR VGND sg13g2_decap_8
XFILLER_41_420 VPWR VGND sg13g2_decap_8
XFILLER_26_494 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_42_987 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_8
XFILLER_41_497 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_6_844 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_17_483 VPWR VGND sg13g2_decap_8
XFILLER_45_770 VPWR VGND sg13g2_decap_8
XFILLER_33_910 VPWR VGND sg13g2_decap_8
XFILLER_18_984 VPWR VGND sg13g2_decap_8
XFILLER_44_280 VPWR VGND sg13g2_decap_8
XFILLER_32_420 VPWR VGND sg13g2_decap_8
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_32_497 VPWR VGND sg13g2_decap_8
XFILLER_20_648 VPWR VGND sg13g2_decap_8
XFILLER_28_704 VPWR VGND sg13g2_decap_8
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_43_707 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_36_770 VPWR VGND sg13g2_decap_8
XFILLER_24_921 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_3_858 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
XFILLER_19_704 VPWR VGND sg13g2_decap_8
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_34_707 VPWR VGND sg13g2_decap_8
XFILLER_15_921 VPWR VGND sg13g2_decap_8
XFILLER_33_217 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_14_431 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
XFILLER_15_998 VPWR VGND sg13g2_decap_8
XFILLER_30_924 VPWR VGND sg13g2_decap_8
XFILLER_18_1026 VPWR VGND sg13g2_fill_2
XFILLER_42_784 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
XFILLER_6_641 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_37_567 VPWR VGND sg13g2_decap_8
XFILLER_25_718 VPWR VGND sg13g2_decap_8
XFILLER_18_781 VPWR VGND sg13g2_decap_8
XFILLER_17_280 VPWR VGND sg13g2_decap_8
XFILLER_24_228 VPWR VGND sg13g2_decap_8
XFILLER_33_784 VPWR VGND sg13g2_decap_8
XFILLER_21_935 VPWR VGND sg13g2_decap_8
XFILLER_32_294 VPWR VGND sg13g2_decap_8
XFILLER_20_445 VPWR VGND sg13g2_decap_8
XFILLER_28_501 VPWR VGND sg13g2_decap_8
XFILLER_16_718 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_28_578 VPWR VGND sg13g2_decap_8
XFILLER_15_228 VPWR VGND sg13g2_decap_8
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_11_445 VPWR VGND sg13g2_decap_8
XFILLER_8_928 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_decap_8
XFILLER_7_427 VPWR VGND sg13g2_decap_8
XFILLER_48_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_19_501 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_34_504 VPWR VGND sg13g2_decap_8
XFILLER_19_578 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_15_795 VPWR VGND sg13g2_decap_8
XFILLER_42_581 VPWR VGND sg13g2_decap_8
XFILLER_30_721 VPWR VGND sg13g2_decap_8
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_31_1001 VPWR VGND sg13g2_decap_8
XFILLER_30_798 VPWR VGND sg13g2_decap_8
XFILLER_7_994 VPWR VGND sg13g2_decap_8
XFILLER_29_0 VPWR VGND sg13g2_decap_8
XFILLER_38_854 VPWR VGND sg13g2_decap_8
XFILLER_37_364 VPWR VGND sg13g2_decap_8
XFILLER_25_515 VPWR VGND sg13g2_decap_8
XFILLER_40_518 VPWR VGND sg13g2_decap_8
XFILLER_33_581 VPWR VGND sg13g2_decap_8
XFILLER_21_732 VPWR VGND sg13g2_decap_8
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_29_854 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_16_515 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_28_375 VPWR VGND sg13g2_decap_8
XFILLER_44_868 VPWR VGND sg13g2_decap_8
XFILLER_31_518 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_decap_8
XFILLER_24_592 VPWR VGND sg13g2_decap_8
XFILLER_11_242 VPWR VGND sg13g2_decap_8
XFILLER_8_725 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_decap_8
XFILLER_4_942 VPWR VGND sg13g2_decap_8
XFILLER_3_452 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_375 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_34_301 VPWR VGND sg13g2_decap_8
XFILLER_35_868 VPWR VGND sg13g2_decap_8
XFILLER_34_378 VPWR VGND sg13g2_decap_8
XFILLER_22_529 VPWR VGND sg13g2_decap_8
XFILLER_15_592 VPWR VGND sg13g2_decap_8
XFILLER_30_595 VPWR VGND sg13g2_decap_8
XFILLER_7_791 VPWR VGND sg13g2_decap_8
XFILLER_38_651 VPWR VGND sg13g2_decap_8
XFILLER_26_802 VPWR VGND sg13g2_decap_8
XFILLER_37_161 VPWR VGND sg13g2_decap_8
XFILLER_25_312 VPWR VGND sg13g2_decap_8
XFILLER_41_805 VPWR VGND sg13g2_decap_8
XFILLER_26_879 VPWR VGND sg13g2_decap_8
XFILLER_13_529 VPWR VGND sg13g2_decap_8
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_25_389 VPWR VGND sg13g2_decap_8
XFILLER_5_739 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_49_938 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_29_63 VPWR VGND sg13g2_decap_8
XFILLER_29_651 VPWR VGND sg13g2_decap_8
XFILLER_16_312 VPWR VGND sg13g2_decap_8
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_44_665 VPWR VGND sg13g2_decap_8
XFILLER_32_805 VPWR VGND sg13g2_decap_8
XFILLER_17_868 VPWR VGND sg13g2_decap_8
XFILLER_16_389 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_31_315 VPWR VGND sg13g2_decap_8
XFILLER_8_522 VPWR VGND sg13g2_decap_8
XFILLER_40_882 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_8_599 VPWR VGND sg13g2_decap_8
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_448 VPWR VGND sg13g2_decap_8
XFILLER_26_109 VPWR VGND sg13g2_decap_8
XFILLER_19_172 VPWR VGND sg13g2_decap_8
XFILLER_35_665 VPWR VGND sg13g2_decap_8
XFILLER_34_175 VPWR VGND sg13g2_decap_8
XFILLER_23_816 VPWR VGND sg13g2_decap_8
XFILLER_22_326 VPWR VGND sg13g2_decap_8
XFILLER_31_882 VPWR VGND sg13g2_decap_8
XFILLER_30_392 VPWR VGND sg13g2_decap_8
XFILLER_44_1022 VPWR VGND sg13g2_decap_8
Xheichips25_template_10 VPWR VGND uo_out[4] sg13g2_tielo
Xheichips25_template_21 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_14_816 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_41_602 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_25_186 VPWR VGND sg13g2_decap_8
XFILLER_9_319 VPWR VGND sg13g2_decap_8
XFILLER_41_679 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_decap_8
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_45_952 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_8
XFILLER_32_602 VPWR VGND sg13g2_decap_8
XFILLER_16_186 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_8
XFILLER_32_679 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_31_189 VPWR VGND sg13g2_decap_8
XFILLER_9_886 VPWR VGND sg13g2_decap_8
XFILLER_8_396 VPWR VGND sg13g2_decap_8
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_245 VPWR VGND sg13g2_decap_8
XFILLER_36_952 VPWR VGND sg13g2_decap_8
XFILLER_35_462 VPWR VGND sg13g2_decap_8
XFILLER_23_613 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_27_952 VPWR VGND sg13g2_decap_8
XFILLER_14_613 VPWR VGND sg13g2_decap_8
XFILLER_26_53 VPWR VGND sg13g2_decap_8
XFILLER_26_473 VPWR VGND sg13g2_decap_8
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_41_476 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_22_690 VPWR VGND sg13g2_decap_8
XFILLER_6_823 VPWR VGND sg13g2_decap_8
XFILLER_5_333 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_37_749 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_18_963 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_decap_8
XFILLER_33_966 VPWR VGND sg13g2_decap_8
XFILLER_32_476 VPWR VGND sg13g2_decap_8
XFILLER_20_627 VPWR VGND sg13g2_decap_8
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_9_683 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
XFILLER_27_259 VPWR VGND sg13g2_decap_8
XFILLER_24_900 VPWR VGND sg13g2_decap_8
XFILLER_23_410 VPWR VGND sg13g2_decap_8
XFILLER_24_977 VPWR VGND sg13g2_decap_8
XFILLER_11_627 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_7_609 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_3_837 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_15_900 VPWR VGND sg13g2_decap_8
XFILLER_14_410 VPWR VGND sg13g2_decap_8
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_15_977 VPWR VGND sg13g2_decap_8
XFILLER_42_763 VPWR VGND sg13g2_decap_8
XFILLER_30_903 VPWR VGND sg13g2_decap_8
XFILLER_18_1005 VPWR VGND sg13g2_decap_8
XFILLER_14_487 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_6_620 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_6_697 VPWR VGND sg13g2_decap_8
XFILLER_37_546 VPWR VGND sg13g2_decap_8
XFILLER_24_207 VPWR VGND sg13g2_decap_8
XFILLER_18_760 VPWR VGND sg13g2_decap_8
XFILLER_33_763 VPWR VGND sg13g2_decap_8
XFILLER_21_914 VPWR VGND sg13g2_decap_8
XFILLER_32_273 VPWR VGND sg13g2_decap_8
XFILLER_20_424 VPWR VGND sg13g2_decap_8
XFILLER_9_480 VPWR VGND sg13g2_decap_8
XFILLER_28_557 VPWR VGND sg13g2_decap_8
XFILLER_15_207 VPWR VGND sg13g2_decap_8
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_11_424 VPWR VGND sg13g2_decap_8
XFILLER_24_774 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_8_907 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_23_284 VPWR VGND sg13g2_decap_8
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_3_634 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_19_557 VPWR VGND sg13g2_decap_8
XFILLER_15_774 VPWR VGND sg13g2_decap_8
XFILLER_42_560 VPWR VGND sg13g2_decap_8
XFILLER_30_700 VPWR VGND sg13g2_decap_8
XFILLER_14_284 VPWR VGND sg13g2_decap_8
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_30_777 VPWR VGND sg13g2_decap_8
XFILLER_11_991 VPWR VGND sg13g2_decap_8
XFILLER_7_973 VPWR VGND sg13g2_decap_8
XFILLER_6_494 VPWR VGND sg13g2_decap_8
XFILLER_38_833 VPWR VGND sg13g2_decap_8
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_33_560 VPWR VGND sg13g2_decap_8
XFILLER_21_711 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_21_788 VPWR VGND sg13g2_decap_8
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_29_833 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_28_354 VPWR VGND sg13g2_decap_8
XFILLER_44_847 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_decap_8
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_24_571 VPWR VGND sg13g2_decap_8
XFILLER_11_221 VPWR VGND sg13g2_decap_8
XFILLER_15_1019 VPWR VGND sg13g2_decap_8
XFILLER_8_704 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_decap_8
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_3_431 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_19_354 VPWR VGND sg13g2_decap_8
XFILLER_35_847 VPWR VGND sg13g2_decap_8
XFILLER_34_357 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_30_574 VPWR VGND sg13g2_decap_8
XFILLER_7_770 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_38_630 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_38_1008 VPWR VGND sg13g2_decap_8
XFILLER_26_858 VPWR VGND sg13g2_decap_8
XFILLER_13_508 VPWR VGND sg13g2_decap_8
XFILLER_25_368 VPWR VGND sg13g2_decap_8
XFILLER_21_585 VPWR VGND sg13g2_decap_8
XFILLER_5_718 VPWR VGND sg13g2_decap_8
XFILLER_4_228 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_42 VPWR VGND sg13g2_decap_8
XFILLER_29_630 VPWR VGND sg13g2_decap_8
XFILLER_21_1012 VPWR VGND sg13g2_decap_8
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_17_847 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_44_644 VPWR VGND sg13g2_decap_8
XFILLER_16_368 VPWR VGND sg13g2_decap_8
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_8_501 VPWR VGND sg13g2_decap_8
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_12_585 VPWR VGND sg13g2_decap_8
XFILLER_8_578 VPWR VGND sg13g2_decap_8
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_4_795 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_39_427 VPWR VGND sg13g2_decap_8
XFILLER_48_994 VPWR VGND sg13g2_decap_8
XFILLER_19_151 VPWR VGND sg13g2_decap_8
XFILLER_35_644 VPWR VGND sg13g2_decap_8
XFILLER_34_154 VPWR VGND sg13g2_decap_8
XFILLER_22_305 VPWR VGND sg13g2_decap_8
XFILLER_31_861 VPWR VGND sg13g2_decap_8
XFILLER_30_371 VPWR VGND sg13g2_decap_8
XFILLER_44_1001 VPWR VGND sg13g2_decap_8
Xheichips25_template_11 VPWR VGND uo_out[5] sg13g2_tielo
Xheichips25_template_22 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_39_994 VPWR VGND sg13g2_decap_8
XFILLER_26_655 VPWR VGND sg13g2_decap_8
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_25_165 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_21_382 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_5_515 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_49_714 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_45_931 VPWR VGND sg13g2_decap_8
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_17_644 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_8
XFILLER_32_658 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_31_168 VPWR VGND sg13g2_decap_8
XFILLER_20_809 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_decap_8
XFILLER_9_865 VPWR VGND sg13g2_decap_8
XFILLER_8_375 VPWR VGND sg13g2_decap_8
XFILLER_4_592 VPWR VGND sg13g2_decap_8
XFILLER_39_224 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_36_931 VPWR VGND sg13g2_decap_8
XFILLER_35_441 VPWR VGND sg13g2_decap_8
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
XFILLER_23_669 VPWR VGND sg13g2_decap_8
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_22_179 VPWR VGND sg13g2_decap_8
XFILLER_2_529 VPWR VGND sg13g2_decap_8
XFILLER_46_728 VPWR VGND sg13g2_decap_8
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_39_791 VPWR VGND sg13g2_decap_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_26_452 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_14_669 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_decap_8
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_6_802 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_511 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_37_728 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_18_942 VPWR VGND sg13g2_decap_8
XFILLER_17_441 VPWR VGND sg13g2_decap_8
XFILLER_33_945 VPWR VGND sg13g2_decap_8
XFILLER_32_455 VPWR VGND sg13g2_decap_8
XFILLER_20_606 VPWR VGND sg13g2_decap_8
XFILLER_34_1022 VPWR VGND sg13g2_decap_8
XFILLER_9_662 VPWR VGND sg13g2_decap_8
XFILLER_8_172 VPWR VGND sg13g2_decap_8
XFILLER_41_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_739 VPWR VGND sg13g2_decap_8
XFILLER_27_238 VPWR VGND sg13g2_decap_8
XFILLER_24_956 VPWR VGND sg13g2_decap_8
XFILLER_11_606 VPWR VGND sg13g2_decap_8
XFILLER_23_466 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_19_739 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_15_956 VPWR VGND sg13g2_decap_8
XFILLER_42_742 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_14_466 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_525 VPWR VGND sg13g2_decap_8
XFILLER_49_385 VPWR VGND sg13g2_decap_8
XFILLER_33_742 VPWR VGND sg13g2_decap_8
XFILLER_32_252 VPWR VGND sg13g2_decap_8
XFILLER_20_403 VPWR VGND sg13g2_decap_8
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_536 VPWR VGND sg13g2_decap_8
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_24_753 VPWR VGND sg13g2_decap_8
XFILLER_11_403 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_3_613 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_19_536 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_34_539 VPWR VGND sg13g2_decap_8
XFILLER_15_753 VPWR VGND sg13g2_decap_8
XFILLER_14_263 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_30_756 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_7_952 VPWR VGND sg13g2_decap_8
XFILLER_6_473 VPWR VGND sg13g2_decap_8
XFILLER_9_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_38_812 VPWR VGND sg13g2_decap_8
XFILLER_49_182 VPWR VGND sg13g2_decap_8
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_38_889 VPWR VGND sg13g2_decap_8
XFILLER_37_399 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
XFILLER_21_767 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_29_812 VPWR VGND sg13g2_decap_8
XFILLER_28_333 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_29_889 VPWR VGND sg13g2_decap_8
XFILLER_44_826 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_24_550 VPWR VGND sg13g2_decap_8
XFILLER_11_200 VPWR VGND sg13g2_decap_8
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_3_410 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_39_609 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_decap_8
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_35_826 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_decap_8
XFILLER_34_336 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
XFILLER_30_553 VPWR VGND sg13g2_decap_8
XFILLER_6_270 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_29_119 VPWR VGND sg13g2_decap_8
XFILLER_38_686 VPWR VGND sg13g2_decap_8
XFILLER_26_837 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_25_347 VPWR VGND sg13g2_decap_8
XFILLER_21_564 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_29_21 VPWR VGND sg13g2_decap_8
XFILLER_29_98 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_44_623 VPWR VGND sg13g2_decap_8
XFILLER_29_686 VPWR VGND sg13g2_decap_8
XFILLER_17_826 VPWR VGND sg13g2_decap_8
XFILLER_16_347 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_8
XFILLER_40_840 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_8_557 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_decap_8
XFILLER_3_284 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_48_973 VPWR VGND sg13g2_decap_8
XFILLER_19_130 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_35_623 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
XFILLER_31_840 VPWR VGND sg13g2_decap_8
XFILLER_30_350 VPWR VGND sg13g2_decap_8
Xheichips25_template_12 VPWR VGND uo_out[6] sg13g2_tielo
Xheichips25_template_23 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_39_973 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_26_634 VPWR VGND sg13g2_decap_8
XFILLER_25_144 VPWR VGND sg13g2_decap_8
XFILLER_41_637 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_22_851 VPWR VGND sg13g2_decap_8
XFILLER_21_361 VPWR VGND sg13g2_decap_8
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_1_700 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_45_910 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_29_483 VPWR VGND sg13g2_decap_8
XFILLER_17_623 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_decap_8
XFILLER_45_987 VPWR VGND sg13g2_decap_8
XFILLER_44_497 VPWR VGND sg13g2_decap_8
XFILLER_32_637 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_31_147 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_9_844 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
XFILLER_4_571 VPWR VGND sg13g2_decap_8
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_203 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_36_910 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_35_420 VPWR VGND sg13g2_decap_8
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_35_497 VPWR VGND sg13g2_decap_8
XFILLER_23_648 VPWR VGND sg13g2_decap_8
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_508 VPWR VGND sg13g2_decap_8
XFILLER_46_707 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_39_770 VPWR VGND sg13g2_decap_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_26_431 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_14_648 VPWR VGND sg13g2_decap_8
XFILLER_42_924 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_6_858 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_37_707 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_18_921 VPWR VGND sg13g2_decap_8
XFILLER_17_420 VPWR VGND sg13g2_decap_8
XFILLER_29_280 VPWR VGND sg13g2_decap_8
XFILLER_17_497 VPWR VGND sg13g2_decap_8
XFILLER_45_784 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_18_998 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_32_434 VPWR VGND sg13g2_decap_8
XFILLER_34_1001 VPWR VGND sg13g2_decap_8
XFILLER_9_641 VPWR VGND sg13g2_decap_8
XFILLER_8_151 VPWR VGND sg13g2_decap_8
XFILLER_28_718 VPWR VGND sg13g2_decap_8
XFILLER_27_217 VPWR VGND sg13g2_decap_8
XFILLER_36_784 VPWR VGND sg13g2_decap_8
XFILLER_24_935 VPWR VGND sg13g2_decap_8
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_19_718 VPWR VGND sg13g2_decap_8
XFILLER_18_228 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_15_935 VPWR VGND sg13g2_decap_8
XFILLER_42_721 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_14_445 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_42_798 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_655 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_49_364 VPWR VGND sg13g2_decap_8
XFILLER_37_504 VPWR VGND sg13g2_decap_8
XFILLER_45_581 VPWR VGND sg13g2_decap_8
XFILLER_33_721 VPWR VGND sg13g2_decap_8
XFILLER_18_795 VPWR VGND sg13g2_decap_8
XFILLER_17_294 VPWR VGND sg13g2_decap_8
XFILLER_32_231 VPWR VGND sg13g2_decap_8
XFILLER_33_798 VPWR VGND sg13g2_decap_8
XFILLER_21_949 VPWR VGND sg13g2_decap_8
XFILLER_20_459 VPWR VGND sg13g2_decap_8
XFILLER_28_515 VPWR VGND sg13g2_decap_8
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_36_581 VPWR VGND sg13g2_decap_8
XFILLER_24_732 VPWR VGND sg13g2_decap_8
XFILLER_23_242 VPWR VGND sg13g2_decap_8
XFILLER_12_949 VPWR VGND sg13g2_decap_8
XFILLER_11_459 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_669 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_19_515 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_34_518 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_15_732 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_42_595 VPWR VGND sg13g2_decap_8
XFILLER_30_735 VPWR VGND sg13g2_decap_8
XFILLER_31_1015 VPWR VGND sg13g2_decap_8
XFILLER_7_931 VPWR VGND sg13g2_decap_8
XFILLER_6_452 VPWR VGND sg13g2_decap_8
XFILLER_9_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_38_868 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_25_529 VPWR VGND sg13g2_decap_8
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_33_595 VPWR VGND sg13g2_decap_8
XFILLER_21_746 VPWR VGND sg13g2_decap_8
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
XFILLER_28_312 VPWR VGND sg13g2_decap_8
XFILLER_44_805 VPWR VGND sg13g2_decap_8
XFILLER_29_868 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_16_529 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_28_389 VPWR VGND sg13g2_decap_8
XFILLER_12_746 VPWR VGND sg13g2_decap_8
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_8_739 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_8
XFILLER_19_312 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_34_315 VPWR VGND sg13g2_decap_8
XFILLER_19_389 VPWR VGND sg13g2_decap_8
XFILLER_43_882 VPWR VGND sg13g2_decap_8
XFILLER_42_392 VPWR VGND sg13g2_decap_8
XFILLER_30_532 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_38_665 VPWR VGND sg13g2_decap_8
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_26_816 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_25_326 VPWR VGND sg13g2_decap_8
XFILLER_41_819 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_34_882 VPWR VGND sg13g2_decap_8
XFILLER_33_392 VPWR VGND sg13g2_decap_8
XFILLER_21_543 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_29_77 VPWR VGND sg13g2_decap_8
XFILLER_29_665 VPWR VGND sg13g2_decap_8
XFILLER_17_805 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_602 VPWR VGND sg13g2_decap_8
XFILLER_16_326 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_44_679 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_decap_8
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_31_329 VPWR VGND sg13g2_decap_8
XFILLER_25_893 VPWR VGND sg13g2_decap_8
XFILLER_12_543 VPWR VGND sg13g2_decap_8
XFILLER_8_536 VPWR VGND sg13g2_decap_8
XFILLER_40_896 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
XFILLER_6_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_952 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_35_602 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_19_186 VPWR VGND sg13g2_decap_8
XFILLER_35_679 VPWR VGND sg13g2_decap_8
XFILLER_16_893 VPWR VGND sg13g2_decap_8
XFILLER_34_189 VPWR VGND sg13g2_decap_8
XFILLER_31_896 VPWR VGND sg13g2_decap_8
Xheichips25_template_13 VPWR VGND uo_out[7] sg13g2_tielo
XFILLER_39_952 VPWR VGND sg13g2_decap_8
XFILLER_38_462 VPWR VGND sg13g2_decap_8
XFILLER_26_613 VPWR VGND sg13g2_decap_8
XFILLER_25_123 VPWR VGND sg13g2_decap_8
XFILLER_41_616 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_22_830 VPWR VGND sg13g2_decap_8
XFILLER_21_340 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_49_749 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_29_462 VPWR VGND sg13g2_decap_8
XFILLER_17_602 VPWR VGND sg13g2_decap_8
XFILLER_16_123 VPWR VGND sg13g2_decap_8
XFILLER_45_966 VPWR VGND sg13g2_decap_8
XFILLER_17_679 VPWR VGND sg13g2_decap_8
XFILLER_44_476 VPWR VGND sg13g2_decap_8
XFILLER_32_616 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_31_126 VPWR VGND sg13g2_decap_8
XFILLER_25_690 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
XFILLER_40_693 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_8
XFILLER_39_259 VPWR VGND sg13g2_decap_8
XFILLER_36_966 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
XFILLER_16_690 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_decap_8
XFILLER_31_693 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_26_410 VPWR VGND sg13g2_decap_8
XFILLER_42_903 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_14_627 VPWR VGND sg13g2_decap_8
XFILLER_41_413 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_6_837 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_45_763 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_18_977 VPWR VGND sg13g2_decap_8
XFILLER_17_476 VPWR VGND sg13g2_decap_8
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_32_413 VPWR VGND sg13g2_decap_8
XFILLER_9_620 VPWR VGND sg13g2_decap_8
XFILLER_41_980 VPWR VGND sg13g2_decap_8
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_40_490 VPWR VGND sg13g2_decap_8
XFILLER_9_697 VPWR VGND sg13g2_decap_8
XFILLER_36_763 VPWR VGND sg13g2_decap_8
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_24_914 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_32_980 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_31_490 VPWR VGND sg13g2_decap_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_15_914 VPWR VGND sg13g2_decap_8
XFILLER_42_700 VPWR VGND sg13g2_decap_8
XFILLER_14_424 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_18_1019 VPWR VGND sg13g2_decap_8
XFILLER_42_777 VPWR VGND sg13g2_decap_8
XFILLER_30_917 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_23_991 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
XFILLER_17_273 VPWR VGND sg13g2_decap_8
XFILLER_45_560 VPWR VGND sg13g2_decap_8
XFILLER_33_700 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_decap_8
XFILLER_32_210 VPWR VGND sg13g2_decap_8
XFILLER_33_777 VPWR VGND sg13g2_decap_8
XFILLER_21_928 VPWR VGND sg13g2_decap_8
XFILLER_14_991 VPWR VGND sg13g2_decap_8
XFILLER_32_287 VPWR VGND sg13g2_decap_8
XFILLER_20_438 VPWR VGND sg13g2_decap_8
XFILLER_9_494 VPWR VGND sg13g2_decap_8
XFILLER_4_81 VPWR VGND sg13g2_decap_8
XFILLER_36_560 VPWR VGND sg13g2_decap_8
XFILLER_24_711 VPWR VGND sg13g2_decap_8
XFILLER_23_221 VPWR VGND sg13g2_decap_8
XFILLER_12_928 VPWR VGND sg13g2_decap_8
XFILLER_24_788 VPWR VGND sg13g2_decap_8
XFILLER_11_438 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_8
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_15_788 VPWR VGND sg13g2_decap_8
XFILLER_42_574 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
XFILLER_14_298 VPWR VGND sg13g2_decap_8
XFILLER_7_910 VPWR VGND sg13g2_decap_8
XFILLER_6_431 VPWR VGND sg13g2_decap_8
XFILLER_7_987 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_140 VPWR VGND sg13g2_decap_8
XFILLER_38_847 VPWR VGND sg13g2_decap_8
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_25_508 VPWR VGND sg13g2_decap_8
XFILLER_18_571 VPWR VGND sg13g2_decap_8
XFILLER_33_574 VPWR VGND sg13g2_decap_8
XFILLER_21_725 VPWR VGND sg13g2_decap_8
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
XFILLER_29_847 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_16_508 VPWR VGND sg13g2_decap_8
XFILLER_28_368 VPWR VGND sg13g2_decap_8
XFILLER_12_725 VPWR VGND sg13g2_decap_8
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_24_585 VPWR VGND sg13g2_decap_8
XFILLER_11_235 VPWR VGND sg13g2_decap_8
XFILLER_8_718 VPWR VGND sg13g2_decap_8
XFILLER_7_217 VPWR VGND sg13g2_decap_8
XFILLER_4_935 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_19_368 VPWR VGND sg13g2_decap_8
XFILLER_43_861 VPWR VGND sg13g2_decap_8
XFILLER_15_585 VPWR VGND sg13g2_decap_8
XFILLER_42_371 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_decap_8
XFILLER_30_588 VPWR VGND sg13g2_decap_8
XFILLER_7_784 VPWR VGND sg13g2_decap_8
XFILLER_38_644 VPWR VGND sg13g2_decap_8
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_25_305 VPWR VGND sg13g2_decap_8
XFILLER_40_308 VPWR VGND sg13g2_decap_8
XFILLER_34_861 VPWR VGND sg13g2_decap_8
XFILLER_33_371 VPWR VGND sg13g2_decap_8
XFILLER_21_522 VPWR VGND sg13g2_decap_8
XFILLER_21_599 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_1_938 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_56 VPWR VGND sg13g2_decap_8
XFILLER_29_644 VPWR VGND sg13g2_decap_8
XFILLER_21_1026 VPWR VGND sg13g2_fill_2
XFILLER_16_305 VPWR VGND sg13g2_decap_8
XFILLER_28_165 VPWR VGND sg13g2_decap_8
XFILLER_44_658 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_31_308 VPWR VGND sg13g2_decap_8
XFILLER_25_872 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_24_382 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_decap_8
XFILLER_40_875 VPWR VGND sg13g2_decap_8
XFILLER_12_599 VPWR VGND sg13g2_decap_8
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_3_242 VPWR VGND sg13g2_decap_8
XFILLER_48_931 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_165 VPWR VGND sg13g2_decap_8
XFILLER_35_658 VPWR VGND sg13g2_decap_8
XFILLER_23_809 VPWR VGND sg13g2_decap_8
XFILLER_16_872 VPWR VGND sg13g2_decap_8
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
XFILLER_34_168 VPWR VGND sg13g2_decap_8
XFILLER_22_319 VPWR VGND sg13g2_decap_8
XFILLER_15_382 VPWR VGND sg13g2_decap_8
XFILLER_31_875 VPWR VGND sg13g2_decap_8
XFILLER_30_385 VPWR VGND sg13g2_decap_8
XFILLER_7_581 VPWR VGND sg13g2_decap_8
XFILLER_44_1015 VPWR VGND sg13g2_decap_8
Xheichips25_template_14 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_39_931 VPWR VGND sg13g2_decap_8
XFILLER_38_441 VPWR VGND sg13g2_decap_8
XFILLER_25_102 VPWR VGND sg13g2_decap_8
XFILLER_14_809 VPWR VGND sg13g2_decap_8
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_25_179 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_decap_8
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_21_396 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_decap_8
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_49_728 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_29_441 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_decap_8
XFILLER_45_945 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_17_658 VPWR VGND sg13g2_decap_8
XFILLER_16_179 VPWR VGND sg13g2_decap_8
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_9_802 VPWR VGND sg13g2_decap_8
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_40_672 VPWR VGND sg13g2_decap_8
XFILLER_12_396 VPWR VGND sg13g2_decap_8
XFILLER_9_879 VPWR VGND sg13g2_decap_8
XFILLER_8_389 VPWR VGND sg13g2_decap_8
XFILLER_39_238 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_36_945 VPWR VGND sg13g2_decap_8
XFILLER_35_455 VPWR VGND sg13g2_decap_8
XFILLER_23_606 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_31_672 VPWR VGND sg13g2_decap_8
XFILLER_30_182 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_decap_8
XFILLER_14_606 VPWR VGND sg13g2_decap_8
XFILLER_26_466 VPWR VGND sg13g2_decap_8
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_6_816 VPWR VGND sg13g2_decap_8
XFILLER_21_193 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_17_455 VPWR VGND sg13g2_decap_8
XFILLER_45_742 VPWR VGND sg13g2_decap_8
XFILLER_18_956 VPWR VGND sg13g2_decap_8
XFILLER_44_252 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_32_469 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_decap_8
XFILLER_9_676 VPWR VGND sg13g2_decap_8
XFILLER_8_186 VPWR VGND sg13g2_decap_8
XFILLER_5_893 VPWR VGND sg13g2_decap_8
XFILLER_36_742 VPWR VGND sg13g2_decap_8
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_23_403 VPWR VGND sg13g2_decap_8
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_14_403 VPWR VGND sg13g2_decap_8
XFILLER_26_263 VPWR VGND sg13g2_decap_8
XFILLER_42_756 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_decap_8
XFILLER_22_480 VPWR VGND sg13g2_decap_8
XFILLER_6_613 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_49_322 VPWR VGND sg13g2_decap_8
XFILLER_49_399 VPWR VGND sg13g2_decap_8
XFILLER_37_539 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_17_252 VPWR VGND sg13g2_decap_8
XFILLER_33_756 VPWR VGND sg13g2_decap_8
XFILLER_32_266 VPWR VGND sg13g2_decap_8
XFILLER_21_907 VPWR VGND sg13g2_decap_8
XFILLER_14_970 VPWR VGND sg13g2_decap_8
XFILLER_20_417 VPWR VGND sg13g2_decap_8
XFILLER_13_480 VPWR VGND sg13g2_decap_8
Xheichips25_template_1 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_9_473 VPWR VGND sg13g2_decap_8
XFILLER_5_690 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_24_767 VPWR VGND sg13g2_decap_8
XFILLER_11_417 VPWR VGND sg13g2_decap_8
XFILLER_23_277 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_20_984 VPWR VGND sg13g2_decap_8
XFILLER_3_627 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_14_200 VPWR VGND sg13g2_decap_8
XFILLER_15_767 VPWR VGND sg13g2_decap_8
XFILLER_42_553 VPWR VGND sg13g2_decap_8
XFILLER_14_277 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_6_410 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_7_966 VPWR VGND sg13g2_decap_8
XFILLER_6_487 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_38_826 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_8
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_18_550 VPWR VGND sg13g2_decap_8
XFILLER_33_553 VPWR VGND sg13g2_decap_8
XFILLER_21_704 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
XFILLER_9_270 VPWR VGND sg13g2_decap_8
XFILLER_29_826 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_decap_8
XFILLER_12_704 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_decap_8
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_20_781 VPWR VGND sg13g2_decap_8
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_3_424 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_19_347 VPWR VGND sg13g2_decap_8
XFILLER_43_840 VPWR VGND sg13g2_decap_8
XFILLER_15_564 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_11_781 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_decap_8
XFILLER_7_763 VPWR VGND sg13g2_decap_8
XFILLER_6_284 VPWR VGND sg13g2_decap_8
XFILLER_3_991 VPWR VGND sg13g2_decap_8
XFILLER_38_623 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_34_840 VPWR VGND sg13g2_decap_8
XFILLER_33_350 VPWR VGND sg13g2_decap_8
XFILLER_21_501 VPWR VGND sg13g2_decap_8
XFILLER_14_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_578 VPWR VGND sg13g2_decap_8
XFILLER_1_917 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_35 VPWR VGND sg13g2_decap_8
XFILLER_29_623 VPWR VGND sg13g2_decap_8
XFILLER_21_1005 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_44_637 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_25_851 VPWR VGND sg13g2_decap_8
XFILLER_12_501 VPWR VGND sg13g2_decap_8
XFILLER_24_361 VPWR VGND sg13g2_decap_8
XFILLER_40_854 VPWR VGND sg13g2_decap_8
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_48_987 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_35_637 VPWR VGND sg13g2_decap_8
XFILLER_16_851 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_34_147 VPWR VGND sg13g2_decap_8
XFILLER_15_361 VPWR VGND sg13g2_decap_8
XFILLER_31_854 VPWR VGND sg13g2_decap_8
XFILLER_30_364 VPWR VGND sg13g2_decap_8
XFILLER_7_560 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_39_910 VPWR VGND sg13g2_decap_8
Xheichips25_template_15 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_38_420 VPWR VGND sg13g2_decap_8
XFILLER_39_987 VPWR VGND sg13g2_decap_8
XFILLER_38_497 VPWR VGND sg13g2_decap_8
XFILLER_26_648 VPWR VGND sg13g2_decap_8
XFILLER_25_158 VPWR VGND sg13g2_decap_8
XFILLER_22_865 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
XFILLER_21_375 VPWR VGND sg13g2_decap_8
XFILLER_5_508 VPWR VGND sg13g2_decap_8
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_29_420 VPWR VGND sg13g2_decap_8
XFILLER_45_924 VPWR VGND sg13g2_decap_8
XFILLER_29_497 VPWR VGND sg13g2_decap_8
XFILLER_17_637 VPWR VGND sg13g2_decap_8
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_16_158 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_40_651 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_decap_8
XFILLER_9_858 VPWR VGND sg13g2_decap_8
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_4_585 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_8
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_36_924 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_35_434 VPWR VGND sg13g2_decap_8
XFILLER_31_651 VPWR VGND sg13g2_decap_8
XFILLER_30_161 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_784 VPWR VGND sg13g2_decap_8
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_26_445 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_42_938 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_22_662 VPWR VGND sg13g2_decap_8
XFILLER_21_172 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_45_721 VPWR VGND sg13g2_decap_8
XFILLER_18_935 VPWR VGND sg13g2_decap_8
XFILLER_17_434 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_29_294 VPWR VGND sg13g2_decap_8
XFILLER_45_798 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_32_448 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_34_1015 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
XFILLER_5_872 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_decap_8
XFILLER_41_1008 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_721 VPWR VGND sg13g2_decap_8
XFILLER_35_231 VPWR VGND sg13g2_decap_8
XFILLER_36_798 VPWR VGND sg13g2_decap_8
XFILLER_24_949 VPWR VGND sg13g2_decap_8
XFILLER_23_459 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_2_319 VPWR VGND sg13g2_decap_8
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_39_581 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_26_242 VPWR VGND sg13g2_decap_8
XFILLER_15_949 VPWR VGND sg13g2_decap_8
XFILLER_42_735 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_14_459 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_6_669 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_49_301 VPWR VGND sg13g2_decap_8
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_49_378 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_decap_8
XFILLER_18_732 VPWR VGND sg13g2_decap_8
XFILLER_17_231 VPWR VGND sg13g2_decap_8
XFILLER_45_595 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_decap_8
XFILLER_32_245 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_decap_8
Xheichips25_template_2 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_28_529 VPWR VGND sg13g2_decap_8
XFILLER_36_595 VPWR VGND sg13g2_decap_8
XFILLER_24_746 VPWR VGND sg13g2_decap_8
XFILLER_23_256 VPWR VGND sg13g2_decap_8
XFILLER_20_963 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_19_529 VPWR VGND sg13g2_decap_8
XFILLER_15_746 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_14_256 VPWR VGND sg13g2_decap_8
XFILLER_42_532 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_7_945 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_9_1019 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_38_805 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_49_175 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
XFILLER_33_532 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_805 VPWR VGND sg13g2_decap_8
XFILLER_28_326 VPWR VGND sg13g2_decap_8
XFILLER_44_819 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_decap_8
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_24_543 VPWR VGND sg13g2_decap_8
XFILLER_20_760 VPWR VGND sg13g2_decap_8
XFILLER_3_403 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_8
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_35_819 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_34_329 VPWR VGND sg13g2_decap_8
XFILLER_28_893 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_27_392 VPWR VGND sg13g2_decap_8
XFILLER_43_896 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_decap_8
XFILLER_11_760 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_7_742 VPWR VGND sg13g2_decap_8
XFILLER_6_263 VPWR VGND sg13g2_decap_8
XFILLER_3_970 VPWR VGND sg13g2_decap_8
XFILLER_2_480 VPWR VGND sg13g2_decap_8
XFILLER_38_602 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_38_679 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_19_893 VPWR VGND sg13g2_decap_8
XFILLER_34_896 VPWR VGND sg13g2_decap_8
XFILLER_21_557 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_29_14 VPWR VGND sg13g2_decap_8
XFILLER_29_602 VPWR VGND sg13g2_decap_8
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_29_679 VPWR VGND sg13g2_decap_8
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_17_819 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_44_616 VPWR VGND sg13g2_decap_8
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_25_830 VPWR VGND sg13g2_decap_8
XFILLER_24_340 VPWR VGND sg13g2_decap_8
XFILLER_40_833 VPWR VGND sg13g2_decap_8
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_3_200 VPWR VGND sg13g2_decap_8
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_48_966 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_35_616 VPWR VGND sg13g2_decap_8
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_decap_8
XFILLER_28_690 VPWR VGND sg13g2_decap_8
XFILLER_15_340 VPWR VGND sg13g2_decap_8
XFILLER_43_693 VPWR VGND sg13g2_decap_8
XFILLER_31_833 VPWR VGND sg13g2_decap_8
XFILLER_30_343 VPWR VGND sg13g2_decap_8
Xheichips25_template_16 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_39_966 VPWR VGND sg13g2_decap_8
XFILLER_38_476 VPWR VGND sg13g2_decap_8
XFILLER_26_627 VPWR VGND sg13g2_decap_8
XFILLER_25_137 VPWR VGND sg13g2_decap_8
XFILLER_19_690 VPWR VGND sg13g2_decap_8
XFILLER_34_693 VPWR VGND sg13g2_decap_8
XFILLER_22_844 VPWR VGND sg13g2_decap_8
XFILLER_21_354 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_45_903 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_29_476 VPWR VGND sg13g2_decap_8
XFILLER_17_616 VPWR VGND sg13g2_decap_8
XFILLER_16_137 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_40_630 VPWR VGND sg13g2_decap_8
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_9_837 VPWR VGND sg13g2_decap_8
XFILLER_8_347 VPWR VGND sg13g2_decap_8
XFILLER_21_81 VPWR VGND sg13g2_decap_8
XFILLER_4_564 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_36_903 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_35_413 VPWR VGND sg13g2_decap_8
XFILLER_44_980 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_31_630 VPWR VGND sg13g2_decap_8
XFILLER_30_140 VPWR VGND sg13g2_decap_8
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_763 VPWR VGND sg13g2_decap_8
XFILLER_27_903 VPWR VGND sg13g2_decap_8
XFILLER_38_273 VPWR VGND sg13g2_decap_8
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_42_917 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_35_980 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_34_490 VPWR VGND sg13g2_decap_8
XFILLER_22_641 VPWR VGND sg13g2_decap_8
XFILLER_21_151 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_decap_8
XFILLER_45_700 VPWR VGND sg13g2_decap_8
XFILLER_29_273 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_45_777 VPWR VGND sg13g2_decap_8
XFILLER_33_917 VPWR VGND sg13g2_decap_8
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_32_427 VPWR VGND sg13g2_decap_8
XFILLER_26_991 VPWR VGND sg13g2_decap_8
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_16_81 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_9_634 VPWR VGND sg13g2_decap_8
XFILLER_41_994 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
XFILLER_32_91 VPWR VGND sg13g2_decap_8
XFILLER_5_851 VPWR VGND sg13g2_decap_8
XFILLER_4_361 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_36_700 VPWR VGND sg13g2_decap_8
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_36_777 VPWR VGND sg13g2_decap_8
XFILLER_24_928 VPWR VGND sg13g2_decap_8
XFILLER_35_287 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_17_980 VPWR VGND sg13g2_decap_8
XFILLER_32_994 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_39_560 VPWR VGND sg13g2_decap_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_15_928 VPWR VGND sg13g2_decap_8
XFILLER_42_714 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_14_438 VPWR VGND sg13g2_decap_8
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_648 VPWR VGND sg13g2_decap_8
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_357 VPWR VGND sg13g2_decap_8
XFILLER_18_711 VPWR VGND sg13g2_decap_8
XFILLER_17_210 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_17_287 VPWR VGND sg13g2_decap_8
XFILLER_45_574 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_32_224 VPWR VGND sg13g2_decap_8
XFILLER_9_431 VPWR VGND sg13g2_decap_8
XFILLER_41_791 VPWR VGND sg13g2_decap_8
Xheichips25_template_3 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_28_508 VPWR VGND sg13g2_decap_8
XFILLER_36_574 VPWR VGND sg13g2_decap_8
XFILLER_24_725 VPWR VGND sg13g2_decap_8
XFILLER_23_235 VPWR VGND sg13g2_decap_8
XFILLER_17_1022 VPWR VGND sg13g2_decap_8
XFILLER_32_791 VPWR VGND sg13g2_decap_8
XFILLER_20_942 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_508 VPWR VGND sg13g2_decap_8
XFILLER_15_725 VPWR VGND sg13g2_decap_8
XFILLER_42_511 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_14_235 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_42_588 VPWR VGND sg13g2_decap_8
XFILLER_30_728 VPWR VGND sg13g2_decap_8
XFILLER_11_942 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_7_924 VPWR VGND sg13g2_decap_8
XFILLER_31_1008 VPWR VGND sg13g2_decap_8
XFILLER_6_445 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_29_7 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_8
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_33_511 VPWR VGND sg13g2_decap_8
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_33_588 VPWR VGND sg13g2_decap_8
XFILLER_21_739 VPWR VGND sg13g2_decap_8
XFILLER_20_249 VPWR VGND sg13g2_decap_8
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_305 VPWR VGND sg13g2_decap_8
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_37_861 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_24_522 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
XFILLER_24_599 VPWR VGND sg13g2_decap_8
XFILLER_11_249 VPWR VGND sg13g2_decap_8
XFILLER_4_949 VPWR VGND sg13g2_decap_8
XFILLER_3_459 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_34_308 VPWR VGND sg13g2_decap_8
XFILLER_28_872 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_43_875 VPWR VGND sg13g2_decap_8
XFILLER_15_599 VPWR VGND sg13g2_decap_8
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_30_525 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_7_721 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_7_798 VPWR VGND sg13g2_decap_8
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_38_658 VPWR VGND sg13g2_decap_8
XFILLER_26_809 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_25_319 VPWR VGND sg13g2_decap_8
XFILLER_19_872 VPWR VGND sg13g2_decap_8
XFILLER_18_382 VPWR VGND sg13g2_decap_8
XFILLER_34_875 VPWR VGND sg13g2_decap_8
XFILLER_33_385 VPWR VGND sg13g2_decap_8
XFILLER_21_536 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_29_658 VPWR VGND sg13g2_decap_8
XFILLER_16_319 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_40_812 VPWR VGND sg13g2_decap_8
XFILLER_25_886 VPWR VGND sg13g2_decap_8
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_24_396 VPWR VGND sg13g2_decap_8
XFILLER_40_889 VPWR VGND sg13g2_decap_8
XFILLER_8_529 VPWR VGND sg13g2_decap_8
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_48_945 VPWR VGND sg13g2_decap_8
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_decap_8
XFILLER_19_179 VPWR VGND sg13g2_decap_8
XFILLER_16_886 VPWR VGND sg13g2_decap_8
XFILLER_43_672 VPWR VGND sg13g2_decap_8
XFILLER_31_812 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_30_322 VPWR VGND sg13g2_decap_8
XFILLER_31_889 VPWR VGND sg13g2_decap_8
XFILLER_30_399 VPWR VGND sg13g2_decap_8
XFILLER_7_595 VPWR VGND sg13g2_decap_8
Xheichips25_template_17 VPWR VGND uio_oe[3] sg13g2_tielo
XFILLER_39_945 VPWR VGND sg13g2_decap_8
XFILLER_38_455 VPWR VGND sg13g2_decap_8
XFILLER_26_606 VPWR VGND sg13g2_decap_8
XFILLER_25_116 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_41_609 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_34_672 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_21_333 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_decap_8
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_5_1012 VPWR VGND sg13g2_decap_8
XFILLER_29_455 VPWR VGND sg13g2_decap_8
XFILLER_16_116 VPWR VGND sg13g2_decap_8
XFILLER_45_959 VPWR VGND sg13g2_decap_8
XFILLER_44_469 VPWR VGND sg13g2_decap_8
XFILLER_32_609 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_31_119 VPWR VGND sg13g2_decap_8
XFILLER_25_683 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_4_543 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_36_959 VPWR VGND sg13g2_decap_8
XFILLER_35_469 VPWR VGND sg13g2_decap_8
XFILLER_16_683 VPWR VGND sg13g2_decap_8
XFILLER_15_193 VPWR VGND sg13g2_decap_8
XFILLER_31_686 VPWR VGND sg13g2_decap_8
XFILLER_30_196 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_392 VPWR VGND sg13g2_decap_8
XFILLER_8_893 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_39_742 VPWR VGND sg13g2_decap_8
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_26_403 VPWR VGND sg13g2_decap_8
XFILLER_27_959 VPWR VGND sg13g2_decap_8
XFILLER_41_406 VPWR VGND sg13g2_decap_8
XFILLER_22_620 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_22_697 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_29_252 VPWR VGND sg13g2_decap_8
XFILLER_17_469 VPWR VGND sg13g2_decap_8
XFILLER_45_756 VPWR VGND sg13g2_decap_8
XFILLER_32_406 VPWR VGND sg13g2_decap_8
XFILLER_16_60 VPWR VGND sg13g2_decap_8
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_26_970 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_25_480 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_9_613 VPWR VGND sg13g2_decap_8
XFILLER_41_973 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_32_70 VPWR VGND sg13g2_decap_8
XFILLER_5_830 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
XFILLER_36_756 VPWR VGND sg13g2_decap_8
XFILLER_24_907 VPWR VGND sg13g2_decap_8
XFILLER_35_266 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
XFILLER_16_480 VPWR VGND sg13g2_decap_8
XFILLER_32_973 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_483 VPWR VGND sg13g2_decap_8
XFILLER_8_690 VPWR VGND sg13g2_decap_8
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_15_907 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_14_417 VPWR VGND sg13g2_decap_8
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_22_494 VPWR VGND sg13g2_decap_8
XFILLER_6_627 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_45_553 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_18_767 VPWR VGND sg13g2_decap_8
XFILLER_17_266 VPWR VGND sg13g2_decap_8
XFILLER_32_203 VPWR VGND sg13g2_decap_8
XFILLER_14_984 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_41_770 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
Xheichips25_template_4 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_9_487 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_decap_8
XFILLER_36_553 VPWR VGND sg13g2_decap_8
XFILLER_24_704 VPWR VGND sg13g2_decap_8
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_17_1001 VPWR VGND sg13g2_decap_8
XFILLER_32_770 VPWR VGND sg13g2_decap_8
XFILLER_31_280 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_20_921 VPWR VGND sg13g2_decap_8
XFILLER_20_998 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_15_704 VPWR VGND sg13g2_decap_8
XFILLER_14_214 VPWR VGND sg13g2_decap_8
XFILLER_42_567 VPWR VGND sg13g2_decap_8
XFILLER_30_707 VPWR VGND sg13g2_decap_8
XFILLER_11_921 VPWR VGND sg13g2_decap_8
XFILLER_23_781 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_7_903 VPWR VGND sg13g2_decap_8
XFILLER_22_291 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_6_424 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_46_840 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_33_567 VPWR VGND sg13g2_decap_8
XFILLER_21_718 VPWR VGND sg13g2_decap_8
XFILLER_14_781 VPWR VGND sg13g2_decap_8
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_13_291 VPWR VGND sg13g2_decap_8
XFILLER_9_284 VPWR VGND sg13g2_decap_8
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
XFILLER_37_840 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_24_501 VPWR VGND sg13g2_decap_8
XFILLER_12_718 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
XFILLER_24_578 VPWR VGND sg13g2_decap_8
XFILLER_11_228 VPWR VGND sg13g2_decap_8
XFILLER_20_795 VPWR VGND sg13g2_decap_8
XFILLER_4_928 VPWR VGND sg13g2_decap_8
XFILLER_3_438 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_28_851 VPWR VGND sg13g2_decap_8
XFILLER_15_501 VPWR VGND sg13g2_decap_8
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_43_854 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_8
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_30_504 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_7_700 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_7_777 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_38_637 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_19_851 VPWR VGND sg13g2_decap_8
XFILLER_18_361 VPWR VGND sg13g2_decap_8
XFILLER_34_854 VPWR VGND sg13g2_decap_8
XFILLER_33_364 VPWR VGND sg13g2_decap_8
XFILLER_21_515 VPWR VGND sg13g2_decap_8
XFILLER_14_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_18 VPWR VGND sg13g2_decap_8
XFILLER_29_49 VPWR VGND sg13g2_decap_8
XFILLER_29_637 VPWR VGND sg13g2_decap_8
XFILLER_21_1019 VPWR VGND sg13g2_decap_8
XFILLER_28_158 VPWR VGND sg13g2_decap_8
XFILLER_25_865 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_decap_8
XFILLER_24_375 VPWR VGND sg13g2_decap_8
XFILLER_8_508 VPWR VGND sg13g2_decap_8
XFILLER_40_868 VPWR VGND sg13g2_decap_8
XFILLER_20_592 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_3_235 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_19_158 VPWR VGND sg13g2_decap_8
XFILLER_16_865 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_decap_8
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_decap_8
XFILLER_31_868 VPWR VGND sg13g2_decap_8
XFILLER_30_378 VPWR VGND sg13g2_decap_8
XFILLER_11_592 VPWR VGND sg13g2_decap_8
XFILLER_7_574 VPWR VGND sg13g2_decap_8
XFILLER_44_1008 VPWR VGND sg13g2_decap_8
Xheichips25_template_18 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_39_924 VPWR VGND sg13g2_decap_8
XFILLER_38_434 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_decap_8
XFILLER_22_802 VPWR VGND sg13g2_decap_8
XFILLER_33_161 VPWR VGND sg13g2_decap_8
XFILLER_21_312 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
XFILLER_21_389 VPWR VGND sg13g2_decap_8
XFILLER_31_28 VPWR VGND sg13g2_decap_8
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_434 VPWR VGND sg13g2_decap_8
XFILLER_45_938 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_25_662 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_24_172 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_40_665 VPWR VGND sg13g2_decap_8
XFILLER_12_389 VPWR VGND sg13g2_decap_8
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_36_938 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_35_448 VPWR VGND sg13g2_decap_8
XFILLER_16_662 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_8
XFILLER_31_665 VPWR VGND sg13g2_decap_8
XFILLER_30_175 VPWR VGND sg13g2_decap_8
XFILLER_8_872 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_7_371 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
XFILLER_39_721 VPWR VGND sg13g2_decap_8
XFILLER_38_231 VPWR VGND sg13g2_decap_8
XFILLER_39_798 VPWR VGND sg13g2_decap_8
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_22_676 VPWR VGND sg13g2_decap_8
XFILLER_6_809 VPWR VGND sg13g2_decap_8
XFILLER_21_186 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
XFILLER_29_231 VPWR VGND sg13g2_decap_8
XFILLER_45_735 VPWR VGND sg13g2_decap_8
XFILLER_18_949 VPWR VGND sg13g2_decap_8
XFILLER_17_448 VPWR VGND sg13g2_decap_8
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_41_952 VPWR VGND sg13g2_decap_8
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_12_186 VPWR VGND sg13g2_decap_8
XFILLER_9_669 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_5_886 VPWR VGND sg13g2_decap_8
XFILLER_4_396 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_36_735 VPWR VGND sg13g2_decap_8
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_32_952 VPWR VGND sg13g2_decap_8
XFILLER_31_462 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_595 VPWR VGND sg13g2_decap_8
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_26_256 VPWR VGND sg13g2_decap_8
XFILLER_42_749 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_23_963 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_22_473 VPWR VGND sg13g2_decap_8
XFILLER_6_606 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_17_245 VPWR VGND sg13g2_decap_8
XFILLER_45_532 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_33_749 VPWR VGND sg13g2_decap_8
XFILLER_14_963 VPWR VGND sg13g2_decap_8
XFILLER_32_259 VPWR VGND sg13g2_decap_8
XFILLER_13_473 VPWR VGND sg13g2_decap_8
XFILLER_43_70 VPWR VGND sg13g2_decap_8
Xheichips25_template_5 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_9_466 VPWR VGND sg13g2_decap_8
XFILLER_5_683 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_49_882 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_36_532 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_20_900 VPWR VGND sg13g2_decap_8
XFILLER_20_977 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_42_546 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_8
XFILLER_23_760 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_22_270 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_6_403 VPWR VGND sg13g2_decap_8
XFILLER_7_959 VPWR VGND sg13g2_decap_8
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
XFILLER_38_819 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_18_543 VPWR VGND sg13g2_decap_8
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_33_546 VPWR VGND sg13g2_decap_8
XFILLER_14_760 VPWR VGND sg13g2_decap_8
XFILLER_13_270 VPWR VGND sg13g2_decap_8
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_9_263 VPWR VGND sg13g2_decap_8
XFILLER_6_970 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
XFILLER_29_819 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_24_557 VPWR VGND sg13g2_decap_8
XFILLER_11_207 VPWR VGND sg13g2_decap_8
XFILLER_20_774 VPWR VGND sg13g2_decap_8
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_28_830 VPWR VGND sg13g2_decap_8
XFILLER_43_833 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_6_200 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_7_756 VPWR VGND sg13g2_decap_8
XFILLER_6_277 VPWR VGND sg13g2_decap_8
XFILLER_3_984 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_38_616 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_19_830 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_8
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_34_833 VPWR VGND sg13g2_decap_8
XFILLER_33_343 VPWR VGND sg13g2_decap_8
XFILLER_14_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_28 VPWR VGND sg13g2_decap_8
XFILLER_29_616 VPWR VGND sg13g2_decap_8
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_37_693 VPWR VGND sg13g2_decap_8
XFILLER_25_844 VPWR VGND sg13g2_decap_8
XFILLER_24_354 VPWR VGND sg13g2_decap_8
XFILLER_40_847 VPWR VGND sg13g2_decap_8
XFILLER_20_571 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_16_844 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_31_847 VPWR VGND sg13g2_decap_8
XFILLER_30_357 VPWR VGND sg13g2_decap_8
XFILLER_11_571 VPWR VGND sg13g2_decap_8
XFILLER_7_553 VPWR VGND sg13g2_decap_8
XFILLER_3_781 VPWR VGND sg13g2_decap_8
XFILLER_39_903 VPWR VGND sg13g2_decap_8
XFILLER_2_291 VPWR VGND sg13g2_decap_8
Xheichips25_template_19 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_38_413 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_34_630 VPWR VGND sg13g2_decap_8
XFILLER_33_140 VPWR VGND sg13g2_decap_8
XFILLER_22_858 VPWR VGND sg13g2_decap_8
XFILLER_21_368 VPWR VGND sg13g2_decap_8
XFILLER_1_707 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_29_413 VPWR VGND sg13g2_decap_8
XFILLER_45_917 VPWR VGND sg13g2_decap_8
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_38_980 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_25_641 VPWR VGND sg13g2_decap_8
XFILLER_24_151 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_40_644 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_decap_8
XFILLER_4_578 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_36_917 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_35_427 VPWR VGND sg13g2_decap_8
XFILLER_29_980 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_44_994 VPWR VGND sg13g2_decap_8
XFILLER_31_644 VPWR VGND sg13g2_decap_8
XFILLER_30_154 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_8_851 VPWR VGND sg13g2_decap_8
XFILLER_39_700 VPWR VGND sg13g2_decap_8
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_39_777 VPWR VGND sg13g2_decap_8
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_38_287 VPWR VGND sg13g2_decap_8
XFILLER_26_438 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_35_994 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_22_655 VPWR VGND sg13g2_decap_8
XFILLER_21_165 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_210 VPWR VGND sg13g2_decap_8
XFILLER_17_427 VPWR VGND sg13g2_decap_8
XFILLER_45_714 VPWR VGND sg13g2_decap_8
XFILLER_29_287 VPWR VGND sg13g2_decap_8
XFILLER_18_928 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_16_95 VPWR VGND sg13g2_decap_8
XFILLER_41_931 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_40_441 VPWR VGND sg13g2_decap_8
XFILLER_34_1008 VPWR VGND sg13g2_decap_8
XFILLER_12_165 VPWR VGND sg13g2_decap_8
XFILLER_9_648 VPWR VGND sg13g2_decap_8
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_5_865 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_36_714 VPWR VGND sg13g2_decap_8
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_44_791 VPWR VGND sg13g2_decap_8
XFILLER_32_931 VPWR VGND sg13g2_decap_8
XFILLER_17_994 VPWR VGND sg13g2_decap_8
XFILLER_31_441 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_39_574 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_26_235 VPWR VGND sg13g2_decap_8
XFILLER_42_728 VPWR VGND sg13g2_decap_8
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_35_791 VPWR VGND sg13g2_decap_8
XFILLER_23_942 VPWR VGND sg13g2_decap_8
XFILLER_22_452 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_45_511 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_decap_8
XFILLER_17_224 VPWR VGND sg13g2_decap_8
XFILLER_45_588 VPWR VGND sg13g2_decap_8
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_14_942 VPWR VGND sg13g2_decap_8
XFILLER_32_238 VPWR VGND sg13g2_decap_8
XFILLER_13_452 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_decap_8
Xheichips25_template_6 VPWR VGND uo_out[0] sg13g2_tielo
XFILLER_5_662 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_49_861 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_36_511 VPWR VGND sg13g2_decap_8
XFILLER_36_588 VPWR VGND sg13g2_decap_8
XFILLER_24_739 VPWR VGND sg13g2_decap_8
XFILLER_17_791 VPWR VGND sg13g2_decap_8
XFILLER_23_249 VPWR VGND sg13g2_decap_8
XFILLER_20_956 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_15_739 VPWR VGND sg13g2_decap_8
XFILLER_42_525 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_14_249 VPWR VGND sg13g2_decap_8
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_7_938 VPWR VGND sg13g2_decap_8
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_49_168 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_18_522 VPWR VGND sg13g2_decap_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_45_385 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_decap_8
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_28_319 VPWR VGND sg13g2_decap_8
XFILLER_37_875 VPWR VGND sg13g2_decap_8
XFILLER_36_385 VPWR VGND sg13g2_decap_8
XFILLER_24_536 VPWR VGND sg13g2_decap_8
XFILLER_20_753 VPWR VGND sg13g2_decap_8
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_1012 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_19_319 VPWR VGND sg13g2_decap_8
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_43_889 VPWR VGND sg13g2_decap_8
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_7_735 VPWR VGND sg13g2_decap_8
XFILLER_6_256 VPWR VGND sg13g2_decap_8
XFILLER_3_963 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_decap_8
XFILLER_34_812 VPWR VGND sg13g2_decap_8
XFILLER_19_886 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_33_322 VPWR VGND sg13g2_decap_8
XFILLER_18_396 VPWR VGND sg13g2_decap_8
XFILLER_34_889 VPWR VGND sg13g2_decap_8
XFILLER_33_399 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_116 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_44_609 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_37_672 VPWR VGND sg13g2_decap_8
XFILLER_25_823 VPWR VGND sg13g2_decap_8
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_24_333 VPWR VGND sg13g2_decap_8
XFILLER_40_826 VPWR VGND sg13g2_decap_8
XFILLER_20_550 VPWR VGND sg13g2_decap_8
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_48_959 VPWR VGND sg13g2_decap_8
Xheichips25_template VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_35_609 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_16_823 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_28_683 VPWR VGND sg13g2_decap_8
XFILLER_15_333 VPWR VGND sg13g2_decap_8
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_43_686 VPWR VGND sg13g2_decap_8
XFILLER_31_826 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_30_336 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_decap_8
XFILLER_7_532 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_39_959 VPWR VGND sg13g2_decap_8
XFILLER_38_469 VPWR VGND sg13g2_decap_8
XFILLER_19_683 VPWR VGND sg13g2_decap_8
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_34_686 VPWR VGND sg13g2_decap_8
XFILLER_33_196 VPWR VGND sg13g2_decap_8
XFILLER_22_837 VPWR VGND sg13g2_decap_8
XFILLER_21_347 VPWR VGND sg13g2_decap_8
XFILLER_5_1026 VPWR VGND sg13g2_fill_2
XFILLER_29_469 VPWR VGND sg13g2_decap_8
XFILLER_17_609 VPWR VGND sg13g2_decap_8
XFILLER_44_406 VPWR VGND sg13g2_decap_8
XFILLER_25_620 VPWR VGND sg13g2_decap_8
XFILLER_24_130 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_40_623 VPWR VGND sg13g2_decap_8
XFILLER_25_697 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_4_557 VPWR VGND sg13g2_decap_8
XFILLER_21_74 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_decap_8
XFILLER_16_620 VPWR VGND sg13g2_decap_8
XFILLER_28_480 VPWR VGND sg13g2_decap_8
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_44_973 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_31_623 VPWR VGND sg13g2_decap_8
XFILLER_30_133 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_830 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_39_756 VPWR VGND sg13g2_decap_8
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_26_417 VPWR VGND sg13g2_decap_8
XFILLER_19_480 VPWR VGND sg13g2_decap_8
XFILLER_35_973 VPWR VGND sg13g2_decap_8
XFILLER_34_483 VPWR VGND sg13g2_decap_8
XFILLER_22_634 VPWR VGND sg13g2_decap_8
XFILLER_21_144 VPWR VGND sg13g2_decap_8
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_17_406 VPWR VGND sg13g2_decap_8
XFILLER_44_203 VPWR VGND sg13g2_decap_8
XFILLER_29_266 VPWR VGND sg13g2_decap_8
XFILLER_41_910 VPWR VGND sg13g2_decap_8
XFILLER_26_984 VPWR VGND sg13g2_decap_8
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_16_74 VPWR VGND sg13g2_decap_8
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_25_494 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_decap_8
XFILLER_41_987 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_40_497 VPWR VGND sg13g2_decap_8
XFILLER_32_84 VPWR VGND sg13g2_decap_8
XFILLER_5_844 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_32_910 VPWR VGND sg13g2_decap_8
XFILLER_17_973 VPWR VGND sg13g2_decap_8
XFILLER_16_494 VPWR VGND sg13g2_decap_8
XFILLER_44_770 VPWR VGND sg13g2_decap_8
XFILLER_31_420 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
XFILLER_32_987 VPWR VGND sg13g2_decap_8
XFILLER_31_497 VPWR VGND sg13g2_decap_8
XFILLER_39_553 VPWR VGND sg13g2_decap_8
XFILLER_26_214 VPWR VGND sg13g2_decap_8
XFILLER_42_707 VPWR VGND sg13g2_decap_8
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_35_770 VPWR VGND sg13g2_decap_8
XFILLER_23_921 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_22_431 VPWR VGND sg13g2_decap_8
XFILLER_23_998 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_17_203 VPWR VGND sg13g2_decap_8
XFILLER_18_704 VPWR VGND sg13g2_decap_8
XFILLER_45_567 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_decap_8
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_14_921 VPWR VGND sg13g2_decap_8
XFILLER_32_217 VPWR VGND sg13g2_decap_8
XFILLER_26_781 VPWR VGND sg13g2_decap_8
XFILLER_13_431 VPWR VGND sg13g2_decap_8
XFILLER_25_291 VPWR VGND sg13g2_decap_8
XFILLER_14_998 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_41_784 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
Xheichips25_template_7 VPWR VGND uo_out[1] sg13g2_tielo
XFILLER_5_641 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_36_567 VPWR VGND sg13g2_decap_8
XFILLER_24_718 VPWR VGND sg13g2_decap_8
XFILLER_23_228 VPWR VGND sg13g2_decap_8
XFILLER_17_770 VPWR VGND sg13g2_decap_8
XFILLER_16_291 VPWR VGND sg13g2_decap_8
XFILLER_17_1015 VPWR VGND sg13g2_decap_8
XFILLER_32_784 VPWR VGND sg13g2_decap_8
XFILLER_20_935 VPWR VGND sg13g2_decap_8
XFILLER_31_294 VPWR VGND sg13g2_decap_8
XFILLER_9_991 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_15_718 VPWR VGND sg13g2_decap_8
XFILLER_42_504 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_decap_8
XFILLER_11_935 VPWR VGND sg13g2_decap_8
XFILLER_7_917 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_6_438 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_18_501 VPWR VGND sg13g2_decap_8
XFILLER_46_854 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_decap_8
XFILLER_18_578 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_14_795 VPWR VGND sg13g2_decap_8
XFILLER_9_221 VPWR VGND sg13g2_decap_8
XFILLER_41_581 VPWR VGND sg13g2_decap_8
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
XFILLER_37_854 VPWR VGND sg13g2_decap_8
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_24_515 VPWR VGND sg13g2_decap_8
XFILLER_32_581 VPWR VGND sg13g2_decap_8
XFILLER_20_732 VPWR VGND sg13g2_decap_8
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_865 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_decap_8
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_30_518 VPWR VGND sg13g2_decap_8
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_23_592 VPWR VGND sg13g2_decap_8
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_7_714 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_19_865 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_decap_8
XFILLER_18_375 VPWR VGND sg13g2_decap_8
XFILLER_34_868 VPWR VGND sg13g2_decap_8
XFILLER_33_378 VPWR VGND sg13g2_decap_8
XFILLER_14_592 VPWR VGND sg13g2_decap_8
XFILLER_21_529 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_37_651 VPWR VGND sg13g2_decap_8
XFILLER_25_802 VPWR VGND sg13g2_decap_8
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_24_312 VPWR VGND sg13g2_decap_8
XFILLER_40_805 VPWR VGND sg13g2_decap_8
XFILLER_25_879 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_8
XFILLER_24_389 VPWR VGND sg13g2_decap_8
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_249 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_938 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_16_802 VPWR VGND sg13g2_decap_8
XFILLER_28_662 VPWR VGND sg13g2_decap_8
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_decap_8
XFILLER_16_879 VPWR VGND sg13g2_decap_8
XFILLER_43_665 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_31_805 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_decap_8
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_30_315 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_decap_8
XFILLER_7_588 VPWR VGND sg13g2_decap_8
XFILLER_39_938 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_38_448 VPWR VGND sg13g2_decap_8
XFILLER_25_109 VPWR VGND sg13g2_decap_8
XFILLER_19_662 VPWR VGND sg13g2_decap_8
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_34_665 VPWR VGND sg13g2_decap_8
XFILLER_22_816 VPWR VGND sg13g2_decap_8
XFILLER_33_175 VPWR VGND sg13g2_decap_8
XFILLER_21_326 VPWR VGND sg13g2_decap_8
XFILLER_30_882 VPWR VGND sg13g2_decap_8
XFILLER_5_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_448 VPWR VGND sg13g2_decap_8
XFILLER_16_109 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_40_602 VPWR VGND sg13g2_decap_8
XFILLER_25_676 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_40_679 VPWR VGND sg13g2_decap_8
XFILLER_21_893 VPWR VGND sg13g2_decap_8
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_43_1022 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_44_952 VPWR VGND sg13g2_decap_8
XFILLER_16_676 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_31_602 VPWR VGND sg13g2_decap_8
XFILLER_15_186 VPWR VGND sg13g2_decap_8
XFILLER_30_112 VPWR VGND sg13g2_decap_8
XFILLER_31_679 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
XFILLER_30_189 VPWR VGND sg13g2_decap_8
XFILLER_8_886 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_7_385 VPWR VGND sg13g2_decap_8
XFILLER_39_735 VPWR VGND sg13g2_decap_8
XFILLER_38_245 VPWR VGND sg13g2_decap_8
XFILLER_35_952 VPWR VGND sg13g2_decap_8
XFILLER_34_462 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_8
XFILLER_21_123 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_29_245 VPWR VGND sg13g2_decap_8
XFILLER_45_749 VPWR VGND sg13g2_decap_8
XFILLER_16_53 VPWR VGND sg13g2_decap_8
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_26_963 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_25_473 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_41_966 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_40_476 VPWR VGND sg13g2_decap_8
XFILLER_32_63 VPWR VGND sg13g2_decap_8
XFILLER_21_690 VPWR VGND sg13g2_decap_8
XFILLER_5_823 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_36_749 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_17_952 VPWR VGND sg13g2_decap_8
XFILLER_16_473 VPWR VGND sg13g2_decap_8
XFILLER_32_966 VPWR VGND sg13g2_decap_8
XFILLER_31_476 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_decap_8
XFILLER_8_683 VPWR VGND sg13g2_decap_8
XFILLER_7_182 VPWR VGND sg13g2_decap_8
XFILLER_39_532 VPWR VGND sg13g2_decap_8
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_23_900 VPWR VGND sg13g2_decap_8
XFILLER_22_410 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_23_977 VPWR VGND sg13g2_decap_8
XFILLER_22_487 VPWR VGND sg13g2_decap_8
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_45_546 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_14_900 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_8
XFILLER_13_410 VPWR VGND sg13g2_decap_8
XFILLER_26_760 VPWR VGND sg13g2_decap_8
XFILLER_25_270 VPWR VGND sg13g2_decap_8
XFILLER_14_977 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_41_763 VPWR VGND sg13g2_decap_8
XFILLER_13_487 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
Xheichips25_template_8 VPWR VGND uo_out[2] sg13g2_tielo
XFILLER_5_620 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_5_697 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_49_896 VPWR VGND sg13g2_decap_8
XFILLER_36_546 VPWR VGND sg13g2_decap_8
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_16_270 VPWR VGND sg13g2_decap_8
XFILLER_32_763 VPWR VGND sg13g2_decap_8
XFILLER_20_914 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_decap_8
XFILLER_9_970 VPWR VGND sg13g2_decap_8
XFILLER_8_480 VPWR VGND sg13g2_decap_8
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_14_207 VPWR VGND sg13g2_decap_8
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_23_774 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_22_284 VPWR VGND sg13g2_decap_8
XFILLER_6_417 VPWR VGND sg13g2_decap_8
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_46_833 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_18_557 VPWR VGND sg13g2_decap_8
XFILLER_14_774 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
XFILLER_41_560 VPWR VGND sg13g2_decap_8
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_9_277 VPWR VGND sg13g2_decap_8
XFILLER_10_991 VPWR VGND sg13g2_decap_8
XFILLER_6_984 VPWR VGND sg13g2_decap_8
XFILLER_5_494 VPWR VGND sg13g2_decap_8
XFILLER_49_693 VPWR VGND sg13g2_decap_8
XFILLER_37_833 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_32_560 VPWR VGND sg13g2_decap_8
XFILLER_20_711 VPWR VGND sg13g2_decap_8
XFILLER_20_788 VPWR VGND sg13g2_decap_8
XFILLER_28_844 VPWR VGND sg13g2_decap_8
XFILLER_27_343 VPWR VGND sg13g2_decap_8
XFILLER_43_847 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_3_921 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_46_630 VPWR VGND sg13g2_decap_8
XFILLER_19_844 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_decap_8
XFILLER_34_847 VPWR VGND sg13g2_decap_8
XFILLER_33_357 VPWR VGND sg13g2_decap_8
XFILLER_21_508 VPWR VGND sg13g2_decap_8
XFILLER_14_571 VPWR VGND sg13g2_decap_8
XFILLER_14_1019 VPWR VGND sg13g2_decap_8
XFILLER_6_781 VPWR VGND sg13g2_decap_8
XFILLER_5_291 VPWR VGND sg13g2_decap_8
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_49_490 VPWR VGND sg13g2_decap_8
XFILLER_37_630 VPWR VGND sg13g2_decap_8
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_25_858 VPWR VGND sg13g2_decap_8
XFILLER_12_508 VPWR VGND sg13g2_decap_8
XFILLER_24_368 VPWR VGND sg13g2_decap_8
XFILLER_20_585 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_3_228 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_28_641 VPWR VGND sg13g2_decap_8
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_16_858 VPWR VGND sg13g2_decap_8
XFILLER_43_644 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_11_585 VPWR VGND sg13g2_decap_8
XFILLER_7_567 VPWR VGND sg13g2_decap_8
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_decap_8
XFILLER_39_917 VPWR VGND sg13g2_decap_8
XFILLER_38_427 VPWR VGND sg13g2_decap_8
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_19_641 VPWR VGND sg13g2_decap_8
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_18_151 VPWR VGND sg13g2_decap_8
XFILLER_34_644 VPWR VGND sg13g2_decap_8
XFILLER_33_154 VPWR VGND sg13g2_decap_8
XFILLER_21_305 VPWR VGND sg13g2_decap_8
XFILLER_30_861 VPWR VGND sg13g2_decap_8
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_427 VPWR VGND sg13g2_decap_8
XFILLER_38_994 VPWR VGND sg13g2_decap_8
XFILLER_25_655 VPWR VGND sg13g2_decap_8
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_decap_8
XFILLER_40_658 VPWR VGND sg13g2_decap_8
XFILLER_21_872 VPWR VGND sg13g2_decap_8
XFILLER_20_382 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_44_931 VPWR VGND sg13g2_decap_8
XFILLER_29_994 VPWR VGND sg13g2_decap_8
XFILLER_16_655 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_31_658 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
XFILLER_30_168 VPWR VGND sg13g2_decap_8
XFILLER_11_382 VPWR VGND sg13g2_decap_8
XFILLER_8_865 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_3_592 VPWR VGND sg13g2_decap_8
XFILLER_39_714 VPWR VGND sg13g2_decap_8
XFILLER_38_224 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_35_931 VPWR VGND sg13g2_decap_8
XFILLER_34_441 VPWR VGND sg13g2_decap_8
XFILLER_21_102 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_22_669 VPWR VGND sg13g2_decap_8
XFILLER_21_179 VPWR VGND sg13g2_decap_8
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_29_224 VPWR VGND sg13g2_decap_8
XFILLER_45_728 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_38_791 VPWR VGND sg13g2_decap_8
XFILLER_26_942 VPWR VGND sg13g2_decap_8
XFILLER_16_32 VPWR VGND sg13g2_decap_8
XFILLER_25_452 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_40_455 VPWR VGND sg13g2_decap_8
XFILLER_12_179 VPWR VGND sg13g2_decap_8
XFILLER_32_42 VPWR VGND sg13g2_decap_8
XFILLER_5_802 VPWR VGND sg13g2_decap_8
XFILLER_4_312 VPWR VGND sg13g2_decap_8
XFILLER_5_879 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_36_728 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_29_791 VPWR VGND sg13g2_decap_8
XFILLER_17_931 VPWR VGND sg13g2_decap_8
XFILLER_16_452 VPWR VGND sg13g2_decap_8
XFILLER_32_945 VPWR VGND sg13g2_decap_8
XFILLER_31_455 VPWR VGND sg13g2_decap_8
XFILLER_8_662 VPWR VGND sg13g2_decap_8
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_39_511 VPWR VGND sg13g2_decap_8
XFILLER_39_588 VPWR VGND sg13g2_decap_8
XFILLER_27_728 VPWR VGND sg13g2_decap_8
XFILLER_26_249 VPWR VGND sg13g2_decap_8
XFILLER_23_956 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_22_466 VPWR VGND sg13g2_decap_8
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_308 VPWR VGND sg13g2_decap_8
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_45_525 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_18_739 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_decap_8
XFILLER_14_956 VPWR VGND sg13g2_decap_8
XFILLER_41_742 VPWR VGND sg13g2_decap_8
XFILLER_13_466 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
Xheichips25_template_9 VPWR VGND uo_out[3] sg13g2_tielo
XFILLER_5_676 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_49_875 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_36_525 VPWR VGND sg13g2_decap_8
XFILLER_32_742 VPWR VGND sg13g2_decap_8
XFILLER_31_252 VPWR VGND sg13g2_decap_8
XFILLER_39_385 VPWR VGND sg13g2_decap_8
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_42_539 VPWR VGND sg13g2_decap_8
XFILLER_23_753 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_22_263 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_18_536 VPWR VGND sg13g2_decap_8
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_decap_8
XFILLER_14_753 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_9_256 VPWR VGND sg13g2_decap_8
XFILLER_10_970 VPWR VGND sg13g2_decap_8
XFILLER_6_963 VPWR VGND sg13g2_decap_8
XFILLER_5_473 VPWR VGND sg13g2_decap_8
XFILLER_49_672 VPWR VGND sg13g2_decap_8
XFILLER_37_812 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_36_399 VPWR VGND sg13g2_decap_8
XFILLER_20_767 VPWR VGND sg13g2_decap_8
XFILLER_8_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_28_823 VPWR VGND sg13g2_decap_8
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_27_322 VPWR VGND sg13g2_decap_8
XFILLER_43_826 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_27_399 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_23_550 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_7_749 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_38_609 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_19_823 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_decap_8
XFILLER_34_826 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
XFILLER_33_336 VPWR VGND sg13g2_decap_8
XFILLER_14_550 VPWR VGND sg13g2_decap_8
XFILLER_6_760 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_8
XFILLER_29_609 VPWR VGND sg13g2_decap_8
XFILLER_37_686 VPWR VGND sg13g2_decap_8
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_25_837 VPWR VGND sg13g2_decap_8
XFILLER_24_347 VPWR VGND sg13g2_decap_8
XFILLER_20_564 VPWR VGND sg13g2_decap_8
XFILLER_3_207 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_28_620 VPWR VGND sg13g2_decap_8
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_43_623 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_28_697 VPWR VGND sg13g2_decap_8
XFILLER_15_347 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_11_564 VPWR VGND sg13g2_decap_8
XFILLER_7_546 VPWR VGND sg13g2_decap_8
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_38_406 VPWR VGND sg13g2_decap_8
XFILLER_19_620 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_34_623 VPWR VGND sg13g2_decap_8
XFILLER_19_697 VPWR VGND sg13g2_decap_8
XFILLER_33_133 VPWR VGND sg13g2_decap_8
XFILLER_30_840 VPWR VGND sg13g2_decap_8
XFILLER_29_406 VPWR VGND sg13g2_decap_8
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_37_483 VPWR VGND sg13g2_decap_8
XFILLER_25_634 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_decap_8
XFILLER_40_637 VPWR VGND sg13g2_decap_8
XFILLER_21_851 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_20_361 VPWR VGND sg13g2_decap_8
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_29_973 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_44_910 VPWR VGND sg13g2_decap_8
XFILLER_28_494 VPWR VGND sg13g2_decap_8
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_44_987 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_31_637 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_30_147 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_8_844 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_decap_8
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_35_910 VPWR VGND sg13g2_decap_8
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_34_420 VPWR VGND sg13g2_decap_8
XFILLER_19_494 VPWR VGND sg13g2_decap_8
XFILLER_35_987 VPWR VGND sg13g2_decap_8
XFILLER_34_497 VPWR VGND sg13g2_decap_8
XFILLER_22_648 VPWR VGND sg13g2_decap_8
XFILLER_21_158 VPWR VGND sg13g2_decap_8
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_203 VPWR VGND sg13g2_decap_8
XFILLER_45_707 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_44_217 VPWR VGND sg13g2_decap_8
XFILLER_38_770 VPWR VGND sg13g2_decap_8
XFILLER_26_921 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_25_431 VPWR VGND sg13g2_decap_8
XFILLER_41_924 VPWR VGND sg13g2_decap_8
XFILLER_26_998 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_16_88 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_32_21 VPWR VGND sg13g2_decap_8
XFILLER_32_98 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_5_858 VPWR VGND sg13g2_decap_8
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_36_707 VPWR VGND sg13g2_decap_8
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_29_770 VPWR VGND sg13g2_decap_8
XFILLER_17_910 VPWR VGND sg13g2_decap_8
XFILLER_16_431 VPWR VGND sg13g2_decap_8
XFILLER_28_291 VPWR VGND sg13g2_decap_8
XFILLER_44_784 VPWR VGND sg13g2_decap_8
XFILLER_32_924 VPWR VGND sg13g2_decap_8
XFILLER_17_987 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_31_434 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_8_641 VPWR VGND sg13g2_decap_8
XFILLER_39_567 VPWR VGND sg13g2_decap_8
XFILLER_27_707 VPWR VGND sg13g2_decap_8
XFILLER_26_228 VPWR VGND sg13g2_decap_8
XFILLER_19_291 VPWR VGND sg13g2_decap_8
XFILLER_35_784 VPWR VGND sg13g2_decap_8
XFILLER_34_294 VPWR VGND sg13g2_decap_8
XFILLER_23_935 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
XFILLER_22_445 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_decap_8
XFILLER_17_217 VPWR VGND sg13g2_decap_8
XFILLER_45_504 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
XFILLER_14_935 VPWR VGND sg13g2_decap_8
XFILLER_41_721 VPWR VGND sg13g2_decap_8
XFILLER_26_795 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_41_798 VPWR VGND sg13g2_decap_8
XFILLER_5_655 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_36_504 VPWR VGND sg13g2_decap_8
XFILLER_44_581 VPWR VGND sg13g2_decap_8
XFILLER_32_721 VPWR VGND sg13g2_decap_8
XFILLER_17_784 VPWR VGND sg13g2_decap_8
XFILLER_31_231 VPWR VGND sg13g2_decap_8
XFILLER_32_798 VPWR VGND sg13g2_decap_8
XFILLER_20_949 VPWR VGND sg13g2_decap_8
XFILLER_39_364 VPWR VGND sg13g2_decap_8
XFILLER_27_504 VPWR VGND sg13g2_decap_8
XFILLER_42_518 VPWR VGND sg13g2_decap_8
XFILLER_35_581 VPWR VGND sg13g2_decap_8
XFILLER_23_732 VPWR VGND sg13g2_decap_8
XFILLER_22_242 VPWR VGND sg13g2_decap_8
XFILLER_11_949 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_18_515 VPWR VGND sg13g2_decap_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_33_518 VPWR VGND sg13g2_decap_8
XFILLER_14_732 VPWR VGND sg13g2_decap_8
XFILLER_26_592 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_41_595 VPWR VGND sg13g2_decap_8
XFILLER_6_942 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
XFILLER_49_651 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_24_529 VPWR VGND sg13g2_decap_8
XFILLER_17_581 VPWR VGND sg13g2_decap_8
XFILLER_32_595 VPWR VGND sg13g2_decap_8
XFILLER_20_746 VPWR VGND sg13g2_decap_8
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_161 VPWR VGND sg13g2_decap_8
XFILLER_28_802 VPWR VGND sg13g2_decap_8
XFILLER_27_301 VPWR VGND sg13g2_decap_8
XFILLER_43_805 VPWR VGND sg13g2_decap_8
XFILLER_28_879 VPWR VGND sg13g2_decap_8
XFILLER_27_378 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_7_728 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_3_956 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_19_802 VPWR VGND sg13g2_decap_8
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_34_805 VPWR VGND sg13g2_decap_8
XFILLER_19_879 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_33_315 VPWR VGND sg13g2_decap_8
XFILLER_18_389 VPWR VGND sg13g2_decap_8
XFILLER_42_882 VPWR VGND sg13g2_decap_8
XFILLER_41_392 VPWR VGND sg13g2_decap_8
XFILLER_28_109 VPWR VGND sg13g2_decap_8
XFILLER_37_665 VPWR VGND sg13g2_decap_8
XFILLER_25_816 VPWR VGND sg13g2_decap_8
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_24_326 VPWR VGND sg13g2_decap_8
XFILLER_40_819 VPWR VGND sg13g2_decap_8
XFILLER_33_882 VPWR VGND sg13g2_decap_8
XFILLER_32_392 VPWR VGND sg13g2_decap_8
XFILLER_20_543 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_16_816 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_28_676 VPWR VGND sg13g2_decap_8
XFILLER_15_326 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_43_679 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_31_819 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_30_329 VPWR VGND sg13g2_decap_8
XFILLER_24_893 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_7_525 VPWR VGND sg13g2_decap_8
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_19_676 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_34_602 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_33_112 VPWR VGND sg13g2_decap_8
XFILLER_34_679 VPWR VGND sg13g2_decap_8
XFILLER_15_893 VPWR VGND sg13g2_decap_8
XFILLER_33_189 VPWR VGND sg13g2_decap_8
XFILLER_30_896 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
XFILLER_5_1019 VPWR VGND sg13g2_decap_8
XFILLER_38_952 VPWR VGND sg13g2_decap_8
XFILLER_37_462 VPWR VGND sg13g2_decap_8
XFILLER_25_613 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_decap_8
XFILLER_40_616 VPWR VGND sg13g2_decap_8
XFILLER_21_830 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_decap_8
XFILLER_28_473 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_44_966 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_31_616 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_8
XFILLER_30_126 VPWR VGND sg13g2_decap_8
XFILLER_24_690 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_decap_8
XFILLER_8_823 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_399 VPWR VGND sg13g2_decap_8
XFILLER_3_550 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_39_749 VPWR VGND sg13g2_decap_8
XFILLER_38_259 VPWR VGND sg13g2_decap_8
XFILLER_19_473 VPWR VGND sg13g2_decap_8
XFILLER_35_966 VPWR VGND sg13g2_decap_8
XFILLER_34_476 VPWR VGND sg13g2_decap_8
XFILLER_15_690 VPWR VGND sg13g2_decap_8
XFILLER_22_627 VPWR VGND sg13g2_decap_8
XFILLER_21_137 VPWR VGND sg13g2_decap_8
XFILLER_30_693 VPWR VGND sg13g2_decap_8
XFILLER_29_259 VPWR VGND sg13g2_decap_8
XFILLER_26_900 VPWR VGND sg13g2_decap_8
XFILLER_25_410 VPWR VGND sg13g2_decap_8
XFILLER_16_67 VPWR VGND sg13g2_decap_8
XFILLER_41_903 VPWR VGND sg13g2_decap_8
XFILLER_26_977 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_40_413 VPWR VGND sg13g2_decap_8
XFILLER_25_487 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_32_77 VPWR VGND sg13g2_decap_8
XFILLER_5_837 VPWR VGND sg13g2_decap_8
XFILLER_4_347 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_16_410 VPWR VGND sg13g2_decap_8
XFILLER_28_270 VPWR VGND sg13g2_decap_8
XFILLER_17_966 VPWR VGND sg13g2_decap_8
XFILLER_44_763 VPWR VGND sg13g2_decap_8
XFILLER_32_903 VPWR VGND sg13g2_decap_8
XFILLER_16_487 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_31_413 VPWR VGND sg13g2_decap_8
XFILLER_8_620 VPWR VGND sg13g2_decap_8
XFILLER_40_980 VPWR VGND sg13g2_decap_8
XFILLER_8_697 VPWR VGND sg13g2_decap_8
XFILLER_7_196 VPWR VGND sg13g2_decap_8
XFILLER_39_546 VPWR VGND sg13g2_decap_8
XFILLER_26_207 VPWR VGND sg13g2_decap_8
XFILLER_19_270 VPWR VGND sg13g2_decap_8
XFILLER_35_763 VPWR VGND sg13g2_decap_8
XFILLER_23_914 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_22_424 VPWR VGND sg13g2_decap_8
XFILLER_31_980 VPWR VGND sg13g2_decap_8
XFILLER_30_490 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_14_914 VPWR VGND sg13g2_decap_8
XFILLER_41_700 VPWR VGND sg13g2_decap_8
XFILLER_26_774 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_25_284 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_41_777 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_22_991 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
XFILLER_44_560 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_decap_8
XFILLER_17_763 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_decap_8
XFILLER_17_1008 VPWR VGND sg13g2_decap_8
XFILLER_32_777 VPWR VGND sg13g2_decap_8
XFILLER_20_928 VPWR VGND sg13g2_decap_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_31_287 VPWR VGND sg13g2_decap_8
XFILLER_9_984 VPWR VGND sg13g2_decap_8
XFILLER_8_494 VPWR VGND sg13g2_decap_8
XFILLER_39_343 VPWR VGND sg13g2_decap_8
XFILLER_35_560 VPWR VGND sg13g2_decap_8
XFILLER_23_711 VPWR VGND sg13g2_decap_8
XFILLER_22_221 VPWR VGND sg13g2_decap_8
XFILLER_11_928 VPWR VGND sg13g2_decap_8
XFILLER_23_788 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_22_298 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_46_847 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_14_711 VPWR VGND sg13g2_decap_8
XFILLER_26_571 VPWR VGND sg13g2_decap_8
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_14_788 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_41_574 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_5_431 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_49_630 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_37_847 VPWR VGND sg13g2_decap_8
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_24_508 VPWR VGND sg13g2_decap_8
XFILLER_17_560 VPWR VGND sg13g2_decap_8
XFILLER_32_574 VPWR VGND sg13g2_decap_8
XFILLER_20_725 VPWR VGND sg13g2_decap_8
XFILLER_9_781 VPWR VGND sg13g2_decap_8
XFILLER_8_291 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_140 VPWR VGND sg13g2_decap_8
XFILLER_28_858 VPWR VGND sg13g2_decap_8
XFILLER_15_508 VPWR VGND sg13g2_decap_8
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_7_707 VPWR VGND sg13g2_decap_8
XFILLER_23_585 VPWR VGND sg13g2_decap_8
XFILLER_10_235 VPWR VGND sg13g2_decap_8
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_3_935 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_858 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_18_368 VPWR VGND sg13g2_decap_8
XFILLER_42_861 VPWR VGND sg13g2_decap_8
XFILLER_14_585 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_decap_8
XFILLER_6_795 VPWR VGND sg13g2_decap_8
XFILLER_37_644 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_24_305 VPWR VGND sg13g2_decap_8
XFILLER_33_861 VPWR VGND sg13g2_decap_8
XFILLER_32_371 VPWR VGND sg13g2_decap_8
XFILLER_20_522 VPWR VGND sg13g2_decap_8
XFILLER_20_599 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_28_655 VPWR VGND sg13g2_decap_8
XFILLER_15_305 VPWR VGND sg13g2_decap_8
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_43_658 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_30_308 VPWR VGND sg13g2_decap_8
XFILLER_24_872 VPWR VGND sg13g2_decap_8
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_23_382 VPWR VGND sg13g2_decap_8
XFILLER_7_504 VPWR VGND sg13g2_decap_8
XFILLER_11_599 VPWR VGND sg13g2_decap_8
XFILLER_3_732 VPWR VGND sg13g2_decap_8
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_655 VPWR VGND sg13g2_decap_8
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_34_658 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_decap_8
XFILLER_33_168 VPWR VGND sg13g2_decap_8
XFILLER_21_319 VPWR VGND sg13g2_decap_8
XFILLER_14_382 VPWR VGND sg13g2_decap_8
XFILLER_30_875 VPWR VGND sg13g2_decap_8
XFILLER_6_592 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_38_931 VPWR VGND sg13g2_decap_8
XFILLER_37_441 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_25_669 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
XFILLER_24_179 VPWR VGND sg13g2_decap_8
XFILLER_21_886 VPWR VGND sg13g2_decap_8
XFILLER_21_46 VPWR VGND sg13g2_decap_8
XFILLER_20_396 VPWR VGND sg13g2_decap_8
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_43_1015 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_29_931 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_28_452 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_44_945 VPWR VGND sg13g2_decap_8
XFILLER_16_669 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_15_179 VPWR VGND sg13g2_decap_8
XFILLER_30_105 VPWR VGND sg13g2_decap_8
XFILLER_8_802 VPWR VGND sg13g2_decap_8
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_decap_8
XFILLER_11_396 VPWR VGND sg13g2_decap_8
XFILLER_8_879 VPWR VGND sg13g2_decap_8
XFILLER_7_378 VPWR VGND sg13g2_decap_8
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_39_728 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
XFILLER_19_452 VPWR VGND sg13g2_decap_8
XFILLER_35_945 VPWR VGND sg13g2_decap_8
XFILLER_34_455 VPWR VGND sg13g2_decap_8
XFILLER_22_606 VPWR VGND sg13g2_decap_8
XFILLER_21_116 VPWR VGND sg13g2_decap_8
XFILLER_30_672 VPWR VGND sg13g2_decap_8
XFILLER_29_238 VPWR VGND sg13g2_decap_8
XFILLER_26_956 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_16_46 VPWR VGND sg13g2_decap_8
XFILLER_25_466 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_41_959 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_32_56 VPWR VGND sg13g2_decap_8
XFILLER_21_683 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_5_816 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_44_742 VPWR VGND sg13g2_decap_8
XFILLER_17_945 VPWR VGND sg13g2_decap_8
XFILLER_16_466 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_32_959 VPWR VGND sg13g2_decap_8
XFILLER_31_469 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_decap_8
XFILLER_11_193 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_8_676 VPWR VGND sg13g2_decap_8
XFILLER_4_893 VPWR VGND sg13g2_decap_8
XFILLER_39_525 VPWR VGND sg13g2_decap_8
XFILLER_35_742 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
XFILLER_22_403 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_45_539 VPWR VGND sg13g2_decap_8
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_26_753 VPWR VGND sg13g2_decap_8
XFILLER_13_403 VPWR VGND sg13g2_decap_8
XFILLER_25_263 VPWR VGND sg13g2_decap_8
XFILLER_41_756 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_22_970 VPWR VGND sg13g2_decap_8
XFILLER_21_480 VPWR VGND sg13g2_decap_8
XFILLER_5_613 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_49_812 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_36_539 VPWR VGND sg13g2_decap_8
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_742 VPWR VGND sg13g2_decap_8
XFILLER_16_263 VPWR VGND sg13g2_decap_8
XFILLER_32_756 VPWR VGND sg13g2_decap_8
XFILLER_20_907 VPWR VGND sg13g2_decap_8
XFILLER_13_970 VPWR VGND sg13g2_decap_8
XFILLER_31_266 VPWR VGND sg13g2_decap_8
XFILLER_12_480 VPWR VGND sg13g2_decap_8
XFILLER_9_963 VPWR VGND sg13g2_decap_8
XFILLER_8_473 VPWR VGND sg13g2_decap_8
XFILLER_4_690 VPWR VGND sg13g2_decap_8
XFILLER_39_322 VPWR VGND sg13g2_decap_8
XFILLER_39_399 VPWR VGND sg13g2_decap_8
XFILLER_27_539 VPWR VGND sg13g2_decap_8
XFILLER_22_200 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_23_767 VPWR VGND sg13g2_decap_8
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_22_277 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_49_119 VPWR VGND sg13g2_decap_8
XFILLER_46_826 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_26_550 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_14_767 VPWR VGND sg13g2_decap_8
XFILLER_41_553 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_37_826 VPWR VGND sg13g2_decap_8
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_32_553 VPWR VGND sg13g2_decap_8
XFILLER_20_704 VPWR VGND sg13g2_decap_8
XFILLER_9_760 VPWR VGND sg13g2_decap_8
XFILLER_8_270 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_28_837 VPWR VGND sg13g2_decap_8
XFILLER_39_196 VPWR VGND sg13g2_decap_8
XFILLER_27_336 VPWR VGND sg13g2_decap_8
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_23_564 VPWR VGND sg13g2_decap_8
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_46_623 VPWR VGND sg13g2_decap_8
XFILLER_19_837 VPWR VGND sg13g2_decap_8
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_18_347 VPWR VGND sg13g2_decap_8
XFILLER_42_840 VPWR VGND sg13g2_decap_8
XFILLER_14_564 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_6_774 VPWR VGND sg13g2_decap_8
XFILLER_5_284 VPWR VGND sg13g2_decap_8
XFILLER_2_991 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_49_483 VPWR VGND sg13g2_decap_8
XFILLER_37_623 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_33_840 VPWR VGND sg13g2_decap_8
XFILLER_32_350 VPWR VGND sg13g2_decap_8
XFILLER_20_501 VPWR VGND sg13g2_decap_8
XFILLER_20_578 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_28_634 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_decap_8
XFILLER_43_637 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_23_361 VPWR VGND sg13g2_decap_8
XFILLER_11_578 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_711 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
XFILLER_19_634 VPWR VGND sg13g2_decap_8
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
XFILLER_34_637 VPWR VGND sg13g2_decap_8
XFILLER_15_851 VPWR VGND sg13g2_decap_8
XFILLER_33_147 VPWR VGND sg13g2_decap_8
XFILLER_14_361 VPWR VGND sg13g2_decap_8
XFILLER_30_854 VPWR VGND sg13g2_decap_8
XFILLER_6_571 VPWR VGND sg13g2_decap_8
XFILLER_38_910 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_49_280 VPWR VGND sg13g2_decap_8
XFILLER_37_420 VPWR VGND sg13g2_decap_8
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_37_497 VPWR VGND sg13g2_decap_8
XFILLER_25_648 VPWR VGND sg13g2_decap_8
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
XFILLER_24_158 VPWR VGND sg13g2_decap_8
XFILLER_21_865 VPWR VGND sg13g2_decap_8
XFILLER_20_375 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_4_508 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_29_910 VPWR VGND sg13g2_decap_8
XFILLER_28_431 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_44_924 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_decap_8
XFILLER_16_648 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_8_858 VPWR VGND sg13g2_decap_8
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_39_707 VPWR VGND sg13g2_decap_8
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_19_431 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_35_924 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_434 VPWR VGND sg13g2_decap_8
XFILLER_30_651 VPWR VGND sg13g2_decap_8
XFILLER_29_217 VPWR VGND sg13g2_decap_8
XFILLER_38_784 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_26_935 VPWR VGND sg13g2_decap_8
XFILLER_25_445 VPWR VGND sg13g2_decap_8
XFILLER_41_938 VPWR VGND sg13g2_decap_8
XFILLER_40_448 VPWR VGND sg13g2_decap_8
XFILLER_32_35 VPWR VGND sg13g2_decap_8
XFILLER_21_662 VPWR VGND sg13g2_decap_8
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_44_721 VPWR VGND sg13g2_decap_8
XFILLER_29_784 VPWR VGND sg13g2_decap_8
XFILLER_17_924 VPWR VGND sg13g2_decap_8
XFILLER_16_445 VPWR VGND sg13g2_decap_8
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_44_798 VPWR VGND sg13g2_decap_8
XFILLER_32_938 VPWR VGND sg13g2_decap_8
XFILLER_31_448 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_decap_8
XFILLER_8_655 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
XFILLER_4_872 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_35_721 VPWR VGND sg13g2_decap_8
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_35_798 VPWR VGND sg13g2_decap_8
XFILLER_23_949 VPWR VGND sg13g2_decap_8
XFILLER_22_459 VPWR VGND sg13g2_decap_8
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_2_809 VPWR VGND sg13g2_decap_8
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
XFILLER_45_518 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_38_581 VPWR VGND sg13g2_decap_8
XFILLER_26_732 VPWR VGND sg13g2_decap_8
XFILLER_25_242 VPWR VGND sg13g2_decap_8
XFILLER_14_949 VPWR VGND sg13g2_decap_8
XFILLER_13_459 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_49_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_669 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_49_868 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_36_518 VPWR VGND sg13g2_decap_8
XFILLER_29_581 VPWR VGND sg13g2_decap_8
XFILLER_17_721 VPWR VGND sg13g2_decap_8
XFILLER_16_242 VPWR VGND sg13g2_decap_8
XFILLER_17_798 VPWR VGND sg13g2_decap_8
XFILLER_44_595 VPWR VGND sg13g2_decap_8
XFILLER_32_735 VPWR VGND sg13g2_decap_8
XFILLER_31_245 VPWR VGND sg13g2_decap_8
XFILLER_9_942 VPWR VGND sg13g2_decap_8
XFILLER_8_452 VPWR VGND sg13g2_decap_8
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_27_518 VPWR VGND sg13g2_decap_8
XFILLER_39_378 VPWR VGND sg13g2_decap_8
XFILLER_35_595 VPWR VGND sg13g2_decap_8
XFILLER_23_746 VPWR VGND sg13g2_decap_8
XFILLER_22_256 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_46_805 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_18_529 VPWR VGND sg13g2_decap_8
XFILLER_14_746 VPWR VGND sg13g2_decap_8
XFILLER_41_532 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_49_665 VPWR VGND sg13g2_decap_8
XFILLER_37_805 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_45_882 VPWR VGND sg13g2_decap_8
XFILLER_44_392 VPWR VGND sg13g2_decap_8
XFILLER_32_532 VPWR VGND sg13g2_decap_8
XFILLER_17_595 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
XFILLER_8_1019 VPWR VGND sg13g2_decap_8
XFILLER_28_816 VPWR VGND sg13g2_decap_8
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_27_315 VPWR VGND sg13g2_decap_8
XFILLER_43_819 VPWR VGND sg13g2_decap_8
XFILLER_36_882 VPWR VGND sg13g2_decap_8
XFILLER_42_329 VPWR VGND sg13g2_decap_8
XFILLER_35_392 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_23_543 VPWR VGND sg13g2_decap_8
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_19_816 VPWR VGND sg13g2_decap_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_46_679 VPWR VGND sg13g2_decap_8
XFILLER_34_819 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_33_329 VPWR VGND sg13g2_decap_8
XFILLER_14_543 VPWR VGND sg13g2_decap_8
XFILLER_42_896 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_6_753 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
XFILLER_49_462 VPWR VGND sg13g2_decap_8
XFILLER_37_602 VPWR VGND sg13g2_decap_8
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_37_679 VPWR VGND sg13g2_decap_8
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_18_893 VPWR VGND sg13g2_decap_8
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_33_896 VPWR VGND sg13g2_decap_8
XFILLER_20_557 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_613 VPWR VGND sg13g2_decap_8
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_24_830 VPWR VGND sg13g2_decap_8
XFILLER_23_340 VPWR VGND sg13g2_decap_8
XFILLER_11_557 VPWR VGND sg13g2_decap_8
XFILLER_7_539 VPWR VGND sg13g2_decap_8
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_19_613 VPWR VGND sg13g2_decap_8
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_34_616 VPWR VGND sg13g2_decap_8
XFILLER_15_830 VPWR VGND sg13g2_decap_8
XFILLER_33_126 VPWR VGND sg13g2_decap_8
XFILLER_14_340 VPWR VGND sg13g2_decap_8
XFILLER_42_693 VPWR VGND sg13g2_decap_8
XFILLER_30_833 VPWR VGND sg13g2_decap_8
XFILLER_6_550 VPWR VGND sg13g2_decap_8
XFILLER_38_966 VPWR VGND sg13g2_decap_8
XFILLER_37_476 VPWR VGND sg13g2_decap_8
XFILLER_25_627 VPWR VGND sg13g2_decap_8
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_24_137 VPWR VGND sg13g2_decap_8
XFILLER_33_693 VPWR VGND sg13g2_decap_8
XFILLER_21_844 VPWR VGND sg13g2_decap_8
XFILLER_20_354 VPWR VGND sg13g2_decap_8
XFILLER_29_966 VPWR VGND sg13g2_decap_8
XFILLER_28_410 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_44_903 VPWR VGND sg13g2_decap_8
XFILLER_16_627 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_28_487 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_8_837 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_3_564 VPWR VGND sg13g2_decap_8
XFILLER_19_410 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_35_903 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_34_413 VPWR VGND sg13g2_decap_8
XFILLER_19_487 VPWR VGND sg13g2_decap_8
XFILLER_43_980 VPWR VGND sg13g2_decap_8
XFILLER_42_490 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_38_763 VPWR VGND sg13g2_decap_8
XFILLER_26_914 VPWR VGND sg13g2_decap_8
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_25_424 VPWR VGND sg13g2_decap_8
XFILLER_41_917 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_decap_8
XFILLER_34_980 VPWR VGND sg13g2_decap_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
XFILLER_32_14 VPWR VGND sg13g2_decap_8
XFILLER_21_641 VPWR VGND sg13g2_decap_8
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_44_700 VPWR VGND sg13g2_decap_8
XFILLER_29_763 VPWR VGND sg13g2_decap_8
XFILLER_17_903 VPWR VGND sg13g2_decap_8
XFILLER_16_424 VPWR VGND sg13g2_decap_8
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_44_777 VPWR VGND sg13g2_decap_8
XFILLER_32_917 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_31_427 VPWR VGND sg13g2_decap_8
XFILLER_25_991 VPWR VGND sg13g2_decap_8
XFILLER_12_641 VPWR VGND sg13g2_decap_8
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_8_634 VPWR VGND sg13g2_decap_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_4_851 VPWR VGND sg13g2_decap_8
XFILLER_3_361 VPWR VGND sg13g2_decap_8
XFILLER_26_1012 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_35_700 VPWR VGND sg13g2_decap_8
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_35_777 VPWR VGND sg13g2_decap_8
XFILLER_23_928 VPWR VGND sg13g2_decap_8
XFILLER_16_991 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_8
XFILLER_22_438 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_31_994 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_38_560 VPWR VGND sg13g2_decap_8
XFILLER_26_711 VPWR VGND sg13g2_decap_8
XFILLER_25_221 VPWR VGND sg13g2_decap_8
XFILLER_14_928 VPWR VGND sg13g2_decap_8
XFILLER_41_714 VPWR VGND sg13g2_decap_8
XFILLER_26_788 VPWR VGND sg13g2_decap_8
XFILLER_13_438 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_25_298 VPWR VGND sg13g2_decap_8
XFILLER_5_648 VPWR VGND sg13g2_decap_8
XFILLER_49_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_29_560 VPWR VGND sg13g2_decap_8
XFILLER_17_700 VPWR VGND sg13g2_decap_8
XFILLER_16_221 VPWR VGND sg13g2_decap_8
XFILLER_44_574 VPWR VGND sg13g2_decap_8
XFILLER_32_714 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_17_777 VPWR VGND sg13g2_decap_8
XFILLER_16_298 VPWR VGND sg13g2_decap_8
XFILLER_31_224 VPWR VGND sg13g2_decap_8
XFILLER_9_921 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_decap_8
XFILLER_40_791 VPWR VGND sg13g2_decap_8
XFILLER_9_998 VPWR VGND sg13g2_decap_8
XFILLER_39_357 VPWR VGND sg13g2_decap_8
XFILLER_35_574 VPWR VGND sg13g2_decap_8
XFILLER_23_725 VPWR VGND sg13g2_decap_8
XFILLER_22_235 VPWR VGND sg13g2_decap_8
XFILLER_31_791 VPWR VGND sg13g2_decap_8
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_18_508 VPWR VGND sg13g2_decap_8
XFILLER_14_725 VPWR VGND sg13g2_decap_8
XFILLER_41_511 VPWR VGND sg13g2_decap_8
XFILLER_26_585 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_41_588 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_644 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_45_861 VPWR VGND sg13g2_decap_8
XFILLER_17_574 VPWR VGND sg13g2_decap_8
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_32_511 VPWR VGND sg13g2_decap_8
XFILLER_32_588 VPWR VGND sg13g2_decap_8
XFILLER_20_739 VPWR VGND sg13g2_decap_8
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
XFILLER_9_795 VPWR VGND sg13g2_decap_8
XFILLER_39_154 VPWR VGND sg13g2_decap_8
XFILLER_42_308 VPWR VGND sg13g2_decap_8
XFILLER_36_861 VPWR VGND sg13g2_decap_8
XFILLER_39_1022 VPWR VGND sg13g2_decap_8
XFILLER_35_371 VPWR VGND sg13g2_decap_8
XFILLER_23_522 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_23_599 VPWR VGND sg13g2_decap_8
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_949 VPWR VGND sg13g2_decap_8
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_33_308 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_14_522 VPWR VGND sg13g2_decap_8
XFILLER_26_382 VPWR VGND sg13g2_decap_8
XFILLER_42_875 VPWR VGND sg13g2_decap_8
XFILLER_14_599 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_14_81 VPWR VGND sg13g2_decap_8
XFILLER_6_732 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_30_91 VPWR VGND sg13g2_decap_8
XFILLER_49_441 VPWR VGND sg13g2_decap_8
XFILLER_37_658 VPWR VGND sg13g2_decap_8
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_25_809 VPWR VGND sg13g2_decap_8
XFILLER_18_872 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_decap_8
XFILLER_24_319 VPWR VGND sg13g2_decap_8
XFILLER_33_875 VPWR VGND sg13g2_decap_8
XFILLER_32_385 VPWR VGND sg13g2_decap_8
XFILLER_20_536 VPWR VGND sg13g2_decap_8
XFILLER_9_592 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_16_809 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_28_669 VPWR VGND sg13g2_decap_8
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_15_319 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_24_886 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_23_396 VPWR VGND sg13g2_decap_8
XFILLER_7_518 VPWR VGND sg13g2_decap_8
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_19_669 VPWR VGND sg13g2_decap_8
XFILLER_33_105 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_decap_8
XFILLER_15_886 VPWR VGND sg13g2_decap_8
XFILLER_42_672 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_decap_8
XFILLER_14_396 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
XFILLER_30_889 VPWR VGND sg13g2_decap_8
XFILLER_38_945 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_37_455 VPWR VGND sg13g2_decap_8
XFILLER_25_606 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_40_609 VPWR VGND sg13g2_decap_8
XFILLER_33_672 VPWR VGND sg13g2_decap_8
XFILLER_21_823 VPWR VGND sg13g2_decap_8
XFILLER_32_182 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_29_945 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_28_466 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_44_959 VPWR VGND sg13g2_decap_8
XFILLER_31_609 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_8
XFILLER_12_823 VPWR VGND sg13g2_decap_8
XFILLER_24_683 VPWR VGND sg13g2_decap_8
XFILLER_11_333 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_8_816 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_543 VPWR VGND sg13g2_decap_8
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_19_466 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_35_959 VPWR VGND sg13g2_decap_8
XFILLER_34_469 VPWR VGND sg13g2_decap_8
XFILLER_15_683 VPWR VGND sg13g2_decap_8
XFILLER_14_193 VPWR VGND sg13g2_decap_8
XFILLER_30_686 VPWR VGND sg13g2_decap_8
XFILLER_7_882 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_38_742 VPWR VGND sg13g2_decap_8
XFILLER_37_252 VPWR VGND sg13g2_decap_8
XFILLER_25_403 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_8
XFILLER_21_620 VPWR VGND sg13g2_decap_8
XFILLER_20_130 VPWR VGND sg13g2_decap_8
XFILLER_21_697 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_29_742 VPWR VGND sg13g2_decap_8
XFILLER_16_403 VPWR VGND sg13g2_decap_8
XFILLER_28_263 VPWR VGND sg13g2_decap_8
XFILLER_44_756 VPWR VGND sg13g2_decap_8
XFILLER_17_959 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_31_406 VPWR VGND sg13g2_decap_8
XFILLER_25_970 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_8
XFILLER_24_480 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_8_613 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_3_340 VPWR VGND sg13g2_decap_8
XFILLER_39_539 VPWR VGND sg13g2_decap_8
XFILLER_19_263 VPWR VGND sg13g2_decap_8
XFILLER_35_756 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_decap_8
XFILLER_16_970 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_22_417 VPWR VGND sg13g2_decap_8
XFILLER_15_480 VPWR VGND sg13g2_decap_8
XFILLER_31_973 VPWR VGND sg13g2_decap_8
XFILLER_30_483 VPWR VGND sg13g2_decap_8
XFILLER_25_200 VPWR VGND sg13g2_decap_8
XFILLER_14_907 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_26_767 VPWR VGND sg13g2_decap_8
XFILLER_13_417 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_25_277 VPWR VGND sg13g2_decap_8
XFILLER_22_984 VPWR VGND sg13g2_decap_8
XFILLER_21_494 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_16_200 VPWR VGND sg13g2_decap_8
XFILLER_17_756 VPWR VGND sg13g2_decap_8
XFILLER_44_553 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_16_277 VPWR VGND sg13g2_decap_8
XFILLER_31_203 VPWR VGND sg13g2_decap_8
XFILLER_9_900 VPWR VGND sg13g2_decap_8
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_40_770 VPWR VGND sg13g2_decap_8
XFILLER_12_494 VPWR VGND sg13g2_decap_8
XFILLER_9_977 VPWR VGND sg13g2_decap_8
XFILLER_33_91 VPWR VGND sg13g2_decap_8
XFILLER_8_487 VPWR VGND sg13g2_decap_8
XFILLER_39_336 VPWR VGND sg13g2_decap_8
XFILLER_35_553 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_31_770 VPWR VGND sg13g2_decap_8
XFILLER_30_280 VPWR VGND sg13g2_decap_8
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_14_704 VPWR VGND sg13g2_decap_8
XFILLER_26_564 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_41_567 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
XFILLER_22_781 VPWR VGND sg13g2_decap_8
XFILLER_21_291 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_45_840 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_17_553 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_decap_8
XFILLER_20_718 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
XFILLER_9_774 VPWR VGND sg13g2_decap_8
XFILLER_8_284 VPWR VGND sg13g2_decap_8
XFILLER_5_991 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
XFILLER_39_133 VPWR VGND sg13g2_decap_8
XFILLER_36_840 VPWR VGND sg13g2_decap_8
XFILLER_39_1001 VPWR VGND sg13g2_decap_8
XFILLER_35_350 VPWR VGND sg13g2_decap_8
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_11_718 VPWR VGND sg13g2_decap_8
XFILLER_23_578 VPWR VGND sg13g2_decap_8
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_3_928 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_46_637 VPWR VGND sg13g2_decap_8
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_14_501 VPWR VGND sg13g2_decap_8
XFILLER_26_361 VPWR VGND sg13g2_decap_8
XFILLER_42_854 VPWR VGND sg13g2_decap_8
XFILLER_14_578 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_14_60 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_6_788 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_30_70 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_420 VPWR VGND sg13g2_decap_8
XFILLER_49_497 VPWR VGND sg13g2_decap_8
XFILLER_37_637 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_18_851 VPWR VGND sg13g2_decap_8
XFILLER_17_350 VPWR VGND sg13g2_decap_8
XFILLER_33_854 VPWR VGND sg13g2_decap_8
XFILLER_32_364 VPWR VGND sg13g2_decap_8
XFILLER_20_515 VPWR VGND sg13g2_decap_8
XFILLER_9_571 VPWR VGND sg13g2_decap_8
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_28_648 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_decap_8
XFILLER_24_865 VPWR VGND sg13g2_decap_8
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_23_375 VPWR VGND sg13g2_decap_8
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_725 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_648 VPWR VGND sg13g2_decap_8
XFILLER_18_158 VPWR VGND sg13g2_decap_8
XFILLER_15_865 VPWR VGND sg13g2_decap_8
XFILLER_42_651 VPWR VGND sg13g2_decap_8
XFILLER_25_81 VPWR VGND sg13g2_decap_8
XFILLER_14_375 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_30_868 VPWR VGND sg13g2_decap_8
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_585 VPWR VGND sg13g2_decap_8
XFILLER_29_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_924 VPWR VGND sg13g2_decap_8
XFILLER_37_434 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
XFILLER_33_651 VPWR VGND sg13g2_decap_8
XFILLER_21_802 VPWR VGND sg13g2_decap_8
XFILLER_32_161 VPWR VGND sg13g2_decap_8
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XFILLER_21_879 VPWR VGND sg13g2_decap_8
XFILLER_20_389 VPWR VGND sg13g2_decap_8
XFILLER_21_39 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_43_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_924 VPWR VGND sg13g2_decap_8
XFILLER_28_445 VPWR VGND sg13g2_decap_8
XFILLER_44_938 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_12_802 VPWR VGND sg13g2_decap_8
XFILLER_24_662 VPWR VGND sg13g2_decap_8
XFILLER_11_312 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_12_879 VPWR VGND sg13g2_decap_8
XFILLER_11_389 VPWR VGND sg13g2_decap_8
XFILLER_3_522 VPWR VGND sg13g2_decap_8
XFILLER_3_599 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_19_445 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_35_938 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_34_448 VPWR VGND sg13g2_decap_8
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_21_109 VPWR VGND sg13g2_decap_8
XFILLER_14_172 VPWR VGND sg13g2_decap_8
XFILLER_30_665 VPWR VGND sg13g2_decap_8
XFILLER_7_861 VPWR VGND sg13g2_decap_8
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_38_721 VPWR VGND sg13g2_decap_8
XFILLER_37_231 VPWR VGND sg13g2_decap_8
XFILLER_38_798 VPWR VGND sg13g2_decap_8
XFILLER_16_39 VPWR VGND sg13g2_decap_8
XFILLER_26_949 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
XFILLER_25_459 VPWR VGND sg13g2_decap_8
XFILLER_32_49 VPWR VGND sg13g2_decap_8
XFILLER_21_676 VPWR VGND sg13g2_decap_8
XFILLER_5_809 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_29_721 VPWR VGND sg13g2_decap_8
XFILLER_29_798 VPWR VGND sg13g2_decap_8
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_17_938 VPWR VGND sg13g2_decap_8
XFILLER_44_735 VPWR VGND sg13g2_decap_8
XFILLER_16_459 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_40_952 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_8
XFILLER_11_186 VPWR VGND sg13g2_decap_8
XFILLER_8_669 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_decap_8
XFILLER_39_518 VPWR VGND sg13g2_decap_8
XFILLER_19_242 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_31_952 VPWR VGND sg13g2_decap_8
XFILLER_30_462 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_27_49 VPWR VGND sg13g2_decap_8
XFILLER_38_595 VPWR VGND sg13g2_decap_8
XFILLER_26_746 VPWR VGND sg13g2_decap_8
XFILLER_25_256 VPWR VGND sg13g2_decap_8
XFILLER_41_749 VPWR VGND sg13g2_decap_8
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_22_963 VPWR VGND sg13g2_decap_8
XFILLER_21_473 VPWR VGND sg13g2_decap_8
XFILLER_5_606 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_44_532 VPWR VGND sg13g2_decap_8
XFILLER_29_595 VPWR VGND sg13g2_decap_8
XFILLER_17_735 VPWR VGND sg13g2_decap_8
XFILLER_16_256 VPWR VGND sg13g2_decap_8
XFILLER_32_749 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_31_259 VPWR VGND sg13g2_decap_8
XFILLER_12_473 VPWR VGND sg13g2_decap_8
XFILLER_33_70 VPWR VGND sg13g2_decap_8
XFILLER_9_956 VPWR VGND sg13g2_decap_8
XFILLER_8_466 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
XFILLER_3_193 VPWR VGND sg13g2_decap_8
XFILLER_39_315 VPWR VGND sg13g2_decap_8
XFILLER_48_882 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_35_532 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_46_819 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_39_882 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_26_543 VPWR VGND sg13g2_decap_8
XFILLER_41_546 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_22_760 VPWR VGND sg13g2_decap_8
XFILLER_21_270 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_37_819 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_29_392 VPWR VGND sg13g2_decap_8
XFILLER_17_532 VPWR VGND sg13g2_decap_8
XFILLER_45_896 VPWR VGND sg13g2_decap_8
XFILLER_32_546 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_12_270 VPWR VGND sg13g2_decap_8
XFILLER_9_753 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
XFILLER_5_970 VPWR VGND sg13g2_decap_8
XFILLER_4_480 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_27_329 VPWR VGND sg13g2_decap_8
XFILLER_36_896 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_23_557 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_3_907 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_616 VPWR VGND sg13g2_decap_8
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_26_340 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_14_557 VPWR VGND sg13g2_decap_8
XFILLER_42_833 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_6_767 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_7_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_37_616 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
XFILLER_45_693 VPWR VGND sg13g2_decap_8
XFILLER_33_833 VPWR VGND sg13g2_decap_8
XFILLER_32_343 VPWR VGND sg13g2_decap_8
XFILLER_9_550 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_28_627 VPWR VGND sg13g2_decap_8
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
XFILLER_36_693 VPWR VGND sg13g2_decap_8
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_23_354 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_704 VPWR VGND sg13g2_decap_8
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_19_627 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_15_844 VPWR VGND sg13g2_decap_8
XFILLER_42_630 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_14_354 VPWR VGND sg13g2_decap_8
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
XFILLER_30_847 VPWR VGND sg13g2_decap_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_564 VPWR VGND sg13g2_decap_8
XFILLER_29_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
XFILLER_38_903 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_49_273 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_decap_8
XFILLER_46_980 VPWR VGND sg13g2_decap_8
XFILLER_45_490 VPWR VGND sg13g2_decap_8
XFILLER_33_630 VPWR VGND sg13g2_decap_8
XFILLER_32_140 VPWR VGND sg13g2_decap_8
XFILLER_21_858 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_20_368 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_29_903 VPWR VGND sg13g2_decap_8
XFILLER_28_424 VPWR VGND sg13g2_decap_8
XFILLER_44_917 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_36_490 VPWR VGND sg13g2_decap_8
XFILLER_24_641 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_decap_8
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_3_501 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_8
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_19_424 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_35_917 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_34_427 VPWR VGND sg13g2_decap_8
XFILLER_28_991 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_15_641 VPWR VGND sg13g2_decap_8
XFILLER_14_151 VPWR VGND sg13g2_decap_8
XFILLER_43_994 VPWR VGND sg13g2_decap_8
XFILLER_30_644 VPWR VGND sg13g2_decap_8
XFILLER_7_840 VPWR VGND sg13g2_decap_8
XFILLER_6_361 VPWR VGND sg13g2_decap_8
XFILLER_38_700 VPWR VGND sg13g2_decap_8
XFILLER_37_210 VPWR VGND sg13g2_decap_8
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_26_928 VPWR VGND sg13g2_decap_8
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_25_438 VPWR VGND sg13g2_decap_8
XFILLER_19_991 VPWR VGND sg13g2_decap_8
XFILLER_34_994 VPWR VGND sg13g2_decap_8
XFILLER_32_28 VPWR VGND sg13g2_decap_8
XFILLER_21_655 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_700 VPWR VGND sg13g2_decap_8
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_44_714 VPWR VGND sg13g2_decap_8
XFILLER_29_777 VPWR VGND sg13g2_decap_8
XFILLER_17_917 VPWR VGND sg13g2_decap_8
XFILLER_16_438 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_8_648 VPWR VGND sg13g2_decap_8
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_26_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_221 VPWR VGND sg13g2_decap_8
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_35_714 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_43_791 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
XFILLER_31_931 VPWR VGND sg13g2_decap_8
XFILLER_30_441 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_38_574 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_26_725 VPWR VGND sg13g2_decap_8
XFILLER_25_235 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_34_791 VPWR VGND sg13g2_decap_8
XFILLER_22_942 VPWR VGND sg13g2_decap_8
XFILLER_21_452 VPWR VGND sg13g2_decap_8
XFILLER_49_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_17_714 VPWR VGND sg13g2_decap_8
XFILLER_44_511 VPWR VGND sg13g2_decap_8
XFILLER_29_574 VPWR VGND sg13g2_decap_8
XFILLER_16_235 VPWR VGND sg13g2_decap_8
XFILLER_44_588 VPWR VGND sg13g2_decap_8
XFILLER_32_728 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_decap_8
XFILLER_9_935 VPWR VGND sg13g2_decap_8
XFILLER_8_445 VPWR VGND sg13g2_decap_8
XFILLER_4_662 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_48_861 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_35_511 VPWR VGND sg13g2_decap_8
XFILLER_35_588 VPWR VGND sg13g2_decap_8
XFILLER_23_739 VPWR VGND sg13g2_decap_8
XFILLER_22_249 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_39_861 VPWR VGND sg13g2_decap_8
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_26_522 VPWR VGND sg13g2_decap_8
XFILLER_14_739 VPWR VGND sg13g2_decap_8
XFILLER_41_525 VPWR VGND sg13g2_decap_8
XFILLER_26_599 VPWR VGND sg13g2_decap_8
XFILLER_13_249 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_49_658 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_17_511 VPWR VGND sg13g2_decap_8
XFILLER_29_371 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_45_875 VPWR VGND sg13g2_decap_8
XFILLER_17_588 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_8
XFILLER_8_242 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_39_168 VPWR VGND sg13g2_decap_8
XFILLER_28_809 VPWR VGND sg13g2_decap_8
XFILLER_27_308 VPWR VGND sg13g2_decap_8
XFILLER_36_875 VPWR VGND sg13g2_decap_8
XFILLER_35_385 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
XFILLER_19_809 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_42_812 VPWR VGND sg13g2_decap_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_14_536 VPWR VGND sg13g2_decap_8
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_26_396 VPWR VGND sg13g2_decap_8
XFILLER_42_889 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_14_95 VPWR VGND sg13g2_decap_8
XFILLER_6_746 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_7_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_49_455 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_decap_8
XFILLER_33_812 VPWR VGND sg13g2_decap_8
XFILLER_18_886 VPWR VGND sg13g2_decap_8
XFILLER_17_385 VPWR VGND sg13g2_decap_8
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_32_322 VPWR VGND sg13g2_decap_8
XFILLER_33_889 VPWR VGND sg13g2_decap_8
XFILLER_32_399 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_28_606 VPWR VGND sg13g2_decap_8
XFILLER_27_105 VPWR VGND sg13g2_decap_8
XFILLER_43_609 VPWR VGND sg13g2_decap_8
XFILLER_36_672 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_23_333 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_606 VPWR VGND sg13g2_decap_8
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_34_609 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_15_823 VPWR VGND sg13g2_decap_8
XFILLER_33_119 VPWR VGND sg13g2_decap_8
XFILLER_14_333 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_decap_8
XFILLER_42_686 VPWR VGND sg13g2_decap_8
XFILLER_30_826 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_543 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_37_469 VPWR VGND sg13g2_decap_8
XFILLER_17_182 VPWR VGND sg13g2_decap_8
XFILLER_18_683 VPWR VGND sg13g2_decap_8
XFILLER_33_686 VPWR VGND sg13g2_decap_8
XFILLER_21_837 VPWR VGND sg13g2_decap_8
XFILLER_32_196 VPWR VGND sg13g2_decap_8
XFILLER_20_347 VPWR VGND sg13g2_decap_8
XFILLER_28_403 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_29_959 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_24_620 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_decap_8
XFILLER_24_697 VPWR VGND sg13g2_decap_8
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_7_329 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_557 VPWR VGND sg13g2_decap_8
XFILLER_19_403 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_4_1026 VPWR VGND sg13g2_fill_2
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_34_406 VPWR VGND sg13g2_decap_8
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_decap_8
XFILLER_15_697 VPWR VGND sg13g2_decap_8
XFILLER_30_623 VPWR VGND sg13g2_decap_8
XFILLER_42_483 VPWR VGND sg13g2_decap_8
XFILLER_6_340 VPWR VGND sg13g2_decap_8
XFILLER_7_896 VPWR VGND sg13g2_decap_8
XFILLER_38_756 VPWR VGND sg13g2_decap_8
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_26_907 VPWR VGND sg13g2_decap_8
XFILLER_19_970 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_decap_8
XFILLER_18_480 VPWR VGND sg13g2_decap_8
XFILLER_34_973 VPWR VGND sg13g2_decap_8
XFILLER_33_483 VPWR VGND sg13g2_decap_8
XFILLER_21_634 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_29_756 VPWR VGND sg13g2_decap_8
XFILLER_28_200 VPWR VGND sg13g2_decap_8
XFILLER_16_417 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_28_277 VPWR VGND sg13g2_decap_8
XFILLER_40_910 VPWR VGND sg13g2_decap_8
XFILLER_25_984 VPWR VGND sg13g2_decap_8
XFILLER_19_1012 VPWR VGND sg13g2_decap_8
XFILLER_12_634 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_decap_8
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_8_627 VPWR VGND sg13g2_decap_8
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_354 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1005 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_34_203 VPWR VGND sg13g2_decap_8
XFILLER_19_277 VPWR VGND sg13g2_decap_8
XFILLER_16_984 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_8
XFILLER_31_910 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_42_280 VPWR VGND sg13g2_decap_8
XFILLER_30_420 VPWR VGND sg13g2_decap_8
XFILLER_31_987 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_30_497 VPWR VGND sg13g2_decap_8
XFILLER_7_693 VPWR VGND sg13g2_decap_8
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_38_553 VPWR VGND sg13g2_decap_8
XFILLER_26_704 VPWR VGND sg13g2_decap_8
XFILLER_25_214 VPWR VGND sg13g2_decap_8
XFILLER_41_707 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_34_770 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_decap_8
XFILLER_33_280 VPWR VGND sg13g2_decap_8
XFILLER_21_431 VPWR VGND sg13g2_decap_8
XFILLER_22_998 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_29_553 VPWR VGND sg13g2_decap_8
XFILLER_16_214 VPWR VGND sg13g2_decap_8
XFILLER_32_707 VPWR VGND sg13g2_decap_8
XFILLER_44_567 VPWR VGND sg13g2_decap_8
XFILLER_31_217 VPWR VGND sg13g2_decap_8
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_25_781 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_decap_8
XFILLER_9_914 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_decap_8
XFILLER_40_784 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_35_567 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_8
XFILLER_16_781 VPWR VGND sg13g2_decap_8
XFILLER_22_228 VPWR VGND sg13g2_decap_8
XFILLER_15_291 VPWR VGND sg13g2_decap_8
XFILLER_31_784 VPWR VGND sg13g2_decap_8
XFILLER_30_294 VPWR VGND sg13g2_decap_8
XFILLER_8_991 VPWR VGND sg13g2_decap_8
XFILLER_7_490 VPWR VGND sg13g2_decap_8
XFILLER_38_28 VPWR VGND sg13g2_decap_8
XFILLER_39_840 VPWR VGND sg13g2_decap_8
XFILLER_38_350 VPWR VGND sg13g2_decap_8
XFILLER_26_501 VPWR VGND sg13g2_decap_8
XFILLER_14_718 VPWR VGND sg13g2_decap_8
XFILLER_41_504 VPWR VGND sg13g2_decap_8
XFILLER_26_578 VPWR VGND sg13g2_decap_8
XFILLER_13_228 VPWR VGND sg13g2_decap_8
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_22_795 VPWR VGND sg13g2_decap_8
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_decap_8
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_637 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_29_350 VPWR VGND sg13g2_decap_8
XFILLER_45_854 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_32_504 VPWR VGND sg13g2_decap_8
XFILLER_17_567 VPWR VGND sg13g2_decap_8
XFILLER_9_711 VPWR VGND sg13g2_decap_8
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
XFILLER_40_581 VPWR VGND sg13g2_decap_8
XFILLER_9_788 VPWR VGND sg13g2_decap_8
XFILLER_8_298 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_39_147 VPWR VGND sg13g2_decap_8
XFILLER_36_854 VPWR VGND sg13g2_decap_8
XFILLER_39_1015 VPWR VGND sg13g2_decap_8
XFILLER_35_364 VPWR VGND sg13g2_decap_8
XFILLER_23_515 VPWR VGND sg13g2_decap_8
XFILLER_31_581 VPWR VGND sg13g2_decap_8
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_14_515 VPWR VGND sg13g2_decap_8
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_26_375 VPWR VGND sg13g2_decap_8
XFILLER_42_868 VPWR VGND sg13g2_decap_8
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_14_74 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_decap_8
XFILLER_6_725 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_8
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_49_434 VPWR VGND sg13g2_decap_8
XFILLER_17_364 VPWR VGND sg13g2_decap_8
XFILLER_45_651 VPWR VGND sg13g2_decap_8
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_44_161 VPWR VGND sg13g2_decap_8
XFILLER_32_301 VPWR VGND sg13g2_decap_8
XFILLER_33_868 VPWR VGND sg13g2_decap_8
XFILLER_32_378 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_decap_8
XFILLER_13_592 VPWR VGND sg13g2_decap_8
XFILLER_9_585 VPWR VGND sg13g2_decap_8
XFILLER_36_651 VPWR VGND sg13g2_decap_8
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_24_879 VPWR VGND sg13g2_decap_8
XFILLER_11_529 VPWR VGND sg13g2_decap_8
XFILLER_23_389 VPWR VGND sg13g2_decap_8
XFILLER_3_739 VPWR VGND sg13g2_decap_8
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_15_802 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_14_312 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_42_665 VPWR VGND sg13g2_decap_8
XFILLER_30_805 VPWR VGND sg13g2_decap_8
XFILLER_14_389 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_decap_8
XFILLER_6_522 VPWR VGND sg13g2_decap_8
XFILLER_6_599 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_38_938 VPWR VGND sg13g2_decap_8
XFILLER_37_448 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_decap_8
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XFILLER_33_665 VPWR VGND sg13g2_decap_8
XFILLER_21_816 VPWR VGND sg13g2_decap_8
XFILLER_32_175 VPWR VGND sg13g2_decap_8
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XFILLER_9_382 VPWR VGND sg13g2_decap_8
XFILLER_29_938 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_28_459 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_24_676 VPWR VGND sg13g2_decap_8
XFILLER_11_326 VPWR VGND sg13g2_decap_8
XFILLER_8_809 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_20_893 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_19_459 VPWR VGND sg13g2_decap_8
XFILLER_43_952 VPWR VGND sg13g2_decap_8
XFILLER_15_676 VPWR VGND sg13g2_decap_8
XFILLER_42_462 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_14_186 VPWR VGND sg13g2_decap_8
XFILLER_30_679 VPWR VGND sg13g2_decap_8
XFILLER_11_893 VPWR VGND sg13g2_decap_8
XFILLER_7_875 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_decap_8
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_735 VPWR VGND sg13g2_decap_8
XFILLER_37_245 VPWR VGND sg13g2_decap_8
XFILLER_34_952 VPWR VGND sg13g2_decap_8
XFILLER_33_462 VPWR VGND sg13g2_decap_8
XFILLER_21_613 VPWR VGND sg13g2_decap_8
XFILLER_20_123 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_29_735 VPWR VGND sg13g2_decap_8
XFILLER_28_256 VPWR VGND sg13g2_decap_8
XFILLER_44_749 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_decap_8
XFILLER_25_963 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_24_473 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_8_606 VPWR VGND sg13g2_decap_8
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_19_256 VPWR VGND sg13g2_decap_8
XFILLER_35_749 VPWR VGND sg13g2_decap_8
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_31_966 VPWR VGND sg13g2_decap_8
XFILLER_30_476 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
XFILLER_7_672 VPWR VGND sg13g2_decap_8
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_38_532 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_21_410 VPWR VGND sg13g2_decap_8
XFILLER_22_977 VPWR VGND sg13g2_decap_8
XFILLER_21_487 VPWR VGND sg13g2_decap_8
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_29_532 VPWR VGND sg13g2_decap_8
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_44_546 VPWR VGND sg13g2_decap_8
XFILLER_17_749 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_25_760 VPWR VGND sg13g2_decap_8
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_24_270 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_40_763 VPWR VGND sg13g2_decap_8
XFILLER_12_487 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_decap_8
XFILLER_4_620 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_39_329 VPWR VGND sg13g2_decap_8
XFILLER_48_896 VPWR VGND sg13g2_decap_8
XFILLER_35_546 VPWR VGND sg13g2_decap_8
XFILLER_16_760 VPWR VGND sg13g2_decap_8
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_15_270 VPWR VGND sg13g2_decap_8
XFILLER_31_763 VPWR VGND sg13g2_decap_8
XFILLER_30_273 VPWR VGND sg13g2_decap_8
XFILLER_8_970 VPWR VGND sg13g2_decap_8
XFILLER_39_896 VPWR VGND sg13g2_decap_8
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_26_557 VPWR VGND sg13g2_decap_8
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_21_284 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_45_833 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_17_546 VPWR VGND sg13g2_decap_8
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_40_560 VPWR VGND sg13g2_decap_8
XFILLER_12_284 VPWR VGND sg13g2_decap_8
XFILLER_9_767 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_984 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_36_833 VPWR VGND sg13g2_decap_8
XFILLER_35_343 VPWR VGND sg13g2_decap_8
XFILLER_31_560 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_39_693 VPWR VGND sg13g2_decap_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_decap_8
XFILLER_42_847 VPWR VGND sg13g2_decap_8
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_53 VPWR VGND sg13g2_decap_8
XFILLER_22_571 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_49_413 VPWR VGND sg13g2_decap_8
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_45_630 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_17_343 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_33_847 VPWR VGND sg13g2_decap_8
XFILLER_32_357 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_decap_8
XFILLER_20_508 VPWR VGND sg13g2_decap_8
XFILLER_9_564 VPWR VGND sg13g2_decap_8
XFILLER_5_781 VPWR VGND sg13g2_decap_8
XFILLER_4_291 VPWR VGND sg13g2_decap_8
XFILLER_49_980 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_36_630 VPWR VGND sg13g2_decap_8
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_8
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_718 VPWR VGND sg13g2_decap_8
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_39_490 VPWR VGND sg13g2_decap_8
XFILLER_26_151 VPWR VGND sg13g2_decap_8
XFILLER_15_858 VPWR VGND sg13g2_decap_8
XFILLER_42_644 VPWR VGND sg13g2_decap_8
XFILLER_14_368 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_25_74 VPWR VGND sg13g2_decap_8
XFILLER_6_501 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_decap_8
XFILLER_29_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_38_917 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_49_287 VPWR VGND sg13g2_decap_8
XFILLER_37_427 VPWR VGND sg13g2_decap_8
XFILLER_18_641 VPWR VGND sg13g2_decap_8
XFILLER_17_140 VPWR VGND sg13g2_decap_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
XFILLER_33_644 VPWR VGND sg13g2_decap_8
XFILLER_32_154 VPWR VGND sg13g2_decap_8
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XFILLER_9_361 VPWR VGND sg13g2_decap_8
XFILLER_29_917 VPWR VGND sg13g2_decap_8
XFILLER_28_438 VPWR VGND sg13g2_decap_8
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_24_655 VPWR VGND sg13g2_decap_8
XFILLER_11_305 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_20_872 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_decap_8
XFILLER_3_515 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_438 VPWR VGND sg13g2_decap_8
XFILLER_43_931 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_decap_8
XFILLER_42_441 VPWR VGND sg13g2_decap_8
XFILLER_14_165 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_decap_8
XFILLER_11_872 VPWR VGND sg13g2_decap_8
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_7_854 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_38_714 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_34_931 VPWR VGND sg13g2_decap_8
XFILLER_33_441 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_8
XFILLER_21_669 VPWR VGND sg13g2_decap_8
XFILLER_20_179 VPWR VGND sg13g2_decap_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_29_714 VPWR VGND sg13g2_decap_8
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_44_728 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_37_791 VPWR VGND sg13g2_decap_8
XFILLER_25_942 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_11_102 VPWR VGND sg13g2_decap_8
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_3_389 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_19_235 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_35_728 VPWR VGND sg13g2_decap_8
XFILLER_16_942 VPWR VGND sg13g2_decap_8
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_8
XFILLER_31_945 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_30_455 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
XFILLER_7_651 VPWR VGND sg13g2_decap_8
XFILLER_6_172 VPWR VGND sg13g2_decap_8
XFILLER_38_511 VPWR VGND sg13g2_decap_8
XFILLER_38_588 VPWR VGND sg13g2_decap_8
XFILLER_26_739 VPWR VGND sg13g2_decap_8
XFILLER_25_249 VPWR VGND sg13g2_decap_8
XFILLER_22_956 VPWR VGND sg13g2_decap_8
XFILLER_21_466 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_29_511 VPWR VGND sg13g2_decap_8
XFILLER_29_588 VPWR VGND sg13g2_decap_8
XFILLER_17_728 VPWR VGND sg13g2_decap_8
XFILLER_17_42 VPWR VGND sg13g2_decap_8
XFILLER_44_525 VPWR VGND sg13g2_decap_8
XFILLER_16_249 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_40_742 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_decap_8
XFILLER_9_949 VPWR VGND sg13g2_decap_8
XFILLER_33_63 VPWR VGND sg13g2_decap_8
XFILLER_32_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_459 VPWR VGND sg13g2_decap_8
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_35_525 VPWR VGND sg13g2_decap_8
XFILLER_31_742 VPWR VGND sg13g2_decap_8
XFILLER_30_252 VPWR VGND sg13g2_decap_8
XFILLER_39_875 VPWR VGND sg13g2_decap_8
XFILLER_38_385 VPWR VGND sg13g2_decap_8
XFILLER_26_536 VPWR VGND sg13g2_decap_8
XFILLER_41_539 VPWR VGND sg13g2_decap_8
XFILLER_22_753 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_263 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_45_812 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_29_385 VPWR VGND sg13g2_decap_8
XFILLER_17_525 VPWR VGND sg13g2_decap_8
XFILLER_45_889 VPWR VGND sg13g2_decap_8
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_32_539 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_12_263 VPWR VGND sg13g2_decap_8
XFILLER_9_746 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_8
XFILLER_5_963 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_36_812 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_36_889 VPWR VGND sg13g2_decap_8
XFILLER_35_399 VPWR VGND sg13g2_decap_8
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_39_672 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
XFILLER_42_826 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_30_42 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_7_1015 VPWR VGND sg13g2_decap_8
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_49_469 VPWR VGND sg13g2_decap_8
XFILLER_37_609 VPWR VGND sg13g2_decap_8
XFILLER_17_322 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_29_182 VPWR VGND sg13g2_decap_8
XFILLER_45_686 VPWR VGND sg13g2_decap_8
XFILLER_33_826 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
XFILLER_32_336 VPWR VGND sg13g2_decap_8
XFILLER_13_550 VPWR VGND sg13g2_decap_8
XFILLER_9_543 VPWR VGND sg13g2_decap_8
XFILLER_5_760 VPWR VGND sg13g2_decap_8
XFILLER_4_270 VPWR VGND sg13g2_decap_8
XFILLER_27_119 VPWR VGND sg13g2_decap_8
XFILLER_36_686 VPWR VGND sg13g2_decap_8
XFILLER_24_837 VPWR VGND sg13g2_decap_8
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_23_347 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_26_130 VPWR VGND sg13g2_decap_8
XFILLER_15_837 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_14_347 VPWR VGND sg13g2_decap_8
XFILLER_42_623 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_6_557 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_49_266 VPWR VGND sg13g2_decap_8
XFILLER_37_406 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_18_620 VPWR VGND sg13g2_decap_8
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_17_196 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_decap_8
XFILLER_33_623 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_decap_8
XFILLER_32_133 VPWR VGND sg13g2_decap_8
XFILLER_9_340 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_28_417 VPWR VGND sg13g2_decap_8
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_36_483 VPWR VGND sg13g2_decap_8
XFILLER_24_634 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_20_851 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_19_417 VPWR VGND sg13g2_decap_8
XFILLER_43_910 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_15_634 VPWR VGND sg13g2_decap_8
XFILLER_42_420 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_43_987 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_decap_8
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_7_833 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_46_770 VPWR VGND sg13g2_decap_8
XFILLER_34_910 VPWR VGND sg13g2_decap_8
XFILLER_19_984 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_33_420 VPWR VGND sg13g2_decap_8
XFILLER_18_494 VPWR VGND sg13g2_decap_8
XFILLER_34_987 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_decap_8
XFILLER_21_648 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_8
XFILLER_28_214 VPWR VGND sg13g2_decap_8
XFILLER_44_707 VPWR VGND sg13g2_decap_8
XFILLER_37_770 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_25_921 VPWR VGND sg13g2_decap_8
XFILLER_24_431 VPWR VGND sg13g2_decap_8
XFILLER_19_1026 VPWR VGND sg13g2_fill_2
XFILLER_40_924 VPWR VGND sg13g2_decap_8
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_12_648 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_26_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_214 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_35_707 VPWR VGND sg13g2_decap_8
XFILLER_16_921 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_28_781 VPWR VGND sg13g2_decap_8
XFILLER_27_280 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_16_998 VPWR VGND sg13g2_decap_8
XFILLER_43_784 VPWR VGND sg13g2_decap_8
XFILLER_31_924 VPWR VGND sg13g2_decap_8
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_30_434 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_7_630 VPWR VGND sg13g2_decap_8
XFILLER_6_151 VPWR VGND sg13g2_decap_8
XFILLER_38_567 VPWR VGND sg13g2_decap_8
XFILLER_26_718 VPWR VGND sg13g2_decap_8
XFILLER_25_228 VPWR VGND sg13g2_decap_8
XFILLER_19_781 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
XFILLER_34_784 VPWR VGND sg13g2_decap_8
XFILLER_22_935 VPWR VGND sg13g2_decap_8
XFILLER_33_294 VPWR VGND sg13g2_decap_8
XFILLER_21_445 VPWR VGND sg13g2_decap_8
XFILLER_49_1008 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_decap_8
XFILLER_44_504 VPWR VGND sg13g2_decap_8
XFILLER_29_567 VPWR VGND sg13g2_decap_8
XFILLER_17_707 VPWR VGND sg13g2_decap_8
XFILLER_16_228 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_40_721 VPWR VGND sg13g2_decap_8
XFILLER_25_795 VPWR VGND sg13g2_decap_8
XFILLER_12_445 VPWR VGND sg13g2_decap_8
XFILLER_33_42 VPWR VGND sg13g2_decap_8
XFILLER_9_928 VPWR VGND sg13g2_decap_8
XFILLER_32_1001 VPWR VGND sg13g2_decap_8
XFILLER_8_438 VPWR VGND sg13g2_decap_8
XFILLER_40_798 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_35_504 VPWR VGND sg13g2_decap_8
XFILLER_16_795 VPWR VGND sg13g2_decap_8
XFILLER_31_721 VPWR VGND sg13g2_decap_8
XFILLER_43_581 VPWR VGND sg13g2_decap_8
XFILLER_30_231 VPWR VGND sg13g2_decap_8
XFILLER_31_798 VPWR VGND sg13g2_decap_8
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_38_364 VPWR VGND sg13g2_decap_8
XFILLER_26_515 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_decap_8
XFILLER_34_581 VPWR VGND sg13g2_decap_8
XFILLER_22_732 VPWR VGND sg13g2_decap_8
XFILLER_21_242 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_17_504 VPWR VGND sg13g2_decap_8
XFILLER_29_364 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_45_868 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
XFILLER_32_518 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_25_592 VPWR VGND sg13g2_decap_8
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
XFILLER_40_595 VPWR VGND sg13g2_decap_8
XFILLER_5_942 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_36_868 VPWR VGND sg13g2_decap_8
XFILLER_35_378 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_decap_8
XFILLER_16_592 VPWR VGND sg13g2_decap_8
XFILLER_31_595 VPWR VGND sg13g2_decap_8
XFILLER_39_651 VPWR VGND sg13g2_decap_8
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_decap_8
XFILLER_42_805 VPWR VGND sg13g2_decap_8
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_14_529 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
XFILLER_26_389 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_14_88 VPWR VGND sg13g2_decap_8
XFILLER_6_739 VPWR VGND sg13g2_decap_8
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_30_98 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_decap_8
XFILLER_17_301 VPWR VGND sg13g2_decap_8
XFILLER_29_161 VPWR VGND sg13g2_decap_8
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_17_378 VPWR VGND sg13g2_decap_8
XFILLER_45_665 VPWR VGND sg13g2_decap_8
XFILLER_33_805 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_32_315 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_41_882 VPWR VGND sg13g2_decap_8
XFILLER_40_392 VPWR VGND sg13g2_decap_8
XFILLER_9_599 VPWR VGND sg13g2_decap_8
XFILLER_45_1022 VPWR VGND sg13g2_decap_8
XFILLER_36_665 VPWR VGND sg13g2_decap_8
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_23_326 VPWR VGND sg13g2_decap_8
XFILLER_32_882 VPWR VGND sg13g2_decap_8
XFILLER_31_392 VPWR VGND sg13g2_decap_8
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_15_816 VPWR VGND sg13g2_decap_8
XFILLER_42_602 VPWR VGND sg13g2_decap_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_14_326 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_42_679 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_23_893 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_536 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_245 VPWR VGND sg13g2_decap_8
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_33_602 VPWR VGND sg13g2_decap_8
XFILLER_18_676 VPWR VGND sg13g2_decap_8
XFILLER_17_175 VPWR VGND sg13g2_decap_8
XFILLER_32_112 VPWR VGND sg13g2_decap_8
XFILLER_33_679 VPWR VGND sg13g2_decap_8
XFILLER_14_893 VPWR VGND sg13g2_decap_8
XFILLER_32_189 VPWR VGND sg13g2_decap_8
XFILLER_9_396 VPWR VGND sg13g2_decap_8
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_36_462 VPWR VGND sg13g2_decap_8
XFILLER_24_613 VPWR VGND sg13g2_decap_8
XFILLER_23_123 VPWR VGND sg13g2_decap_8
XFILLER_20_830 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_decap_8
XFILLER_4_1019 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_27_462 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_decap_8
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_43_966 VPWR VGND sg13g2_decap_8
XFILLER_42_476 VPWR VGND sg13g2_decap_8
XFILLER_30_616 VPWR VGND sg13g2_decap_8
XFILLER_11_830 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_decap_8
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_7_812 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_7_889 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_38_749 VPWR VGND sg13g2_decap_8
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_19_963 VPWR VGND sg13g2_decap_8
XFILLER_18_473 VPWR VGND sg13g2_decap_8
XFILLER_34_966 VPWR VGND sg13g2_decap_8
XFILLER_33_476 VPWR VGND sg13g2_decap_8
XFILLER_21_627 VPWR VGND sg13g2_decap_8
XFILLER_14_690 VPWR VGND sg13g2_decap_8
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_9_193 VPWR VGND sg13g2_decap_8
XFILLER_29_749 VPWR VGND sg13g2_decap_8
XFILLER_25_900 VPWR VGND sg13g2_decap_8
XFILLER_24_410 VPWR VGND sg13g2_decap_8
XFILLER_40_903 VPWR VGND sg13g2_decap_8
XFILLER_25_977 VPWR VGND sg13g2_decap_8
XFILLER_19_1005 VPWR VGND sg13g2_decap_8
XFILLER_12_627 VPWR VGND sg13g2_decap_8
XFILLER_24_487 VPWR VGND sg13g2_decap_8
XFILLER_11_137 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_3_347 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_16_900 VPWR VGND sg13g2_decap_8
XFILLER_28_760 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_31_903 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_30_413 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_6_130 VPWR VGND sg13g2_decap_8
XFILLER_7_686 VPWR VGND sg13g2_decap_8
XFILLER_38_546 VPWR VGND sg13g2_decap_8
XFILLER_19_760 VPWR VGND sg13g2_decap_8
XFILLER_25_207 VPWR VGND sg13g2_decap_8
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_34_763 VPWR VGND sg13g2_decap_8
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_33_273 VPWR VGND sg13g2_decap_8
XFILLER_21_424 VPWR VGND sg13g2_decap_8
XFILLER_30_980 VPWR VGND sg13g2_decap_8
XFILLER_29_546 VPWR VGND sg13g2_decap_8
XFILLER_16_207 VPWR VGND sg13g2_decap_8
XFILLER_17_77 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_40_700 VPWR VGND sg13g2_decap_8
XFILLER_25_774 VPWR VGND sg13g2_decap_8
XFILLER_12_424 VPWR VGND sg13g2_decap_8
XFILLER_9_907 VPWR VGND sg13g2_decap_8
XFILLER_33_21 VPWR VGND sg13g2_decap_8
XFILLER_24_284 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_40_777 VPWR VGND sg13g2_decap_8
XFILLER_33_98 VPWR VGND sg13g2_decap_8
XFILLER_21_991 VPWR VGND sg13g2_decap_8
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_16_774 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
XFILLER_31_700 VPWR VGND sg13g2_decap_8
XFILLER_15_284 VPWR VGND sg13g2_decap_8
XFILLER_30_210 VPWR VGND sg13g2_decap_8
XFILLER_31_777 VPWR VGND sg13g2_decap_8
XFILLER_12_991 VPWR VGND sg13g2_decap_8
XFILLER_30_287 VPWR VGND sg13g2_decap_8
XFILLER_8_984 VPWR VGND sg13g2_decap_8
XFILLER_7_483 VPWR VGND sg13g2_decap_8
XFILLER_39_833 VPWR VGND sg13g2_decap_8
XFILLER_38_343 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_34_560 VPWR VGND sg13g2_decap_8
XFILLER_22_711 VPWR VGND sg13g2_decap_8
XFILLER_21_221 VPWR VGND sg13g2_decap_8
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
XFILLER_22_788 VPWR VGND sg13g2_decap_8
XFILLER_21_298 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_343 VPWR VGND sg13g2_decap_8
XFILLER_45_847 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_12_221 VPWR VGND sg13g2_decap_8
XFILLER_25_571 VPWR VGND sg13g2_decap_8
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_40_574 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_921 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_5_998 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_39_1008 VPWR VGND sg13g2_decap_8
XFILLER_36_847 VPWR VGND sg13g2_decap_8
XFILLER_35_357 VPWR VGND sg13g2_decap_8
XFILLER_23_508 VPWR VGND sg13g2_decap_8
XFILLER_16_571 VPWR VGND sg13g2_decap_8
XFILLER_31_574 VPWR VGND sg13g2_decap_8
XFILLER_8_781 VPWR VGND sg13g2_decap_8
XFILLER_7_280 VPWR VGND sg13g2_decap_8
XFILLER_39_630 VPWR VGND sg13g2_decap_8
XFILLER_22_1012 VPWR VGND sg13g2_decap_8
XFILLER_38_140 VPWR VGND sg13g2_decap_8
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_14_508 VPWR VGND sg13g2_decap_8
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_14_67 VPWR VGND sg13g2_decap_8
XFILLER_22_585 VPWR VGND sg13g2_decap_8
XFILLER_6_718 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_49_427 VPWR VGND sg13g2_decap_8
XFILLER_29_140 VPWR VGND sg13g2_decap_8
XFILLER_45_644 VPWR VGND sg13g2_decap_8
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_17_357 VPWR VGND sg13g2_decap_8
XFILLER_44_154 VPWR VGND sg13g2_decap_8
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_41_861 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_9_578 VPWR VGND sg13g2_decap_8
XFILLER_5_795 VPWR VGND sg13g2_decap_8
XFILLER_45_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_994 VPWR VGND sg13g2_decap_8
XFILLER_36_644 VPWR VGND sg13g2_decap_8
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_decap_8
XFILLER_32_861 VPWR VGND sg13g2_decap_8
XFILLER_31_371 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_14_305 VPWR VGND sg13g2_decap_8
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_42_658 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_23_872 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_22_382 VPWR VGND sg13g2_decap_8
XFILLER_6_515 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_33_658 VPWR VGND sg13g2_decap_8
XFILLER_21_809 VPWR VGND sg13g2_decap_8
XFILLER_14_872 VPWR VGND sg13g2_decap_8
XFILLER_32_168 VPWR VGND sg13g2_decap_8
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_9_375 VPWR VGND sg13g2_decap_8
XFILLER_5_592 VPWR VGND sg13g2_decap_8
XFILLER_49_791 VPWR VGND sg13g2_decap_8
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_24_669 VPWR VGND sg13g2_decap_8
XFILLER_11_319 VPWR VGND sg13g2_decap_8
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_20_886 VPWR VGND sg13g2_decap_8
XFILLER_11_46 VPWR VGND sg13g2_decap_8
XFILLER_3_529 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_28_942 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_14_102 VPWR VGND sg13g2_decap_8
XFILLER_43_945 VPWR VGND sg13g2_decap_8
XFILLER_15_669 VPWR VGND sg13g2_decap_8
XFILLER_42_455 VPWR VGND sg13g2_decap_8
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_decap_8
XFILLER_35_1022 VPWR VGND sg13g2_decap_8
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_7_868 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_38_728 VPWR VGND sg13g2_decap_8
XFILLER_37_238 VPWR VGND sg13g2_decap_8
XFILLER_19_942 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_decap_8
XFILLER_34_945 VPWR VGND sg13g2_decap_8
XFILLER_33_455 VPWR VGND sg13g2_decap_8
XFILLER_21_606 VPWR VGND sg13g2_decap_8
XFILLER_20_116 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_decap_8
XFILLER_29_728 VPWR VGND sg13g2_decap_8
XFILLER_28_249 VPWR VGND sg13g2_decap_8
XFILLER_25_956 VPWR VGND sg13g2_decap_8
XFILLER_12_606 VPWR VGND sg13g2_decap_8
XFILLER_24_466 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_116 VPWR VGND sg13g2_decap_8
XFILLER_40_959 VPWR VGND sg13g2_decap_8
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_20_683 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_43_742 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_31_959 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_30_469 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_7_665 VPWR VGND sg13g2_decap_8
XFILLER_6_186 VPWR VGND sg13g2_decap_8
XFILLER_3_893 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_525 VPWR VGND sg13g2_decap_8
XFILLER_34_742 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_decap_8
XFILLER_21_403 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_525 VPWR VGND sg13g2_decap_8
XFILLER_44_539 VPWR VGND sg13g2_decap_8
XFILLER_17_56 VPWR VGND sg13g2_decap_8
XFILLER_25_753 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_24_263 VPWR VGND sg13g2_decap_8
XFILLER_40_756 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_decap_8
XFILLER_21_970 VPWR VGND sg13g2_decap_8
XFILLER_20_480 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_35_539 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_16_753 VPWR VGND sg13g2_decap_8
XFILLER_15_263 VPWR VGND sg13g2_decap_8
XFILLER_31_756 VPWR VGND sg13g2_decap_8
XFILLER_12_970 VPWR VGND sg13g2_decap_8
XFILLER_30_266 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_decap_8
XFILLER_8_963 VPWR VGND sg13g2_decap_8
XFILLER_7_462 VPWR VGND sg13g2_decap_8
XFILLER_3_690 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_889 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_38_399 VPWR VGND sg13g2_decap_8
XFILLER_21_200 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_22_767 VPWR VGND sg13g2_decap_8
XFILLER_21_277 VPWR VGND sg13g2_decap_8
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_29_322 VPWR VGND sg13g2_decap_8
XFILLER_45_826 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_29_399 VPWR VGND sg13g2_decap_8
XFILLER_17_539 VPWR VGND sg13g2_decap_8
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_25_550 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_40_553 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_decap_8
XFILLER_5_900 VPWR VGND sg13g2_decap_8
XFILLER_4_410 VPWR VGND sg13g2_decap_8
XFILLER_5_977 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_36_826 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_16_550 VPWR VGND sg13g2_decap_8
XFILLER_31_553 VPWR VGND sg13g2_decap_8
XFILLER_8_760 VPWR VGND sg13g2_decap_8
XFILLER_39_686 VPWR VGND sg13g2_decap_8
XFILLER_27_826 VPWR VGND sg13g2_decap_8
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_26_347 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_14_46 VPWR VGND sg13g2_decap_8
XFILLER_22_564 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_49_406 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_17_336 VPWR VGND sg13g2_decap_8
XFILLER_45_623 VPWR VGND sg13g2_decap_8
XFILLER_29_196 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_41_840 VPWR VGND sg13g2_decap_8
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_5_774 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_49_973 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_36_623 VPWR VGND sg13g2_decap_8
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_32_840 VPWR VGND sg13g2_decap_8
XFILLER_31_350 VPWR VGND sg13g2_decap_8
XFILLER_39_483 VPWR VGND sg13g2_decap_8
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_26_144 VPWR VGND sg13g2_decap_8
XFILLER_42_637 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_23_851 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_22_361 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_29_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_8
XFILLER_17_133 VPWR VGND sg13g2_decap_8
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_45_497 VPWR VGND sg13g2_decap_8
XFILLER_33_637 VPWR VGND sg13g2_decap_8
XFILLER_14_851 VPWR VGND sg13g2_decap_8
XFILLER_32_147 VPWR VGND sg13g2_decap_8
XFILLER_13_361 VPWR VGND sg13g2_decap_8
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
XFILLER_9_354 VPWR VGND sg13g2_decap_8
XFILLER_5_571 VPWR VGND sg13g2_decap_8
XFILLER_49_770 VPWR VGND sg13g2_decap_8
XFILLER_37_910 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_420 VPWR VGND sg13g2_decap_8
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_36_497 VPWR VGND sg13g2_decap_8
XFILLER_24_648 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_20_865 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
XFILLER_3_508 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_28_921 VPWR VGND sg13g2_decap_8
XFILLER_27_420 VPWR VGND sg13g2_decap_8
XFILLER_43_924 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_42_434 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_14_158 VPWR VGND sg13g2_decap_8
XFILLER_35_1001 VPWR VGND sg13g2_decap_8
XFILLER_11_865 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_7_847 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_38_707 VPWR VGND sg13g2_decap_8
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_19_921 VPWR VGND sg13g2_decap_8
XFILLER_18_431 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_34_924 VPWR VGND sg13g2_decap_8
XFILLER_19_998 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_decap_8
XFILLER_33_434 VPWR VGND sg13g2_decap_8
XFILLER_9_151 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_29_707 VPWR VGND sg13g2_decap_8
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_37_784 VPWR VGND sg13g2_decap_8
XFILLER_25_935 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_24_445 VPWR VGND sg13g2_decap_8
XFILLER_40_938 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_20_662 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_19_228 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_16_935 VPWR VGND sg13g2_decap_8
XFILLER_28_795 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_8
XFILLER_27_294 VPWR VGND sg13g2_decap_8
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_43_798 VPWR VGND sg13g2_decap_8
XFILLER_31_938 VPWR VGND sg13g2_decap_8
XFILLER_30_448 VPWR VGND sg13g2_decap_8
XFILLER_11_662 VPWR VGND sg13g2_decap_8
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_7_644 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_3_872 VPWR VGND sg13g2_decap_8
XFILLER_2_382 VPWR VGND sg13g2_decap_8
XFILLER_38_504 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_34_721 VPWR VGND sg13g2_decap_8
XFILLER_19_795 VPWR VGND sg13g2_decap_8
XFILLER_33_231 VPWR VGND sg13g2_decap_8
XFILLER_34_798 VPWR VGND sg13g2_decap_8
XFILLER_22_949 VPWR VGND sg13g2_decap_8
XFILLER_21_459 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_29_504 VPWR VGND sg13g2_decap_8
XFILLER_17_35 VPWR VGND sg13g2_decap_8
XFILLER_44_518 VPWR VGND sg13g2_decap_8
XFILLER_37_581 VPWR VGND sg13g2_decap_8
XFILLER_25_732 VPWR VGND sg13g2_decap_8
XFILLER_24_242 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_40_735 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_decap_8
XFILLER_33_56 VPWR VGND sg13g2_decap_8
XFILLER_32_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_35_518 VPWR VGND sg13g2_decap_8
XFILLER_16_732 VPWR VGND sg13g2_decap_8
XFILLER_28_592 VPWR VGND sg13g2_decap_8
XFILLER_15_242 VPWR VGND sg13g2_decap_8
XFILLER_43_595 VPWR VGND sg13g2_decap_8
XFILLER_31_735 VPWR VGND sg13g2_decap_8
XFILLER_30_245 VPWR VGND sg13g2_decap_8
XFILLER_7_441 VPWR VGND sg13g2_decap_8
XFILLER_8_942 VPWR VGND sg13g2_decap_8
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
XFILLER_38_301 VPWR VGND sg13g2_decap_8
XFILLER_39_868 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_decap_8
XFILLER_26_529 VPWR VGND sg13g2_decap_8
XFILLER_19_592 VPWR VGND sg13g2_decap_8
XFILLER_34_595 VPWR VGND sg13g2_decap_8
XFILLER_22_746 VPWR VGND sg13g2_decap_8
XFILLER_21_256 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_29_301 VPWR VGND sg13g2_decap_8
XFILLER_17_518 VPWR VGND sg13g2_decap_8
XFILLER_45_805 VPWR VGND sg13g2_decap_8
XFILLER_29_378 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_40_532 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_5_956 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
XFILLER_36_805 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_44_882 VPWR VGND sg13g2_decap_8
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_31_532 VPWR VGND sg13g2_decap_8
XFILLER_39_665 VPWR VGND sg13g2_decap_8
XFILLER_27_805 VPWR VGND sg13g2_decap_8
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_26_326 VPWR VGND sg13g2_decap_8
XFILLER_42_819 VPWR VGND sg13g2_decap_8
XFILLER_41_329 VPWR VGND sg13g2_decap_8
XFILLER_35_882 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_34_392 VPWR VGND sg13g2_decap_8
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_7_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_45_602 VPWR VGND sg13g2_decap_8
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_17_315 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_29_175 VPWR VGND sg13g2_decap_8
XFILLER_45_679 VPWR VGND sg13g2_decap_8
XFILLER_33_819 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_32_329 VPWR VGND sg13g2_decap_8
XFILLER_26_893 VPWR VGND sg13g2_decap_8
XFILLER_13_543 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
XFILLER_41_896 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_8
XFILLER_4_263 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_36_602 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_36_679 VPWR VGND sg13g2_decap_8
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_17_882 VPWR VGND sg13g2_decap_8
XFILLER_32_896 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_39_462 VPWR VGND sg13g2_decap_8
XFILLER_27_602 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_42_616 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_23_830 VPWR VGND sg13g2_decap_8
XFILLER_22_340 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_17_112 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_decap_8
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_decap_8
XFILLER_33_616 VPWR VGND sg13g2_decap_8
XFILLER_14_830 VPWR VGND sg13g2_decap_8
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_32_126 VPWR VGND sg13g2_decap_8
XFILLER_26_690 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
XFILLER_41_693 VPWR VGND sg13g2_decap_8
XFILLER_5_550 VPWR VGND sg13g2_decap_8
XFILLER_37_966 VPWR VGND sg13g2_decap_8
XFILLER_36_476 VPWR VGND sg13g2_decap_8
XFILLER_24_627 VPWR VGND sg13g2_decap_8
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_32_693 VPWR VGND sg13g2_decap_8
XFILLER_20_844 VPWR VGND sg13g2_decap_8
XFILLER_28_900 VPWR VGND sg13g2_decap_8
XFILLER_43_903 VPWR VGND sg13g2_decap_8
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_decap_8
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_7_826 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_19_900 VPWR VGND sg13g2_decap_8
XFILLER_18_410 VPWR VGND sg13g2_decap_8
XFILLER_19_977 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_decap_8
XFILLER_34_903 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_33_413 VPWR VGND sg13g2_decap_8
XFILLER_42_980 VPWR VGND sg13g2_decap_8
XFILLER_9_130 VPWR VGND sg13g2_decap_8
XFILLER_41_490 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_28_207 VPWR VGND sg13g2_decap_8
XFILLER_37_763 VPWR VGND sg13g2_decap_8
XFILLER_25_914 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_40_917 VPWR VGND sg13g2_decap_8
XFILLER_19_1019 VPWR VGND sg13g2_decap_8
XFILLER_33_980 VPWR VGND sg13g2_decap_8
XFILLER_32_490 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_20_641 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_207 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_16_914 VPWR VGND sg13g2_decap_8
XFILLER_43_700 VPWR VGND sg13g2_decap_8
XFILLER_28_774 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_27_273 VPWR VGND sg13g2_decap_8
XFILLER_43_777 VPWR VGND sg13g2_decap_8
XFILLER_31_917 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_30_427 VPWR VGND sg13g2_decap_8
XFILLER_24_991 VPWR VGND sg13g2_decap_8
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_7_623 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
XFILLER_3_851 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_34_700 VPWR VGND sg13g2_decap_8
XFILLER_19_774 VPWR VGND sg13g2_decap_8
XFILLER_33_210 VPWR VGND sg13g2_decap_8
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_34_777 VPWR VGND sg13g2_decap_8
XFILLER_15_991 VPWR VGND sg13g2_decap_8
XFILLER_33_287 VPWR VGND sg13g2_decap_8
XFILLER_22_928 VPWR VGND sg13g2_decap_8
XFILLER_21_438 VPWR VGND sg13g2_decap_8
XFILLER_30_994 VPWR VGND sg13g2_decap_8
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_37_560 VPWR VGND sg13g2_decap_8
XFILLER_25_711 VPWR VGND sg13g2_decap_8
XFILLER_24_221 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_40_714 VPWR VGND sg13g2_decap_8
XFILLER_25_788 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_decap_8
XFILLER_33_35 VPWR VGND sg13g2_decap_8
XFILLER_24_298 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_16_711 VPWR VGND sg13g2_decap_8
XFILLER_28_571 VPWR VGND sg13g2_decap_8
XFILLER_15_221 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_decap_8
XFILLER_15_298 VPWR VGND sg13g2_decap_8
XFILLER_30_224 VPWR VGND sg13g2_decap_8
XFILLER_8_921 VPWR VGND sg13g2_decap_8
XFILLER_7_420 VPWR VGND sg13g2_decap_8
XFILLER_8_998 VPWR VGND sg13g2_decap_8
XFILLER_48_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_497 VPWR VGND sg13g2_decap_8
XFILLER_39_847 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
XFILLER_26_508 VPWR VGND sg13g2_decap_8
XFILLER_19_571 VPWR VGND sg13g2_decap_8
XFILLER_34_574 VPWR VGND sg13g2_decap_8
XFILLER_22_725 VPWR VGND sg13g2_decap_8
XFILLER_21_235 VPWR VGND sg13g2_decap_8
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_30_791 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_357 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_decap_8
XFILLER_25_585 VPWR VGND sg13g2_decap_8
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_9_718 VPWR VGND sg13g2_decap_8
XFILLER_40_588 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_5_935 VPWR VGND sg13g2_decap_8
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_44_861 VPWR VGND sg13g2_decap_8
XFILLER_16_585 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_31_511 VPWR VGND sg13g2_decap_8
XFILLER_31_588 VPWR VGND sg13g2_decap_8
XFILLER_8_795 VPWR VGND sg13g2_decap_8
XFILLER_7_294 VPWR VGND sg13g2_decap_8
XFILLER_39_644 VPWR VGND sg13g2_decap_8
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_22_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_305 VPWR VGND sg13g2_decap_8
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_35_861 VPWR VGND sg13g2_decap_8
XFILLER_34_371 VPWR VGND sg13g2_decap_8
XFILLER_22_522 VPWR VGND sg13g2_decap_8
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_30_14 VPWR VGND sg13g2_decap_8
XFILLER_2_949 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_29_154 VPWR VGND sg13g2_decap_8
XFILLER_45_658 VPWR VGND sg13g2_decap_8
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_38_1022 VPWR VGND sg13g2_decap_8
XFILLER_32_308 VPWR VGND sg13g2_decap_8
XFILLER_26_872 VPWR VGND sg13g2_decap_8
XFILLER_13_522 VPWR VGND sg13g2_decap_8
XFILLER_25_382 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_41_875 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_732 VPWR VGND sg13g2_decap_8
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_45_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_931 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_36_658 VPWR VGND sg13g2_decap_8
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_23_319 VPWR VGND sg13g2_decap_8
XFILLER_17_861 VPWR VGND sg13g2_decap_8
XFILLER_16_382 VPWR VGND sg13g2_decap_8
XFILLER_32_875 VPWR VGND sg13g2_decap_8
XFILLER_31_385 VPWR VGND sg13g2_decap_8
XFILLER_8_592 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_39_441 VPWR VGND sg13g2_decap_8
XFILLER_26_102 VPWR VGND sg13g2_decap_8
XFILLER_15_809 VPWR VGND sg13g2_decap_8
XFILLER_27_658 VPWR VGND sg13g2_decap_8
XFILLER_14_319 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_23_886 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_22_396 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_49_238 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_46_945 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_decap_8
XFILLER_17_168 VPWR VGND sg13g2_decap_8
XFILLER_32_105 VPWR VGND sg13g2_decap_8
XFILLER_14_886 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
XFILLER_41_672 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_9_389 VPWR VGND sg13g2_decap_8
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_36_455 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_32_672 VPWR VGND sg13g2_decap_8
XFILLER_20_823 VPWR VGND sg13g2_decap_8
XFILLER_31_182 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_15_606 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_decap_8
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_42_469 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_7_805 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_19_956 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_18_466 VPWR VGND sg13g2_decap_8
XFILLER_34_959 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_decap_8
XFILLER_14_683 VPWR VGND sg13g2_decap_8
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_9_186 VPWR VGND sg13g2_decap_8
XFILLER_6_893 VPWR VGND sg13g2_decap_8
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_742 VPWR VGND sg13g2_decap_8
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_24_403 VPWR VGND sg13g2_decap_8
XFILLER_20_620 VPWR VGND sg13g2_decap_8
XFILLER_20_697 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_753 VPWR VGND sg13g2_decap_8
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_42_266 VPWR VGND sg13g2_decap_8
XFILLER_30_406 VPWR VGND sg13g2_decap_8
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_11_620 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_7_602 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_7_679 VPWR VGND sg13g2_decap_8
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_38_539 VPWR VGND sg13g2_decap_8
XFILLER_19_753 VPWR VGND sg13g2_decap_8
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_34_756 VPWR VGND sg13g2_decap_8
XFILLER_22_907 VPWR VGND sg13g2_decap_8
XFILLER_15_970 VPWR VGND sg13g2_decap_8
XFILLER_33_266 VPWR VGND sg13g2_decap_8
XFILLER_21_417 VPWR VGND sg13g2_decap_8
XFILLER_14_480 VPWR VGND sg13g2_decap_8
XFILLER_30_973 VPWR VGND sg13g2_decap_8
XFILLER_6_690 VPWR VGND sg13g2_decap_8
XFILLER_29_539 VPWR VGND sg13g2_decap_8
XFILLER_24_200 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_25_767 VPWR VGND sg13g2_decap_8
XFILLER_12_417 VPWR VGND sg13g2_decap_8
XFILLER_33_14 VPWR VGND sg13g2_decap_8
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_21_984 VPWR VGND sg13g2_decap_8
XFILLER_20_494 VPWR VGND sg13g2_decap_8
XFILLER_4_627 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_28_550 VPWR VGND sg13g2_decap_8
XFILLER_15_200 VPWR VGND sg13g2_decap_8
XFILLER_16_767 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_decap_8
XFILLER_15_277 VPWR VGND sg13g2_decap_8
XFILLER_30_203 VPWR VGND sg13g2_decap_8
XFILLER_8_900 VPWR VGND sg13g2_decap_8
XFILLER_12_984 VPWR VGND sg13g2_decap_8
XFILLER_11_494 VPWR VGND sg13g2_decap_8
XFILLER_7_476 VPWR VGND sg13g2_decap_8
XFILLER_8_977 VPWR VGND sg13g2_decap_8
XFILLER_39_826 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_38_336 VPWR VGND sg13g2_decap_8
XFILLER_19_550 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_553 VPWR VGND sg13g2_decap_8
XFILLER_22_704 VPWR VGND sg13g2_decap_8
XFILLER_21_214 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_decap_8
XFILLER_30_770 VPWR VGND sg13g2_decap_8
XFILLER_29_336 VPWR VGND sg13g2_decap_8
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_25_564 VPWR VGND sg13g2_decap_8
XFILLER_12_214 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_40_567 VPWR VGND sg13g2_decap_8
XFILLER_21_781 VPWR VGND sg13g2_decap_8
XFILLER_5_914 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_4_424 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_44_840 VPWR VGND sg13g2_decap_8
XFILLER_16_564 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
XFILLER_15_1012 VPWR VGND sg13g2_decap_8
XFILLER_31_567 VPWR VGND sg13g2_decap_8
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_11_291 VPWR VGND sg13g2_decap_8
XFILLER_8_774 VPWR VGND sg13g2_decap_8
XFILLER_7_273 VPWR VGND sg13g2_decap_8
XFILLER_4_991 VPWR VGND sg13g2_decap_8
XFILLER_39_623 VPWR VGND sg13g2_decap_8
XFILLER_22_1005 VPWR VGND sg13g2_decap_8
XFILLER_38_133 VPWR VGND sg13g2_decap_8
XFILLER_35_840 VPWR VGND sg13g2_decap_8
XFILLER_34_350 VPWR VGND sg13g2_decap_8
XFILLER_22_501 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_decap_8
XFILLER_2_928 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_29_133 VPWR VGND sg13g2_decap_8
XFILLER_45_637 VPWR VGND sg13g2_decap_8
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_26_851 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_8
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_25_361 VPWR VGND sg13g2_decap_8
XFILLER_41_854 VPWR VGND sg13g2_decap_8
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_decap_8
XFILLER_4_221 VPWR VGND sg13g2_decap_8
XFILLER_5_788 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
XFILLER_49_987 VPWR VGND sg13g2_decap_8
XFILLER_36_637 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_17_840 VPWR VGND sg13g2_decap_8
XFILLER_16_361 VPWR VGND sg13g2_decap_8
XFILLER_32_854 VPWR VGND sg13g2_decap_8
XFILLER_31_364 VPWR VGND sg13g2_decap_8
XFILLER_8_571 VPWR VGND sg13g2_decap_8
XFILLER_39_420 VPWR VGND sg13g2_decap_8
XFILLER_39_497 VPWR VGND sg13g2_decap_8
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_26_158 VPWR VGND sg13g2_decap_8
XFILLER_23_865 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_6_508 VPWR VGND sg13g2_decap_8
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_decap_8
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_18_648 VPWR VGND sg13g2_decap_8
XFILLER_17_147 VPWR VGND sg13g2_decap_8
XFILLER_14_865 VPWR VGND sg13g2_decap_8
XFILLER_41_651 VPWR VGND sg13g2_decap_8
XFILLER_13_375 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
XFILLER_31_91 VPWR VGND sg13g2_decap_8
XFILLER_5_585 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_49_784 VPWR VGND sg13g2_decap_8
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_36_434 VPWR VGND sg13g2_decap_8
XFILLER_32_651 VPWR VGND sg13g2_decap_8
XFILLER_31_161 VPWR VGND sg13g2_decap_8
XFILLER_20_802 VPWR VGND sg13g2_decap_8
XFILLER_20_879 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
XFILLER_28_935 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_43_938 VPWR VGND sg13g2_decap_8
XFILLER_42_448 VPWR VGND sg13g2_decap_8
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_35_1015 VPWR VGND sg13g2_decap_8
XFILLER_23_662 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_8
XFILLER_19_935 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_18_445 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_decap_8
XFILLER_34_938 VPWR VGND sg13g2_decap_8
XFILLER_33_448 VPWR VGND sg13g2_decap_8
XFILLER_14_662 VPWR VGND sg13g2_decap_8
XFILLER_20_109 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_decap_8
XFILLER_9_165 VPWR VGND sg13g2_decap_8
XFILLER_6_872 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_49_581 VPWR VGND sg13g2_decap_8
XFILLER_37_721 VPWR VGND sg13g2_decap_8
XFILLER_36_231 VPWR VGND sg13g2_decap_8
XFILLER_37_798 VPWR VGND sg13g2_decap_8
XFILLER_25_949 VPWR VGND sg13g2_decap_8
XFILLER_24_459 VPWR VGND sg13g2_decap_8
XFILLER_11_109 VPWR VGND sg13g2_decap_8
XFILLER_20_676 VPWR VGND sg13g2_decap_8
XFILLER_4_809 VPWR VGND sg13g2_decap_8
XFILLER_3_319 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_28_732 VPWR VGND sg13g2_decap_8
XFILLER_27_231 VPWR VGND sg13g2_decap_8
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_43_735 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_decap_8
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_7_658 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_3_886 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_38_518 VPWR VGND sg13g2_decap_8
XFILLER_19_732 VPWR VGND sg13g2_decap_8
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_34_735 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_decap_8
XFILLER_30_952 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_29_518 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_37_595 VPWR VGND sg13g2_decap_8
XFILLER_25_746 VPWR VGND sg13g2_decap_8
XFILLER_24_256 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_decap_8
XFILLER_21_963 VPWR VGND sg13g2_decap_8
XFILLER_20_473 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_16_746 VPWR VGND sg13g2_decap_8
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_15_256 VPWR VGND sg13g2_decap_8
XFILLER_31_749 VPWR VGND sg13g2_decap_8
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_30_259 VPWR VGND sg13g2_decap_8
XFILLER_11_473 VPWR VGND sg13g2_decap_8
XFILLER_8_956 VPWR VGND sg13g2_decap_8
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_7_455 VPWR VGND sg13g2_decap_8
XFILLER_3_683 VPWR VGND sg13g2_decap_8
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
XFILLER_34_532 VPWR VGND sg13g2_decap_8
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_315 VPWR VGND sg13g2_decap_8
XFILLER_45_819 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_38_882 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_25_543 VPWR VGND sg13g2_decap_8
XFILLER_40_546 VPWR VGND sg13g2_decap_8
XFILLER_21_760 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_36_819 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_29_882 VPWR VGND sg13g2_decap_8
XFILLER_16_543 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_44_896 VPWR VGND sg13g2_decap_8
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_31_546 VPWR VGND sg13g2_decap_8
XFILLER_12_760 VPWR VGND sg13g2_decap_8
XFILLER_11_270 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_decap_8
XFILLER_4_970 VPWR VGND sg13g2_decap_8
XFILLER_3_480 VPWR VGND sg13g2_decap_8
XFILLER_39_602 VPWR VGND sg13g2_decap_8
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_679 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
XFILLER_35_896 VPWR VGND sg13g2_decap_8
XFILLER_14_39 VPWR VGND sg13g2_decap_8
XFILLER_22_557 VPWR VGND sg13g2_decap_8
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_29_112 VPWR VGND sg13g2_decap_8
XFILLER_45_616 VPWR VGND sg13g2_decap_8
XFILLER_17_329 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_29_189 VPWR VGND sg13g2_decap_8
XFILLER_26_830 VPWR VGND sg13g2_decap_8
XFILLER_25_340 VPWR VGND sg13g2_decap_8
XFILLER_41_833 VPWR VGND sg13g2_decap_8
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_49_966 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_36_616 VPWR VGND sg13g2_decap_8
XFILLER_29_91 VPWR VGND sg13g2_decap_8
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_16_340 VPWR VGND sg13g2_decap_8
XFILLER_44_693 VPWR VGND sg13g2_decap_8
XFILLER_32_833 VPWR VGND sg13g2_decap_8
XFILLER_17_896 VPWR VGND sg13g2_decap_8
XFILLER_31_343 VPWR VGND sg13g2_decap_8
XFILLER_8_550 VPWR VGND sg13g2_decap_8
XFILLER_6_95 VPWR VGND sg13g2_decap_8
XFILLER_39_476 VPWR VGND sg13g2_decap_8
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_35_693 VPWR VGND sg13g2_decap_8
XFILLER_23_844 VPWR VGND sg13g2_decap_8
XFILLER_22_354 VPWR VGND sg13g2_decap_8
XFILLER_2_704 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_46_903 VPWR VGND sg13g2_decap_8
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_17_126 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_14_844 VPWR VGND sg13g2_decap_8
XFILLER_41_630 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_decap_8
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_5_564 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_413 VPWR VGND sg13g2_decap_8
XFILLER_45_980 VPWR VGND sg13g2_decap_8
XFILLER_44_490 VPWR VGND sg13g2_decap_8
XFILLER_32_630 VPWR VGND sg13g2_decap_8
XFILLER_17_693 VPWR VGND sg13g2_decap_8
XFILLER_31_140 VPWR VGND sg13g2_decap_8
XFILLER_20_858 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
XFILLER_28_914 VPWR VGND sg13g2_decap_8
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_27_413 VPWR VGND sg13g2_decap_8
XFILLER_43_917 VPWR VGND sg13g2_decap_8
XFILLER_42_427 VPWR VGND sg13g2_decap_8
XFILLER_36_980 VPWR VGND sg13g2_decap_8
XFILLER_35_490 VPWR VGND sg13g2_decap_8
XFILLER_23_641 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
XFILLER_19_914 VPWR VGND sg13g2_decap_8
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_18_424 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_8
XFILLER_34_917 VPWR VGND sg13g2_decap_8
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_33_427 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_14_641 VPWR VGND sg13g2_decap_8
XFILLER_26_81 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
XFILLER_42_91 VPWR VGND sg13g2_decap_8
XFILLER_6_851 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_decap_8
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_49_560 VPWR VGND sg13g2_decap_8
XFILLER_37_700 VPWR VGND sg13g2_decap_8
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_37_777 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_25_928 VPWR VGND sg13g2_decap_8
XFILLER_18_991 VPWR VGND sg13g2_decap_8
XFILLER_17_490 VPWR VGND sg13g2_decap_8
XFILLER_24_438 VPWR VGND sg13g2_decap_8
XFILLER_33_994 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_20_655 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_711 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_16_928 VPWR VGND sg13g2_decap_8
XFILLER_43_714 VPWR VGND sg13g2_decap_8
XFILLER_28_788 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_27_287 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_7_637 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_decap_8
XFILLER_3_865 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_19_711 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_46_574 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_34_714 VPWR VGND sg13g2_decap_8
XFILLER_19_788 VPWR VGND sg13g2_decap_8
XFILLER_33_224 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_42_791 VPWR VGND sg13g2_decap_8
XFILLER_30_931 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
XFILLER_17_28 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_decap_8
XFILLER_25_725 VPWR VGND sg13g2_decap_8
XFILLER_24_235 VPWR VGND sg13g2_decap_8
XFILLER_40_728 VPWR VGND sg13g2_decap_8
XFILLER_33_791 VPWR VGND sg13g2_decap_8
XFILLER_33_49 VPWR VGND sg13g2_decap_8
XFILLER_32_1008 VPWR VGND sg13g2_decap_8
XFILLER_21_942 VPWR VGND sg13g2_decap_8
XFILLER_20_452 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_16_725 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_28_585 VPWR VGND sg13g2_decap_8
XFILLER_15_235 VPWR VGND sg13g2_decap_8
XFILLER_43_588 VPWR VGND sg13g2_decap_8
XFILLER_31_728 VPWR VGND sg13g2_decap_8
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_30_238 VPWR VGND sg13g2_decap_8
XFILLER_11_452 VPWR VGND sg13g2_decap_8
XFILLER_8_935 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_7_434 VPWR VGND sg13g2_decap_8
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
XFILLER_34_511 VPWR VGND sg13g2_decap_8
XFILLER_19_585 VPWR VGND sg13g2_decap_8
XFILLER_34_588 VPWR VGND sg13g2_decap_8
XFILLER_22_739 VPWR VGND sg13g2_decap_8
XFILLER_21_249 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_44_308 VPWR VGND sg13g2_decap_8
XFILLER_38_861 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_25_522 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_40_525 VPWR VGND sg13g2_decap_8
XFILLER_25_599 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_5_949 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_29_861 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_16_522 VPWR VGND sg13g2_decap_8
XFILLER_28_382 VPWR VGND sg13g2_decap_8
XFILLER_44_875 VPWR VGND sg13g2_decap_8
XFILLER_16_599 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_31_525 VPWR VGND sg13g2_decap_8
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_8_732 VPWR VGND sg13g2_decap_8
XFILLER_7_231 VPWR VGND sg13g2_decap_8
XFILLER_39_658 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_decap_8
XFILLER_19_382 VPWR VGND sg13g2_decap_8
XFILLER_35_875 VPWR VGND sg13g2_decap_8
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_34_385 VPWR VGND sg13g2_decap_8
XFILLER_22_536 VPWR VGND sg13g2_decap_8
XFILLER_30_28 VPWR VGND sg13g2_decap_8
XFILLER_18_809 VPWR VGND sg13g2_decap_8
XFILLER_17_308 VPWR VGND sg13g2_decap_8
XFILLER_29_168 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_41_812 VPWR VGND sg13g2_decap_8
XFILLER_26_886 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_25_396 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_41_889 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_5_746 VPWR VGND sg13g2_decap_8
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_49_945 VPWR VGND sg13g2_decap_8
XFILLER_29_70 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_17_875 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_44_672 VPWR VGND sg13g2_decap_8
XFILLER_32_812 VPWR VGND sg13g2_decap_8
XFILLER_16_396 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_31_322 VPWR VGND sg13g2_decap_8
XFILLER_32_889 VPWR VGND sg13g2_decap_8
XFILLER_31_399 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_455 VPWR VGND sg13g2_decap_8
XFILLER_26_116 VPWR VGND sg13g2_decap_8
XFILLER_42_609 VPWR VGND sg13g2_decap_8
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_35_672 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_23_823 VPWR VGND sg13g2_decap_8
XFILLER_34_182 VPWR VGND sg13g2_decap_8
XFILLER_22_333 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_18_606 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_8
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_33_609 VPWR VGND sg13g2_decap_8
XFILLER_14_823 VPWR VGND sg13g2_decap_8
XFILLER_32_119 VPWR VGND sg13g2_decap_8
XFILLER_26_683 VPWR VGND sg13g2_decap_8
XFILLER_13_333 VPWR VGND sg13g2_decap_8
XFILLER_25_193 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_543 VPWR VGND sg13g2_decap_8
XFILLER_49_742 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_36_469 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_decap_8
XFILLER_16_193 VPWR VGND sg13g2_decap_8
XFILLER_32_686 VPWR VGND sg13g2_decap_8
XFILLER_20_837 VPWR VGND sg13g2_decap_8
XFILLER_31_196 VPWR VGND sg13g2_decap_8
XFILLER_9_893 VPWR VGND sg13g2_decap_8
XFILLER_39_252 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_27_469 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
XFILLER_7_819 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_18_403 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_decap_8
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_33_406 VPWR VGND sg13g2_decap_8
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_14_620 VPWR VGND sg13g2_decap_8
XFILLER_26_480 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_14_697 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_41_483 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_6_830 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
XFILLER_37_756 VPWR VGND sg13g2_decap_8
XFILLER_25_907 VPWR VGND sg13g2_decap_8
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_24_417 VPWR VGND sg13g2_decap_8
XFILLER_18_970 VPWR VGND sg13g2_decap_8
XFILLER_33_973 VPWR VGND sg13g2_decap_8
XFILLER_32_483 VPWR VGND sg13g2_decap_8
XFILLER_20_634 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_9_690 VPWR VGND sg13g2_decap_8
XFILLER_16_907 VPWR VGND sg13g2_decap_8
XFILLER_28_767 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_27_266 VPWR VGND sg13g2_decap_8
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_7_616 VPWR VGND sg13g2_decap_8
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_6_137 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_844 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_19_767 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_33_203 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_18_1012 VPWR VGND sg13g2_decap_8
XFILLER_15_984 VPWR VGND sg13g2_decap_8
XFILLER_42_770 VPWR VGND sg13g2_decap_8
XFILLER_30_910 VPWR VGND sg13g2_decap_8
XFILLER_14_494 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
XFILLER_30_987 VPWR VGND sg13g2_decap_8
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
XFILLER_37_553 VPWR VGND sg13g2_decap_8
XFILLER_25_704 VPWR VGND sg13g2_decap_8
XFILLER_24_214 VPWR VGND sg13g2_decap_8
XFILLER_40_707 VPWR VGND sg13g2_decap_8
XFILLER_33_770 VPWR VGND sg13g2_decap_8
XFILLER_33_28 VPWR VGND sg13g2_decap_8
XFILLER_21_921 VPWR VGND sg13g2_decap_8
XFILLER_32_280 VPWR VGND sg13g2_decap_8
XFILLER_20_431 VPWR VGND sg13g2_decap_8
XFILLER_21_998 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_16_704 VPWR VGND sg13g2_decap_8
XFILLER_28_564 VPWR VGND sg13g2_decap_8
XFILLER_15_214 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_31_707 VPWR VGND sg13g2_decap_8
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_30_217 VPWR VGND sg13g2_decap_8
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_11_431 VPWR VGND sg13g2_decap_8
XFILLER_8_914 VPWR VGND sg13g2_decap_8
XFILLER_23_291 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
XFILLER_7_413 VPWR VGND sg13g2_decap_8
XFILLER_3_641 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_19_564 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_34_567 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_decap_8
XFILLER_15_781 VPWR VGND sg13g2_decap_8
XFILLER_21_228 VPWR VGND sg13g2_decap_8
XFILLER_14_291 VPWR VGND sg13g2_decap_8
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_30_784 VPWR VGND sg13g2_decap_8
XFILLER_7_980 VPWR VGND sg13g2_decap_8
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_38_840 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
XFILLER_25_501 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_40_504 VPWR VGND sg13g2_decap_8
XFILLER_25_578 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_21_795 VPWR VGND sg13g2_decap_8
XFILLER_5_928 VPWR VGND sg13g2_decap_8
XFILLER_4_438 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_29_840 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_16_501 VPWR VGND sg13g2_decap_8
XFILLER_28_361 VPWR VGND sg13g2_decap_8
XFILLER_44_854 VPWR VGND sg13g2_decap_8
XFILLER_16_578 VPWR VGND sg13g2_decap_8
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_31_504 VPWR VGND sg13g2_decap_8
XFILLER_15_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_711 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_8_788 VPWR VGND sg13g2_decap_8
XFILLER_7_287 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_decap_8
XFILLER_22_1019 VPWR VGND sg13g2_decap_8
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_19_361 VPWR VGND sg13g2_decap_8
XFILLER_35_854 VPWR VGND sg13g2_decap_8
XFILLER_34_364 VPWR VGND sg13g2_decap_8
XFILLER_22_515 VPWR VGND sg13g2_decap_8
XFILLER_30_581 VPWR VGND sg13g2_decap_8
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_29_147 VPWR VGND sg13g2_decap_8
XFILLER_26_865 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_38_1015 VPWR VGND sg13g2_decap_8
XFILLER_25_375 VPWR VGND sg13g2_decap_8
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_41_868 VPWR VGND sg13g2_decap_8
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_21_592 VPWR VGND sg13g2_decap_8
XFILLER_5_725 VPWR VGND sg13g2_decap_8
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_45_1008 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_44_651 VPWR VGND sg13g2_decap_8
XFILLER_17_854 VPWR VGND sg13g2_decap_8
XFILLER_16_375 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_decap_8
XFILLER_32_868 VPWR VGND sg13g2_decap_8
XFILLER_31_378 VPWR VGND sg13g2_decap_8
XFILLER_12_592 VPWR VGND sg13g2_decap_8
XFILLER_8_585 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
XFILLER_39_434 VPWR VGND sg13g2_decap_8
XFILLER_35_651 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_34_161 VPWR VGND sg13g2_decap_8
XFILLER_23_802 VPWR VGND sg13g2_decap_8
XFILLER_22_312 VPWR VGND sg13g2_decap_8
XFILLER_23_879 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_22_389 VPWR VGND sg13g2_decap_8
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_46_938 VPWR VGND sg13g2_decap_8
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_14_802 VPWR VGND sg13g2_decap_8
XFILLER_26_662 VPWR VGND sg13g2_decap_8
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_25_172 VPWR VGND sg13g2_decap_8
XFILLER_14_879 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_41_665 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_599 VPWR VGND sg13g2_decap_8
XFILLER_49_721 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_49_798 VPWR VGND sg13g2_decap_8
XFILLER_37_938 VPWR VGND sg13g2_decap_8
XFILLER_36_448 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_17_651 VPWR VGND sg13g2_decap_8
XFILLER_16_172 VPWR VGND sg13g2_decap_8
XFILLER_32_665 VPWR VGND sg13g2_decap_8
XFILLER_20_816 VPWR VGND sg13g2_decap_8
XFILLER_31_175 VPWR VGND sg13g2_decap_8
XFILLER_9_872 VPWR VGND sg13g2_decap_8
XFILLER_8_382 VPWR VGND sg13g2_decap_8
XFILLER_39_231 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_28_949 VPWR VGND sg13g2_decap_8
XFILLER_27_448 VPWR VGND sg13g2_decap_8
XFILLER_14_109 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_decap_8
XFILLER_19_949 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_18_459 VPWR VGND sg13g2_decap_8
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_14_676 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_41_462 VPWR VGND sg13g2_decap_8
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_5_396 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_37_735 VPWR VGND sg13g2_decap_8
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_33_952 VPWR VGND sg13g2_decap_8
XFILLER_32_462 VPWR VGND sg13g2_decap_8
XFILLER_20_613 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_41_1022 VPWR VGND sg13g2_decap_8
XFILLER_28_746 VPWR VGND sg13g2_decap_8
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_43_749 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_19_746 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_34_749 VPWR VGND sg13g2_decap_8
XFILLER_15_963 VPWR VGND sg13g2_decap_8
XFILLER_33_259 VPWR VGND sg13g2_decap_8
XFILLER_14_473 VPWR VGND sg13g2_decap_8
XFILLER_30_966 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_decap_8
XFILLER_6_683 VPWR VGND sg13g2_decap_8
XFILLER_5_193 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_392 VPWR VGND sg13g2_decap_8
XFILLER_37_532 VPWR VGND sg13g2_decap_8
XFILLER_21_900 VPWR VGND sg13g2_decap_8
XFILLER_20_410 VPWR VGND sg13g2_decap_8
XFILLER_21_977 VPWR VGND sg13g2_decap_8
XFILLER_20_487 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_28_543 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_24_760 VPWR VGND sg13g2_decap_8
XFILLER_11_410 VPWR VGND sg13g2_decap_8
XFILLER_23_270 VPWR VGND sg13g2_decap_8
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_7_469 VPWR VGND sg13g2_decap_8
XFILLER_3_620 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_3_697 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_19_543 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_34_546 VPWR VGND sg13g2_decap_8
XFILLER_15_760 VPWR VGND sg13g2_decap_8
XFILLER_21_207 VPWR VGND sg13g2_decap_8
XFILLER_14_270 VPWR VGND sg13g2_decap_8
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_30_763 VPWR VGND sg13g2_decap_8
XFILLER_6_480 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_29_329 VPWR VGND sg13g2_decap_8
XFILLER_38_896 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_8
XFILLER_25_557 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_decap_8
XFILLER_21_774 VPWR VGND sg13g2_decap_8
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_5_907 VPWR VGND sg13g2_decap_8
XFILLER_4_417 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_28_340 VPWR VGND sg13g2_decap_8
XFILLER_44_833 VPWR VGND sg13g2_decap_8
XFILLER_29_896 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_16_557 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
XFILLER_15_1005 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
XFILLER_8_767 VPWR VGND sg13g2_decap_8
XFILLER_4_984 VPWR VGND sg13g2_decap_8
XFILLER_3_494 VPWR VGND sg13g2_decap_8
XFILLER_39_616 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_38_126 VPWR VGND sg13g2_decap_8
XFILLER_19_340 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_35_833 VPWR VGND sg13g2_decap_8
XFILLER_34_343 VPWR VGND sg13g2_decap_8
XFILLER_30_560 VPWR VGND sg13g2_decap_8
XFILLER_39_28 VPWR VGND sg13g2_decap_8
XFILLER_29_126 VPWR VGND sg13g2_decap_8
XFILLER_38_693 VPWR VGND sg13g2_decap_8
XFILLER_26_844 VPWR VGND sg13g2_decap_8
XFILLER_25_354 VPWR VGND sg13g2_decap_8
XFILLER_41_847 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_21_571 VPWR VGND sg13g2_decap_8
XFILLER_5_704 VPWR VGND sg13g2_decap_8
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_49_903 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_44_630 VPWR VGND sg13g2_decap_8
XFILLER_29_693 VPWR VGND sg13g2_decap_8
XFILLER_17_833 VPWR VGND sg13g2_decap_8
XFILLER_16_354 VPWR VGND sg13g2_decap_8
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_32_847 VPWR VGND sg13g2_decap_8
XFILLER_31_357 VPWR VGND sg13g2_decap_8
XFILLER_12_571 VPWR VGND sg13g2_decap_8
XFILLER_8_564 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
XFILLER_4_781 VPWR VGND sg13g2_decap_8
XFILLER_3_291 VPWR VGND sg13g2_decap_8
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_48_980 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_35_630 VPWR VGND sg13g2_decap_8
XFILLER_34_140 VPWR VGND sg13g2_decap_8
XFILLER_23_858 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_22_368 VPWR VGND sg13g2_decap_8
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_46_917 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_39_980 VPWR VGND sg13g2_decap_8
XFILLER_38_490 VPWR VGND sg13g2_decap_8
XFILLER_26_641 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_decap_8
XFILLER_14_858 VPWR VGND sg13g2_decap_8
XFILLER_13_368 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_decap_8
XFILLER_5_578 VPWR VGND sg13g2_decap_8
XFILLER_49_700 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_36_427 VPWR VGND sg13g2_decap_8
XFILLER_29_490 VPWR VGND sg13g2_decap_8
XFILLER_17_630 VPWR VGND sg13g2_decap_8
XFILLER_16_151 VPWR VGND sg13g2_decap_8
XFILLER_45_994 VPWR VGND sg13g2_decap_8
XFILLER_32_644 VPWR VGND sg13g2_decap_8
XFILLER_31_154 VPWR VGND sg13g2_decap_8
XFILLER_9_851 VPWR VGND sg13g2_decap_8
XFILLER_8_361 VPWR VGND sg13g2_decap_8
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_28_928 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
XFILLER_27_427 VPWR VGND sg13g2_decap_8
XFILLER_36_994 VPWR VGND sg13g2_decap_8
XFILLER_35_1008 VPWR VGND sg13g2_decap_8
XFILLER_23_655 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_decap_8
XFILLER_19_928 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_decap_8
XFILLER_42_931 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_14_655 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_9_158 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_6_865 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_574 VPWR VGND sg13g2_decap_8
XFILLER_37_714 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_45_791 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_8
XFILLER_32_441 VPWR VGND sg13g2_decap_8
XFILLER_20_669 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_41_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_725 VPWR VGND sg13g2_decap_8
XFILLER_27_224 VPWR VGND sg13g2_decap_8
XFILLER_43_728 VPWR VGND sg13g2_decap_8
XFILLER_36_791 VPWR VGND sg13g2_decap_8
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_24_942 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_3_879 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_19_725 VPWR VGND sg13g2_decap_8
XFILLER_18_235 VPWR VGND sg13g2_decap_8
XFILLER_46_588 VPWR VGND sg13g2_decap_8
XFILLER_34_728 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_15_942 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_decap_8
XFILLER_14_452 VPWR VGND sg13g2_decap_8
XFILLER_30_945 VPWR VGND sg13g2_decap_8
XFILLER_6_662 VPWR VGND sg13g2_decap_8
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_49_371 VPWR VGND sg13g2_decap_8
XFILLER_37_511 VPWR VGND sg13g2_decap_8
XFILLER_37_588 VPWR VGND sg13g2_decap_8
XFILLER_25_739 VPWR VGND sg13g2_decap_8
XFILLER_24_249 VPWR VGND sg13g2_decap_8
XFILLER_21_956 VPWR VGND sg13g2_decap_8
XFILLER_20_466 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_28_522 VPWR VGND sg13g2_decap_8
XFILLER_16_739 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_28_599 VPWR VGND sg13g2_decap_8
XFILLER_15_249 VPWR VGND sg13g2_decap_8
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_11_466 VPWR VGND sg13g2_decap_8
XFILLER_7_448 VPWR VGND sg13g2_decap_8
XFILLER_8_949 VPWR VGND sg13g2_decap_8
XFILLER_23_74 VPWR VGND sg13g2_decap_8
XFILLER_3_676 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_19_522 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_34_525 VPWR VGND sg13g2_decap_8
XFILLER_19_599 VPWR VGND sg13g2_decap_8
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_30_742 VPWR VGND sg13g2_decap_8
XFILLER_31_1022 VPWR VGND sg13g2_decap_8
XFILLER_9_1012 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_29_308 VPWR VGND sg13g2_decap_8
XFILLER_38_875 VPWR VGND sg13g2_decap_8
XFILLER_37_385 VPWR VGND sg13g2_decap_8
XFILLER_25_536 VPWR VGND sg13g2_decap_8
XFILLER_40_539 VPWR VGND sg13g2_decap_8
XFILLER_21_753 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_44_812 VPWR VGND sg13g2_decap_8
XFILLER_29_875 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_16_536 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_28_396 VPWR VGND sg13g2_decap_8
XFILLER_44_889 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_31_539 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_7_245 VPWR VGND sg13g2_decap_8
XFILLER_4_963 VPWR VGND sg13g2_decap_8
XFILLER_3_473 VPWR VGND sg13g2_decap_8
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
XFILLER_34_322 VPWR VGND sg13g2_decap_8
XFILLER_19_396 VPWR VGND sg13g2_decap_8
XFILLER_35_889 VPWR VGND sg13g2_decap_8
XFILLER_34_399 VPWR VGND sg13g2_decap_8
XFILLER_29_105 VPWR VGND sg13g2_decap_8
XFILLER_45_609 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_38_672 VPWR VGND sg13g2_decap_8
XFILLER_26_823 VPWR VGND sg13g2_decap_8
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_25_333 VPWR VGND sg13g2_decap_8
XFILLER_41_826 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_21_550 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_49_959 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_36_609 VPWR VGND sg13g2_decap_8
XFILLER_29_84 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_29_672 VPWR VGND sg13g2_decap_8
XFILLER_17_812 VPWR VGND sg13g2_decap_8
XFILLER_16_333 VPWR VGND sg13g2_decap_8
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_17_889 VPWR VGND sg13g2_decap_8
XFILLER_44_686 VPWR VGND sg13g2_decap_8
XFILLER_32_826 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_31_336 VPWR VGND sg13g2_decap_8
XFILLER_12_550 VPWR VGND sg13g2_decap_8
XFILLER_8_543 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_4_760 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
XFILLER_6_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_469 VPWR VGND sg13g2_decap_8
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_19_193 VPWR VGND sg13g2_decap_8
XFILLER_35_686 VPWR VGND sg13g2_decap_8
XFILLER_23_837 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_decap_8
XFILLER_22_347 VPWR VGND sg13g2_decap_8
Xheichips25_template_20 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_17_119 VPWR VGND sg13g2_decap_8
XFILLER_26_620 VPWR VGND sg13g2_decap_8
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_14_837 VPWR VGND sg13g2_decap_8
XFILLER_41_623 VPWR VGND sg13g2_decap_8
XFILLER_26_697 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_31_63 VPWR VGND sg13g2_decap_8
XFILLER_5_557 VPWR VGND sg13g2_decap_8
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_756 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_406 VPWR VGND sg13g2_decap_8
XFILLER_16_130 VPWR VGND sg13g2_decap_8
XFILLER_45_973 VPWR VGND sg13g2_decap_8
XFILLER_44_483 VPWR VGND sg13g2_decap_8
XFILLER_32_623 VPWR VGND sg13g2_decap_8
XFILLER_17_686 VPWR VGND sg13g2_decap_8
XFILLER_31_133 VPWR VGND sg13g2_decap_8
XFILLER_9_830 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
.ends

