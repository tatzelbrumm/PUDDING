** sch_path: /home/user/PUDDING/tb/DC_sim.sch
**.subckt DC_sim
DAC_TOP net1 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3
+ net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 net3 Vout GND net2 DAC_TOP
V1 net1 GND 1.5
.save i(v1)
V2 Vout GND 0.4
.save i(v2)
Iref net2 GND 100n
V3 net3 GND 0
.save i(v3)
**** begin user architecture code


*.include dc_dac.save
.param temp=27
.control
save all
op
write dc_dac.raw
set appendwrite
dc VON 0 1.2 1.2
write dc_dac.raw.raw
.endc


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  /home/user/PUDDING/schematic/DAC_TOP.sym # of pins=5
** sym_path: /home/user/PUDDING/schematic/DAC_TOP.sym
** sch_path: /home/user/PUDDING/schematic/DAC_TOP.sch
.subckt DAC_TOP VDD ON[255] ON[254] ON[253] ON[252] ON[251] ON[250] ON[249] ON[248] ON[247] ON[246] ON[245] ON[244] ON[243]
+ ON[242] ON[241] ON[240] ON[239] ON[238] ON[237] ON[236] ON[235] ON[234] ON[233] ON[232] ON[231] ON[230] ON[229] ON[228] ON[227] ON[226]
+ ON[225] ON[224] ON[223] ON[222] ON[221] ON[220] ON[219] ON[218] ON[217] ON[216] ON[215] ON[214] ON[213] ON[212] ON[211] ON[210] ON[209]
+ ON[208] ON[207] ON[206] ON[205] ON[204] ON[203] ON[202] ON[201] ON[200] ON[199] ON[198] ON[197] ON[196] ON[195] ON[194] ON[193] ON[192]
+ ON[191] ON[190] ON[189] ON[188] ON[187] ON[186] ON[185] ON[184] ON[183] ON[182] ON[181] ON[180] ON[179] ON[178] ON[177] ON[176] ON[175]
+ ON[174] ON[173] ON[172] ON[171] ON[170] ON[169] ON[168] ON[167] ON[166] ON[165] ON[164] ON[163] ON[162] ON[161] ON[160] ON[159] ON[158]
+ ON[157] ON[156] ON[155] ON[154] ON[153] ON[152] ON[151] ON[150] ON[149] ON[148] ON[147] ON[146] ON[145] ON[144] ON[143] ON[142] ON[141]
+ ON[140] ON[139] ON[138] ON[137] ON[136] ON[135] ON[134] ON[133] ON[132] ON[131] ON[130] ON[129] ON[128] ON[127] ON[126] ON[125] ON[124]
+ ON[123] ON[122] ON[121] ON[120] ON[119] ON[118] ON[117] ON[116] ON[115] ON[114] ON[113] ON[112] ON[111] ON[110] ON[109] ON[108] ON[107]
+ ON[106] ON[105] ON[104] ON[103] ON[102] ON[101] ON[100] ON[99] ON[98] ON[97] ON[96] ON[95] ON[94] ON[93] ON[92] ON[91] ON[90] ON[89]
+ ON[88] ON[87] ON[86] ON[85] ON[84] ON[83] ON[82] ON[81] ON[80] ON[79] ON[78] ON[77] ON[76] ON[75] ON[74] ON[73] ON[72] ON[71] ON[70]
+ ON[69] ON[68] ON[67] ON[66] ON[65] ON[64] ON[63] ON[62] ON[61] ON[60] ON[59] ON[58] ON[57] ON[56] ON[55] ON[54] ON[53] ON[52] ON[51]
+ ON[50] ON[49] ON[48] ON[47] ON[46] ON[45] ON[44] ON[43] ON[42] ON[41] ON[40] ON[39] ON[38] ON[37] ON[36] ON[35] ON[34] ON[33] ON[32]
+ ON[31] ON[30] ON[29] ON[28] ON[27] ON[26] ON[25] ON[24] ON[23] ON[22] ON[21] ON[20] ON[19] ON[18] ON[17] ON[16] ON[15] ON[14] ON[13]
+ ON[12] ON[11] ON[10] ON[9] ON[8] ON[7] ON[6] ON[5] ON[4] ON[3] ON[2] ON[1] ON[0] Iout ESDGND Iref
*.ipin VDD
*.opin Iout
*.ipin ESDGND
*.ipin
*+ ON[255],ON[254],ON[253],ON[252],ON[251],ON[250],ON[249],ON[248],ON[247],ON[246],ON[245],ON[244],ON[243],ON[242],ON[241],ON[240],ON[239],ON[238],ON[237],ON[236],ON[235],ON[234],ON[233],ON[232],ON[231],ON[230],ON[229],ON[228],ON[227],ON[226],ON[225],ON[224],ON[223],ON[222],ON[221],ON[220],ON[219],ON[218],ON[217],ON[216],ON[215],ON[214],ON[213],ON[212],ON[211],ON[210],ON[209],ON[208],ON[207],ON[206],ON[205],ON[204],ON[203],ON[202],ON[201],ON[200],ON[199],ON[198],ON[197],ON[196],ON[195],ON[194],ON[193],ON[192],ON[191],ON[190],ON[189],ON[188],ON[187],ON[186],ON[185],ON[184],ON[183],ON[182],ON[181],ON[180],ON[179],ON[178],ON[177],ON[176],ON[175],ON[174],ON[173],ON[172],ON[171],ON[170],ON[169],ON[168],ON[167],ON[166],ON[165],ON[164],ON[163],ON[162],ON[161],ON[160],ON[159],ON[158],ON[157],ON[156],ON[155],ON[154],ON[153],ON[152],ON[151],ON[150],ON[149],ON[148],ON[147],ON[146],ON[145],ON[144],ON[143],ON[142],ON[141],ON[140],ON[139],ON[138],ON[137],ON[136],ON[135],ON[134],ON[133],ON[132],ON[131],ON[130],ON[129],ON[128],ON[127],ON[126],ON[125],ON[124],ON[123],ON[122],ON[121],ON[120],ON[119],ON[118],ON[117],ON[116],ON[115],ON[114],ON[113],ON[112],ON[111],ON[110],ON[109],ON[108],ON[107],ON[106],ON[105],ON[104],ON[103],ON[102],ON[101],ON[100],ON[99],ON[98],ON[97],ON[96],ON[95],ON[94],ON[93],ON[92],ON[91],ON[90],ON[89],ON[88],ON[87],ON[86],ON[85],ON[84],ON[83],ON[82],ON[81],ON[80],ON[79],ON[78],ON[77],ON[76],ON[75],ON[74],ON[73],ON[72],ON[71],ON[70],ON[69],ON[68],ON[67],ON[66],ON[65],ON[64],ON[63],ON[62],ON[61],ON[60],ON[59],ON[58],ON[57],ON[56],ON[55],ON[54],ON[53],ON[52],ON[51],ON[50],ON[49],ON[48],ON[47],ON[46],ON[45],ON[44],ON[43],ON[42],ON[41],ON[40],ON[39],ON[38],ON[37],ON[36],ON[35],ON[34],ON[33],ON[32],ON[31],ON[30],ON[29],ON[28],ON[27],ON[26],ON[25],ON[24],ON[23],ON[22],ON[21],ON[20],ON[19],ON[18],ON[17],ON[16],ON[15],ON[14],ON[13],ON[12],ON[11],ON[10],ON[9],ON[8],ON[7],ON[6],ON[5],ON[4],ON[3],ON[2],ON[1],ON[0]
*.ipin Iref
x1 VDD Iout Vbias CASCODE_SW[255] CASCODE_SW[254] CASCODE_SW[253] CASCODE_SW[252] CASCODE_SW[251] CASCODE_SW[250] CASCODE_SW[249]
+ CASCODE_SW[248] CASCODE_SW[247] CASCODE_SW[246] CASCODE_SW[245] CASCODE_SW[244] CASCODE_SW[243] CASCODE_SW[242] CASCODE_SW[241] CASCODE_SW[240]
+ CASCODE_SW[239] CASCODE_SW[238] CASCODE_SW[237] CASCODE_SW[236] CASCODE_SW[235] CASCODE_SW[234] CASCODE_SW[233] CASCODE_SW[232] CASCODE_SW[231]
+ CASCODE_SW[230] CASCODE_SW[229] CASCODE_SW[228] CASCODE_SW[227] CASCODE_SW[226] CASCODE_SW[225] CASCODE_SW[224] CASCODE_SW[223] CASCODE_SW[222]
+ CASCODE_SW[221] CASCODE_SW[220] CASCODE_SW[219] CASCODE_SW[218] CASCODE_SW[217] CASCODE_SW[216] CASCODE_SW[215] CASCODE_SW[214] CASCODE_SW[213]
+ CASCODE_SW[212] CASCODE_SW[211] CASCODE_SW[210] CASCODE_SW[209] CASCODE_SW[208] CASCODE_SW[207] CASCODE_SW[206] CASCODE_SW[205] CASCODE_SW[204]
+ CASCODE_SW[203] CASCODE_SW[202] CASCODE_SW[201] CASCODE_SW[200] CASCODE_SW[199] CASCODE_SW[198] CASCODE_SW[197] CASCODE_SW[196] CASCODE_SW[195]
+ CASCODE_SW[194] CASCODE_SW[193] CASCODE_SW[192] CASCODE_SW[191] CASCODE_SW[190] CASCODE_SW[189] CASCODE_SW[188] CASCODE_SW[187] CASCODE_SW[186]
+ CASCODE_SW[185] CASCODE_SW[184] CASCODE_SW[183] CASCODE_SW[182] CASCODE_SW[181] CASCODE_SW[180] CASCODE_SW[179] CASCODE_SW[178] CASCODE_SW[177]
+ CASCODE_SW[176] CASCODE_SW[175] CASCODE_SW[174] CASCODE_SW[173] CASCODE_SW[172] CASCODE_SW[171] CASCODE_SW[170] CASCODE_SW[169] CASCODE_SW[168]
+ CASCODE_SW[167] CASCODE_SW[166] CASCODE_SW[165] CASCODE_SW[164] CASCODE_SW[163] CASCODE_SW[162] CASCODE_SW[161] CASCODE_SW[160] CASCODE_SW[159]
+ CASCODE_SW[158] CASCODE_SW[157] CASCODE_SW[156] CASCODE_SW[155] CASCODE_SW[154] CASCODE_SW[153] CASCODE_SW[152] CASCODE_SW[151] CASCODE_SW[150]
+ CASCODE_SW[149] CASCODE_SW[148] CASCODE_SW[147] CASCODE_SW[146] CASCODE_SW[145] CASCODE_SW[144] CASCODE_SW[143] CASCODE_SW[142] CASCODE_SW[141]
+ CASCODE_SW[140] CASCODE_SW[139] CASCODE_SW[138] CASCODE_SW[137] CASCODE_SW[136] CASCODE_SW[135] CASCODE_SW[134] CASCODE_SW[133] CASCODE_SW[132]
+ CASCODE_SW[131] CASCODE_SW[130] CASCODE_SW[129] CASCODE_SW[128] CASCODE_SW[127] CASCODE_SW[126] CASCODE_SW[125] CASCODE_SW[124] CASCODE_SW[123]
+ CASCODE_SW[122] CASCODE_SW[121] CASCODE_SW[120] CASCODE_SW[119] CASCODE_SW[118] CASCODE_SW[117] CASCODE_SW[116] CASCODE_SW[115] CASCODE_SW[114]
+ CASCODE_SW[113] CASCODE_SW[112] CASCODE_SW[111] CASCODE_SW[110] CASCODE_SW[109] CASCODE_SW[108] CASCODE_SW[107] CASCODE_SW[106] CASCODE_SW[105]
+ CASCODE_SW[104] CASCODE_SW[103] CASCODE_SW[102] CASCODE_SW[101] CASCODE_SW[100] CASCODE_SW[99] CASCODE_SW[98] CASCODE_SW[97] CASCODE_SW[96]
+ CASCODE_SW[95] CASCODE_SW[94] CASCODE_SW[93] CASCODE_SW[92] CASCODE_SW[91] CASCODE_SW[90] CASCODE_SW[89] CASCODE_SW[88] CASCODE_SW[87]
+ CASCODE_SW[86] CASCODE_SW[85] CASCODE_SW[84] CASCODE_SW[83] CASCODE_SW[82] CASCODE_SW[81] CASCODE_SW[80] CASCODE_SW[79] CASCODE_SW[78]
+ CASCODE_SW[77] CASCODE_SW[76] CASCODE_SW[75] CASCODE_SW[74] CASCODE_SW[73] CASCODE_SW[72] CASCODE_SW[71] CASCODE_SW[70] CASCODE_SW[69]
+ CASCODE_SW[68] CASCODE_SW[67] CASCODE_SW[66] CASCODE_SW[65] CASCODE_SW[64] CASCODE_SW[63] CASCODE_SW[62] CASCODE_SW[61] CASCODE_SW[60]
+ CASCODE_SW[59] CASCODE_SW[58] CASCODE_SW[57] CASCODE_SW[56] CASCODE_SW[55] CASCODE_SW[54] CASCODE_SW[53] CASCODE_SW[52] CASCODE_SW[51]
+ CASCODE_SW[50] CASCODE_SW[49] CASCODE_SW[48] CASCODE_SW[47] CASCODE_SW[46] CASCODE_SW[45] CASCODE_SW[44] CASCODE_SW[43] CASCODE_SW[42]
+ CASCODE_SW[41] CASCODE_SW[40] CASCODE_SW[39] CASCODE_SW[38] CASCODE_SW[37] CASCODE_SW[36] CASCODE_SW[35] CASCODE_SW[34] CASCODE_SW[33]
+ CASCODE_SW[32] CASCODE_SW[31] CASCODE_SW[30] CASCODE_SW[29] CASCODE_SW[28] CASCODE_SW[27] CASCODE_SW[26] CASCODE_SW[25] CASCODE_SW[24]
+ CASCODE_SW[23] CASCODE_SW[22] CASCODE_SW[21] CASCODE_SW[20] CASCODE_SW[19] CASCODE_SW[18] CASCODE_SW[17] CASCODE_SW[16] CASCODE_SW[15]
+ CASCODE_SW[14] CASCODE_SW[13] CASCODE_SW[12] CASCODE_SW[11] CASCODE_SW[10] CASCODE_SW[9] CASCODE_SW[8] CASCODE_SW[7] CASCODE_SW[6] CASCODE_SW[5]
+ CASCODE_SW[4] CASCODE_SW[3] CASCODE_SW[2] CASCODE_SW[1] CASCODE_SW[0] Pmirrors_top
SW VDD ON[255] CASCODE_SW[255] Iref ESDGND DAC_SW
XM2 Vbias Vbias VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 Iref Iref Vbias VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/user/PUDDING/schematic/Pmirrors_top.sym # of pins=4
** sym_path: /home/user/PUDDING/schematic/Pmirrors_top.sym
** sch_path: /home/user/PUDDING/schematic/Pmirrors_top.sch
.subckt Pmirrors_top VDD Iout Vbiasp VcascodeP[255] VcascodeP[254] VcascodeP[253] VcascodeP[252] VcascodeP[251] VcascodeP[250]
+ VcascodeP[249] VcascodeP[248] VcascodeP[247] VcascodeP[246] VcascodeP[245] VcascodeP[244] VcascodeP[243] VcascodeP[242] VcascodeP[241]
+ VcascodeP[240] VcascodeP[239] VcascodeP[238] VcascodeP[237] VcascodeP[236] VcascodeP[235] VcascodeP[234] VcascodeP[233] VcascodeP[232]
+ VcascodeP[231] VcascodeP[230] VcascodeP[229] VcascodeP[228] VcascodeP[227] VcascodeP[226] VcascodeP[225] VcascodeP[224] VcascodeP[223]
+ VcascodeP[222] VcascodeP[221] VcascodeP[220] VcascodeP[219] VcascodeP[218] VcascodeP[217] VcascodeP[216] VcascodeP[215] VcascodeP[214]
+ VcascodeP[213] VcascodeP[212] VcascodeP[211] VcascodeP[210] VcascodeP[209] VcascodeP[208] VcascodeP[207] VcascodeP[206] VcascodeP[205]
+ VcascodeP[204] VcascodeP[203] VcascodeP[202] VcascodeP[201] VcascodeP[200] VcascodeP[199] VcascodeP[198] VcascodeP[197] VcascodeP[196]
+ VcascodeP[195] VcascodeP[194] VcascodeP[193] VcascodeP[192] VcascodeP[191] VcascodeP[190] VcascodeP[189] VcascodeP[188] VcascodeP[187]
+ VcascodeP[186] VcascodeP[185] VcascodeP[184] VcascodeP[183] VcascodeP[182] VcascodeP[181] VcascodeP[180] VcascodeP[179] VcascodeP[178]
+ VcascodeP[177] VcascodeP[176] VcascodeP[175] VcascodeP[174] VcascodeP[173] VcascodeP[172] VcascodeP[171] VcascodeP[170] VcascodeP[169]
+ VcascodeP[168] VcascodeP[167] VcascodeP[166] VcascodeP[165] VcascodeP[164] VcascodeP[163] VcascodeP[162] VcascodeP[161] VcascodeP[160]
+ VcascodeP[159] VcascodeP[158] VcascodeP[157] VcascodeP[156] VcascodeP[155] VcascodeP[154] VcascodeP[153] VcascodeP[152] VcascodeP[151]
+ VcascodeP[150] VcascodeP[149] VcascodeP[148] VcascodeP[147] VcascodeP[146] VcascodeP[145] VcascodeP[144] VcascodeP[143] VcascodeP[142]
+ VcascodeP[141] VcascodeP[140] VcascodeP[139] VcascodeP[138] VcascodeP[137] VcascodeP[136] VcascodeP[135] VcascodeP[134] VcascodeP[133]
+ VcascodeP[132] VcascodeP[131] VcascodeP[130] VcascodeP[129] VcascodeP[128] VcascodeP[127] VcascodeP[126] VcascodeP[125] VcascodeP[124]
+ VcascodeP[123] VcascodeP[122] VcascodeP[121] VcascodeP[120] VcascodeP[119] VcascodeP[118] VcascodeP[117] VcascodeP[116] VcascodeP[115]
+ VcascodeP[114] VcascodeP[113] VcascodeP[112] VcascodeP[111] VcascodeP[110] VcascodeP[109] VcascodeP[108] VcascodeP[107] VcascodeP[106]
+ VcascodeP[105] VcascodeP[104] VcascodeP[103] VcascodeP[102] VcascodeP[101] VcascodeP[100] VcascodeP[99] VcascodeP[98] VcascodeP[97]
+ VcascodeP[96] VcascodeP[95] VcascodeP[94] VcascodeP[93] VcascodeP[92] VcascodeP[91] VcascodeP[90] VcascodeP[89] VcascodeP[88] VcascodeP[87]
+ VcascodeP[86] VcascodeP[85] VcascodeP[84] VcascodeP[83] VcascodeP[82] VcascodeP[81] VcascodeP[80] VcascodeP[79] VcascodeP[78] VcascodeP[77]
+ VcascodeP[76] VcascodeP[75] VcascodeP[74] VcascodeP[73] VcascodeP[72] VcascodeP[71] VcascodeP[70] VcascodeP[69] VcascodeP[68] VcascodeP[67]
+ VcascodeP[66] VcascodeP[65] VcascodeP[64] VcascodeP[63] VcascodeP[62] VcascodeP[61] VcascodeP[60] VcascodeP[59] VcascodeP[58] VcascodeP[57]
+ VcascodeP[56] VcascodeP[55] VcascodeP[54] VcascodeP[53] VcascodeP[52] VcascodeP[51] VcascodeP[50] VcascodeP[49] VcascodeP[48] VcascodeP[47]
+ VcascodeP[46] VcascodeP[45] VcascodeP[44] VcascodeP[43] VcascodeP[42] VcascodeP[41] VcascodeP[40] VcascodeP[39] VcascodeP[38] VcascodeP[37]
+ VcascodeP[36] VcascodeP[35] VcascodeP[34] VcascodeP[33] VcascodeP[32] VcascodeP[31] VcascodeP[30] VcascodeP[29] VcascodeP[28] VcascodeP[27]
+ VcascodeP[26] VcascodeP[25] VcascodeP[24] VcascodeP[23] VcascodeP[22] VcascodeP[21] VcascodeP[20] VcascodeP[19] VcascodeP[18] VcascodeP[17]
+ VcascodeP[16] VcascodeP[15] VcascodeP[14] VcascodeP[13] VcascodeP[12] VcascodeP[11] VcascodeP[10] VcascodeP[9] VcascodeP[8] VcascodeP[7]
+ VcascodeP[6] VcascodeP[5] VcascodeP[4] VcascodeP[3] VcascodeP[2] VcascodeP[1] VcascodeP[0]
*.ipin Vbiasp
*.ipin VDD
*.ipin
*+ VcascodeP[255],VcascodeP[254],VcascodeP[253],VcascodeP[252],VcascodeP[251],VcascodeP[250],VcascodeP[249],VcascodeP[248],VcascodeP[247],VcascodeP[246],VcascodeP[245],VcascodeP[244],VcascodeP[243],VcascodeP[242],VcascodeP[241],VcascodeP[240],VcascodeP[239],VcascodeP[238],VcascodeP[237],VcascodeP[236],VcascodeP[235],VcascodeP[234],VcascodeP[233],VcascodeP[232],VcascodeP[231],VcascodeP[230],VcascodeP[229],VcascodeP[228],VcascodeP[227],VcascodeP[226],VcascodeP[225],VcascodeP[224],VcascodeP[223],VcascodeP[222],VcascodeP[221],VcascodeP[220],VcascodeP[219],VcascodeP[218],VcascodeP[217],VcascodeP[216],VcascodeP[215],VcascodeP[214],VcascodeP[213],VcascodeP[212],VcascodeP[211],VcascodeP[210],VcascodeP[209],VcascodeP[208],VcascodeP[207],VcascodeP[206],VcascodeP[205],VcascodeP[204],VcascodeP[203],VcascodeP[202],VcascodeP[201],VcascodeP[200],VcascodeP[199],VcascodeP[198],VcascodeP[197],VcascodeP[196],VcascodeP[195],VcascodeP[194],VcascodeP[193],VcascodeP[192],VcascodeP[191],VcascodeP[190],VcascodeP[189],VcascodeP[188],VcascodeP[187],VcascodeP[186],VcascodeP[185],VcascodeP[184],VcascodeP[183],VcascodeP[182],VcascodeP[181],VcascodeP[180],VcascodeP[179],VcascodeP[178],VcascodeP[177],VcascodeP[176],VcascodeP[175],VcascodeP[174],VcascodeP[173],VcascodeP[172],VcascodeP[171],VcascodeP[170],VcascodeP[169],VcascodeP[168],VcascodeP[167],VcascodeP[166],VcascodeP[165],VcascodeP[164],VcascodeP[163],VcascodeP[162],VcascodeP[161],VcascodeP[160],VcascodeP[159],VcascodeP[158],VcascodeP[157],VcascodeP[156],VcascodeP[155],VcascodeP[154],VcascodeP[153],VcascodeP[152],VcascodeP[151],VcascodeP[150],VcascodeP[149],VcascodeP[148],VcascodeP[147],VcascodeP[146],VcascodeP[145],VcascodeP[144],VcascodeP[143],VcascodeP[142],VcascodeP[141],VcascodeP[140],VcascodeP[139],VcascodeP[138],VcascodeP[137],VcascodeP[136],VcascodeP[135],VcascodeP[134],VcascodeP[133],VcascodeP[132],VcascodeP[131],VcascodeP[130],VcascodeP[129],VcascodeP[128],VcascodeP[127],VcascodeP[126],VcascodeP[125],VcascodeP[124],VcascodeP[123],VcascodeP[122],VcascodeP[121],VcascodeP[120],VcascodeP[119],VcascodeP[118],VcascodeP[117],VcascodeP[116],VcascodeP[115],VcascodeP[114],VcascodeP[113],VcascodeP[112],VcascodeP[111],VcascodeP[110],VcascodeP[109],VcascodeP[108],VcascodeP[107],VcascodeP[106],VcascodeP[105],VcascodeP[104],VcascodeP[103],VcascodeP[102],VcascodeP[101],VcascodeP[100],VcascodeP[99],VcascodeP[98],VcascodeP[97],VcascodeP[96],VcascodeP[95],VcascodeP[94],VcascodeP[93],VcascodeP[92],VcascodeP[91],VcascodeP[90],VcascodeP[89],VcascodeP[88],VcascodeP[87],VcascodeP[86],VcascodeP[85],VcascodeP[84],VcascodeP[83],VcascodeP[82],VcascodeP[81],VcascodeP[80],VcascodeP[79],VcascodeP[78],VcascodeP[77],VcascodeP[76],VcascodeP[75],VcascodeP[74],VcascodeP[73],VcascodeP[72],VcascodeP[71],VcascodeP[70],VcascodeP[69],VcascodeP[68],VcascodeP[67],VcascodeP[66],VcascodeP[65],VcascodeP[64],VcascodeP[63],VcascodeP[62],VcascodeP[61],VcascodeP[60],VcascodeP[59],VcascodeP[58],VcascodeP[57],VcascodeP[56],VcascodeP[55],VcascodeP[54],VcascodeP[53],VcascodeP[52],VcascodeP[51],VcascodeP[50],VcascodeP[49],VcascodeP[48],VcascodeP[47],VcascodeP[46],VcascodeP[45],VcascodeP[44],VcascodeP[43],VcascodeP[42],VcascodeP[41],VcascodeP[40],VcascodeP[39],VcascodeP[38],VcascodeP[37],VcascodeP[36],VcascodeP[35],VcascodeP[34],VcascodeP[33],VcascodeP[32],VcascodeP[31],VcascodeP[30],VcascodeP[29],VcascodeP[28],VcascodeP[27],VcascodeP[26],VcascodeP[25],VcascodeP[24],VcascodeP[23],VcascodeP[22],VcascodeP[21],VcascodeP[20],VcascodeP[19],VcascodeP[18],VcascodeP[17],VcascodeP[16],VcascodeP[15],VcascodeP[14],VcascodeP[13],VcascodeP[12],VcascodeP[11],VcascodeP[10],VcascodeP[9],VcascodeP[8],VcascodeP[7],VcascodeP[6],VcascodeP[5],VcascodeP[4],VcascodeP[3],VcascodeP[2],VcascodeP[1],VcascodeP[0]
*.opin Iout
I_MIRROR[255] VDD Vbiasp VcascodeP[255] Iout Pmirror_StdCell
I_MIRROR[254] VDD Vbiasp VcascodeP[254] Iout Pmirror_StdCell
I_MIRROR[253] VDD Vbiasp VcascodeP[253] Iout Pmirror_StdCell
I_MIRROR[252] VDD Vbiasp VcascodeP[252] Iout Pmirror_StdCell
I_MIRROR[251] VDD Vbiasp VcascodeP[251] Iout Pmirror_StdCell
I_MIRROR[250] VDD Vbiasp VcascodeP[250] Iout Pmirror_StdCell
I_MIRROR[249] VDD Vbiasp VcascodeP[249] Iout Pmirror_StdCell
I_MIRROR[248] VDD Vbiasp VcascodeP[248] Iout Pmirror_StdCell
I_MIRROR[247] VDD Vbiasp VcascodeP[247] Iout Pmirror_StdCell
I_MIRROR[246] VDD Vbiasp VcascodeP[246] Iout Pmirror_StdCell
I_MIRROR[245] VDD Vbiasp VcascodeP[245] Iout Pmirror_StdCell
I_MIRROR[244] VDD Vbiasp VcascodeP[244] Iout Pmirror_StdCell
I_MIRROR[243] VDD Vbiasp VcascodeP[243] Iout Pmirror_StdCell
I_MIRROR[242] VDD Vbiasp VcascodeP[242] Iout Pmirror_StdCell
I_MIRROR[241] VDD Vbiasp VcascodeP[241] Iout Pmirror_StdCell
I_MIRROR[240] VDD Vbiasp VcascodeP[240] Iout Pmirror_StdCell
I_MIRROR[239] VDD Vbiasp VcascodeP[239] Iout Pmirror_StdCell
I_MIRROR[238] VDD Vbiasp VcascodeP[238] Iout Pmirror_StdCell
I_MIRROR[237] VDD Vbiasp VcascodeP[237] Iout Pmirror_StdCell
I_MIRROR[236] VDD Vbiasp VcascodeP[236] Iout Pmirror_StdCell
I_MIRROR[235] VDD Vbiasp VcascodeP[235] Iout Pmirror_StdCell
I_MIRROR[234] VDD Vbiasp VcascodeP[234] Iout Pmirror_StdCell
I_MIRROR[233] VDD Vbiasp VcascodeP[233] Iout Pmirror_StdCell
I_MIRROR[232] VDD Vbiasp VcascodeP[232] Iout Pmirror_StdCell
I_MIRROR[231] VDD Vbiasp VcascodeP[231] Iout Pmirror_StdCell
I_MIRROR[230] VDD Vbiasp VcascodeP[230] Iout Pmirror_StdCell
I_MIRROR[229] VDD Vbiasp VcascodeP[229] Iout Pmirror_StdCell
I_MIRROR[228] VDD Vbiasp VcascodeP[228] Iout Pmirror_StdCell
I_MIRROR[227] VDD Vbiasp VcascodeP[227] Iout Pmirror_StdCell
I_MIRROR[226] VDD Vbiasp VcascodeP[226] Iout Pmirror_StdCell
I_MIRROR[225] VDD Vbiasp VcascodeP[225] Iout Pmirror_StdCell
I_MIRROR[224] VDD Vbiasp VcascodeP[224] Iout Pmirror_StdCell
I_MIRROR[223] VDD Vbiasp VcascodeP[223] Iout Pmirror_StdCell
I_MIRROR[222] VDD Vbiasp VcascodeP[222] Iout Pmirror_StdCell
I_MIRROR[221] VDD Vbiasp VcascodeP[221] Iout Pmirror_StdCell
I_MIRROR[220] VDD Vbiasp VcascodeP[220] Iout Pmirror_StdCell
I_MIRROR[219] VDD Vbiasp VcascodeP[219] Iout Pmirror_StdCell
I_MIRROR[218] VDD Vbiasp VcascodeP[218] Iout Pmirror_StdCell
I_MIRROR[217] VDD Vbiasp VcascodeP[217] Iout Pmirror_StdCell
I_MIRROR[216] VDD Vbiasp VcascodeP[216] Iout Pmirror_StdCell
I_MIRROR[215] VDD Vbiasp VcascodeP[215] Iout Pmirror_StdCell
I_MIRROR[214] VDD Vbiasp VcascodeP[214] Iout Pmirror_StdCell
I_MIRROR[213] VDD Vbiasp VcascodeP[213] Iout Pmirror_StdCell
I_MIRROR[212] VDD Vbiasp VcascodeP[212] Iout Pmirror_StdCell
I_MIRROR[211] VDD Vbiasp VcascodeP[211] Iout Pmirror_StdCell
I_MIRROR[210] VDD Vbiasp VcascodeP[210] Iout Pmirror_StdCell
I_MIRROR[209] VDD Vbiasp VcascodeP[209] Iout Pmirror_StdCell
I_MIRROR[208] VDD Vbiasp VcascodeP[208] Iout Pmirror_StdCell
I_MIRROR[207] VDD Vbiasp VcascodeP[207] Iout Pmirror_StdCell
I_MIRROR[206] VDD Vbiasp VcascodeP[206] Iout Pmirror_StdCell
I_MIRROR[205] VDD Vbiasp VcascodeP[205] Iout Pmirror_StdCell
I_MIRROR[204] VDD Vbiasp VcascodeP[204] Iout Pmirror_StdCell
I_MIRROR[203] VDD Vbiasp VcascodeP[203] Iout Pmirror_StdCell
I_MIRROR[202] VDD Vbiasp VcascodeP[202] Iout Pmirror_StdCell
I_MIRROR[201] VDD Vbiasp VcascodeP[201] Iout Pmirror_StdCell
I_MIRROR[200] VDD Vbiasp VcascodeP[200] Iout Pmirror_StdCell
I_MIRROR[199] VDD Vbiasp VcascodeP[199] Iout Pmirror_StdCell
I_MIRROR[198] VDD Vbiasp VcascodeP[198] Iout Pmirror_StdCell
I_MIRROR[197] VDD Vbiasp VcascodeP[197] Iout Pmirror_StdCell
I_MIRROR[196] VDD Vbiasp VcascodeP[196] Iout Pmirror_StdCell
I_MIRROR[195] VDD Vbiasp VcascodeP[195] Iout Pmirror_StdCell
I_MIRROR[194] VDD Vbiasp VcascodeP[194] Iout Pmirror_StdCell
I_MIRROR[193] VDD Vbiasp VcascodeP[193] Iout Pmirror_StdCell
I_MIRROR[192] VDD Vbiasp VcascodeP[192] Iout Pmirror_StdCell
I_MIRROR[191] VDD Vbiasp VcascodeP[191] Iout Pmirror_StdCell
I_MIRROR[190] VDD Vbiasp VcascodeP[190] Iout Pmirror_StdCell
I_MIRROR[189] VDD Vbiasp VcascodeP[189] Iout Pmirror_StdCell
I_MIRROR[188] VDD Vbiasp VcascodeP[188] Iout Pmirror_StdCell
I_MIRROR[187] VDD Vbiasp VcascodeP[187] Iout Pmirror_StdCell
I_MIRROR[186] VDD Vbiasp VcascodeP[186] Iout Pmirror_StdCell
I_MIRROR[185] VDD Vbiasp VcascodeP[185] Iout Pmirror_StdCell
I_MIRROR[184] VDD Vbiasp VcascodeP[184] Iout Pmirror_StdCell
I_MIRROR[183] VDD Vbiasp VcascodeP[183] Iout Pmirror_StdCell
I_MIRROR[182] VDD Vbiasp VcascodeP[182] Iout Pmirror_StdCell
I_MIRROR[181] VDD Vbiasp VcascodeP[181] Iout Pmirror_StdCell
I_MIRROR[180] VDD Vbiasp VcascodeP[180] Iout Pmirror_StdCell
I_MIRROR[179] VDD Vbiasp VcascodeP[179] Iout Pmirror_StdCell
I_MIRROR[178] VDD Vbiasp VcascodeP[178] Iout Pmirror_StdCell
I_MIRROR[177] VDD Vbiasp VcascodeP[177] Iout Pmirror_StdCell
I_MIRROR[176] VDD Vbiasp VcascodeP[176] Iout Pmirror_StdCell
I_MIRROR[175] VDD Vbiasp VcascodeP[175] Iout Pmirror_StdCell
I_MIRROR[174] VDD Vbiasp VcascodeP[174] Iout Pmirror_StdCell
I_MIRROR[173] VDD Vbiasp VcascodeP[173] Iout Pmirror_StdCell
I_MIRROR[172] VDD Vbiasp VcascodeP[172] Iout Pmirror_StdCell
I_MIRROR[171] VDD Vbiasp VcascodeP[171] Iout Pmirror_StdCell
I_MIRROR[170] VDD Vbiasp VcascodeP[170] Iout Pmirror_StdCell
I_MIRROR[169] VDD Vbiasp VcascodeP[169] Iout Pmirror_StdCell
I_MIRROR[168] VDD Vbiasp VcascodeP[168] Iout Pmirror_StdCell
I_MIRROR[167] VDD Vbiasp VcascodeP[167] Iout Pmirror_StdCell
I_MIRROR[166] VDD Vbiasp VcascodeP[166] Iout Pmirror_StdCell
I_MIRROR[165] VDD Vbiasp VcascodeP[165] Iout Pmirror_StdCell
I_MIRROR[164] VDD Vbiasp VcascodeP[164] Iout Pmirror_StdCell
I_MIRROR[163] VDD Vbiasp VcascodeP[163] Iout Pmirror_StdCell
I_MIRROR[162] VDD Vbiasp VcascodeP[162] Iout Pmirror_StdCell
I_MIRROR[161] VDD Vbiasp VcascodeP[161] Iout Pmirror_StdCell
I_MIRROR[160] VDD Vbiasp VcascodeP[160] Iout Pmirror_StdCell
I_MIRROR[159] VDD Vbiasp VcascodeP[159] Iout Pmirror_StdCell
I_MIRROR[158] VDD Vbiasp VcascodeP[158] Iout Pmirror_StdCell
I_MIRROR[157] VDD Vbiasp VcascodeP[157] Iout Pmirror_StdCell
I_MIRROR[156] VDD Vbiasp VcascodeP[156] Iout Pmirror_StdCell
I_MIRROR[155] VDD Vbiasp VcascodeP[155] Iout Pmirror_StdCell
I_MIRROR[154] VDD Vbiasp VcascodeP[154] Iout Pmirror_StdCell
I_MIRROR[153] VDD Vbiasp VcascodeP[153] Iout Pmirror_StdCell
I_MIRROR[152] VDD Vbiasp VcascodeP[152] Iout Pmirror_StdCell
I_MIRROR[151] VDD Vbiasp VcascodeP[151] Iout Pmirror_StdCell
I_MIRROR[150] VDD Vbiasp VcascodeP[150] Iout Pmirror_StdCell
I_MIRROR[149] VDD Vbiasp VcascodeP[149] Iout Pmirror_StdCell
I_MIRROR[148] VDD Vbiasp VcascodeP[148] Iout Pmirror_StdCell
I_MIRROR[147] VDD Vbiasp VcascodeP[147] Iout Pmirror_StdCell
I_MIRROR[146] VDD Vbiasp VcascodeP[146] Iout Pmirror_StdCell
I_MIRROR[145] VDD Vbiasp VcascodeP[145] Iout Pmirror_StdCell
I_MIRROR[144] VDD Vbiasp VcascodeP[144] Iout Pmirror_StdCell
I_MIRROR[143] VDD Vbiasp VcascodeP[143] Iout Pmirror_StdCell
I_MIRROR[142] VDD Vbiasp VcascodeP[142] Iout Pmirror_StdCell
I_MIRROR[141] VDD Vbiasp VcascodeP[141] Iout Pmirror_StdCell
I_MIRROR[140] VDD Vbiasp VcascodeP[140] Iout Pmirror_StdCell
I_MIRROR[139] VDD Vbiasp VcascodeP[139] Iout Pmirror_StdCell
I_MIRROR[138] VDD Vbiasp VcascodeP[138] Iout Pmirror_StdCell
I_MIRROR[137] VDD Vbiasp VcascodeP[137] Iout Pmirror_StdCell
I_MIRROR[136] VDD Vbiasp VcascodeP[136] Iout Pmirror_StdCell
I_MIRROR[135] VDD Vbiasp VcascodeP[135] Iout Pmirror_StdCell
I_MIRROR[134] VDD Vbiasp VcascodeP[134] Iout Pmirror_StdCell
I_MIRROR[133] VDD Vbiasp VcascodeP[133] Iout Pmirror_StdCell
I_MIRROR[132] VDD Vbiasp VcascodeP[132] Iout Pmirror_StdCell
I_MIRROR[131] VDD Vbiasp VcascodeP[131] Iout Pmirror_StdCell
I_MIRROR[130] VDD Vbiasp VcascodeP[130] Iout Pmirror_StdCell
I_MIRROR[129] VDD Vbiasp VcascodeP[129] Iout Pmirror_StdCell
I_MIRROR[128] VDD Vbiasp VcascodeP[128] Iout Pmirror_StdCell
I_MIRROR[127] VDD Vbiasp VcascodeP[127] Iout Pmirror_StdCell
I_MIRROR[126] VDD Vbiasp VcascodeP[126] Iout Pmirror_StdCell
I_MIRROR[125] VDD Vbiasp VcascodeP[125] Iout Pmirror_StdCell
I_MIRROR[124] VDD Vbiasp VcascodeP[124] Iout Pmirror_StdCell
I_MIRROR[123] VDD Vbiasp VcascodeP[123] Iout Pmirror_StdCell
I_MIRROR[122] VDD Vbiasp VcascodeP[122] Iout Pmirror_StdCell
I_MIRROR[121] VDD Vbiasp VcascodeP[121] Iout Pmirror_StdCell
I_MIRROR[120] VDD Vbiasp VcascodeP[120] Iout Pmirror_StdCell
I_MIRROR[119] VDD Vbiasp VcascodeP[119] Iout Pmirror_StdCell
I_MIRROR[118] VDD Vbiasp VcascodeP[118] Iout Pmirror_StdCell
I_MIRROR[117] VDD Vbiasp VcascodeP[117] Iout Pmirror_StdCell
I_MIRROR[116] VDD Vbiasp VcascodeP[116] Iout Pmirror_StdCell
I_MIRROR[115] VDD Vbiasp VcascodeP[115] Iout Pmirror_StdCell
I_MIRROR[114] VDD Vbiasp VcascodeP[114] Iout Pmirror_StdCell
I_MIRROR[113] VDD Vbiasp VcascodeP[113] Iout Pmirror_StdCell
I_MIRROR[112] VDD Vbiasp VcascodeP[112] Iout Pmirror_StdCell
I_MIRROR[111] VDD Vbiasp VcascodeP[111] Iout Pmirror_StdCell
I_MIRROR[110] VDD Vbiasp VcascodeP[110] Iout Pmirror_StdCell
I_MIRROR[109] VDD Vbiasp VcascodeP[109] Iout Pmirror_StdCell
I_MIRROR[108] VDD Vbiasp VcascodeP[108] Iout Pmirror_StdCell
I_MIRROR[107] VDD Vbiasp VcascodeP[107] Iout Pmirror_StdCell
I_MIRROR[106] VDD Vbiasp VcascodeP[106] Iout Pmirror_StdCell
I_MIRROR[105] VDD Vbiasp VcascodeP[105] Iout Pmirror_StdCell
I_MIRROR[104] VDD Vbiasp VcascodeP[104] Iout Pmirror_StdCell
I_MIRROR[103] VDD Vbiasp VcascodeP[103] Iout Pmirror_StdCell
I_MIRROR[102] VDD Vbiasp VcascodeP[102] Iout Pmirror_StdCell
I_MIRROR[101] VDD Vbiasp VcascodeP[101] Iout Pmirror_StdCell
I_MIRROR[100] VDD Vbiasp VcascodeP[100] Iout Pmirror_StdCell
I_MIRROR[99] VDD Vbiasp VcascodeP[99] Iout Pmirror_StdCell
I_MIRROR[98] VDD Vbiasp VcascodeP[98] Iout Pmirror_StdCell
I_MIRROR[97] VDD Vbiasp VcascodeP[97] Iout Pmirror_StdCell
I_MIRROR[96] VDD Vbiasp VcascodeP[96] Iout Pmirror_StdCell
I_MIRROR[95] VDD Vbiasp VcascodeP[95] Iout Pmirror_StdCell
I_MIRROR[94] VDD Vbiasp VcascodeP[94] Iout Pmirror_StdCell
I_MIRROR[93] VDD Vbiasp VcascodeP[93] Iout Pmirror_StdCell
I_MIRROR[92] VDD Vbiasp VcascodeP[92] Iout Pmirror_StdCell
I_MIRROR[91] VDD Vbiasp VcascodeP[91] Iout Pmirror_StdCell
I_MIRROR[90] VDD Vbiasp VcascodeP[90] Iout Pmirror_StdCell
I_MIRROR[89] VDD Vbiasp VcascodeP[89] Iout Pmirror_StdCell
I_MIRROR[88] VDD Vbiasp VcascodeP[88] Iout Pmirror_StdCell
I_MIRROR[87] VDD Vbiasp VcascodeP[87] Iout Pmirror_StdCell
I_MIRROR[86] VDD Vbiasp VcascodeP[86] Iout Pmirror_StdCell
I_MIRROR[85] VDD Vbiasp VcascodeP[85] Iout Pmirror_StdCell
I_MIRROR[84] VDD Vbiasp VcascodeP[84] Iout Pmirror_StdCell
I_MIRROR[83] VDD Vbiasp VcascodeP[83] Iout Pmirror_StdCell
I_MIRROR[82] VDD Vbiasp VcascodeP[82] Iout Pmirror_StdCell
I_MIRROR[81] VDD Vbiasp VcascodeP[81] Iout Pmirror_StdCell
I_MIRROR[80] VDD Vbiasp VcascodeP[80] Iout Pmirror_StdCell
I_MIRROR[79] VDD Vbiasp VcascodeP[79] Iout Pmirror_StdCell
I_MIRROR[78] VDD Vbiasp VcascodeP[78] Iout Pmirror_StdCell
I_MIRROR[77] VDD Vbiasp VcascodeP[77] Iout Pmirror_StdCell
I_MIRROR[76] VDD Vbiasp VcascodeP[76] Iout Pmirror_StdCell
I_MIRROR[75] VDD Vbiasp VcascodeP[75] Iout Pmirror_StdCell
I_MIRROR[74] VDD Vbiasp VcascodeP[74] Iout Pmirror_StdCell
I_MIRROR[73] VDD Vbiasp VcascodeP[73] Iout Pmirror_StdCell
I_MIRROR[72] VDD Vbiasp VcascodeP[72] Iout Pmirror_StdCell
I_MIRROR[71] VDD Vbiasp VcascodeP[71] Iout Pmirror_StdCell
I_MIRROR[70] VDD Vbiasp VcascodeP[70] Iout Pmirror_StdCell
I_MIRROR[69] VDD Vbiasp VcascodeP[69] Iout Pmirror_StdCell
I_MIRROR[68] VDD Vbiasp VcascodeP[68] Iout Pmirror_StdCell
I_MIRROR[67] VDD Vbiasp VcascodeP[67] Iout Pmirror_StdCell
I_MIRROR[66] VDD Vbiasp VcascodeP[66] Iout Pmirror_StdCell
I_MIRROR[65] VDD Vbiasp VcascodeP[65] Iout Pmirror_StdCell
I_MIRROR[64] VDD Vbiasp VcascodeP[64] Iout Pmirror_StdCell
I_MIRROR[63] VDD Vbiasp VcascodeP[63] Iout Pmirror_StdCell
I_MIRROR[62] VDD Vbiasp VcascodeP[62] Iout Pmirror_StdCell
I_MIRROR[61] VDD Vbiasp VcascodeP[61] Iout Pmirror_StdCell
I_MIRROR[60] VDD Vbiasp VcascodeP[60] Iout Pmirror_StdCell
I_MIRROR[59] VDD Vbiasp VcascodeP[59] Iout Pmirror_StdCell
I_MIRROR[58] VDD Vbiasp VcascodeP[58] Iout Pmirror_StdCell
I_MIRROR[57] VDD Vbiasp VcascodeP[57] Iout Pmirror_StdCell
I_MIRROR[56] VDD Vbiasp VcascodeP[56] Iout Pmirror_StdCell
I_MIRROR[55] VDD Vbiasp VcascodeP[55] Iout Pmirror_StdCell
I_MIRROR[54] VDD Vbiasp VcascodeP[54] Iout Pmirror_StdCell
I_MIRROR[53] VDD Vbiasp VcascodeP[53] Iout Pmirror_StdCell
I_MIRROR[52] VDD Vbiasp VcascodeP[52] Iout Pmirror_StdCell
I_MIRROR[51] VDD Vbiasp VcascodeP[51] Iout Pmirror_StdCell
I_MIRROR[50] VDD Vbiasp VcascodeP[50] Iout Pmirror_StdCell
I_MIRROR[49] VDD Vbiasp VcascodeP[49] Iout Pmirror_StdCell
I_MIRROR[48] VDD Vbiasp VcascodeP[48] Iout Pmirror_StdCell
I_MIRROR[47] VDD Vbiasp VcascodeP[47] Iout Pmirror_StdCell
I_MIRROR[46] VDD Vbiasp VcascodeP[46] Iout Pmirror_StdCell
I_MIRROR[45] VDD Vbiasp VcascodeP[45] Iout Pmirror_StdCell
I_MIRROR[44] VDD Vbiasp VcascodeP[44] Iout Pmirror_StdCell
I_MIRROR[43] VDD Vbiasp VcascodeP[43] Iout Pmirror_StdCell
I_MIRROR[42] VDD Vbiasp VcascodeP[42] Iout Pmirror_StdCell
I_MIRROR[41] VDD Vbiasp VcascodeP[41] Iout Pmirror_StdCell
I_MIRROR[40] VDD Vbiasp VcascodeP[40] Iout Pmirror_StdCell
I_MIRROR[39] VDD Vbiasp VcascodeP[39] Iout Pmirror_StdCell
I_MIRROR[38] VDD Vbiasp VcascodeP[38] Iout Pmirror_StdCell
I_MIRROR[37] VDD Vbiasp VcascodeP[37] Iout Pmirror_StdCell
I_MIRROR[36] VDD Vbiasp VcascodeP[36] Iout Pmirror_StdCell
I_MIRROR[35] VDD Vbiasp VcascodeP[35] Iout Pmirror_StdCell
I_MIRROR[34] VDD Vbiasp VcascodeP[34] Iout Pmirror_StdCell
I_MIRROR[33] VDD Vbiasp VcascodeP[33] Iout Pmirror_StdCell
I_MIRROR[32] VDD Vbiasp VcascodeP[32] Iout Pmirror_StdCell
I_MIRROR[31] VDD Vbiasp VcascodeP[31] Iout Pmirror_StdCell
I_MIRROR[30] VDD Vbiasp VcascodeP[30] Iout Pmirror_StdCell
I_MIRROR[29] VDD Vbiasp VcascodeP[29] Iout Pmirror_StdCell
I_MIRROR[28] VDD Vbiasp VcascodeP[28] Iout Pmirror_StdCell
I_MIRROR[27] VDD Vbiasp VcascodeP[27] Iout Pmirror_StdCell
I_MIRROR[26] VDD Vbiasp VcascodeP[26] Iout Pmirror_StdCell
I_MIRROR[25] VDD Vbiasp VcascodeP[25] Iout Pmirror_StdCell
I_MIRROR[24] VDD Vbiasp VcascodeP[24] Iout Pmirror_StdCell
I_MIRROR[23] VDD Vbiasp VcascodeP[23] Iout Pmirror_StdCell
I_MIRROR[22] VDD Vbiasp VcascodeP[22] Iout Pmirror_StdCell
I_MIRROR[21] VDD Vbiasp VcascodeP[21] Iout Pmirror_StdCell
I_MIRROR[20] VDD Vbiasp VcascodeP[20] Iout Pmirror_StdCell
I_MIRROR[19] VDD Vbiasp VcascodeP[19] Iout Pmirror_StdCell
I_MIRROR[18] VDD Vbiasp VcascodeP[18] Iout Pmirror_StdCell
I_MIRROR[17] VDD Vbiasp VcascodeP[17] Iout Pmirror_StdCell
I_MIRROR[16] VDD Vbiasp VcascodeP[16] Iout Pmirror_StdCell
I_MIRROR[15] VDD Vbiasp VcascodeP[15] Iout Pmirror_StdCell
I_MIRROR[14] VDD Vbiasp VcascodeP[14] Iout Pmirror_StdCell
I_MIRROR[13] VDD Vbiasp VcascodeP[13] Iout Pmirror_StdCell
I_MIRROR[12] VDD Vbiasp VcascodeP[12] Iout Pmirror_StdCell
I_MIRROR[11] VDD Vbiasp VcascodeP[11] Iout Pmirror_StdCell
I_MIRROR[10] VDD Vbiasp VcascodeP[10] Iout Pmirror_StdCell
I_MIRROR[9] VDD Vbiasp VcascodeP[9] Iout Pmirror_StdCell
I_MIRROR[8] VDD Vbiasp VcascodeP[8] Iout Pmirror_StdCell
I_MIRROR[7] VDD Vbiasp VcascodeP[7] Iout Pmirror_StdCell
I_MIRROR[6] VDD Vbiasp VcascodeP[6] Iout Pmirror_StdCell
I_MIRROR[5] VDD Vbiasp VcascodeP[5] Iout Pmirror_StdCell
I_MIRROR[4] VDD Vbiasp VcascodeP[4] Iout Pmirror_StdCell
I_MIRROR[3] VDD Vbiasp VcascodeP[3] Iout Pmirror_StdCell
I_MIRROR[2] VDD Vbiasp VcascodeP[2] Iout Pmirror_StdCell
I_MIRROR[1] VDD Vbiasp VcascodeP[1] Iout Pmirror_StdCell
I_MIRROR[0] VDD Vbiasp VcascodeP[0] Iout Pmirror_StdCell
.ends


* expanding   symbol:  /home/user/PUDDING/schematic/DAC_SW.sym # of pins=5
** sym_path: /home/user/PUDDING/schematic/DAC_SW.sym
** sch_path: /home/user/PUDDING/schematic/DAC_SW.sch
.subckt DAC_SW VDD ON Pcascode_sw Pcascode ESDGND
*.ipin ON
*.ipin Pcascode
*.ipin ESDGND
*.ipin VDD
*.opin Pcascode_sw
XM1 VDD ON Pcascode_sw VDD sg13_lv_pmos w=0.5u l=0.13u ng=1 m=1
XM2 net1 ON VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 Pcascode net1 Pcascode_sw VDD sg13_lv_pmos w=0.5u l=0.13u ng=1 m=1
XM4 net1 ON ESDGND ESDGND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/user/PUDDING/schematic/Pmirror_StdCell.sym # of pins=4
** sym_path: /home/user/PUDDING/schematic/Pmirror_StdCell.sym
** sch_path: /home/user/PUDDING/schematic/Pmirror_StdCell.sch
.subckt Pmirror_StdCell VDD VbiasP VcascodeP Iout
*.ipin VcascodeP
*.ipin VbiasP
*.opin Iout
*.ipin VDD
XM2 net1 VbiasP VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 Iout VcascodeP net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
