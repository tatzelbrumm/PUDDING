VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO analog_wires
  CLASS BLOCK ;
  ORIGIN 0.35 0.35 ;
  SIZE 100.35 BY 200.35 ;
  SYMMETRY X Y R90 ;
END analog_wires

END LIBRARY
