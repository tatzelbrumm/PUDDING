magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771125512
<< nwell >>
rect -124 -124 6660 6524
<< hvpmos >>
rect 68 0 6468 6400
<< hvpdiff >>
rect 0 6386 68 6400
rect 0 6354 14 6386
rect 46 6354 68 6386
rect 0 6317 68 6354
rect 0 6285 14 6317
rect 46 6285 68 6317
rect 0 6249 68 6285
rect 0 6217 14 6249
rect 46 6217 68 6249
rect 0 6181 68 6217
rect 0 6149 14 6181
rect 46 6149 68 6181
rect 0 6113 68 6149
rect 0 6081 14 6113
rect 46 6081 68 6113
rect 0 6045 68 6081
rect 0 6013 14 6045
rect 46 6013 68 6045
rect 0 5976 68 6013
rect 0 5944 14 5976
rect 46 5944 68 5976
rect 0 5908 68 5944
rect 0 5876 14 5908
rect 46 5876 68 5908
rect 0 5840 68 5876
rect 0 5808 14 5840
rect 46 5808 68 5840
rect 0 5772 68 5808
rect 0 5740 14 5772
rect 46 5740 68 5772
rect 0 5704 68 5740
rect 0 5672 14 5704
rect 46 5672 68 5704
rect 0 5636 68 5672
rect 0 5604 14 5636
rect 46 5604 68 5636
rect 0 5567 68 5604
rect 0 5535 14 5567
rect 46 5535 68 5567
rect 0 5499 68 5535
rect 0 5467 14 5499
rect 46 5467 68 5499
rect 0 5431 68 5467
rect 0 5399 14 5431
rect 46 5399 68 5431
rect 0 5363 68 5399
rect 0 5331 14 5363
rect 46 5331 68 5363
rect 0 5295 68 5331
rect 0 5263 14 5295
rect 46 5263 68 5295
rect 0 5227 68 5263
rect 0 5195 14 5227
rect 46 5195 68 5227
rect 0 5158 68 5195
rect 0 5126 14 5158
rect 46 5126 68 5158
rect 0 5090 68 5126
rect 0 5058 14 5090
rect 46 5058 68 5090
rect 0 5022 68 5058
rect 0 4990 14 5022
rect 46 4990 68 5022
rect 0 4954 68 4990
rect 0 4922 14 4954
rect 46 4922 68 4954
rect 0 4886 68 4922
rect 0 4854 14 4886
rect 46 4854 68 4886
rect 0 4818 68 4854
rect 0 4786 14 4818
rect 46 4786 68 4818
rect 0 4749 68 4786
rect 0 4717 14 4749
rect 46 4717 68 4749
rect 0 4681 68 4717
rect 0 4649 14 4681
rect 46 4649 68 4681
rect 0 4613 68 4649
rect 0 4581 14 4613
rect 46 4581 68 4613
rect 0 4545 68 4581
rect 0 4513 14 4545
rect 46 4513 68 4545
rect 0 4477 68 4513
rect 0 4445 14 4477
rect 46 4445 68 4477
rect 0 4409 68 4445
rect 0 4377 14 4409
rect 46 4377 68 4409
rect 0 4340 68 4377
rect 0 4308 14 4340
rect 46 4308 68 4340
rect 0 4272 68 4308
rect 0 4240 14 4272
rect 46 4240 68 4272
rect 0 4204 68 4240
rect 0 4172 14 4204
rect 46 4172 68 4204
rect 0 4136 68 4172
rect 0 4104 14 4136
rect 46 4104 68 4136
rect 0 4068 68 4104
rect 0 4036 14 4068
rect 46 4036 68 4068
rect 0 3999 68 4036
rect 0 3967 14 3999
rect 46 3967 68 3999
rect 0 3931 68 3967
rect 0 3899 14 3931
rect 46 3899 68 3931
rect 0 3863 68 3899
rect 0 3831 14 3863
rect 46 3831 68 3863
rect 0 3795 68 3831
rect 0 3763 14 3795
rect 46 3763 68 3795
rect 0 3727 68 3763
rect 0 3695 14 3727
rect 46 3695 68 3727
rect 0 3659 68 3695
rect 0 3627 14 3659
rect 46 3627 68 3659
rect 0 3590 68 3627
rect 0 3558 14 3590
rect 46 3558 68 3590
rect 0 3522 68 3558
rect 0 3490 14 3522
rect 46 3490 68 3522
rect 0 3454 68 3490
rect 0 3422 14 3454
rect 46 3422 68 3454
rect 0 3386 68 3422
rect 0 3354 14 3386
rect 46 3354 68 3386
rect 0 3318 68 3354
rect 0 3286 14 3318
rect 46 3286 68 3318
rect 0 3250 68 3286
rect 0 3218 14 3250
rect 46 3218 68 3250
rect 0 3181 68 3218
rect 0 3149 14 3181
rect 46 3149 68 3181
rect 0 3113 68 3149
rect 0 3081 14 3113
rect 46 3081 68 3113
rect 0 3045 68 3081
rect 0 3013 14 3045
rect 46 3013 68 3045
rect 0 2977 68 3013
rect 0 2945 14 2977
rect 46 2945 68 2977
rect 0 2909 68 2945
rect 0 2877 14 2909
rect 46 2877 68 2909
rect 0 2841 68 2877
rect 0 2809 14 2841
rect 46 2809 68 2841
rect 0 2772 68 2809
rect 0 2740 14 2772
rect 46 2740 68 2772
rect 0 2704 68 2740
rect 0 2672 14 2704
rect 46 2672 68 2704
rect 0 2636 68 2672
rect 0 2604 14 2636
rect 46 2604 68 2636
rect 0 2568 68 2604
rect 0 2536 14 2568
rect 46 2536 68 2568
rect 0 2500 68 2536
rect 0 2468 14 2500
rect 46 2468 68 2500
rect 0 2432 68 2468
rect 0 2400 14 2432
rect 46 2400 68 2432
rect 0 2363 68 2400
rect 0 2331 14 2363
rect 46 2331 68 2363
rect 0 2295 68 2331
rect 0 2263 14 2295
rect 46 2263 68 2295
rect 0 2227 68 2263
rect 0 2195 14 2227
rect 46 2195 68 2227
rect 0 2159 68 2195
rect 0 2127 14 2159
rect 46 2127 68 2159
rect 0 2091 68 2127
rect 0 2059 14 2091
rect 46 2059 68 2091
rect 0 2022 68 2059
rect 0 1990 14 2022
rect 46 1990 68 2022
rect 0 1954 68 1990
rect 0 1922 14 1954
rect 46 1922 68 1954
rect 0 1886 68 1922
rect 0 1854 14 1886
rect 46 1854 68 1886
rect 0 1818 68 1854
rect 0 1786 14 1818
rect 46 1786 68 1818
rect 0 1750 68 1786
rect 0 1718 14 1750
rect 46 1718 68 1750
rect 0 1682 68 1718
rect 0 1650 14 1682
rect 46 1650 68 1682
rect 0 1613 68 1650
rect 0 1581 14 1613
rect 46 1581 68 1613
rect 0 1545 68 1581
rect 0 1513 14 1545
rect 46 1513 68 1545
rect 0 1477 68 1513
rect 0 1445 14 1477
rect 46 1445 68 1477
rect 0 1409 68 1445
rect 0 1377 14 1409
rect 46 1377 68 1409
rect 0 1341 68 1377
rect 0 1309 14 1341
rect 46 1309 68 1341
rect 0 1273 68 1309
rect 0 1241 14 1273
rect 46 1241 68 1273
rect 0 1204 68 1241
rect 0 1172 14 1204
rect 46 1172 68 1204
rect 0 1136 68 1172
rect 0 1104 14 1136
rect 46 1104 68 1136
rect 0 1068 68 1104
rect 0 1036 14 1068
rect 46 1036 68 1068
rect 0 1000 68 1036
rect 0 968 14 1000
rect 46 968 68 1000
rect 0 932 68 968
rect 0 900 14 932
rect 46 900 68 932
rect 0 864 68 900
rect 0 832 14 864
rect 46 832 68 864
rect 0 795 68 832
rect 0 763 14 795
rect 46 763 68 795
rect 0 727 68 763
rect 0 695 14 727
rect 46 695 68 727
rect 0 659 68 695
rect 0 627 14 659
rect 46 627 68 659
rect 0 591 68 627
rect 0 559 14 591
rect 46 559 68 591
rect 0 523 68 559
rect 0 491 14 523
rect 46 491 68 523
rect 0 455 68 491
rect 0 423 14 455
rect 46 423 68 455
rect 0 386 68 423
rect 0 354 14 386
rect 46 354 68 386
rect 0 318 68 354
rect 0 286 14 318
rect 46 286 68 318
rect 0 250 68 286
rect 0 218 14 250
rect 46 218 68 250
rect 0 182 68 218
rect 0 150 14 182
rect 46 150 68 182
rect 0 114 68 150
rect 0 82 14 114
rect 46 82 68 114
rect 0 46 68 82
rect 0 14 14 46
rect 46 14 68 46
rect 0 0 68 14
rect 6468 6386 6536 6400
rect 6468 6354 6490 6386
rect 6522 6354 6536 6386
rect 6468 6317 6536 6354
rect 6468 6285 6490 6317
rect 6522 6285 6536 6317
rect 6468 6249 6536 6285
rect 6468 6217 6490 6249
rect 6522 6217 6536 6249
rect 6468 6181 6536 6217
rect 6468 6149 6490 6181
rect 6522 6149 6536 6181
rect 6468 6113 6536 6149
rect 6468 6081 6490 6113
rect 6522 6081 6536 6113
rect 6468 6045 6536 6081
rect 6468 6013 6490 6045
rect 6522 6013 6536 6045
rect 6468 5976 6536 6013
rect 6468 5944 6490 5976
rect 6522 5944 6536 5976
rect 6468 5908 6536 5944
rect 6468 5876 6490 5908
rect 6522 5876 6536 5908
rect 6468 5840 6536 5876
rect 6468 5808 6490 5840
rect 6522 5808 6536 5840
rect 6468 5772 6536 5808
rect 6468 5740 6490 5772
rect 6522 5740 6536 5772
rect 6468 5704 6536 5740
rect 6468 5672 6490 5704
rect 6522 5672 6536 5704
rect 6468 5636 6536 5672
rect 6468 5604 6490 5636
rect 6522 5604 6536 5636
rect 6468 5567 6536 5604
rect 6468 5535 6490 5567
rect 6522 5535 6536 5567
rect 6468 5499 6536 5535
rect 6468 5467 6490 5499
rect 6522 5467 6536 5499
rect 6468 5431 6536 5467
rect 6468 5399 6490 5431
rect 6522 5399 6536 5431
rect 6468 5363 6536 5399
rect 6468 5331 6490 5363
rect 6522 5331 6536 5363
rect 6468 5295 6536 5331
rect 6468 5263 6490 5295
rect 6522 5263 6536 5295
rect 6468 5227 6536 5263
rect 6468 5195 6490 5227
rect 6522 5195 6536 5227
rect 6468 5158 6536 5195
rect 6468 5126 6490 5158
rect 6522 5126 6536 5158
rect 6468 5090 6536 5126
rect 6468 5058 6490 5090
rect 6522 5058 6536 5090
rect 6468 5022 6536 5058
rect 6468 4990 6490 5022
rect 6522 4990 6536 5022
rect 6468 4954 6536 4990
rect 6468 4922 6490 4954
rect 6522 4922 6536 4954
rect 6468 4886 6536 4922
rect 6468 4854 6490 4886
rect 6522 4854 6536 4886
rect 6468 4818 6536 4854
rect 6468 4786 6490 4818
rect 6522 4786 6536 4818
rect 6468 4749 6536 4786
rect 6468 4717 6490 4749
rect 6522 4717 6536 4749
rect 6468 4681 6536 4717
rect 6468 4649 6490 4681
rect 6522 4649 6536 4681
rect 6468 4613 6536 4649
rect 6468 4581 6490 4613
rect 6522 4581 6536 4613
rect 6468 4545 6536 4581
rect 6468 4513 6490 4545
rect 6522 4513 6536 4545
rect 6468 4477 6536 4513
rect 6468 4445 6490 4477
rect 6522 4445 6536 4477
rect 6468 4409 6536 4445
rect 6468 4377 6490 4409
rect 6522 4377 6536 4409
rect 6468 4340 6536 4377
rect 6468 4308 6490 4340
rect 6522 4308 6536 4340
rect 6468 4272 6536 4308
rect 6468 4240 6490 4272
rect 6522 4240 6536 4272
rect 6468 4204 6536 4240
rect 6468 4172 6490 4204
rect 6522 4172 6536 4204
rect 6468 4136 6536 4172
rect 6468 4104 6490 4136
rect 6522 4104 6536 4136
rect 6468 4068 6536 4104
rect 6468 4036 6490 4068
rect 6522 4036 6536 4068
rect 6468 3999 6536 4036
rect 6468 3967 6490 3999
rect 6522 3967 6536 3999
rect 6468 3931 6536 3967
rect 6468 3899 6490 3931
rect 6522 3899 6536 3931
rect 6468 3863 6536 3899
rect 6468 3831 6490 3863
rect 6522 3831 6536 3863
rect 6468 3795 6536 3831
rect 6468 3763 6490 3795
rect 6522 3763 6536 3795
rect 6468 3727 6536 3763
rect 6468 3695 6490 3727
rect 6522 3695 6536 3727
rect 6468 3659 6536 3695
rect 6468 3627 6490 3659
rect 6522 3627 6536 3659
rect 6468 3590 6536 3627
rect 6468 3558 6490 3590
rect 6522 3558 6536 3590
rect 6468 3522 6536 3558
rect 6468 3490 6490 3522
rect 6522 3490 6536 3522
rect 6468 3454 6536 3490
rect 6468 3422 6490 3454
rect 6522 3422 6536 3454
rect 6468 3386 6536 3422
rect 6468 3354 6490 3386
rect 6522 3354 6536 3386
rect 6468 3318 6536 3354
rect 6468 3286 6490 3318
rect 6522 3286 6536 3318
rect 6468 3250 6536 3286
rect 6468 3218 6490 3250
rect 6522 3218 6536 3250
rect 6468 3181 6536 3218
rect 6468 3149 6490 3181
rect 6522 3149 6536 3181
rect 6468 3113 6536 3149
rect 6468 3081 6490 3113
rect 6522 3081 6536 3113
rect 6468 3045 6536 3081
rect 6468 3013 6490 3045
rect 6522 3013 6536 3045
rect 6468 2977 6536 3013
rect 6468 2945 6490 2977
rect 6522 2945 6536 2977
rect 6468 2909 6536 2945
rect 6468 2877 6490 2909
rect 6522 2877 6536 2909
rect 6468 2841 6536 2877
rect 6468 2809 6490 2841
rect 6522 2809 6536 2841
rect 6468 2772 6536 2809
rect 6468 2740 6490 2772
rect 6522 2740 6536 2772
rect 6468 2704 6536 2740
rect 6468 2672 6490 2704
rect 6522 2672 6536 2704
rect 6468 2636 6536 2672
rect 6468 2604 6490 2636
rect 6522 2604 6536 2636
rect 6468 2568 6536 2604
rect 6468 2536 6490 2568
rect 6522 2536 6536 2568
rect 6468 2500 6536 2536
rect 6468 2468 6490 2500
rect 6522 2468 6536 2500
rect 6468 2432 6536 2468
rect 6468 2400 6490 2432
rect 6522 2400 6536 2432
rect 6468 2363 6536 2400
rect 6468 2331 6490 2363
rect 6522 2331 6536 2363
rect 6468 2295 6536 2331
rect 6468 2263 6490 2295
rect 6522 2263 6536 2295
rect 6468 2227 6536 2263
rect 6468 2195 6490 2227
rect 6522 2195 6536 2227
rect 6468 2159 6536 2195
rect 6468 2127 6490 2159
rect 6522 2127 6536 2159
rect 6468 2091 6536 2127
rect 6468 2059 6490 2091
rect 6522 2059 6536 2091
rect 6468 2022 6536 2059
rect 6468 1990 6490 2022
rect 6522 1990 6536 2022
rect 6468 1954 6536 1990
rect 6468 1922 6490 1954
rect 6522 1922 6536 1954
rect 6468 1886 6536 1922
rect 6468 1854 6490 1886
rect 6522 1854 6536 1886
rect 6468 1818 6536 1854
rect 6468 1786 6490 1818
rect 6522 1786 6536 1818
rect 6468 1750 6536 1786
rect 6468 1718 6490 1750
rect 6522 1718 6536 1750
rect 6468 1682 6536 1718
rect 6468 1650 6490 1682
rect 6522 1650 6536 1682
rect 6468 1613 6536 1650
rect 6468 1581 6490 1613
rect 6522 1581 6536 1613
rect 6468 1545 6536 1581
rect 6468 1513 6490 1545
rect 6522 1513 6536 1545
rect 6468 1477 6536 1513
rect 6468 1445 6490 1477
rect 6522 1445 6536 1477
rect 6468 1409 6536 1445
rect 6468 1377 6490 1409
rect 6522 1377 6536 1409
rect 6468 1341 6536 1377
rect 6468 1309 6490 1341
rect 6522 1309 6536 1341
rect 6468 1273 6536 1309
rect 6468 1241 6490 1273
rect 6522 1241 6536 1273
rect 6468 1204 6536 1241
rect 6468 1172 6490 1204
rect 6522 1172 6536 1204
rect 6468 1136 6536 1172
rect 6468 1104 6490 1136
rect 6522 1104 6536 1136
rect 6468 1068 6536 1104
rect 6468 1036 6490 1068
rect 6522 1036 6536 1068
rect 6468 1000 6536 1036
rect 6468 968 6490 1000
rect 6522 968 6536 1000
rect 6468 932 6536 968
rect 6468 900 6490 932
rect 6522 900 6536 932
rect 6468 864 6536 900
rect 6468 832 6490 864
rect 6522 832 6536 864
rect 6468 795 6536 832
rect 6468 763 6490 795
rect 6522 763 6536 795
rect 6468 727 6536 763
rect 6468 695 6490 727
rect 6522 695 6536 727
rect 6468 659 6536 695
rect 6468 627 6490 659
rect 6522 627 6536 659
rect 6468 591 6536 627
rect 6468 559 6490 591
rect 6522 559 6536 591
rect 6468 523 6536 559
rect 6468 491 6490 523
rect 6522 491 6536 523
rect 6468 455 6536 491
rect 6468 423 6490 455
rect 6522 423 6536 455
rect 6468 386 6536 423
rect 6468 354 6490 386
rect 6522 354 6536 386
rect 6468 318 6536 354
rect 6468 286 6490 318
rect 6522 286 6536 318
rect 6468 250 6536 286
rect 6468 218 6490 250
rect 6522 218 6536 250
rect 6468 182 6536 218
rect 6468 150 6490 182
rect 6522 150 6536 182
rect 6468 114 6536 150
rect 6468 82 6490 114
rect 6522 82 6536 114
rect 6468 46 6536 82
rect 6468 14 6490 46
rect 6522 14 6536 46
rect 6468 0 6536 14
<< hvpdiffc >>
rect 14 6354 46 6386
rect 14 6285 46 6317
rect 14 6217 46 6249
rect 14 6149 46 6181
rect 14 6081 46 6113
rect 14 6013 46 6045
rect 14 5944 46 5976
rect 14 5876 46 5908
rect 14 5808 46 5840
rect 14 5740 46 5772
rect 14 5672 46 5704
rect 14 5604 46 5636
rect 14 5535 46 5567
rect 14 5467 46 5499
rect 14 5399 46 5431
rect 14 5331 46 5363
rect 14 5263 46 5295
rect 14 5195 46 5227
rect 14 5126 46 5158
rect 14 5058 46 5090
rect 14 4990 46 5022
rect 14 4922 46 4954
rect 14 4854 46 4886
rect 14 4786 46 4818
rect 14 4717 46 4749
rect 14 4649 46 4681
rect 14 4581 46 4613
rect 14 4513 46 4545
rect 14 4445 46 4477
rect 14 4377 46 4409
rect 14 4308 46 4340
rect 14 4240 46 4272
rect 14 4172 46 4204
rect 14 4104 46 4136
rect 14 4036 46 4068
rect 14 3967 46 3999
rect 14 3899 46 3931
rect 14 3831 46 3863
rect 14 3763 46 3795
rect 14 3695 46 3727
rect 14 3627 46 3659
rect 14 3558 46 3590
rect 14 3490 46 3522
rect 14 3422 46 3454
rect 14 3354 46 3386
rect 14 3286 46 3318
rect 14 3218 46 3250
rect 14 3149 46 3181
rect 14 3081 46 3113
rect 14 3013 46 3045
rect 14 2945 46 2977
rect 14 2877 46 2909
rect 14 2809 46 2841
rect 14 2740 46 2772
rect 14 2672 46 2704
rect 14 2604 46 2636
rect 14 2536 46 2568
rect 14 2468 46 2500
rect 14 2400 46 2432
rect 14 2331 46 2363
rect 14 2263 46 2295
rect 14 2195 46 2227
rect 14 2127 46 2159
rect 14 2059 46 2091
rect 14 1990 46 2022
rect 14 1922 46 1954
rect 14 1854 46 1886
rect 14 1786 46 1818
rect 14 1718 46 1750
rect 14 1650 46 1682
rect 14 1581 46 1613
rect 14 1513 46 1545
rect 14 1445 46 1477
rect 14 1377 46 1409
rect 14 1309 46 1341
rect 14 1241 46 1273
rect 14 1172 46 1204
rect 14 1104 46 1136
rect 14 1036 46 1068
rect 14 968 46 1000
rect 14 900 46 932
rect 14 832 46 864
rect 14 763 46 795
rect 14 695 46 727
rect 14 627 46 659
rect 14 559 46 591
rect 14 491 46 523
rect 14 423 46 455
rect 14 354 46 386
rect 14 286 46 318
rect 14 218 46 250
rect 14 150 46 182
rect 14 82 46 114
rect 14 14 46 46
rect 6490 6354 6522 6386
rect 6490 6285 6522 6317
rect 6490 6217 6522 6249
rect 6490 6149 6522 6181
rect 6490 6081 6522 6113
rect 6490 6013 6522 6045
rect 6490 5944 6522 5976
rect 6490 5876 6522 5908
rect 6490 5808 6522 5840
rect 6490 5740 6522 5772
rect 6490 5672 6522 5704
rect 6490 5604 6522 5636
rect 6490 5535 6522 5567
rect 6490 5467 6522 5499
rect 6490 5399 6522 5431
rect 6490 5331 6522 5363
rect 6490 5263 6522 5295
rect 6490 5195 6522 5227
rect 6490 5126 6522 5158
rect 6490 5058 6522 5090
rect 6490 4990 6522 5022
rect 6490 4922 6522 4954
rect 6490 4854 6522 4886
rect 6490 4786 6522 4818
rect 6490 4717 6522 4749
rect 6490 4649 6522 4681
rect 6490 4581 6522 4613
rect 6490 4513 6522 4545
rect 6490 4445 6522 4477
rect 6490 4377 6522 4409
rect 6490 4308 6522 4340
rect 6490 4240 6522 4272
rect 6490 4172 6522 4204
rect 6490 4104 6522 4136
rect 6490 4036 6522 4068
rect 6490 3967 6522 3999
rect 6490 3899 6522 3931
rect 6490 3831 6522 3863
rect 6490 3763 6522 3795
rect 6490 3695 6522 3727
rect 6490 3627 6522 3659
rect 6490 3558 6522 3590
rect 6490 3490 6522 3522
rect 6490 3422 6522 3454
rect 6490 3354 6522 3386
rect 6490 3286 6522 3318
rect 6490 3218 6522 3250
rect 6490 3149 6522 3181
rect 6490 3081 6522 3113
rect 6490 3013 6522 3045
rect 6490 2945 6522 2977
rect 6490 2877 6522 2909
rect 6490 2809 6522 2841
rect 6490 2740 6522 2772
rect 6490 2672 6522 2704
rect 6490 2604 6522 2636
rect 6490 2536 6522 2568
rect 6490 2468 6522 2500
rect 6490 2400 6522 2432
rect 6490 2331 6522 2363
rect 6490 2263 6522 2295
rect 6490 2195 6522 2227
rect 6490 2127 6522 2159
rect 6490 2059 6522 2091
rect 6490 1990 6522 2022
rect 6490 1922 6522 1954
rect 6490 1854 6522 1886
rect 6490 1786 6522 1818
rect 6490 1718 6522 1750
rect 6490 1650 6522 1682
rect 6490 1581 6522 1613
rect 6490 1513 6522 1545
rect 6490 1445 6522 1477
rect 6490 1377 6522 1409
rect 6490 1309 6522 1341
rect 6490 1241 6522 1273
rect 6490 1172 6522 1204
rect 6490 1104 6522 1136
rect 6490 1036 6522 1068
rect 6490 968 6522 1000
rect 6490 900 6522 932
rect 6490 832 6522 864
rect 6490 763 6522 795
rect 6490 695 6522 727
rect 6490 627 6522 659
rect 6490 559 6522 591
rect 6490 491 6522 523
rect 6490 423 6522 455
rect 6490 354 6522 386
rect 6490 286 6522 318
rect 6490 218 6522 250
rect 6490 150 6522 182
rect 6490 82 6522 114
rect 6490 14 6522 46
<< poly >>
rect 68 6400 6468 6436
rect 68 -36 6468 0
<< metal1 >>
rect 14 6386 46 6400
rect 14 6317 46 6354
rect 14 6249 46 6285
rect 14 6181 46 6217
rect 14 6113 46 6149
rect 14 6045 46 6081
rect 14 5976 46 6013
rect 14 5908 46 5944
rect 14 5840 46 5876
rect 14 5772 46 5808
rect 14 5704 46 5740
rect 14 5636 46 5672
rect 14 5567 46 5604
rect 14 5499 46 5535
rect 14 5431 46 5467
rect 14 5363 46 5399
rect 14 5295 46 5331
rect 14 5227 46 5263
rect 14 5158 46 5195
rect 14 5090 46 5126
rect 14 5022 46 5058
rect 14 4954 46 4990
rect 14 4886 46 4922
rect 14 4818 46 4854
rect 14 4749 46 4786
rect 14 4681 46 4717
rect 14 4613 46 4649
rect 14 4545 46 4581
rect 14 4477 46 4513
rect 14 4409 46 4445
rect 14 4340 46 4377
rect 14 4272 46 4308
rect 14 4204 46 4240
rect 14 4136 46 4172
rect 14 4068 46 4104
rect 14 3999 46 4036
rect 14 3931 46 3967
rect 14 3863 46 3899
rect 14 3795 46 3831
rect 14 3727 46 3763
rect 14 3659 46 3695
rect 14 3590 46 3627
rect 14 3522 46 3558
rect 14 3454 46 3490
rect 14 3386 46 3422
rect 14 3318 46 3354
rect 14 3250 46 3286
rect 14 3181 46 3218
rect 14 3113 46 3149
rect 14 3045 46 3081
rect 14 2977 46 3013
rect 14 2909 46 2945
rect 14 2841 46 2877
rect 14 2772 46 2809
rect 14 2704 46 2740
rect 14 2636 46 2672
rect 14 2568 46 2604
rect 14 2500 46 2536
rect 14 2432 46 2468
rect 14 2363 46 2400
rect 14 2295 46 2331
rect 14 2227 46 2263
rect 14 2159 46 2195
rect 14 2091 46 2127
rect 14 2022 46 2059
rect 14 1954 46 1990
rect 14 1886 46 1922
rect 14 1818 46 1854
rect 14 1750 46 1786
rect 14 1682 46 1718
rect 14 1613 46 1650
rect 14 1545 46 1581
rect 14 1477 46 1513
rect 14 1409 46 1445
rect 14 1341 46 1377
rect 14 1273 46 1309
rect 14 1204 46 1241
rect 14 1136 46 1172
rect 14 1068 46 1104
rect 14 1000 46 1036
rect 14 932 46 968
rect 14 864 46 900
rect 14 795 46 832
rect 14 727 46 763
rect 14 659 46 695
rect 14 591 46 627
rect 14 523 46 559
rect 14 455 46 491
rect 14 386 46 423
rect 14 318 46 354
rect 14 250 46 286
rect 14 182 46 218
rect 14 114 46 150
rect 14 46 46 82
rect 14 0 46 14
rect 6490 6386 6522 6400
rect 6490 6317 6522 6354
rect 6490 6249 6522 6285
rect 6490 6181 6522 6217
rect 6490 6113 6522 6149
rect 6490 6045 6522 6081
rect 6490 5976 6522 6013
rect 6490 5908 6522 5944
rect 6490 5840 6522 5876
rect 6490 5772 6522 5808
rect 6490 5704 6522 5740
rect 6490 5636 6522 5672
rect 6490 5567 6522 5604
rect 6490 5499 6522 5535
rect 6490 5431 6522 5467
rect 6490 5363 6522 5399
rect 6490 5295 6522 5331
rect 6490 5227 6522 5263
rect 6490 5158 6522 5195
rect 6490 5090 6522 5126
rect 6490 5022 6522 5058
rect 6490 4954 6522 4990
rect 6490 4886 6522 4922
rect 6490 4818 6522 4854
rect 6490 4749 6522 4786
rect 6490 4681 6522 4717
rect 6490 4613 6522 4649
rect 6490 4545 6522 4581
rect 6490 4477 6522 4513
rect 6490 4409 6522 4445
rect 6490 4340 6522 4377
rect 6490 4272 6522 4308
rect 6490 4204 6522 4240
rect 6490 4136 6522 4172
rect 6490 4068 6522 4104
rect 6490 3999 6522 4036
rect 6490 3931 6522 3967
rect 6490 3863 6522 3899
rect 6490 3795 6522 3831
rect 6490 3727 6522 3763
rect 6490 3659 6522 3695
rect 6490 3590 6522 3627
rect 6490 3522 6522 3558
rect 6490 3454 6522 3490
rect 6490 3386 6522 3422
rect 6490 3318 6522 3354
rect 6490 3250 6522 3286
rect 6490 3181 6522 3218
rect 6490 3113 6522 3149
rect 6490 3045 6522 3081
rect 6490 2977 6522 3013
rect 6490 2909 6522 2945
rect 6490 2841 6522 2877
rect 6490 2772 6522 2809
rect 6490 2704 6522 2740
rect 6490 2636 6522 2672
rect 6490 2568 6522 2604
rect 6490 2500 6522 2536
rect 6490 2432 6522 2468
rect 6490 2363 6522 2400
rect 6490 2295 6522 2331
rect 6490 2227 6522 2263
rect 6490 2159 6522 2195
rect 6490 2091 6522 2127
rect 6490 2022 6522 2059
rect 6490 1954 6522 1990
rect 6490 1886 6522 1922
rect 6490 1818 6522 1854
rect 6490 1750 6522 1786
rect 6490 1682 6522 1718
rect 6490 1613 6522 1650
rect 6490 1545 6522 1581
rect 6490 1477 6522 1513
rect 6490 1409 6522 1445
rect 6490 1341 6522 1377
rect 6490 1273 6522 1309
rect 6490 1204 6522 1241
rect 6490 1136 6522 1172
rect 6490 1068 6522 1104
rect 6490 1000 6522 1036
rect 6490 932 6522 968
rect 6490 864 6522 900
rect 6490 795 6522 832
rect 6490 727 6522 763
rect 6490 659 6522 695
rect 6490 591 6522 627
rect 6490 523 6522 559
rect 6490 455 6522 491
rect 6490 386 6522 423
rect 6490 318 6522 354
rect 6490 250 6522 286
rect 6490 182 6522 218
rect 6490 114 6522 150
rect 6490 46 6522 82
rect 6490 0 6522 14
<< labels >>
flabel comment s 3268 3200 3268 3200 0 FreeSans 200 90 0 0 pmosHV
<< end >>
