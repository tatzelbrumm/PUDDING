* NGSPICE file created from heichips25_pudding.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for analog_wires abstract view
.subckt analog_wires Iout VcascP[1] VcascP[0] VbiasP[1] VbiasP[0] VDDA[1] VDDA[0]
+ i_in i_out
.ends

* Black-box entry subcircuit for dac128module abstract view
.subckt dac128module VbiasP[1] Iout VbiasP[0] VcascP[1] VcascP[0] ON[64] ONB[64] ON[65]
+ ONB[65] ON[66] ONB[66] ON[67] ONB[67] ON[68] ONB[68] ON[69] ONB[69] ON[70] ONB[70]
+ ON[71] ONB[71] ON[72] ONB[72] EN[2] ENB[2] ON[73] ONB[73] ON[74] ONB[74] ON[75]
+ ONB[75] ON[76] ONB[76] ON[77] ONB[77] ON[78] ONB[78] ON[79] ONB[79] ON[80] ONB[80]
+ ON[81] ONB[81] ON[82] ONB[82] ON[83] ONB[83] ON[84] ONB[84] ON[85] ONB[85] ON[86]
+ ONB[86] ON[87] ONB[87] ON[88] ONB[88] ON[89] ONB[89] ON[90] ONB[90] ON[91] ONB[91]
+ ON[92] ONB[92] ON[93] ONB[93] ON[94] ONB[94] ON[95] ONB[95] ON[96] ONB[96] ON[97]
+ ONB[97] ON[98] ONB[98] ON[99] ONB[99] ON[100] ONB[100] ON[101] ONB[101] ON[102]
+ ONB[102] ON[103] ONB[103] ON[104] ONB[104] ON[105] ONB[105] ON[106] ONB[106] ON[107]
+ ONB[107] ON[108] ONB[108] ON[109] ONB[109] ON[110] ONB[110] ON[111] ONB[111] ON[112]
+ ONB[112] ON[113] ONB[113] ON[114] ONB[114] ON[115] ONB[115] ON[116] ONB[116] ON[117]
+ ONB[117] ON[118] ONB[118] ON[119] ONB[119] ON[120] ONB[120] ON[121] ONB[121] ON[122]
+ ONB[122] EN[3] ENB[3] ON[123] ONB[123] ON[124] ONB[124] ON[125] ONB[125] ON[126]
+ ONB[126] ON[127] ONB[127] ON[0] ONB[0] ON[1] ONB[1] ON[2] ONB[2] ON[3] ONB[3] ON[4]
+ ONB[4] ON[5] ONB[5] ON[6] EN[0] ENB[0] ONB[6] ON[7] ONB[7] ON[8] ONB[8] ON[9] ONB[9]
+ ON[10] ONB[10] ON[11] ONB[11] ON[12] ONB[12] ON[13] ONB[13] ON[14] ONB[14] ON[15]
+ ONB[15] ON[16] ONB[16] ON[17] ONB[17] ON[18] ONB[18] ON[19] ONB[19] ON[20] ONB[20]
+ ON[21] ONB[21] ON[22] ONB[22] ON[23] ONB[23] ON[24] ONB[24] ON[25] ONB[25] ON[26]
+ ONB[26] ON[27] ONB[27] ON[28] ONB[28] ON[29] ONB[29] ON[30] ONB[30] ON[31] ONB[31]
+ ON[33] ONB[33] ON[32] ONB[32] ON[34] ONB[34] ON[35] ONB[35] ON[36] ONB[36] ON[37]
+ ONB[37] ON[38] ONB[38] ON[39] ONB[39] ON[40] ONB[40] ON[41] ONB[41] ON[42] ONB[42]
+ ON[43] ONB[43] ON[44] ONB[44] ON[45] ONB[45] ON[46] ONB[46] ON[47] ONB[47] ON[48]
+ ONB[48] ON[49] ONB[49] ON[50] ONB[50] ON[51] ONB[51] ON[52] ONB[52] ON[53] ONB[53]
+ ON[54] ONB[54] ON[55] ONB[55] ON[56] ONB[56] ON[57] ONB[57] ON[58] ONB[58] ON[59]
+ ONB[59] ON[60] ONB[60] ON[61] ONB[61] ON[62] ONB[62] ON[63] ONB[63] EN[1] ENB[1]
+ VSS VDD
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

.subckt heichips25_pudding VGND VPWR clk ena i_in i_out rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_266 VPWR VGND sg13g2_decap_8
X_2106_ _0743_ net100 state\[25\] VPWR VGND sg13g2_nand2_1
X_2037_ _0703_ net157 _0702_ VPWR VGND sg13g2_nand2_1
XFILLER_10_339 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_13_111 VPWR VGND sg13g2_decap_8
XFILLER_26_472 VPWR VGND sg13g2_decap_4
XFILLER_26_85 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_13_188 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_4
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_5_321 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_5_398 VPWR VGND sg13g2_decap_8
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_3_78 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_17_494 VPWR VGND sg13g2_decap_8
XFILLER_44_280 VPWR VGND sg13g2_decap_8
X_2488__394 VPWR VGND net393 sg13g2_tiehi
X_1606_ state\[38\] daisychain\[38\] net139 _1002_ VPWR VGND sg13g2_mux2_1
X_1399_ VPWR _0032_ state\[13\] VGND sg13g2_inv_1
X_1468_ VGND VPWR net92 daisychain\[9\] _0892_ net45 sg13g2_a21oi_1
X_1537_ _0947_ net163 _0946_ VPWR VGND sg13g2_nand2_1
Xfanout105 net106 net105 VPWR VGND sg13g2_buf_1
Xfanout116 net117 net116 VPWR VGND sg13g2_buf_1
Xfanout127 net131 net127 VPWR VGND sg13g2_buf_1
Xfanout138 net141 net138 VPWR VGND sg13g2_buf_1
Xfanout149 net150 net149 VPWR VGND sg13g2_buf_1
XFILLER_27_258 VPWR VGND sg13g2_fill_1
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_10_136 VPWR VGND sg13g2_decap_8
XFILLER_6_107 VPWR VGND sg13g2_decap_8
XFILLER_7_608 VPWR VGND sg13g2_fill_2
XFILLER_7_619 VPWR VGND sg13g2_fill_1
XFILLER_12_98 VPWR VGND sg13g2_decap_8
XFILLER_2_357 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_fill_2
XFILLER_18_236 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_46_534 VPWR VGND sg13g2_fill_1
XFILLER_26_280 VPWR VGND sg13g2_fill_2
XFILLER_33_228 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
X_2440_ net328 VGND VPWR _0256_ state\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_5_195 VPWR VGND sg13g2_decap_8
X_1322_ VPWR _0117_ state\[90\] VGND sg13g2_inv_1
X_2371_ net210 VGND VPWR _0187_ daisychain\[59\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2340__273 VPWR VGND net272 sg13g2_tiehi
XFILLER_49_361 VPWR VGND sg13g2_decap_8
X_2555__248 VPWR VGND net247 sg13g2_tiehi
X_2416__377 VPWR VGND net376 sg13g2_tiehi
XFILLER_9_490 VPWR VGND sg13g2_fill_2
XFILLER_23_20 VPWR VGND sg13g2_decap_8
XFILLER_23_97 VPWR VGND sg13g2_decap_4
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_14_261 VPWR VGND sg13g2_decap_8
XFILLER_15_784 VPWR VGND sg13g2_fill_1
XFILLER_30_710 VPWR VGND sg13g2_fill_1
XFILLER_30_743 VPWR VGND sg13g2_fill_1
XFILLER_30_776 VPWR VGND sg13g2_fill_1
XFILLER_9_77 VPWR VGND sg13g2_decap_8
X_2450__290 VPWR VGND net289 sg13g2_tiehi
X_1940_ VGND VPWR _0623_ _0624_ _0232_ _0625_ sg13g2_a21oi_1
X_1871_ state\[91\] daisychain\[91\] net151 _0570_ VPWR VGND sg13g2_mux2_1
XFILLER_6_471 VPWR VGND sg13g2_decap_4
X_2561__296 VPWR VGND net295 sg13g2_tiehi
X_2423_ net362 VGND VPWR _0239_ daisychain\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1305_ VPWR _0008_ state\[107\] VGND sg13g2_inv_1
X_2354_ net244 VGND VPWR _0170_ daisychain\[42\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2285_ VGND VPWR _0663_ _0832_ _0370_ net76 sg13g2_a21oi_1
XFILLER_25_526 VPWR VGND sg13g2_decap_8
XFILLER_37_364 VPWR VGND sg13g2_decap_8
XFILLER_20_264 VPWR VGND sg13g2_decap_8
XFILLER_18_75 VPWR VGND sg13g2_decap_8
XFILLER_28_364 VPWR VGND sg13g2_fill_1
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_48_629 VPWR VGND sg13g2_fill_1
X_2319__315 VPWR VGND net314 sg13g2_tiehi
XFILLER_11_220 VPWR VGND sg13g2_decap_8
XFILLER_34_96 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_11_297 VPWR VGND sg13g2_decap_8
XFILLER_3_463 VPWR VGND sg13g2_decap_8
XFILLER_7_257 VPWR VGND sg13g2_decap_8
XFILLER_8_758 VPWR VGND sg13g2_decap_8
XFILLER_19_320 VPWR VGND sg13g2_fill_2
XFILLER_19_331 VPWR VGND sg13g2_decap_8
X_2070_ _0725_ net101 state\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_22_507 VPWR VGND sg13g2_fill_1
XFILLER_34_334 VPWR VGND sg13g2_fill_1
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_47_673 VPWR VGND sg13g2_decap_8
XFILLER_47_684 VPWR VGND sg13g2_fill_2
X_1923_ VGND VPWR net112 daisychain\[100\] _0612_ net54 sg13g2_a21oi_1
X_1854_ net196 VPWR _0557_ VGND daisychain\[87\] net39 sg13g2_o21ai_1
X_1785_ VGND VPWR _0499_ _0500_ _0201_ _0501_ sg13g2_a21oi_1
XFILLER_7_780 VPWR VGND sg13g2_fill_1
X_2406_ net396 VGND VPWR _0222_ daisychain\[94\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_37_161 VPWR VGND sg13g2_decap_8
X_2337_ net278 VGND VPWR _0153_ daisychain\[25\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2268_ _0824_ net107 state\[106\] VPWR VGND sg13g2_nand2_1
X_2199_ VGND VPWR _0491_ _0789_ _0327_ net87 sg13g2_a21oi_1
XFILLER_25_345 VPWR VGND sg13g2_decap_8
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_4_227 VPWR VGND sg13g2_decap_8
X_2464__234 VPWR VGND net233 sg13g2_tiehi
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_29_52 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_16_356 VPWR VGND sg13g2_fill_1
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_fill_2
XFILLER_45_84 VPWR VGND sg13g2_decap_8
X_2512__268 VPWR VGND net267 sg13g2_tiehi
XFILLER_3_260 VPWR VGND sg13g2_decap_8
X_2443__318 VPWR VGND net317 sg13g2_tiehi
X_1570_ VGND VPWR _0971_ _0972_ _0158_ _0973_ sg13g2_a21oi_1
XFILLER_19_183 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_4
X_2122_ _0751_ net117 state\[33\] VPWR VGND sg13g2_nand2_1
X_2053_ VGND VPWR net91 daisychain\[126\] _0716_ net48 sg13g2_a21oi_1
XFILLER_22_348 VPWR VGND sg13g2_fill_1
XFILLER_34_131 VPWR VGND sg13g2_decap_8
XFILLER_35_687 VPWR VGND sg13g2_decap_8
X_1906_ state\[98\] daisychain\[98\] net142 _0598_ VPWR VGND sg13g2_mux2_1
X_1837_ _0543_ net173 _0542_ VPWR VGND sg13g2_nand2_1
X_1768_ VGND VPWR net129 daisychain\[69\] _0488_ net64 sg13g2_a21oi_1
X_1699_ net194 VPWR _0433_ VGND daisychain\[56\] net37 sg13g2_o21ai_1
XFILLER_15_65 VPWR VGND sg13g2_decap_8
XFILLER_25_186 VPWR VGND sg13g2_decap_8
XFILLER_31_53 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_41_668 VPWR VGND sg13g2_decap_8
XFILLER_5_514 VPWR VGND sg13g2_fill_2
XFILLER_9_308 VPWR VGND sg13g2_decap_8
XFILLER_5_569 VPWR VGND sg13g2_decap_4
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_1_775 VPWR VGND sg13g2_fill_1
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_49_779 VPWR VGND sg13g2_decap_4
XFILLER_16_153 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_fill_1
XFILLER_31_123 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_8
XFILLER_44_473 VPWR VGND sg13g2_fill_1
XFILLER_8_341 VPWR VGND sg13g2_decap_8
X_1622_ _1015_ net169 _1014_ VPWR VGND sg13g2_nand2_1
X_1484_ net180 VPWR _0905_ VGND daisychain\[13\] net23 sg13g2_o21ai_1
X_1553_ VGND VPWR net100 daisychain\[26\] _0960_ net52 sg13g2_a21oi_1
X_2380__449 VPWR VGND net448 sg13g2_tiehi
XFILLER_39_245 VPWR VGND sg13g2_decap_8
X_2105_ VGND VPWR _0947_ _0742_ _0280_ net73 sg13g2_a21oi_1
X_2036_ state\[124\] daisychain\[124\] net135 _0702_ VPWR VGND sg13g2_mux2_1
XFILLER_10_318 VPWR VGND sg13g2_decap_8
XFILLER_11_819 VPWR VGND sg13g2_decap_4
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_31_690 VPWR VGND sg13g2_decap_8
X_2350__253 VPWR VGND net252 sg13g2_tiehi
XFILLER_2_539 VPWR VGND sg13g2_decap_8
X_2426__357 VPWR VGND net356 sg13g2_tiehi
XFILLER_13_167 VPWR VGND sg13g2_decap_8
XFILLER_14_646 VPWR VGND sg13g2_fill_1
XFILLER_14_657 VPWR VGND sg13g2_fill_1
XFILLER_26_42 VPWR VGND sg13g2_decap_4
XFILLER_26_64 VPWR VGND sg13g2_decap_8
XFILLER_41_421 VPWR VGND sg13g2_decap_8
XFILLER_41_432 VPWR VGND sg13g2_fill_2
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_9_105 VPWR VGND sg13g2_decap_8
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_5_300 VPWR VGND sg13g2_decap_8
XFILLER_6_812 VPWR VGND sg13g2_decap_8
XFILLER_1_550 VPWR VGND sg13g2_fill_1
XFILLER_3_35 VPWR VGND sg13g2_fill_2
XFILLER_3_57 VPWR VGND sg13g2_decap_8
XFILLER_5_377 VPWR VGND sg13g2_decap_8
X_2327__299 VPWR VGND net298 sg13g2_tiehi
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_fill_2
X_1536_ state\[24\] daisychain\[24\] net139 _0946_ VPWR VGND sg13g2_mux2_1
X_1605_ VGND VPWR _0999_ _1000_ _0165_ _1001_ sg13g2_a21oi_1
X_1398_ VPWR _0033_ state\[14\] VGND sg13g2_inv_1
X_1467_ _0891_ net158 _0890_ VPWR VGND sg13g2_nand2_1
Xfanout106 net114 net106 VPWR VGND sg13g2_buf_1
Xfanout117 net123 net117 VPWR VGND sg13g2_buf_1
Xfanout128 net130 net128 VPWR VGND sg13g2_buf_1
Xfanout139 net141 net139 VPWR VGND sg13g2_buf_1
X_2495__366 VPWR VGND net365 sg13g2_tiehi
XFILLER_27_237 VPWR VGND sg13g2_decap_8
XFILLER_36_771 VPWR VGND sg13g2_decap_4
XFILLER_36_782 VPWR VGND sg13g2_decap_8
X_2019_ net179 VPWR _0689_ VGND daisychain\[120\] net25 sg13g2_o21ai_1
XFILLER_10_115 VPWR VGND sg13g2_decap_8
XFILLER_12_77 VPWR VGND sg13g2_decap_8
XFILLER_2_336 VPWR VGND sg13g2_decap_8
XFILLER_18_215 VPWR VGND sg13g2_decap_8
XFILLER_19_749 VPWR VGND sg13g2_fill_1
XFILLER_33_207 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_5_174 VPWR VGND sg13g2_decap_8
XFILLER_6_697 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
X_1321_ VPWR _0118_ state\[91\] VGND sg13g2_inv_1
X_2379__451 VPWR VGND net450 sg13g2_tiehi
X_2370_ net212 VGND VPWR _0186_ daisychain\[58\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_17_281 VPWR VGND sg13g2_decap_8
XFILLER_24_218 VPWR VGND sg13g2_fill_2
XFILLER_33_752 VPWR VGND sg13g2_decap_4
XFILLER_37_579 VPWR VGND sg13g2_fill_1
XFILLER_20_479 VPWR VGND sg13g2_fill_1
XFILLER_32_284 VPWR VGND sg13g2_decap_8
X_1519_ net185 VPWR _0933_ VGND daisychain\[20\] net28 sg13g2_o21ai_1
X_2499_ net349 VGND VPWR _0315_ state\[59\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_28_513 VPWR VGND sg13g2_fill_2
XFILLER_28_524 VPWR VGND sg13g2_decap_8
XFILLER_11_457 VPWR VGND sg13g2_fill_1
XFILLER_23_76 VPWR VGND sg13g2_decap_8
XFILLER_7_439 VPWR VGND sg13g2_decap_8
XFILLER_19_502 VPWR VGND sg13g2_fill_2
XFILLER_19_513 VPWR VGND sg13g2_fill_1
XFILLER_2_133 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_14_240 VPWR VGND sg13g2_decap_8
XFILLER_34_549 VPWR VGND sg13g2_fill_1
XFILLER_46_343 VPWR VGND sg13g2_decap_8
X_2515__244 VPWR VGND net243 sg13g2_tiehi
XFILLER_30_722 VPWR VGND sg13g2_fill_2
XFILLER_30_755 VPWR VGND sg13g2_fill_2
X_1870_ VGND VPWR _0567_ _0568_ _0218_ _0569_ sg13g2_a21oi_1
XFILLER_6_450 VPWR VGND sg13g2_decap_8
X_2422_ net364 VGND VPWR _0238_ daisychain\[110\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2353_ net246 VGND VPWR _0169_ daisychain\[41\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_38_822 VPWR VGND sg13g2_fill_1
X_1304_ VPWR _0009_ state\[108\] VGND sg13g2_inv_1
X_2284_ _0832_ net108 state\[114\] VPWR VGND sg13g2_nand2_1
XFILLER_40_508 VPWR VGND sg13g2_fill_2
XFILLER_20_243 VPWR VGND sg13g2_decap_8
XFILLER_4_409 VPWR VGND sg13g2_decap_8
X_1999_ net181 VPWR _0673_ VGND daisychain\[116\] net24 sg13g2_o21ai_1
XFILLER_16_505 VPWR VGND sg13g2_fill_1
XFILLER_16_538 VPWR VGND sg13g2_fill_2
XFILLER_18_54 VPWR VGND sg13g2_decap_8
XFILLER_28_310 VPWR VGND sg13g2_fill_2
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_11_276 VPWR VGND sg13g2_decap_8
XFILLER_12_755 VPWR VGND sg13g2_decap_4
XFILLER_34_75 VPWR VGND sg13g2_decap_8
XFILLER_7_236 VPWR VGND sg13g2_decap_8
X_2549__384 VPWR VGND net383 sg13g2_tiehi
XFILLER_3_442 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_19_387 VPWR VGND sg13g2_fill_1
XFILLER_34_313 VPWR VGND sg13g2_decap_8
XFILLER_34_346 VPWR VGND sg13g2_decap_8
X_1922_ _0611_ net166 _0610_ VPWR VGND sg13g2_nand2_1
XFILLER_30_563 VPWR VGND sg13g2_fill_1
X_1853_ VGND VPWR net124 daisychain\[86\] _0556_ net64 sg13g2_a21oi_1
X_1784_ net198 VPWR _0501_ VGND daisychain\[73\] net41 sg13g2_o21ai_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_2405_ net398 VGND VPWR _0221_ daisychain\[93\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2336_ net280 VGND VPWR _0152_ daisychain\[24\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_29_129 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
X_2390__429 VPWR VGND net428 sg13g2_tiehi
X_2267_ VGND VPWR _0627_ _0823_ _0361_ net76 sg13g2_a21oi_1
X_2198_ _0789_ net130 state\[71\] VPWR VGND sg13g2_nand2_1
XFILLER_4_206 VPWR VGND sg13g2_decap_8
X_2360__233 VPWR VGND net232 sg13g2_tiehi
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_29_31 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
X_2471__206 VPWR VGND net205 sg13g2_tiehi
XFILLER_24_390 VPWR VGND sg13g2_fill_1
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_31_305 VPWR VGND sg13g2_fill_2
XFILLER_31_338 VPWR VGND sg13g2_fill_1
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_44_633 VPWR VGND sg13g2_fill_1
XFILLER_44_644 VPWR VGND sg13g2_fill_2
XFILLER_45_63 VPWR VGND sg13g2_decap_8
X_2436__337 VPWR VGND net336 sg13g2_tiehi
XFILLER_12_541 VPWR VGND sg13g2_fill_1
XFILLER_12_585 VPWR VGND sg13g2_decap_4
XFILLER_6_79 VPWR VGND sg13g2_decap_8
XFILLER_19_162 VPWR VGND sg13g2_decap_8
XFILLER_34_110 VPWR VGND sg13g2_decap_8
XFILLER_35_622 VPWR VGND sg13g2_fill_1
X_2337__279 VPWR VGND net278 sg13g2_tiehi
X_2121_ VGND VPWR _0979_ _0750_ _0288_ net74 sg13g2_a21oi_1
X_2052_ _0715_ net157 _0714_ VPWR VGND sg13g2_nand2_1
XFILLER_34_187 VPWR VGND sg13g2_decap_8
XFILLER_35_699 VPWR VGND sg13g2_decap_8
X_1905_ VGND VPWR _0595_ _0596_ _0225_ _0597_ sg13g2_a21oi_1
XFILLER_30_393 VPWR VGND sg13g2_decap_4
X_1836_ state\[84\] daisychain\[84\] net152 _0542_ VPWR VGND sg13g2_mux2_1
X_1767_ _0487_ net176 _0486_ VPWR VGND sg13g2_nand2_1
X_1698_ VGND VPWR net119 daisychain\[55\] _0432_ net59 sg13g2_a21oi_1
X_2319_ net314 VGND VPWR _0135_ daisychain\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_13_349 VPWR VGND sg13g2_decap_8
XFILLER_14_817 VPWR VGND sg13g2_decap_4
XFILLER_25_165 VPWR VGND sg13g2_decap_8
XFILLER_31_32 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_5_548 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_16_132 VPWR VGND sg13g2_decap_8
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_12_371 VPWR VGND sg13g2_fill_2
XFILLER_17_699 VPWR VGND sg13g2_fill_2
XFILLER_31_102 VPWR VGND sg13g2_decap_8
XFILLER_31_179 VPWR VGND sg13g2_decap_8
XFILLER_40_680 VPWR VGND sg13g2_decap_4
XFILLER_8_320 VPWR VGND sg13g2_decap_8
XFILLER_4_570 VPWR VGND sg13g2_fill_2
XFILLER_8_397 VPWR VGND sg13g2_decap_8
X_1552_ _0959_ net161 _0958_ VPWR VGND sg13g2_nand2_1
X_1621_ state\[41\] daisychain\[41\] net146 _1014_ VPWR VGND sg13g2_mux2_1
XFILLER_27_408 VPWR VGND sg13g2_decap_8
XFILLER_39_224 VPWR VGND sg13g2_decap_8
X_1483_ VGND VPWR net92 daisychain\[12\] _0904_ net45 sg13g2_a21oi_1
X_2104_ _0742_ net105 state\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_22_102 VPWR VGND sg13g2_decap_8
X_2035_ VGND VPWR _0699_ _0700_ _0251_ _0701_ sg13g2_a21oi_1
XFILLER_22_179 VPWR VGND sg13g2_decap_8
X_2389__431 VPWR VGND net430 sg13g2_tiehi
XFILLER_2_518 VPWR VGND sg13g2_decap_8
X_1819_ net199 VPWR _0529_ VGND daisychain\[80\] net42 sg13g2_o21ai_1
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_13_146 VPWR VGND sg13g2_decap_8
XFILLER_41_444 VPWR VGND sg13g2_fill_1
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_5_356 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_45_761 VPWR VGND sg13g2_decap_4
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_49_599 VPWR VGND sg13g2_fill_2
X_2518__220 VPWR VGND net219 sg13g2_tiehi
XFILLER_20_606 VPWR VGND sg13g2_fill_1
XFILLER_8_194 VPWR VGND sg13g2_decap_8
X_1535_ VGND VPWR _0943_ _0944_ _0151_ _0945_ sg13g2_a21oi_1
Xfanout107 net108 net107 VPWR VGND sg13g2_buf_1
Xfanout118 net121 net118 VPWR VGND sg13g2_buf_1
Xfanout129 net130 net129 VPWR VGND sg13g2_buf_1
X_1604_ net185 VPWR _1001_ VGND daisychain\[37\] net28 sg13g2_o21ai_1
XFILLER_27_216 VPWR VGND sg13g2_decap_8
XFILLER_43_709 VPWR VGND sg13g2_decap_8
X_1397_ VPWR _0034_ state\[15\] VGND sg13g2_inv_1
X_1466_ state\[10\] daisychain\[10\] net133 _0890_ VPWR VGND sg13g2_mux2_1
XFILLER_23_444 VPWR VGND sg13g2_fill_2
X_2018_ VGND VPWR net97 daisychain\[119\] _0688_ net46 sg13g2_a21oi_1
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_19_706 VPWR VGND sg13g2_fill_2
XFILLER_2_315 VPWR VGND sg13g2_decap_8
XFILLER_5_6 VPWR VGND sg13g2_fill_1
XFILLER_14_411 VPWR VGND sg13g2_decap_8
XFILLER_19_717 VPWR VGND sg13g2_fill_2
XFILLER_26_282 VPWR VGND sg13g2_fill_1
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_46_569 VPWR VGND sg13g2_fill_2
XFILLER_10_672 VPWR VGND sg13g2_decap_8
XFILLER_14_466 VPWR VGND sg13g2_decap_4
XFILLER_14_488 VPWR VGND sg13g2_fill_2
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_153 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_8
X_1320_ VPWR _0119_ state\[92\] VGND sg13g2_inv_1
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_503 VPWR VGND sg13g2_decap_4
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_17_260 VPWR VGND sg13g2_decap_8
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_33_720 VPWR VGND sg13g2_decap_8
XFILLER_33_764 VPWR VGND sg13g2_fill_2
X_1449_ net187 VPWR _0877_ VGND daisychain\[6\] net30 sg13g2_o21ai_1
X_1518_ VGND VPWR net99 daisychain\[19\] _0932_ net50 sg13g2_a21oi_1
X_2567_ net455 VGND VPWR _0383_ state\[127\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2498_ net353 VGND VPWR _0314_ state\[58\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_15_219 VPWR VGND sg13g2_decap_8
XFILLER_11_469 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_fill_2
XFILLER_23_55 VPWR VGND sg13g2_decap_8
XFILLER_7_418 VPWR VGND sg13g2_decap_8
X_2467__222 VPWR VGND net221 sg13g2_tiehi
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_3_602 VPWR VGND sg13g2_decap_8
XFILLER_3_657 VPWR VGND sg13g2_fill_1
XFILLER_3_668 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
X_2521__452 VPWR VGND net451 sg13g2_tiehi
XFILLER_30_701 VPWR VGND sg13g2_fill_2
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_9_13 VPWR VGND sg13g2_fill_1
X_2370__213 VPWR VGND net212 sg13g2_tiehi
XFILLER_10_491 VPWR VGND sg13g2_decap_8
XFILLER_14_296 VPWR VGND sg13g2_decap_8
XFILLER_30_789 VPWR VGND sg13g2_decap_4
X_2446__306 VPWR VGND net305 sg13g2_tiehi
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_6_484 VPWR VGND sg13g2_fill_1
X_1303_ VPWR _0010_ state\[109\] VGND sg13g2_inv_1
X_2421_ net366 VGND VPWR _0237_ daisychain\[109\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2352_ net248 VGND VPWR _0168_ daisychain\[40\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2283_ VGND VPWR _0659_ _0831_ _0369_ net69 sg13g2_a21oi_1
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_38_801 VPWR VGND sg13g2_fill_1
XFILLER_49_193 VPWR VGND sg13g2_decap_8
X_2533__356 VPWR VGND net355 sg13g2_tiehi
XFILLER_20_222 VPWR VGND sg13g2_decap_8
XFILLER_33_561 VPWR VGND sg13g2_fill_2
XFILLER_20_299 VPWR VGND sg13g2_decap_8
X_2347__259 VPWR VGND net258 sg13g2_tiehi
X_1998_ VGND VPWR net96 daisychain\[115\] _0672_ net46 sg13g2_a21oi_1
XFILLER_18_33 VPWR VGND sg13g2_decap_8
XFILLER_28_300 VPWR VGND sg13g2_fill_1
XFILLER_28_333 VPWR VGND sg13g2_fill_2
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_34_54 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_11_255 VPWR VGND sg13g2_decap_8
XFILLER_7_215 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_421 VPWR VGND sg13g2_decap_8
XFILLER_3_498 VPWR VGND sg13g2_decap_8
XFILLER_19_355 VPWR VGND sg13g2_fill_2
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_30_531 VPWR VGND sg13g2_fill_1
XFILLER_46_196 VPWR VGND sg13g2_decap_8
X_1921_ state\[101\] daisychain\[101\] net143 _0610_ VPWR VGND sg13g2_mux2_1
X_1852_ _0555_ net173 _0554_ VPWR VGND sg13g2_nand2_1
XFILLER_30_597 VPWR VGND sg13g2_fill_1
X_1783_ VGND VPWR net128 daisychain\[72\] _0500_ net62 sg13g2_a21oi_1
XFILLER_29_108 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_2404_ net400 VGND VPWR _0220_ daisychain\[92\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2335_ net282 VGND VPWR _0151_ daisychain\[23\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2266_ _0823_ net107 state\[105\] VPWR VGND sg13g2_nand2_1
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
X_2197_ VGND VPWR _0487_ _0788_ _0326_ net87 sg13g2_a21oi_1
XFILLER_5_708 VPWR VGND sg13g2_fill_2
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_20_89 VPWR VGND sg13g2_decap_8
X_2399__411 VPWR VGND net410 sg13g2_tiehi
XFILLER_16_314 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_29_87 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_8
XFILLER_16_347 VPWR VGND sg13g2_decap_8
XFILLER_16_369 VPWR VGND sg13g2_decap_4
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_44_678 VPWR VGND sg13g2_decap_4
XFILLER_44_689 VPWR VGND sg13g2_fill_1
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_8_557 VPWR VGND sg13g2_fill_1
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_3_295 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_fill_2
X_2120_ _0750_ net106 state\[32\] VPWR VGND sg13g2_nand2_1
XFILLER_19_141 VPWR VGND sg13g2_decap_8
XFILLER_34_166 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
X_2051_ state\[127\] daisychain\[127\] net135 _0714_ VPWR VGND sg13g2_mux2_1
X_1904_ net190 VPWR _0597_ VGND daisychain\[97\] net33 sg13g2_o21ai_1
X_1835_ VGND VPWR _0539_ _0540_ _0211_ _0541_ sg13g2_a21oi_1
X_1766_ state\[70\] daisychain\[70\] net154 _0486_ VPWR VGND sg13g2_mux2_1
X_1697_ _0431_ net171 _0430_ VPWR VGND sg13g2_nand2_1
X_2498__354 VPWR VGND net353 sg13g2_tiehi
X_2318_ net316 VGND VPWR _0134_ daisychain\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2249_ VGND VPWR _0591_ _0814_ _0352_ net78 sg13g2_a21oi_1
XFILLER_13_328 VPWR VGND sg13g2_decap_8
XFILLER_15_34 VPWR VGND sg13g2_fill_1
XFILLER_25_144 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_31_11 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_decap_8
XFILLER_5_527 VPWR VGND sg13g2_fill_2
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_49_759 VPWR VGND sg13g2_decap_8
X_2557__440 VPWR VGND net439 sg13g2_tiehi
Xoutput9 net9 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_out[4] VPWR VGND sg13g2_buf_1
X_2477__438 VPWR VGND net437 sg13g2_tiehi
XFILLER_16_111 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_12_350 VPWR VGND sg13g2_decap_8
XFILLER_16_188 VPWR VGND sg13g2_decap_8
XFILLER_31_158 VPWR VGND sg13g2_decap_8
XFILLER_32_648 VPWR VGND sg13g2_fill_2
XFILLER_9_822 VPWR VGND sg13g2_fill_1
XFILLER_4_593 VPWR VGND sg13g2_decap_4
XFILLER_8_376 VPWR VGND sg13g2_decap_8
X_1482_ _0903_ net159 _0902_ VPWR VGND sg13g2_nand2_1
X_1551_ state\[27\] daisychain\[27\] net138 _0958_ VPWR VGND sg13g2_mux2_1
X_1620_ VGND VPWR _1011_ _1012_ _0168_ _1013_ sg13g2_a21oi_1
XFILLER_39_203 VPWR VGND sg13g2_decap_8
X_2103_ VGND VPWR _0943_ _0741_ _0279_ net73 sg13g2_a21oi_1
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_35_442 VPWR VGND sg13g2_decap_4
XFILLER_47_280 VPWR VGND sg13g2_decap_8
X_2034_ net179 VPWR _0701_ VGND daisychain\[123\] net25 sg13g2_o21ai_1
X_1818_ VGND VPWR net127 daisychain\[79\] _0528_ net63 sg13g2_a21oi_1
X_1749_ net198 VPWR _0473_ VGND daisychain\[66\] net41 sg13g2_o21ai_1
XFILLER_14_604 VPWR VGND sg13g2_fill_2
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_13_125 VPWR VGND sg13g2_decap_8
XFILLER_26_99 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_5_335 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_49_578 VPWR VGND sg13g2_decap_4
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_fill_1
XFILLER_20_618 VPWR VGND sg13g2_fill_1
XFILLER_8_173 VPWR VGND sg13g2_decap_8
XFILLER_9_685 VPWR VGND sg13g2_fill_1
X_1465_ VGND VPWR _0887_ _0888_ _0137_ _0889_ sg13g2_a21oi_1
X_1534_ net185 VPWR _0945_ VGND daisychain\[23\] net28 sg13g2_o21ai_1
Xfanout108 net109 net108 VPWR VGND sg13g2_buf_1
Xfanout119 net121 net119 VPWR VGND sg13g2_buf_1
X_2460__250 VPWR VGND net249 sg13g2_tiehi
X_1603_ VGND VPWR net103 daisychain\[36\] _1000_ net57 sg13g2_a21oi_1
X_1396_ VPWR _0035_ state\[16\] VGND sg13g2_inv_1
X_2536__332 VPWR VGND net331 sg13g2_tiehi
X_2017_ _0687_ net157 _0686_ VPWR VGND sg13g2_nand2_1
XFILLER_23_467 VPWR VGND sg13g2_decap_8
XFILLER_23_478 VPWR VGND sg13g2_fill_2
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_12_13 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_46_515 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_42_743 VPWR VGND sg13g2_fill_2
XFILLER_46_526 VPWR VGND sg13g2_fill_2
X_2357__239 VPWR VGND net238 sg13g2_tiehi
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_5_132 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
X_2559__376 VPWR VGND net375 sg13g2_tiehi
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_9_471 VPWR VGND sg13g2_fill_1
XFILLER_28_504 VPWR VGND sg13g2_decap_4
XFILLER_28_515 VPWR VGND sg13g2_fill_1
XFILLER_4_80 VPWR VGND sg13g2_decap_8
X_1448_ VGND VPWR net108 daisychain\[5\] _0876_ net53 sg13g2_a21oi_1
X_1517_ _0931_ net163 _0930_ VPWR VGND sg13g2_nand2_1
X_2566_ net391 VGND VPWR _0382_ state\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2497_ net357 VGND VPWR _0313_ state\[57\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_43_529 VPWR VGND sg13g2_fill_2
X_1379_ VPWR _0054_ state\[33\] VGND sg13g2_inv_1
XFILLER_11_415 VPWR VGND sg13g2_fill_2
XFILLER_23_286 VPWR VGND sg13g2_decap_4
XFILLER_23_297 VPWR VGND sg13g2_decap_4
XFILLER_23_34 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_19_504 VPWR VGND sg13g2_fill_1
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_14_275 VPWR VGND sg13g2_decap_8
XFILLER_15_754 VPWR VGND sg13g2_decap_8
XFILLER_15_765 VPWR VGND sg13g2_fill_2
XFILLER_30_735 VPWR VGND sg13g2_fill_1
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_fill_2
XFILLER_30_768 VPWR VGND sg13g2_fill_1
Xfanout90 net91 net90 VPWR VGND sg13g2_buf_1
X_2420_ net368 VGND VPWR _0236_ daisychain\[108\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_38_813 VPWR VGND sg13g2_decap_8
X_1302_ VPWR _0012_ state\[110\] VGND sg13g2_inv_1
X_2351_ net250 VGND VPWR _0167_ daisychain\[39\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2282_ _0831_ net108 state\[113\] VPWR VGND sg13g2_nand2_1
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_20_201 VPWR VGND sg13g2_decap_8
XFILLER_20_278 VPWR VGND sg13g2_decap_8
X_1997_ _0671_ net159 _0670_ VPWR VGND sg13g2_nand2_1
X_2549_ net383 VGND VPWR _0365_ state\[109\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_18_89 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_11_234 VPWR VGND sg13g2_decap_8
XFILLER_3_400 VPWR VGND sg13g2_decap_8
XFILLER_8_706 VPWR VGND sg13g2_decap_8
XFILLER_8_728 VPWR VGND sg13g2_decap_8
XFILLER_3_477 VPWR VGND sg13g2_decap_8
XFILLER_19_367 VPWR VGND sg13g2_decap_4
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_47_698 VPWR VGND sg13g2_fill_1
X_2491__382 VPWR VGND net381 sg13g2_tiehi
XFILLER_15_562 VPWR VGND sg13g2_fill_2
XFILLER_42_392 VPWR VGND sg13g2_decap_8
X_1920_ VGND VPWR _0607_ _0608_ _0228_ _0609_ sg13g2_a21oi_1
X_1851_ state\[87\] daisychain\[87\] net152 _0554_ VPWR VGND sg13g2_mux2_1
XFILLER_6_282 VPWR VGND sg13g2_decap_8
X_2403_ net402 VGND VPWR _0219_ daisychain\[91\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1782_ _0499_ net175 _0498_ VPWR VGND sg13g2_nand2_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
X_2334_ net284 VGND VPWR _0150_ daisychain\[22\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2265_ VGND VPWR _0623_ _0822_ _0360_ net78 sg13g2_a21oi_1
X_2196_ _0788_ net130 state\[70\] VPWR VGND sg13g2_nand2_1
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_21_510 VPWR VGND sg13g2_fill_1
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_20_68 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_29_66 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_44_624 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv1 VPWR digitalen.g\[2\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_31_307 VPWR VGND sg13g2_fill_1
XFILLER_32_819 VPWR VGND sg13g2_decap_4
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_19_120 VPWR VGND sg13g2_decap_8
XFILLER_3_274 VPWR VGND sg13g2_decap_8
X_2558__408 VPWR VGND net407 sg13g2_tiehi
X_2050_ VGND VPWR _0711_ _0712_ _0254_ _0713_ sg13g2_a21oi_1
XFILLER_19_197 VPWR VGND sg13g2_decap_8
XFILLER_34_145 VPWR VGND sg13g2_decap_8
XFILLER_35_657 VPWR VGND sg13g2_fill_1
XFILLER_47_462 VPWR VGND sg13g2_decap_8
X_1903_ VGND VPWR net112 daisychain\[96\] _0596_ net54 sg13g2_a21oi_1
X_1834_ net196 VPWR _0541_ VGND daisychain\[83\] net39 sg13g2_o21ai_1
X_1765_ VGND VPWR _0483_ _0484_ _0197_ _0485_ sg13g2_a21oi_1
X_1696_ state\[56\] daisychain\[56\] net148 _0430_ VPWR VGND sg13g2_mux2_1
X_2317_ net318 VGND VPWR _0133_ daisychain\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2248_ _0814_ net112 state\[96\] VPWR VGND sg13g2_nand2_1
X_2179_ VGND VPWR _0451_ _0779_ _0317_ net82 sg13g2_a21oi_1
XFILLER_13_307 VPWR VGND sg13g2_decap_8
XFILLER_15_79 VPWR VGND sg13g2_decap_8
XFILLER_21_340 VPWR VGND sg13g2_fill_1
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_31_67 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_16_167 VPWR VGND sg13g2_decap_8
XFILLER_29_451 VPWR VGND sg13g2_decap_8
X_2336__281 VPWR VGND net280 sg13g2_tiehi
XFILLER_31_137 VPWR VGND sg13g2_decap_8
XFILLER_8_355 VPWR VGND sg13g2_decap_8
X_2367__219 VPWR VGND net218 sg13g2_tiehi
XFILLER_4_572 VPWR VGND sg13g2_fill_1
X_1481_ state\[13\] daisychain\[13\] net134 _0902_ VPWR VGND sg13g2_mux2_1
X_1550_ VGND VPWR _0955_ _0956_ _0154_ _0957_ sg13g2_a21oi_1
XFILLER_39_259 VPWR VGND sg13g2_decap_8
X_2102_ _0741_ net104 state\[23\] VPWR VGND sg13g2_nand2_1
X_2033_ VGND VPWR net90 daisychain\[122\] _0700_ net48 sg13g2_a21oi_1
XFILLER_16_690 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_decap_8
X_1817_ _0527_ net174 _0526_ VPWR VGND sg13g2_nand2_1
X_1748_ VGND VPWR net127 daisychain\[65\] _0472_ net63 sg13g2_a21oi_1
X_1679_ net194 VPWR _0417_ VGND daisychain\[52\] net37 sg13g2_o21ai_1
XFILLER_13_104 VPWR VGND sg13g2_decap_8
XFILLER_26_465 VPWR VGND sg13g2_fill_2
XFILLER_26_78 VPWR VGND sg13g2_decap_8
XFILLER_39_771 VPWR VGND sg13g2_fill_2
XFILLER_41_413 VPWR VGND sg13g2_decap_4
XFILLER_21_192 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_5_314 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_17_454 VPWR VGND sg13g2_decap_4
XFILLER_32_413 VPWR VGND sg13g2_fill_1
XFILLER_32_446 VPWR VGND sg13g2_decap_8
XFILLER_32_457 VPWR VGND sg13g2_fill_2
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_13_682 VPWR VGND sg13g2_decap_8
XFILLER_40_490 VPWR VGND sg13g2_decap_8
XFILLER_8_152 VPWR VGND sg13g2_decap_8
XFILLER_9_697 VPWR VGND sg13g2_decap_8
X_1602_ _0999_ net163 _0998_ VPWR VGND sg13g2_nand2_1
X_1395_ VPWR _0036_ state\[17\] VGND sg13g2_inv_1
X_1464_ net183 VPWR _0889_ VGND daisychain\[9\] net26 sg13g2_o21ai_1
X_1533_ VGND VPWR net104 daisychain\[22\] _0944_ net50 sg13g2_a21oi_1
Xfanout109 net114 net109 VPWR VGND sg13g2_buf_1
XFILLER_35_273 VPWR VGND sg13g2_decap_8
X_2016_ state\[120\] daisychain\[120\] net135 _0686_ VPWR VGND sg13g2_mux2_1
XFILLER_10_129 VPWR VGND sg13g2_decap_8
XFILLER_12_36 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_fill_2
XFILLER_23_446 VPWR VGND sg13g2_fill_1
XFILLER_18_229 VPWR VGND sg13g2_decap_8
XFILLER_19_708 VPWR VGND sg13g2_fill_1
XFILLER_26_251 VPWR VGND sg13g2_decap_8
XFILLER_26_262 VPWR VGND sg13g2_fill_2
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_22_490 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_5_111 VPWR VGND sg13g2_decap_8
XFILLER_6_601 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_5_188 VPWR VGND sg13g2_decap_8
XFILLER_18_785 VPWR VGND sg13g2_fill_2
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_17_295 VPWR VGND sg13g2_decap_8
XFILLER_20_405 VPWR VGND sg13g2_fill_2
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_4
XFILLER_33_788 VPWR VGND sg13g2_decap_4
XFILLER_33_799 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_1516_ state\[20\] daisychain\[20\] net139 _0930_ VPWR VGND sg13g2_mux2_1
X_2565_ net263 VGND VPWR _0381_ state\[125\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1378_ VPWR _0055_ state\[34\] VGND sg13g2_inv_1
X_1447_ _0875_ net161 _0874_ VPWR VGND sg13g2_nand2_1
X_2496_ net361 VGND VPWR _0312_ state\[56\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_23_221 VPWR VGND sg13g2_fill_1
XFILLER_23_265 VPWR VGND sg13g2_fill_1
XFILLER_11_438 VPWR VGND sg13g2_fill_1
XFILLER_23_13 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_14_254 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_fill_1
XFILLER_30_747 VPWR VGND sg13g2_fill_1
XFILLER_42_596 VPWR VGND sg13g2_fill_2
XFILLER_9_37 VPWR VGND sg13g2_fill_1
Xfanout91 net98 net91 VPWR VGND sg13g2_buf_1
Xfanout80 net83 net80 VPWR VGND sg13g2_buf_1
XFILLER_13_90 VPWR VGND sg13g2_decap_8
XFILLER_6_464 VPWR VGND sg13g2_decap_8
XFILLER_6_475 VPWR VGND sg13g2_fill_1
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_49_151 VPWR VGND sg13g2_decap_8
X_1301_ VPWR _0013_ state\[111\] VGND sg13g2_inv_1
Xclkbuf_leaf_1_clk clknet_2_1__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_2350_ net252 VGND VPWR _0166_ daisychain\[38\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2281_ VGND VPWR _0655_ _0830_ _0368_ net76 sg13g2_a21oi_1
XFILLER_25_519 VPWR VGND sg13g2_decap_8
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_20_257 VPWR VGND sg13g2_decap_8
XFILLER_9_280 VPWR VGND sg13g2_decap_8
X_1996_ state\[116\] daisychain\[116\] net134 _0670_ VPWR VGND sg13g2_mux2_1
X_2548_ net399 VGND VPWR _0364_ state\[108\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_18_13 VPWR VGND sg13g2_fill_1
XFILLER_18_68 VPWR VGND sg13g2_decap_8
X_2479_ net429 VGND VPWR _0295_ state\[39\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_11_213 VPWR VGND sg13g2_decap_8
XFILLER_34_89 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_2_3__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_19_302 VPWR VGND sg13g2_decap_8
XFILLER_3_456 VPWR VGND sg13g2_decap_8
XFILLER_15_530 VPWR VGND sg13g2_fill_1
XFILLER_34_327 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_47_666 VPWR VGND sg13g2_decap_8
X_2376__457 VPWR VGND net456 sg13g2_tiehi
XFILLER_42_371 VPWR VGND sg13g2_decap_8
X_1850_ VGND VPWR _0551_ _0552_ _0214_ _0553_ sg13g2_a21oi_1
X_1781_ state\[73\] daisychain\[73\] net153 _0498_ VPWR VGND sg13g2_mux2_1
XFILLER_10_290 VPWR VGND sg13g2_decap_8
XFILLER_6_261 VPWR VGND sg13g2_decap_8
XFILLER_7_773 VPWR VGND sg13g2_decap_8
X_2402_ net404 VGND VPWR _0218_ daisychain\[90\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2346__261 VPWR VGND net260 sg13g2_tiehi
X_2333_ net286 VGND VPWR _0149_ daisychain\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_37_154 VPWR VGND sg13g2_decap_8
X_2500__346 VPWR VGND net345 sg13g2_tiehi
X_2264_ _0822_ net110 state\[104\] VPWR VGND sg13g2_nand2_1
X_2195_ VGND VPWR _0483_ _0787_ _0325_ net86 sg13g2_a21oi_1
XFILLER_25_338 VPWR VGND sg13g2_fill_2
XFILLER_33_382 VPWR VGND sg13g2_decap_8
XFILLER_40_308 VPWR VGND sg13g2_decap_8
X_1979_ net187 VPWR _0657_ VGND daisychain\[112\] net30 sg13g2_o21ai_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_45 VPWR VGND sg13g2_decap_8
XFILLER_28_165 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv2 VPWR digitalen.g\[2\].u.OUTP digitalen.g\[2\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_31_319 VPWR VGND sg13g2_decap_4
XFILLER_10_80 VPWR VGND sg13g2_decap_8
XFILLER_3_253 VPWR VGND sg13g2_decap_8
XFILLER_20_8 VPWR VGND sg13g2_fill_2
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_176 VPWR VGND sg13g2_decap_8
XFILLER_34_124 VPWR VGND sg13g2_decap_8
X_1902_ _0595_ net167 _0594_ VPWR VGND sg13g2_nand2_1
X_1833_ VGND VPWR net125 daisychain\[82\] _0540_ net61 sg13g2_a21oi_1
X_1764_ net199 VPWR _0485_ VGND daisychain\[69\] net42 sg13g2_o21ai_1
X_2316_ net320 VGND VPWR _0132_ daisychain\[4\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1695_ VGND VPWR _0427_ _0428_ _0183_ _0429_ sg13g2_a21oi_1
XFILLER_25_102 VPWR VGND sg13g2_decap_4
XFILLER_25_124 VPWR VGND sg13g2_fill_2
X_2247_ VGND VPWR _0587_ _0813_ _0351_ net77 sg13g2_a21oi_1
X_2178_ _0779_ net122 state\[61\] VPWR VGND sg13g2_nand2_1
XFILLER_15_58 VPWR VGND sg13g2_decap_8
XFILLER_25_179 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_31_46 VPWR VGND sg13g2_decap_8
XFILLER_5_507 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_fill_1
Xoutput13 net13 uio_out[6] VPWR VGND sg13g2_buf_1
X_2507__308 VPWR VGND net307 sg13g2_tiehi
X_2442__322 VPWR VGND net321 sg13g2_tiehi
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_29_463 VPWR VGND sg13g2_decap_4
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_13_820 VPWR VGND sg13g2_fill_2
XFILLER_16_146 VPWR VGND sg13g2_decap_8
XFILLER_24_190 VPWR VGND sg13g2_decap_8
XFILLER_31_116 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_8_334 VPWR VGND sg13g2_decap_8
X_1480_ VGND VPWR _0899_ _0900_ _0140_ _0901_ sg13g2_a21oi_1
XFILLER_39_238 VPWR VGND sg13g2_decap_8
XFILLER_48_772 VPWR VGND sg13g2_fill_2
X_2101_ VGND VPWR _0939_ _0740_ _0278_ net73 sg13g2_a21oi_1
X_2032_ _0699_ net157 _0698_ VPWR VGND sg13g2_nand2_1
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_31_683 VPWR VGND sg13g2_decap_8
XFILLER_30_193 VPWR VGND sg13g2_decap_8
X_1816_ state\[80\] daisychain\[80\] net151 _0526_ VPWR VGND sg13g2_mux2_1
X_1747_ _0471_ net175 _0470_ VPWR VGND sg13g2_nand2_1
X_1678_ VGND VPWR net118 daisychain\[51\] _0416_ net59 sg13g2_a21oi_1
XFILLER_26_35 VPWR VGND sg13g2_decap_8
XFILLER_26_488 VPWR VGND sg13g2_fill_2
XFILLER_26_57 VPWR VGND sg13g2_decap_8
XFILLER_39_783 VPWR VGND sg13g2_fill_2
XFILLER_21_171 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_6_805 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_45_753 VPWR VGND sg13g2_decap_4
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_16_90 VPWR VGND sg13g2_decap_8
XFILLER_44_252 VPWR VGND sg13g2_decap_8
XFILLER_12_182 VPWR VGND sg13g2_decap_8
XFILLER_8_131 VPWR VGND sg13g2_decap_8
XFILLER_9_654 VPWR VGND sg13g2_fill_2
X_1532_ _0943_ net163 _0942_ VPWR VGND sg13g2_nand2_1
X_1601_ state\[37\] daisychain\[37\] net139 _0998_ VPWR VGND sg13g2_mux2_1
XFILLER_4_381 VPWR VGND sg13g2_decap_8
X_1394_ VPWR _0037_ state\[18\] VGND sg13g2_inv_1
X_1463_ VGND VPWR net101 daisychain\[8\] _0888_ net49 sg13g2_a21oi_1
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_36_720 VPWR VGND sg13g2_fill_1
XFILLER_36_764 VPWR VGND sg13g2_decap_8
XFILLER_36_775 VPWR VGND sg13g2_fill_2
X_2015_ VGND VPWR _0683_ _0684_ _0247_ _0685_ sg13g2_a21oi_1
XFILLER_10_108 VPWR VGND sg13g2_decap_8
XFILLER_2_329 VPWR VGND sg13g2_decap_8
X_2404__401 VPWR VGND net400 sg13g2_tiehi
XFILLER_18_208 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_5_167 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_17_274 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_712 VPWR VGND sg13g2_fill_2
XFILLER_33_745 VPWR VGND sg13g2_decap_8
X_2494__370 VPWR VGND net369 sg13g2_tiehi
XFILLER_20_439 VPWR VGND sg13g2_fill_2
XFILLER_32_277 VPWR VGND sg13g2_decap_8
X_2386__437 VPWR VGND net436 sg13g2_tiehi
X_1515_ VGND VPWR _0927_ _0928_ _0147_ _0929_ sg13g2_a21oi_1
X_2564_ net359 VGND VPWR _0380_ state\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2495_ net365 VGND VPWR _0311_ state\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1377_ VPWR _0056_ state\[35\] VGND sg13g2_inv_1
X_1446_ state\[6\] daisychain\[6\] net137 _0874_ VPWR VGND sg13g2_mux2_1
X_2473__454 VPWR VGND net453 sg13g2_tiehi
X_2356__241 VPWR VGND net240 sg13g2_tiehi
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_36_583 VPWR VGND sg13g2_fill_2
XFILLER_23_69 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_3_649 VPWR VGND sg13g2_decap_4
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_14_233 VPWR VGND sg13g2_decap_8
XFILLER_15_789 VPWR VGND sg13g2_decap_4
Xfanout92 net94 net92 VPWR VGND sg13g2_buf_1
Xfanout81 net82 net81 VPWR VGND sg13g2_buf_1
Xfanout70 net89 net70 VPWR VGND sg13g2_buf_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_6_443 VPWR VGND sg13g2_decap_8
XFILLER_2_671 VPWR VGND sg13g2_decap_8
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
X_1300_ VPWR _0014_ state\[112\] VGND sg13g2_inv_1
X_2280_ _0830_ net108 state\[112\] VPWR VGND sg13g2_nand2_1
XFILLER_25_509 VPWR VGND sg13g2_decap_4
XFILLER_20_236 VPWR VGND sg13g2_decap_8
X_1995_ VGND VPWR _0667_ _0668_ _0243_ _0669_ sg13g2_a21oi_1
X_1429_ net180 VPWR _0861_ VGND daisychain\[2\] net23 sg13g2_o21ai_1
X_2547_ net415 VGND VPWR _0363_ state\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2478_ net433 VGND VPWR _0294_ state\[38\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_18_47 VPWR VGND sg13g2_decap_8
XFILLER_11_269 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_fill_2
XFILLER_34_68 VPWR VGND sg13g2_decap_8
XFILLER_7_229 VPWR VGND sg13g2_decap_8
Xclkload1 VPWR clkload1/Y clknet_leaf_3_clk VGND sg13g2_inv_1
XFILLER_20_781 VPWR VGND sg13g2_fill_1
XFILLER_3_435 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_34_306 VPWR VGND sg13g2_decap_8
XFILLER_34_339 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_30_567 VPWR VGND sg13g2_fill_1
XFILLER_30_589 VPWR VGND sg13g2_fill_1
XFILLER_6_240 VPWR VGND sg13g2_decap_8
X_1780_ VGND VPWR _0495_ _0496_ _0200_ _0497_ sg13g2_a21oi_1
XFILLER_2_490 VPWR VGND sg13g2_decap_8
X_2401_ net406 VGND VPWR _0217_ daisychain\[89\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2332_ net288 VGND VPWR _0148_ daisychain\[20\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_25_317 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_38_601 VPWR VGND sg13g2_fill_1
X_2263_ VGND VPWR _0619_ _0821_ _0359_ net78 sg13g2_a21oi_1
X_2194_ _0787_ net130 state\[69\] VPWR VGND sg13g2_nand2_1
X_1978_ VGND VPWR net108 daisychain\[111\] _0656_ net53 sg13g2_a21oi_1
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_24 VPWR VGND sg13g2_decap_8
XFILLER_16_328 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_12_556 VPWR VGND sg13g2_decap_4
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_12_589 VPWR VGND sg13g2_fill_2
XFILLER_24_383 VPWR VGND sg13g2_decap_8
XFILLER_8_538 VPWR VGND sg13g2_decap_4
X_2412__385 VPWR VGND net384 sg13g2_tiehi
XFILLER_3_232 VPWR VGND sg13g2_decap_8
XFILLER_19_155 VPWR VGND sg13g2_decap_8
XFILLER_34_103 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_15_394 VPWR VGND sg13g2_decap_8
X_1901_ state\[97\] daisychain\[97\] net144 _0594_ VPWR VGND sg13g2_mux2_1
X_1832_ _0539_ net173 _0538_ VPWR VGND sg13g2_nand2_1
XFILLER_30_386 VPWR VGND sg13g2_decap_8
X_1763_ VGND VPWR net129 daisychain\[68\] _0484_ net62 sg13g2_a21oi_1
X_1694_ net194 VPWR _0429_ VGND daisychain\[55\] net37 sg13g2_o21ai_1
X_2315_ net322 VGND VPWR _0131_ daisychain\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2246_ _0813_ net111 state\[95\] VPWR VGND sg13g2_nand2_1
XFILLER_25_158 VPWR VGND sg13g2_decap_8
XFILLER_34_670 VPWR VGND sg13g2_decap_8
XFILLER_38_442 VPWR VGND sg13g2_decap_4
X_2470__210 VPWR VGND net209 sg13g2_tiehi
X_2177_ VGND VPWR _0447_ _0778_ _0316_ net82 sg13g2_a21oi_1
XFILLER_31_25 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_1_769 VPWR VGND sg13g2_fill_1
Xoutput14 net14 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_17_626 VPWR VGND sg13g2_fill_1
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_16_125 VPWR VGND sg13g2_decap_8
XFILLER_32_618 VPWR VGND sg13g2_fill_2
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_12_364 VPWR VGND sg13g2_decap_8
XFILLER_21_80 VPWR VGND sg13g2_decap_8
XFILLER_40_673 VPWR VGND sg13g2_decap_8
XFILLER_8_313 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_8
X_2100_ _0740_ net104 state\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_47_294 VPWR VGND sg13g2_decap_8
X_2315__323 VPWR VGND net322 sg13g2_tiehi
X_2031_ state\[123\] daisychain\[123\] net135 _0698_ VPWR VGND sg13g2_mux2_1
XFILLER_15_191 VPWR VGND sg13g2_decap_8
XFILLER_30_172 VPWR VGND sg13g2_decap_8
X_1815_ VGND VPWR _0523_ _0524_ _0207_ _0525_ sg13g2_a21oi_1
XFILLER_7_390 VPWR VGND sg13g2_decap_8
XFILLER_7_82 VPWR VGND sg13g2_decap_8
X_1746_ state\[66\] daisychain\[66\] net153 _0470_ VPWR VGND sg13g2_mux2_1
X_1677_ _0415_ net171 _0414_ VPWR VGND sg13g2_nand2_1
X_2396__417 VPWR VGND net416 sg13g2_tiehi
X_2229_ VGND VPWR _0551_ _0804_ _0342_ net85 sg13g2_a21oi_1
XFILLER_13_139 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_4
XFILLER_26_423 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_21_150 VPWR VGND sg13g2_decap_8
XFILLER_5_349 VPWR VGND sg13g2_decap_8
X_2366__221 VPWR VGND net220 sg13g2_tiehi
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_29_283 VPWR VGND sg13g2_decap_4
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_45_721 VPWR VGND sg13g2_decap_4
XFILLER_45_765 VPWR VGND sg13g2_fill_1
XFILLER_12_161 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_fill_2
XFILLER_32_459 VPWR VGND sg13g2_fill_1
XFILLER_8_110 VPWR VGND sg13g2_decap_8
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_8_187 VPWR VGND sg13g2_decap_8
X_1462_ _0887_ net161 _0886_ VPWR VGND sg13g2_nand2_1
X_1531_ state\[23\] daisychain\[23\] net139 _0942_ VPWR VGND sg13g2_mux2_1
X_1600_ VGND VPWR _0995_ _0996_ _0164_ _0997_ sg13g2_a21oi_1
XFILLER_27_209 VPWR VGND sg13g2_decap_8
X_1393_ VPWR _0038_ state\[19\] VGND sg13g2_inv_1
XFILLER_35_231 VPWR VGND sg13g2_decap_8
X_2014_ net181 VPWR _0685_ VGND daisychain\[119\] net24 sg13g2_o21ai_1
XFILLER_31_492 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
X_2847_ daisychain\[127\] net22 VPWR VGND sg13g2_buf_1
XFILLER_2_308 VPWR VGND sg13g2_decap_8
X_1729_ net195 VPWR _0457_ VGND daisychain\[62\] net38 sg13g2_o21ai_1
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_39_581 VPWR VGND sg13g2_fill_2
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_5_146 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_37_507 VPWR VGND sg13g2_fill_2
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_17_253 VPWR VGND sg13g2_decap_8
XFILLER_27_90 VPWR VGND sg13g2_decap_8
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_20_407 VPWR VGND sg13g2_fill_1
XFILLER_9_441 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_fill_1
XFILLER_4_94 VPWR VGND sg13g2_decap_8
X_1445_ VGND VPWR _0871_ _0872_ _0133_ _0873_ sg13g2_a21oi_1
X_1514_ net183 VPWR _0929_ VGND daisychain\[19\] net26 sg13g2_o21ai_1
X_2563_ net423 VGND VPWR _0379_ state\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2503__334 VPWR VGND net333 sg13g2_tiehi
X_2494_ net369 VGND VPWR _0310_ state\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1376_ VPWR _0057_ state\[36\] VGND sg13g2_inv_1
XFILLER_11_407 VPWR VGND sg13g2_fill_2
XFILLER_23_256 VPWR VGND sg13g2_fill_2
XFILLER_23_48 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
X_2480__426 VPWR VGND net425 sg13g2_tiehi
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_14_212 VPWR VGND sg13g2_decap_8
XFILLER_10_484 VPWR VGND sg13g2_decap_8
XFILLER_14_289 VPWR VGND sg13g2_decap_8
XFILLER_30_727 VPWR VGND sg13g2_fill_1
XFILLER_6_422 VPWR VGND sg13g2_decap_8
Xfanout93 net94 net93 VPWR VGND sg13g2_buf_1
Xfanout82 net83 net82 VPWR VGND sg13g2_buf_1
Xfanout71 net75 net71 VPWR VGND sg13g2_buf_1
Xfanout60 net65 net60 VPWR VGND sg13g2_buf_1
XFILLER_36_7 VPWR VGND sg13g2_decap_8
X_2422__365 VPWR VGND net364 sg13g2_tiehi
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_18_595 VPWR VGND sg13g2_decap_8
XFILLER_20_215 VPWR VGND sg13g2_decap_8
XFILLER_33_554 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
X_1994_ net181 VPWR _0669_ VGND daisychain\[115\] net24 sg13g2_o21ai_1
X_1428_ VGND VPWR net94 daisychain\[1\] _0860_ net45 sg13g2_a21oi_1
X_2546_ net431 VGND VPWR _0362_ state\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2477_ net437 VGND VPWR _0293_ state\[37\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
X_1359_ VPWR _0076_ state\[53\] VGND sg13g2_inv_1
XFILLER_11_248 VPWR VGND sg13g2_decap_8
XFILLER_20_760 VPWR VGND sg13g2_fill_1
XFILLER_20_793 VPWR VGND sg13g2_fill_1
XFILLER_34_47 VPWR VGND sg13g2_decap_8
XFILLER_7_208 VPWR VGND sg13g2_decap_8
Xclkload2 clkload2/Y clknet_leaf_10_clk VPWR VGND sg13g2_inv_2
X_2445__310 VPWR VGND net309 sg13g2_tiehi
XFILLER_3_414 VPWR VGND sg13g2_decap_8
XFILLER_35_819 VPWR VGND sg13g2_decap_4
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_47_646 VPWR VGND sg13g2_fill_2
XFILLER_27_392 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_6_296 VPWR VGND sg13g2_decap_8
X_2567__456 VPWR VGND net455 sg13g2_tiehi
X_2400_ net408 VGND VPWR _0216_ daisychain\[88\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2331_ net290 VGND VPWR _0147_ daisychain\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2262_ _0821_ net110 state\[103\] VPWR VGND sg13g2_nand2_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_38_668 VPWR VGND sg13g2_fill_2
X_2193_ VGND VPWR _0479_ _0786_ _0324_ net86 sg13g2_a21oi_1
XFILLER_21_502 VPWR VGND sg13g2_fill_2
XFILLER_21_535 VPWR VGND sg13g2_fill_2
X_1977_ _0655_ net165 _0654_ VPWR VGND sg13g2_nand2_1
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_20_27 VPWR VGND sg13g2_fill_2
X_2529_ net387 VGND VPWR _0345_ state\[89\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2325__303 VPWR VGND net302 sg13g2_tiehi
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_16_307 VPWR VGND sg13g2_decap_8
XFILLER_40_822 VPWR VGND sg13g2_fill_1
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_3_211 VPWR VGND sg13g2_decap_8
XFILLER_8_528 VPWR VGND sg13g2_decap_4
XFILLER_3_288 VPWR VGND sg13g2_decap_8
XFILLER_19_134 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_31_822 VPWR VGND sg13g2_fill_1
XFILLER_34_159 VPWR VGND sg13g2_decap_8
X_1900_ VGND VPWR _0591_ _0592_ _0224_ _0593_ sg13g2_a21oi_1
X_1831_ state\[83\] daisychain\[83\] net151 _0538_ VPWR VGND sg13g2_mux2_1
X_1762_ _0483_ net176 _0482_ VPWR VGND sg13g2_nand2_1
X_1693_ VGND VPWR net118 daisychain\[54\] _0428_ net59 sg13g2_a21oi_1
XFILLER_38_421 VPWR VGND sg13g2_fill_2
X_2314_ net324 VGND VPWR _0130_ daisychain\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2245_ VGND VPWR _0583_ _0812_ _0350_ net77 sg13g2_a21oi_1
X_2176_ _0778_ net120 state\[60\] VPWR VGND sg13g2_nand2_1
XFILLER_15_27 VPWR VGND sg13g2_decap_8
XFILLER_25_137 VPWR VGND sg13g2_decap_8
XFILLER_38_487 VPWR VGND sg13g2_decap_4
XFILLER_41_619 VPWR VGND sg13g2_fill_2
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_49_719 VPWR VGND sg13g2_fill_1
Xoutput15 net15 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_16_104 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_12_343 VPWR VGND sg13g2_decap_8
XFILLER_13_800 VPWR VGND sg13g2_fill_2
XFILLER_13_822 VPWR VGND sg13g2_fill_1
XFILLER_9_815 VPWR VGND sg13g2_decap_8
XFILLER_8_369 VPWR VGND sg13g2_decap_8
XFILLER_48_741 VPWR VGND sg13g2_decap_8
X_2030_ VGND VPWR _0695_ _0696_ _0250_ _0697_ sg13g2_a21oi_1
XFILLER_15_170 VPWR VGND sg13g2_decap_8
XFILLER_35_435 VPWR VGND sg13g2_decap_8
XFILLER_35_446 VPWR VGND sg13g2_fill_1
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_30_151 VPWR VGND sg13g2_decap_8
XFILLER_7_61 VPWR VGND sg13g2_decap_8
X_1814_ net199 VPWR _0525_ VGND daisychain\[79\] net42 sg13g2_o21ai_1
X_1745_ VGND VPWR _0467_ _0468_ _0193_ _0469_ sg13g2_a21oi_1
X_2541__256 VPWR VGND net255 sg13g2_tiehi
X_1676_ state\[52\] daisychain\[52\] net148 _0414_ VPWR VGND sg13g2_mux2_1
XFILLER_38_273 VPWR VGND sg13g2_decap_8
XFILLER_39_785 VPWR VGND sg13g2_fill_1
X_2476__442 VPWR VGND net441 sg13g2_tiehi
X_2228_ _0804_ net131 state\[86\] VPWR VGND sg13g2_nand2_1
X_2159_ VGND VPWR _0411_ _0769_ _0307_ net81 sg13g2_a21oi_1
XFILLER_13_118 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_5_328 VPWR VGND sg13g2_decap_8
XFILLER_29_262 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_12_140 VPWR VGND sg13g2_decap_8
XFILLER_13_674 VPWR VGND sg13g2_decap_4
XFILLER_13_696 VPWR VGND sg13g2_decap_8
XFILLER_8_166 VPWR VGND sg13g2_decap_8
X_1392_ VPWR _0040_ state\[20\] VGND sg13g2_inv_1
X_1461_ state\[9\] daisychain\[9\] net133 _0886_ VPWR VGND sg13g2_mux2_1
X_1530_ VGND VPWR _0939_ _0940_ _0150_ _0941_ sg13g2_a21oi_1
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
X_2013_ VGND VPWR net97 daisychain\[118\] _0684_ net46 sg13g2_a21oi_1
XFILLER_35_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_2_0__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_2432__345 VPWR VGND net344 sg13g2_tiehi
X_2846_ daisychain\[126\] net21 VPWR VGND sg13g2_buf_1
X_1728_ VGND VPWR net122 daisychain\[61\] _0456_ net60 sg13g2_a21oi_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
X_1659_ net195 VPWR _0401_ VGND daisychain\[48\] net38 sg13g2_o21ai_1
XFILLER_26_232 VPWR VGND sg13g2_fill_1
XFILLER_26_298 VPWR VGND sg13g2_decap_4
XFILLER_39_560 VPWR VGND sg13g2_fill_2
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_46_508 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_fill_2
XFILLER_6_626 VPWR VGND sg13g2_fill_1
X_2333__287 VPWR VGND net286 sg13g2_tiehi
XFILLER_2_810 VPWR VGND sg13g2_decap_8
XFILLER_2_821 VPWR VGND sg13g2_fill_2
XFILLER_5_125 VPWR VGND sg13g2_decap_8
XFILLER_6_659 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_17_232 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_fill_1
XFILLER_45_552 VPWR VGND sg13g2_decap_8
XFILLER_45_563 VPWR VGND sg13g2_fill_1
XFILLER_13_493 VPWR VGND sg13g2_fill_2
XFILLER_9_420 VPWR VGND sg13g2_decap_8
XFILLER_9_464 VPWR VGND sg13g2_fill_2
X_2562_ net231 VGND VPWR _0378_ state\[122\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_4_73 VPWR VGND sg13g2_decap_8
X_1375_ VPWR _0058_ state\[37\] VGND sg13g2_inv_1
X_1444_ net187 VPWR _0873_ VGND daisychain\[5\] net30 sg13g2_o21ai_1
X_1513_ VGND VPWR net99 daisychain\[18\] _0928_ net49 sg13g2_a21oi_1
Xclkbuf_leaf_4_clk clknet_2_3__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_2493_ net373 VGND VPWR _0309_ state\[53\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_596 VPWR VGND sg13g2_decap_4
XFILLER_23_27 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_14_268 VPWR VGND sg13g2_decap_8
XFILLER_30_706 VPWR VGND sg13g2_fill_1
XFILLER_30_739 VPWR VGND sg13g2_fill_1
XFILLER_42_544 VPWR VGND sg13g2_decap_4
XFILLER_42_555 VPWR VGND sg13g2_decap_4
XFILLER_6_401 VPWR VGND sg13g2_decap_8
Xfanout94 net98 net94 VPWR VGND sg13g2_buf_1
Xfanout83 net88 net83 VPWR VGND sg13g2_buf_1
Xfanout72 net75 net72 VPWR VGND sg13g2_buf_1
Xfanout61 net64 net61 VPWR VGND sg13g2_buf_1
Xfanout50 net52 net50 VPWR VGND sg13g2_buf_1
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_18_574 VPWR VGND sg13g2_fill_2
XFILLER_38_806 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
X_1993_ VGND VPWR net96 daisychain\[114\] _0668_ net46 sg13g2_a21oi_1
XFILLER_9_294 VPWR VGND sg13g2_decap_8
X_2545_ net447 VGND VPWR _0361_ state\[105\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_28_327 VPWR VGND sg13g2_fill_1
X_1358_ VPWR _0077_ state\[54\] VGND sg13g2_inv_1
X_1427_ _0859_ net158 _0858_ VPWR VGND sg13g2_nand2_1
X_2476_ net441 VGND VPWR _0292_ state\[36\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_44_809 VPWR VGND sg13g2_decap_8
X_1289_ VPWR _0026_ state\[123\] VGND sg13g2_inv_1
XFILLER_11_227 VPWR VGND sg13g2_decap_8
Xclkload3 clkload3/Y clknet_leaf_15_clk VPWR VGND sg13g2_inv_2
XFILLER_19_316 VPWR VGND sg13g2_decap_4
XFILLER_19_338 VPWR VGND sg13g2_fill_2
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_decap_4
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_11_794 VPWR VGND sg13g2_fill_2
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_6_275 VPWR VGND sg13g2_decap_8
X_2330_ net292 VGND VPWR _0146_ daisychain\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2261_ VGND VPWR _0615_ _0820_ _0358_ net78 sg13g2_a21oi_1
X_2192_ _0786_ net129 state\[68\] VPWR VGND sg13g2_nand2_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_33_396 VPWR VGND sg13g2_fill_2
X_1976_ state\[112\] daisychain\[112\] net142 _0654_ VPWR VGND sg13g2_mux2_1
X_2528_ net395 VGND VPWR _0344_ state\[88\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_29_59 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
X_2459_ net253 VGND VPWR _0275_ state\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_24_330 VPWR VGND sg13g2_decap_4
XFILLER_24_363 VPWR VGND sg13g2_fill_2
XFILLER_20_580 VPWR VGND sg13g2_fill_2
XFILLER_10_94 VPWR VGND sg13g2_decap_8
XFILLER_19_113 VPWR VGND sg13g2_decap_8
XFILLER_3_267 VPWR VGND sg13g2_decap_8
XFILLER_15_330 VPWR VGND sg13g2_decap_8
XFILLER_19_92 VPWR VGND sg13g2_decap_8
XFILLER_31_801 VPWR VGND sg13g2_decap_8
XFILLER_34_138 VPWR VGND sg13g2_decap_8
XFILLER_43_661 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
X_1830_ VGND VPWR _0535_ _0536_ _0210_ _0537_ sg13g2_a21oi_1
X_1761_ state\[69\] daisychain\[69\] net154 _0482_ VPWR VGND sg13g2_mux2_1
XFILLER_7_595 VPWR VGND sg13g2_fill_2
X_2313_ net326 VGND VPWR _0129_ daisychain\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1692_ _0427_ net171 _0426_ VPWR VGND sg13g2_nand2_1
X_2244_ _0812_ net111 state\[94\] VPWR VGND sg13g2_nand2_1
X_2175_ VGND VPWR _0443_ _0777_ _0315_ net82 sg13g2_a21oi_1
XFILLER_15_39 VPWR VGND sg13g2_fill_2
XFILLER_21_333 VPWR VGND sg13g2_decap_8
XFILLER_33_193 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_21_377 VPWR VGND sg13g2_fill_1
X_1959_ net187 VPWR _0641_ VGND daisychain\[108\] net30 sg13g2_o21ai_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_29_444 VPWR VGND sg13g2_decap_8
XFILLER_44_469 VPWR VGND sg13g2_decap_4
XFILLER_12_322 VPWR VGND sg13g2_decap_8
XFILLER_40_697 VPWR VGND sg13g2_decap_8
XFILLER_8_348 VPWR VGND sg13g2_decap_8
X_2343__267 VPWR VGND net266 sg13g2_tiehi
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_16_661 VPWR VGND sg13g2_fill_1
XFILLER_16_683 VPWR VGND sg13g2_decap_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
XFILLER_31_653 VPWR VGND sg13g2_decap_4
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_31_697 VPWR VGND sg13g2_fill_1
X_1813_ VGND VPWR net127 daisychain\[78\] _0524_ net63 sg13g2_a21oi_1
X_1744_ net199 VPWR _0469_ VGND daisychain\[65\] net42 sg13g2_o21ai_1
X_1675_ VGND VPWR _0411_ _0412_ _0179_ _0413_ sg13g2_a21oi_1
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_41_406 VPWR VGND sg13g2_decap_8
X_2227_ VGND VPWR _0547_ _0803_ _0341_ net85 sg13g2_a21oi_1
X_2158_ _0769_ net121 state\[51\] VPWR VGND sg13g2_nand2_1
X_2089_ VGND VPWR _0915_ _0734_ _0272_ net71 sg13g2_a21oi_1
XFILLER_21_185 VPWR VGND sg13g2_decap_8
XFILLER_41_428 VPWR VGND sg13g2_decap_4
XFILLER_41_439 VPWR VGND sg13g2_fill_1
XFILLER_6_819 VPWR VGND sg13g2_decap_4
X_2483__414 VPWR VGND net413 sg13g2_tiehi
XFILLER_5_307 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_4
XFILLER_29_241 VPWR VGND sg13g2_decap_8
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_12_196 VPWR VGND sg13g2_decap_8
XFILLER_13_664 VPWR VGND sg13g2_fill_1
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_40_461 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_8_145 VPWR VGND sg13g2_decap_8
X_2529__388 VPWR VGND net387 sg13g2_tiehi
XFILLER_4_395 VPWR VGND sg13g2_decap_8
X_1391_ VPWR _0041_ state\[21\] VGND sg13g2_inv_1
X_1460_ VGND VPWR _0883_ _0884_ _0136_ _0885_ sg13g2_a21oi_1
XFILLER_36_789 VPWR VGND sg13g2_fill_2
XFILLER_48_572 VPWR VGND sg13g2_fill_2
X_2012_ _0683_ net160 _0682_ VPWR VGND sg13g2_nand2_1
XFILLER_35_266 VPWR VGND sg13g2_decap_8
X_2845_ daisychain\[125\] net20 VPWR VGND sg13g2_buf_1
XFILLER_12_29 VPWR VGND sg13g2_decap_8
X_1727_ _0455_ net172 _0454_ VPWR VGND sg13g2_nand2_1
X_1658_ VGND VPWR net117 daisychain\[47\] _0400_ net60 sg13g2_a21oi_1
X_1589_ net192 VPWR _0989_ VGND daisychain\[34\] net35 sg13g2_o21ai_1
XFILLER_26_211 VPWR VGND sg13g2_decap_8
XFILLER_26_244 VPWR VGND sg13g2_decap_8
XFILLER_39_594 VPWR VGND sg13g2_fill_2
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_22_483 VPWR VGND sg13g2_decap_8
XFILLER_5_104 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_17_211 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_17_288 VPWR VGND sg13g2_decap_8
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
X_2312__328 VPWR VGND net327 sg13g2_tiehi
XFILLER_9_476 VPWR VGND sg13g2_decap_4
X_1512_ _0927_ net162 _0926_ VPWR VGND sg13g2_nand2_1
X_2561_ net295 VGND VPWR _0377_ state\[121\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2492_ net377 VGND VPWR _0308_ state\[52\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_4_192 VPWR VGND sg13g2_decap_8
X_1374_ VPWR _0059_ state\[38\] VGND sg13g2_inv_1
X_1443_ VGND VPWR net95 daisychain\[4\] _0872_ net46 sg13g2_a21oi_1
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_36_531 VPWR VGND sg13g2_fill_1
XFILLER_11_409 VPWR VGND sg13g2_fill_1
XFILLER_23_258 VPWR VGND sg13g2_fill_1
XFILLER_31_291 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_19_509 VPWR VGND sg13g2_decap_4
XFILLER_14_247 VPWR VGND sg13g2_decap_8
XFILLER_30_718 VPWR VGND sg13g2_fill_1
XFILLER_9_19 VPWR VGND sg13g2_fill_1
Xfanout73 net75 net73 VPWR VGND sg13g2_buf_1
Xfanout62 net63 net62 VPWR VGND sg13g2_buf_1
Xfanout51 net52 net51 VPWR VGND sg13g2_buf_1
Xfanout40 net43 net40 VPWR VGND sg13g2_buf_1
XFILLER_13_83 VPWR VGND sg13g2_decap_8
XFILLER_6_457 VPWR VGND sg13g2_decap_8
Xfanout95 net97 net95 VPWR VGND sg13g2_buf_1
Xfanout84 net88 net84 VPWR VGND sg13g2_buf_1
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_2_652 VPWR VGND sg13g2_decap_4
XFILLER_2_685 VPWR VGND sg13g2_fill_1
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_18_520 VPWR VGND sg13g2_fill_2
XFILLER_33_534 VPWR VGND sg13g2_fill_1
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_33_567 VPWR VGND sg13g2_fill_2
XFILLER_9_273 VPWR VGND sg13g2_decap_8
Xclkload10 VPWR clkload10/Y clknet_leaf_11_clk VGND sg13g2_inv_1
X_1992_ _0667_ net159 _0666_ VPWR VGND sg13g2_nand2_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2544_ net207 VGND VPWR _0360_ state\[104\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2475_ net445 VGND VPWR _0291_ state\[35\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2401__407 VPWR VGND net406 sg13g2_tiehi
XFILLER_28_306 VPWR VGND sg13g2_decap_4
X_1288_ VPWR _0027_ state\[124\] VGND sg13g2_inv_1
X_1357_ VPWR _0078_ state\[55\] VGND sg13g2_inv_1
X_1426_ state\[2\] daisychain\[2\] net133 _0858_ VPWR VGND sg13g2_mux2_1
XFILLER_11_206 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_20_773 VPWR VGND sg13g2_fill_1
Xclkload4 clkload4/Y clknet_leaf_16_clk VPWR VGND sg13g2_inv_2
XFILLER_3_449 VPWR VGND sg13g2_decap_8
XFILLER_15_523 VPWR VGND sg13g2_fill_1
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_30_559 VPWR VGND sg13g2_decap_4
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_10_283 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_6_254 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
X_2260_ _0820_ net110 state\[102\] VPWR VGND sg13g2_nand2_1
X_2191_ VGND VPWR _0475_ _0785_ _0323_ net86 sg13g2_a21oi_1
XFILLER_21_504 VPWR VGND sg13g2_fill_1
XFILLER_21_537 VPWR VGND sg13g2_fill_1
XFILLER_33_375 VPWR VGND sg13g2_decap_8
X_2353__247 VPWR VGND net246 sg13g2_tiehi
X_1975_ VGND VPWR _0651_ _0652_ _0239_ _0653_ sg13g2_a21oi_1
XFILLER_29_38 VPWR VGND sg13g2_decap_8
X_1409_ VPWR _0061_ state\[3\] VGND sg13g2_inv_1
X_2527_ net403 VGND VPWR _0343_ state\[87\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2479__430 VPWR VGND net429 sg13g2_tiehi
X_2458_ net257 VGND VPWR _0274_ state\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_28_158 VPWR VGND sg13g2_decap_8
X_2389_ net430 VGND VPWR _0205_ daisychain\[77\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_10_73 VPWR VGND sg13g2_decap_8
XFILLER_3_246 VPWR VGND sg13g2_decap_8
XFILLER_19_71 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_169 VPWR VGND sg13g2_decap_8
XFILLER_30_312 VPWR VGND sg13g2_fill_2
XFILLER_34_117 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_43_695 VPWR VGND sg13g2_decap_8
XFILLER_30_334 VPWR VGND sg13g2_fill_2
XFILLER_30_367 VPWR VGND sg13g2_fill_2
X_1760_ VGND VPWR _0479_ _0480_ _0196_ _0481_ sg13g2_a21oi_1
X_1691_ state\[55\] daisychain\[55\] net148 _0426_ VPWR VGND sg13g2_mux2_1
X_2312_ net327 VGND VPWR _0128_ daisychain\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_25_106 VPWR VGND sg13g2_fill_1
XFILLER_25_117 VPWR VGND sg13g2_decap_8
XFILLER_38_423 VPWR VGND sg13g2_fill_1
X_2243_ VGND VPWR _0579_ _0811_ _0349_ net78 sg13g2_a21oi_1
X_2174_ _0777_ net120 state\[59\] VPWR VGND sg13g2_nand2_1
XFILLER_18_180 VPWR VGND sg13g2_decap_8
XFILLER_33_172 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_decap_8
X_2511__276 VPWR VGND net275 sg13g2_tiehi
XFILLER_31_39 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[2] VPWR VGND sg13g2_buf_1
X_1958_ VGND VPWR net107 daisychain\[107\] _0640_ net53 sg13g2_a21oi_1
X_1889_ net189 VPWR _0585_ VGND daisychain\[94\] net32 sg13g2_o21ai_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_12_301 VPWR VGND sg13g2_decap_8
XFILLER_13_813 VPWR VGND sg13g2_decap_8
XFILLER_16_139 VPWR VGND sg13g2_decap_8
XFILLER_31_109 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_24_183 VPWR VGND sg13g2_decap_8
XFILLER_40_643 VPWR VGND sg13g2_fill_1
XFILLER_8_327 VPWR VGND sg13g2_decap_8
XFILLER_21_94 VPWR VGND sg13g2_decap_8
XFILLER_0_783 VPWR VGND sg13g2_fill_1
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_31_632 VPWR VGND sg13g2_decap_8
XFILLER_31_676 VPWR VGND sg13g2_decap_8
XFILLER_43_492 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_30_186 VPWR VGND sg13g2_decap_8
XFILLER_7_96 VPWR VGND sg13g2_decap_8
X_1812_ _0523_ net176 _0522_ VPWR VGND sg13g2_nand2_1
X_1743_ VGND VPWR net127 daisychain\[64\] _0468_ net63 sg13g2_a21oi_1
X_1674_ net194 VPWR _0413_ VGND daisychain\[51\] net37 sg13g2_o21ai_1
X_2226_ _0803_ net125 state\[85\] VPWR VGND sg13g2_nand2_1
XFILLER_38_231 VPWR VGND sg13g2_decap_8
X_2157_ VGND VPWR _0407_ _0768_ _0306_ net81 sg13g2_a21oi_1
X_2088_ _0734_ net99 state\[16\] VPWR VGND sg13g2_nand2_1
XFILLER_21_164 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_29_220 VPWR VGND sg13g2_decap_8
XFILLER_45_746 VPWR VGND sg13g2_fill_2
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_16_83 VPWR VGND sg13g2_decap_8
XFILLER_32_418 VPWR VGND sg13g2_fill_1
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_12_175 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_8_124 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
X_1390_ VPWR _0042_ state\[22\] VGND sg13g2_inv_1
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_36_735 VPWR VGND sg13g2_fill_2
X_2011_ state\[119\] daisychain\[119\] net136 _0682_ VPWR VGND sg13g2_mux2_1
XFILLER_31_473 VPWR VGND sg13g2_decap_8
X_2844_ daisychain\[124\] net19 VPWR VGND sg13g2_buf_1
X_1726_ state\[62\] daisychain\[62\] net149 _0454_ VPWR VGND sg13g2_mux2_1
X_1657_ _0399_ net172 _0398_ VPWR VGND sg13g2_nand2_1
X_1588_ VGND VPWR net103 daisychain\[33\] _0988_ net57 sg13g2_a21oi_1
XFILLER_37_49 VPWR VGND sg13g2_decap_8
X_2209_ VGND VPWR _0511_ _0794_ _0332_ net86 sg13g2_a21oi_1
XFILLER_14_418 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_10_657 VPWR VGND sg13g2_fill_1
XFILLER_10_679 VPWR VGND sg13g2_fill_2
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_17_267 VPWR VGND sg13g2_decap_8
XFILLER_18_724 VPWR VGND sg13g2_fill_2
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_41_760 VPWR VGND sg13g2_decap_4
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_4_171 VPWR VGND sg13g2_decap_8
XFILLER_5_694 VPWR VGND sg13g2_decap_8
X_1442_ _0871_ net159 _0870_ VPWR VGND sg13g2_nand2_1
X_1511_ state\[19\] daisychain\[19\] net137 _0926_ VPWR VGND sg13g2_mux2_1
X_2560_ net343 VGND VPWR _0376_ state\[120\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2491_ net381 VGND VPWR _0307_ state\[51\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1373_ VPWR _0060_ state\[39\] VGND sg13g2_inv_1
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_31_270 VPWR VGND sg13g2_decap_8
XFILLER_3_609 VPWR VGND sg13g2_fill_2
X_2363__227 VPWR VGND net226 sg13g2_tiehi
XFILLER_2_119 VPWR VGND sg13g2_decap_8
X_2408__393 VPWR VGND net392 sg13g2_tiehi
X_1709_ net195 VPWR _0441_ VGND daisychain\[58\] net38 sg13g2_o21ai_1
XFILLER_27_532 VPWR VGND sg13g2_decap_4
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_14_226 VPWR VGND sg13g2_decap_8
Xfanout30 net34 net30 VPWR VGND sg13g2_buf_1
Xfanout96 net97 net96 VPWR VGND sg13g2_buf_1
Xfanout85 net88 net85 VPWR VGND sg13g2_buf_1
Xfanout74 net75 net74 VPWR VGND sg13g2_buf_1
Xfanout63 net64 net63 VPWR VGND sg13g2_buf_1
Xfanout52 net66 net52 VPWR VGND sg13g2_buf_1
Xfanout41 net42 net41 VPWR VGND sg13g2_buf_1
XFILLER_13_62 VPWR VGND sg13g2_decap_8
XFILLER_6_436 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_4
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_20_229 VPWR VGND sg13g2_decap_8
XFILLER_9_252 VPWR VGND sg13g2_decap_8
Xclkload11 clkload11/Y clknet_leaf_4_clk VPWR VGND sg13g2_inv_2
X_1991_ state\[115\] daisychain\[115\] net134 _0666_ VPWR VGND sg13g2_mux2_1
X_1425_ VGND VPWR _0855_ _0856_ _0129_ _0857_ sg13g2_a21oi_1
X_2543_ net223 VGND VPWR _0359_ state\[103\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2474_ net449 VGND VPWR _0290_ state\[34\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_24_502 VPWR VGND sg13g2_fill_1
X_1287_ VPWR _0028_ state\[125\] VGND sg13g2_inv_1
X_1356_ VPWR _0079_ state\[56\] VGND sg13g2_inv_1
XFILLER_20_752 VPWR VGND sg13g2_fill_1
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_36_395 VPWR VGND sg13g2_decap_8
X_2514__252 VPWR VGND net251 sg13g2_tiehi
Xclkload5 clkload5/Y clknet_leaf_0_clk VPWR VGND sg13g2_inv_8
XFILLER_20_785 VPWR VGND sg13g2_decap_4
XFILLER_3_428 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_27_351 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_43_822 VPWR VGND sg13g2_fill_1
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_10_262 VPWR VGND sg13g2_decap_8
XFILLER_11_763 VPWR VGND sg13g2_fill_1
XFILLER_6_233 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_18_351 VPWR VGND sg13g2_decap_4
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
X_2190_ _0785_ net129 state\[67\] VPWR VGND sg13g2_nand2_1
XFILLER_21_516 VPWR VGND sg13g2_fill_1
XFILLER_33_398 VPWR VGND sg13g2_fill_1
X_1974_ net188 VPWR _0653_ VGND daisychain\[111\] net31 sg13g2_o21ai_1
XFILLER_29_17 VPWR VGND sg13g2_decap_8
X_1408_ VPWR _0072_ state\[4\] VGND sg13g2_inv_1
X_2526_ net411 VGND VPWR _0342_ state\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2457_ net261 VGND VPWR _0273_ state\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2388_ net432 VGND VPWR _0204_ daisychain\[76\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_37_682 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
X_1339_ VPWR _0098_ state\[73\] VGND sg13g2_inv_1
X_2486__402 VPWR VGND net401 sg13g2_tiehi
XFILLER_10_52 VPWR VGND sg13g2_decap_8
XFILLER_3_225 VPWR VGND sg13g2_decap_8
XFILLER_19_148 VPWR VGND sg13g2_decap_8
XFILLER_19_50 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_15_387 VPWR VGND sg13g2_decap_8
XFILLER_16_811 VPWR VGND sg13g2_decap_8
XFILLER_16_822 VPWR VGND sg13g2_fill_1
XFILLER_27_181 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_30_379 VPWR VGND sg13g2_decap_8
XFILLER_7_597 VPWR VGND sg13g2_fill_1
X_1690_ VGND VPWR _0423_ _0424_ _0182_ _0425_ sg13g2_a21oi_1
XFILLER_2_280 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_38_402 VPWR VGND sg13g2_decap_4
X_2311_ VGND VPWR _0715_ _0845_ _0383_ net70 sg13g2_a21oi_1
X_2242_ _0811_ net113 state\[93\] VPWR VGND sg13g2_nand2_1
XFILLER_38_435 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
X_2173_ VGND VPWR _0439_ _0776_ _0314_ net82 sg13g2_a21oi_1
XFILLER_31_18 VPWR VGND sg13g2_decap_8
XFILLER_33_151 VPWR VGND sg13g2_decap_8
XFILLER_34_663 VPWR VGND sg13g2_decap_8
X_1957_ _0639_ net165 _0638_ VPWR VGND sg13g2_nand2_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[3] VPWR VGND sg13g2_buf_1
X_2509_ net291 VGND VPWR _0325_ state\[69\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1888_ VGND VPWR net113 daisychain\[93\] _0584_ net55 sg13g2_a21oi_1
XFILLER_29_435 VPWR VGND sg13g2_decap_4
XFILLER_16_118 VPWR VGND sg13g2_decap_8
XFILLER_24_162 VPWR VGND sg13g2_decap_8
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_12_357 VPWR VGND sg13g2_decap_8
XFILLER_21_73 VPWR VGND sg13g2_decap_8
XFILLER_40_666 VPWR VGND sg13g2_decap_8
XFILLER_8_306 VPWR VGND sg13g2_decap_8
XFILLER_48_711 VPWR VGND sg13g2_fill_2
XFILLER_16_652 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_15_184 VPWR VGND sg13g2_decap_8
XFILLER_30_165 VPWR VGND sg13g2_decap_8
X_1811_ state\[79\] daisychain\[79\] net154 _0522_ VPWR VGND sg13g2_mux2_1
XFILLER_7_383 VPWR VGND sg13g2_decap_8
XFILLER_7_75 VPWR VGND sg13g2_decap_8
X_2322__309 VPWR VGND net308 sg13g2_tiehi
X_1742_ _0467_ net176 _0466_ VPWR VGND sg13g2_nand2_1
X_1673_ VGND VPWR net118 daisychain\[50\] _0412_ net59 sg13g2_a21oi_1
XFILLER_38_210 VPWR VGND sg13g2_decap_8
X_2225_ VGND VPWR _0543_ _0802_ _0340_ net85 sg13g2_a21oi_1
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_26_29 VPWR VGND sg13g2_fill_1
XFILLER_38_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_2_1__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_2156_ _0768_ net118 state\[50\] VPWR VGND sg13g2_nand2_1
X_2087_ VGND VPWR _0911_ _0733_ _0271_ net71 sg13g2_a21oi_1
XFILLER_21_143 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_29_276 VPWR VGND sg13g2_decap_8
XFILLER_29_287 VPWR VGND sg13g2_fill_2
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_45_725 VPWR VGND sg13g2_fill_1
X_2418__373 VPWR VGND net372 sg13g2_tiehi
X_2373__207 VPWR VGND net206 sg13g2_tiehi
XFILLER_12_154 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_16_62 VPWR VGND sg13g2_decap_8
XFILLER_25_471 VPWR VGND sg13g2_decap_8
XFILLER_8_103 VPWR VGND sg13g2_decap_8
XFILLER_4_353 VPWR VGND sg13g2_decap_8
X_2010_ VGND VPWR _0679_ _0680_ _0246_ _0681_ sg13g2_a21oi_1
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_31_485 VPWR VGND sg13g2_decap_8
XFILLER_8_681 VPWR VGND sg13g2_fill_2
XFILLER_8_692 VPWR VGND sg13g2_decap_8
X_2843_ daisychain\[123\] net18 VPWR VGND sg13g2_buf_1
X_1725_ VGND VPWR _0451_ _0452_ _0189_ _0453_ sg13g2_a21oi_1
XFILLER_7_180 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_7_clk clknet_2_3__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_1656_ state\[48\] daisychain\[48\] net149 _0398_ VPWR VGND sg13g2_mux2_1
X_1587_ _0987_ net169 _0986_ VPWR VGND sg13g2_nand2_1
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_39_596 VPWR VGND sg13g2_fill_1
X_2208_ _0794_ net128 state\[76\] VPWR VGND sg13g2_nand2_1
X_2139_ VGND VPWR _1015_ _0759_ _0297_ net80 sg13g2_a21oi_1
XFILLER_35_791 VPWR VGND sg13g2_fill_2
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_17_246 VPWR VGND sg13g2_decap_8
XFILLER_27_83 VPWR VGND sg13g2_decap_8
XFILLER_32_249 VPWR VGND sg13g2_decap_8
XFILLER_9_434 VPWR VGND sg13g2_decap_8
XFILLER_4_10 VPWR VGND sg13g2_fill_1
XFILLER_4_150 VPWR VGND sg13g2_decap_8
X_1441_ state\[5\] daisychain\[5\] net134 _0870_ VPWR VGND sg13g2_mux2_1
X_1510_ VGND VPWR _0923_ _0924_ _0146_ _0925_ sg13g2_a21oi_1
X_2490_ net385 VGND VPWR _0306_ state\[50\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_4_87 VPWR VGND sg13g2_decap_8
X_1372_ VPWR _0062_ state\[40\] VGND sg13g2_inv_1
X_1708_ VGND VPWR net119 daisychain\[57\] _0440_ net59 sg13g2_a21oi_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_1639_ net193 VPWR _0385_ VGND daisychain\[44\] net36 sg13g2_o21ai_1
XFILLER_14_205 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_6_415 VPWR VGND sg13g2_decap_8
Xfanout31 net34 net31 VPWR VGND sg13g2_buf_1
Xfanout97 net98 net97 VPWR VGND sg13g2_buf_1
Xfanout86 net87 net86 VPWR VGND sg13g2_buf_1
Xfanout75 net89 net75 VPWR VGND sg13g2_buf_1
Xfanout64 net65 net64 VPWR VGND sg13g2_buf_1
Xfanout53 net56 net53 VPWR VGND sg13g2_buf_1
Xfanout42 net43 net42 VPWR VGND sg13g2_buf_1
XFILLER_2_632 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_20_208 VPWR VGND sg13g2_decap_8
XFILLER_33_547 VPWR VGND sg13g2_decap_8
XFILLER_33_569 VPWR VGND sg13g2_fill_1
XFILLER_45_385 VPWR VGND sg13g2_decap_8
X_1990_ VGND VPWR _0663_ _0664_ _0242_ _0665_ sg13g2_a21oi_1
XFILLER_13_293 VPWR VGND sg13g2_decap_8
XFILLER_41_591 VPWR VGND sg13g2_decap_8
XFILLER_9_231 VPWR VGND sg13g2_decap_8
X_2542_ net239 VGND VPWR _0358_ state\[102\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_5_470 VPWR VGND sg13g2_fill_1
X_1355_ VPWR _0080_ state\[57\] VGND sg13g2_inv_1
X_1424_ net180 VPWR _0857_ VGND daisychain\[1\] net23 sg13g2_o21ai_1
X_2473_ net453 VGND VPWR _0289_ state\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_36_385 VPWR VGND sg13g2_decap_4
XFILLER_49_680 VPWR VGND sg13g2_decap_4
X_1286_ VPWR _0029_ state\[126\] VGND sg13g2_inv_1
XFILLER_20_731 VPWR VGND sg13g2_fill_1
XFILLER_20_764 VPWR VGND sg13g2_fill_2
Xclkload6 VPWR clkload6/Y clknet_leaf_2_clk VGND sg13g2_inv_1
XFILLER_3_407 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
X_2532__364 VPWR VGND net363 sg13g2_tiehi
XFILLER_10_241 VPWR VGND sg13g2_decap_8
XFILLER_11_775 VPWR VGND sg13g2_decap_4
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_6_212 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_2_462 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_6_289 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_decap_8
X_1973_ VGND VPWR net109 daisychain\[110\] _0652_ net56 sg13g2_a21oi_1
X_2525_ net419 VGND VPWR _0341_ state\[85\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_116 VPWR VGND sg13g2_decap_8
X_1338_ VPWR _0099_ state\[74\] VGND sg13g2_inv_1
X_1407_ VPWR _0083_ state\[5\] VGND sg13g2_inv_1
X_2456_ net265 VGND VPWR _0272_ state\[16\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2387_ net434 VGND VPWR _0203_ daisychain\[75\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_40_815 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_12_539 VPWR VGND sg13g2_fill_2
XFILLER_20_572 VPWR VGND sg13g2_fill_1
XFILLER_10_31 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_decap_8
X_2382__445 VPWR VGND net444 sg13g2_tiehi
XFILLER_19_127 VPWR VGND sg13g2_decap_8
XFILLER_27_160 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_15_344 VPWR VGND sg13g2_fill_2
XFILLER_30_314 VPWR VGND sg13g2_fill_1
XFILLER_31_815 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_43_675 VPWR VGND sg13g2_decap_8
XFILLER_11_561 VPWR VGND sg13g2_fill_2
X_2428__353 VPWR VGND net352 sg13g2_tiehi
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_fill_2
X_2310_ _0845_ state\[127\] net91 VPWR VGND sg13g2_nand2_1
X_2241_ VGND VPWR _0575_ _0810_ _0348_ net84 sg13g2_a21oi_1
X_2172_ _0776_ net120 state\[58\] VPWR VGND sg13g2_nand2_1
XFILLER_33_130 VPWR VGND sg13g2_decap_8
X_1956_ state\[108\] daisychain\[108\] net142 _0638_ VPWR VGND sg13g2_mux2_1
X_1887_ _0583_ net166 _0582_ VPWR VGND sg13g2_nand2_1
Xoutput19 net19 uo_out[4] VPWR VGND sg13g2_buf_1
X_2508_ net299 VGND VPWR _0324_ state\[68\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2329__295 VPWR VGND net294 sg13g2_tiehi
XFILLER_44_406 VPWR VGND sg13g2_decap_8
X_2439_ net330 VGND VPWR _0255_ daisychain\[127\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_12_336 VPWR VGND sg13g2_decap_8
XFILLER_40_612 VPWR VGND sg13g2_fill_2
XFILLER_40_623 VPWR VGND sg13g2_fill_2
XFILLER_9_808 VPWR VGND sg13g2_decap_8
XFILLER_20_391 VPWR VGND sg13g2_decap_8
XFILLER_21_30 VPWR VGND sg13g2_decap_8
XFILLER_21_52 VPWR VGND sg13g2_decap_8
XFILLER_35_428 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_15_163 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_decap_8
XFILLER_30_144 VPWR VGND sg13g2_decap_8
XFILLER_7_43 VPWR VGND sg13g2_fill_1
XFILLER_7_54 VPWR VGND sg13g2_decap_8
X_1810_ VGND VPWR _0519_ _0520_ _0206_ _0521_ sg13g2_a21oi_1
X_1741_ state\[65\] daisychain\[65\] net154 _0466_ VPWR VGND sg13g2_mux2_1
XFILLER_7_362 VPWR VGND sg13g2_decap_8
X_1672_ _0411_ net171 _0410_ VPWR VGND sg13g2_nand2_1
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_39_767 VPWR VGND sg13g2_decap_4
X_2224_ _0802_ net124 state\[84\] VPWR VGND sg13g2_nand2_1
X_2155_ VGND VPWR _0403_ _0767_ _0305_ net82 sg13g2_a21oi_1
XFILLER_21_122 VPWR VGND sg13g2_decap_8
XFILLER_26_439 VPWR VGND sg13g2_fill_1
X_2086_ _0733_ net101 state\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_21_199 VPWR VGND sg13g2_decap_8
X_1939_ net189 VPWR _0625_ VGND daisychain\[104\] net32 sg13g2_o21ai_1
XFILLER_17_406 VPWR VGND sg13g2_fill_2
XFILLER_29_255 VPWR VGND sg13g2_decap_8
XFILLER_44_203 VPWR VGND sg13g2_decap_8
XFILLER_45_748 VPWR VGND sg13g2_fill_1
XFILLER_12_133 VPWR VGND sg13g2_decap_8
XFILLER_13_689 VPWR VGND sg13g2_decap_8
XFILLER_25_494 VPWR VGND sg13g2_decap_8
XFILLER_40_475 VPWR VGND sg13g2_decap_4
XFILLER_40_497 VPWR VGND sg13g2_fill_2
XFILLER_8_159 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_5_822 VPWR VGND sg13g2_fill_1
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
X_2842_ daisychain\[122\] net17 VPWR VGND sg13g2_buf_1
X_1724_ net195 VPWR _0453_ VGND daisychain\[61\] net38 sg13g2_o21ai_1
X_1655_ VGND VPWR _0395_ _0396_ _0175_ _0397_ sg13g2_a21oi_1
X_1586_ state\[34\] daisychain\[34\] net139 _0986_ VPWR VGND sg13g2_mux2_1
XFILLER_26_225 VPWR VGND sg13g2_decap_8
XFILLER_26_258 VPWR VGND sg13g2_decap_4
XFILLER_39_553 VPWR VGND sg13g2_decap_8
X_2207_ VGND VPWR _0507_ _0793_ _0331_ net84 sg13g2_a21oi_1
X_2138_ _0759_ net115 state\[41\] VPWR VGND sg13g2_nand2_1
X_2069_ VGND VPWR _0875_ _0724_ _0262_ net71 sg13g2_a21oi_1
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_22_497 VPWR VGND sg13g2_fill_2
XFILLER_35_770 VPWR VGND sg13g2_fill_2
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_6_608 VPWR VGND sg13g2_fill_2
XFILLER_5_118 VPWR VGND sg13g2_decap_8
XFILLER_6_619 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_17_225 VPWR VGND sg13g2_decap_8
XFILLER_27_62 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_fill_1
XFILLER_45_545 VPWR VGND sg13g2_decap_8
X_2535__340 VPWR VGND net339 sg13g2_tiehi
XFILLER_13_486 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_41_795 VPWR VGND sg13g2_fill_1
XFILLER_9_413 VPWR VGND sg13g2_decap_8
X_1371_ VPWR _0063_ state\[41\] VGND sg13g2_inv_1
X_1440_ VGND VPWR _0867_ _0868_ _0132_ _0869_ sg13g2_a21oi_1
XFILLER_36_523 VPWR VGND sg13g2_fill_2
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_17_781 VPWR VGND sg13g2_fill_2
XFILLER_36_589 VPWR VGND sg13g2_decap_8
X_1707_ _0439_ net172 _0438_ VPWR VGND sg13g2_nand2_1
X_1638_ VGND VPWR net115 daisychain\[43\] _0384_ net58 sg13g2_a21oi_1
XFILLER_27_501 VPWR VGND sg13g2_fill_1
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_1569_ net186 VPWR _0973_ VGND daisychain\[30\] net29 sg13g2_o21ai_1
XFILLER_42_548 VPWR VGND sg13g2_fill_2
XFILLER_42_559 VPWR VGND sg13g2_fill_1
XFILLER_10_423 VPWR VGND sg13g2_fill_2
XFILLER_13_42 VPWR VGND sg13g2_fill_2
XFILLER_13_97 VPWR VGND sg13g2_decap_8
Xfanout32 net34 net32 VPWR VGND sg13g2_buf_1
Xfanout98 net132 net98 VPWR VGND sg13g2_buf_1
Xfanout87 net88 net87 VPWR VGND sg13g2_buf_1
Xfanout76 net79 net76 VPWR VGND sg13g2_buf_1
Xfanout65 net66 net65 VPWR VGND sg13g2_buf_1
Xfanout54 net55 net54 VPWR VGND sg13g2_buf_1
Xfanout43 net44 net43 VPWR VGND sg13g2_buf_1
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
X_2392__425 VPWR VGND net424 sg13g2_tiehi
XFILLER_13_272 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_9_210 VPWR VGND sg13g2_decap_8
XFILLER_9_287 VPWR VGND sg13g2_decap_8
X_2541_ net255 VGND VPWR _0357_ state\[101\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2472_ net VGND VPWR _0288_ state\[32\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1285_ VPWR _0846_ net160 VGND sg13g2_inv_1
X_1354_ VPWR _0081_ state\[58\] VGND sg13g2_inv_1
X_1423_ VGND VPWR net94 daisychain\[0\] _0856_ net45 sg13g2_a21oi_1
X_2438__333 VPWR VGND net332 sg13g2_tiehi
XFILLER_24_537 VPWR VGND sg13g2_decap_8
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_20_710 VPWR VGND sg13g2_fill_1
Xclkload7 clknet_leaf_17_clk clkload7/Y VPWR VGND sg13g2_inv_4
Xfanout200 net201 net200 VPWR VGND sg13g2_buf_1
XFILLER_19_309 VPWR VGND sg13g2_decap_8
X_2339__275 VPWR VGND net274 sg13g2_tiehi
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_24_85 VPWR VGND sg13g2_fill_1
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_10_220 VPWR VGND sg13g2_decap_8
XFILLER_10_297 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_6_268 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_19_810 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_33_312 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_46_662 VPWR VGND sg13g2_fill_2
XFILLER_33_389 VPWR VGND sg13g2_decap_8
X_1972_ _0651_ net168 _0650_ VPWR VGND sg13g2_nand2_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2524_ net427 VGND VPWR _0340_ state\[84\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2455_ net269 VGND VPWR _0271_ state\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_37_651 VPWR VGND sg13g2_fill_2
X_1337_ VPWR _0100_ state\[75\] VGND sg13g2_inv_1
X_1406_ VPWR _0094_ state\[6\] VGND sg13g2_inv_1
X_2386_ net436 VGND VPWR _0202_ daisychain\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_24_334 VPWR VGND sg13g2_fill_1
XFILLER_24_356 VPWR VGND sg13g2_decap_8
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_10_87 VPWR VGND sg13g2_decap_8
XFILLER_15_323 VPWR VGND sg13g2_decap_8
XFILLER_19_106 VPWR VGND sg13g2_decap_8
XFILLER_19_85 VPWR VGND sg13g2_decap_8
XFILLER_43_621 VPWR VGND sg13g2_decap_8
XFILLER_43_654 VPWR VGND sg13g2_fill_2
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_11_551 VPWR VGND sg13g2_fill_1
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_fill_1
XFILLER_19_651 VPWR VGND sg13g2_decap_8
XFILLER_3_794 VPWR VGND sg13g2_fill_2
X_2240_ _0810_ net126 state\[92\] VPWR VGND sg13g2_nand2_1
X_2171_ VGND VPWR _0435_ _0775_ _0313_ net81 sg13g2_a21oi_1
XFILLER_18_194 VPWR VGND sg13g2_decap_8
XFILLER_19_673 VPWR VGND sg13g2_fill_2
XFILLER_21_326 VPWR VGND sg13g2_decap_8
XFILLER_33_186 VPWR VGND sg13g2_decap_8
XFILLER_34_610 VPWR VGND sg13g2_fill_2
X_1955_ VGND VPWR _0635_ _0636_ _0235_ _0637_ sg13g2_a21oi_1
X_1886_ state\[94\] daisychain\[94\] net143 _0582_ VPWR VGND sg13g2_mux2_1
X_2507_ net307 VGND VPWR _0323_ state\[67\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2438_ net332 VGND VPWR _0254_ daisychain\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_37_470 VPWR VGND sg13g2_fill_2
X_2369_ net214 VGND VPWR _0185_ daisychain\[57\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_12_315 VPWR VGND sg13g2_decap_8
XFILLER_24_197 VPWR VGND sg13g2_decap_8
XFILLER_0_753 VPWR VGND sg13g2_fill_2
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_48_713 VPWR VGND sg13g2_fill_1
XFILLER_15_142 VPWR VGND sg13g2_decap_8
XFILLER_16_676 VPWR VGND sg13g2_decap_8
XFILLER_28_481 VPWR VGND sg13g2_decap_8
XFILLER_35_418 VPWR VGND sg13g2_fill_2
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_11_381 VPWR VGND sg13g2_decap_8
XFILLER_30_123 VPWR VGND sg13g2_decap_8
XFILLER_31_646 VPWR VGND sg13g2_decap_8
XFILLER_31_657 VPWR VGND sg13g2_fill_2
XFILLER_7_341 VPWR VGND sg13g2_decap_8
X_1740_ VGND VPWR _0463_ _0464_ _0192_ _0465_ sg13g2_a21oi_1
X_1671_ state\[51\] daisychain\[51\] net148 _0410_ VPWR VGND sg13g2_mux2_1
XFILLER_38_245 VPWR VGND sg13g2_decap_8
X_2223_ VGND VPWR _0539_ _0801_ _0339_ net84 sg13g2_a21oi_1
X_2154_ _0767_ net122 state\[49\] VPWR VGND sg13g2_nand2_1
X_2085_ VGND VPWR _0907_ _0732_ _0270_ net68 sg13g2_a21oi_1
XFILLER_21_101 VPWR VGND sg13g2_decap_8
XFILLER_21_178 VPWR VGND sg13g2_decap_8
XFILLER_34_473 VPWR VGND sg13g2_fill_2
X_1938_ VGND VPWR net107 daisychain\[103\] _0624_ net55 sg13g2_a21oi_1
X_1869_ net196 VPWR _0569_ VGND daisychain\[90\] net39 sg13g2_o21ai_1
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_29_234 VPWR VGND sg13g2_decap_8
XFILLER_25_484 VPWR VGND sg13g2_fill_2
XFILLER_40_410 VPWR VGND sg13g2_fill_2
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_12_112 VPWR VGND sg13g2_decap_8
XFILLER_12_189 VPWR VGND sg13g2_decap_8
XFILLER_16_97 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_40_454 VPWR VGND sg13g2_decap_8
XFILLER_8_138 VPWR VGND sg13g2_decap_8
XFILLER_4_311 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_decap_8
X_2540__272 VPWR VGND net271 sg13g2_tiehi
X_2321__311 VPWR VGND net310 sg13g2_tiehi
XFILLER_0_594 VPWR VGND sg13g2_decap_8
XFILLER_36_716 VPWR VGND sg13g2_decap_4
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_31_432 VPWR VGND sg13g2_fill_2
XFILLER_35_259 VPWR VGND sg13g2_decap_8
X_2841_ daisychain\[121\] net16 VPWR VGND sg13g2_buf_1
X_1723_ VGND VPWR net120 daisychain\[60\] _0452_ net60 sg13g2_a21oi_1
X_1654_ net193 VPWR _0397_ VGND daisychain\[47\] net36 sg13g2_o21ai_1
XFILLER_39_543 VPWR VGND sg13g2_decap_4
X_2206_ _0793_ net125 state\[75\] VPWR VGND sg13g2_nand2_1
X_1585_ VGND VPWR _0983_ _0984_ _0161_ _0985_ sg13g2_a21oi_1
XFILLER_26_204 VPWR VGND sg13g2_decap_8
XFILLER_26_237 VPWR VGND sg13g2_decap_8
XFILLER_39_587 VPWR VGND sg13g2_decap_8
X_2137_ VGND VPWR _1011_ _0758_ _0296_ net80 sg13g2_a21oi_1
X_2068_ _0724_ net101 state\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_34_292 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_17_204 VPWR VGND sg13g2_decap_8
XFILLER_27_41 VPWR VGND sg13g2_decap_8
XFILLER_25_292 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_9_458 VPWR VGND sg13g2_fill_1
X_2349__255 VPWR VGND net254 sg13g2_tiehi
XFILLER_4_185 VPWR VGND sg13g2_decap_8
X_1370_ VPWR _0064_ state\[42\] VGND sg13g2_inv_1
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_31_284 VPWR VGND sg13g2_decap_8
X_1706_ state\[58\] daisychain\[58\] net149 _0438_ VPWR VGND sg13g2_mux2_1
X_1637_ _1027_ net170 _1026_ VPWR VGND sg13g2_nand2_1
X_1499_ net183 VPWR _0917_ VGND daisychain\[16\] net26 sg13g2_o21ai_1
X_1568_ VGND VPWR net105 daisychain\[29\] _0972_ net51 sg13g2_a21oi_1
XFILLER_10_402 VPWR VGND sg13g2_decap_8
Xfanout33 net34 net33 VPWR VGND sg13g2_buf_1
Xfanout55 net56 net55 VPWR VGND sg13g2_buf_1
Xfanout44 _0851_ net44 VPWR VGND sg13g2_buf_1
XFILLER_13_76 VPWR VGND sg13g2_decap_8
Xfanout99 net102 net99 VPWR VGND sg13g2_buf_1
Xfanout88 net89 net88 VPWR VGND sg13g2_buf_1
Xfanout77 net78 net77 VPWR VGND sg13g2_buf_1
Xfanout66 _0850_ net66 VPWR VGND sg13g2_buf_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_645 VPWR VGND sg13g2_decap_8
XFILLER_2_656 VPWR VGND sg13g2_fill_1
XFILLER_2_678 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_fill_1
XFILLER_13_251 VPWR VGND sg13g2_decap_8
XFILLER_9_266 VPWR VGND sg13g2_decap_8
XFILLER_5_461 VPWR VGND sg13g2_decap_8
X_1422_ _0855_ net158 _0854_ VPWR VGND sg13g2_nand2_1
X_2540_ net271 VGND VPWR _0356_ state\[100\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2471_ net205 VGND VPWR _0287_ state\[31\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1284_ VPWR _0030_ state\[127\] VGND sg13g2_inv_1
X_1353_ VPWR _0082_ state\[59\] VGND sg13g2_inv_1
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_20_744 VPWR VGND sg13g2_fill_1
XFILLER_20_777 VPWR VGND sg13g2_fill_1
XFILLER_32_582 VPWR VGND sg13g2_decap_8
Xclkload8 clkload8/Y clknet_leaf_18_clk VPWR VGND sg13g2_inv_8
Xfanout201 net1 net201 VPWR VGND sg13g2_buf_1
XFILLER_43_803 VPWR VGND sg13g2_fill_1
XFILLER_11_744 VPWR VGND sg13g2_fill_1
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_10_276 VPWR VGND sg13g2_decap_8
XFILLER_2_420 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_fill_2
XFILLER_6_247 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_2_497 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_46_696 VPWR VGND sg13g2_decap_8
X_1971_ state\[111\] daisychain\[111\] net145 _0650_ VPWR VGND sg13g2_mux2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_6_792 VPWR VGND sg13g2_decap_4
X_1405_ VPWR _0105_ state\[7\] VGND sg13g2_inv_1
X_2523_ net435 VGND VPWR _0339_ state\[83\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2454_ net273 VGND VPWR _0270_ state\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2405__399 VPWR VGND net398 sg13g2_tiehi
X_2385_ net438 VGND VPWR _0201_ daisychain\[73\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_37_641 VPWR VGND sg13g2_fill_2
XFILLER_37_663 VPWR VGND sg13g2_decap_8
XFILLER_37_674 VPWR VGND sg13g2_fill_2
X_1336_ VPWR _0101_ state\[76\] VGND sg13g2_inv_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
XFILLER_12_508 VPWR VGND sg13g2_decap_4
XFILLER_37_696 VPWR VGND sg13g2_fill_2
XFILLER_20_585 VPWR VGND sg13g2_fill_1
XFILLER_3_239 VPWR VGND sg13g2_decap_8
XFILLER_10_66 VPWR VGND sg13g2_decap_8
XFILLER_19_64 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_27_195 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_fill_1
XFILLER_11_563 VPWR VGND sg13g2_fill_1
XFILLER_11_585 VPWR VGND sg13g2_decap_4
XFILLER_30_305 VPWR VGND sg13g2_decap_8
XFILLER_7_556 VPWR VGND sg13g2_fill_1
XFILLER_7_589 VPWR VGND sg13g2_fill_2
XFILLER_2_294 VPWR VGND sg13g2_decap_8
X_2170_ _0775_ net119 state\[57\] VPWR VGND sg13g2_nand2_1
XFILLER_14_390 VPWR VGND sg13g2_decap_8
XFILLER_18_173 VPWR VGND sg13g2_decap_8
XFILLER_33_165 VPWR VGND sg13g2_decap_8
XFILLER_34_644 VPWR VGND sg13g2_decap_8
XFILLER_34_677 VPWR VGND sg13g2_fill_1
X_1954_ net187 VPWR _0637_ VGND daisychain\[107\] net30 sg13g2_o21ai_1
X_1885_ VGND VPWR _0579_ _0580_ _0221_ _0581_ sg13g2_a21oi_1
X_2506_ net315 VGND VPWR _0322_ state\[66\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2437_ net334 VGND VPWR _0253_ daisychain\[125\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2368_ net216 VGND VPWR _0184_ daisychain\[56\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_13_806 VPWR VGND sg13g2_decap_8
XFILLER_37_460 VPWR VGND sg13g2_fill_1
X_1319_ VPWR _0120_ state\[93\] VGND sg13g2_inv_1
X_2299_ VGND VPWR _0691_ _0839_ _0377_ net70 sg13g2_a21oi_1
XFILLER_24_176 VPWR VGND sg13g2_decap_8
XFILLER_40_636 VPWR VGND sg13g2_decap_8
XFILLER_21_87 VPWR VGND sg13g2_decap_8
XFILLER_4_537 VPWR VGND sg13g2_fill_2
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_15_121 VPWR VGND sg13g2_decap_8
XFILLER_15_198 VPWR VGND sg13g2_decap_8
XFILLER_30_102 VPWR VGND sg13g2_decap_8
XFILLER_31_603 VPWR VGND sg13g2_fill_2
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_43_485 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_11_360 VPWR VGND sg13g2_decap_8
XFILLER_30_179 VPWR VGND sg13g2_decap_8
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_7_397 VPWR VGND sg13g2_decap_8
XFILLER_7_89 VPWR VGND sg13g2_decap_8
X_2506__316 VPWR VGND net315 sg13g2_tiehi
X_1670_ VGND VPWR _0407_ _0408_ _0178_ _0409_ sg13g2_a21oi_1
XFILLER_30_4 VPWR VGND sg13g2_decap_4
X_2222_ _0801_ net131 state\[83\] VPWR VGND sg13g2_nand2_1
XFILLER_38_224 VPWR VGND sg13g2_decap_8
X_2552__336 VPWR VGND net335 sg13g2_tiehi
X_2359__235 VPWR VGND net234 sg13g2_tiehi
X_2153_ VGND VPWR _0399_ _0766_ _0304_ net82 sg13g2_a21oi_1
X_2084_ _0732_ net93 state\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_21_157 VPWR VGND sg13g2_decap_8
X_1937_ _0623_ net166 _0622_ VPWR VGND sg13g2_nand2_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
X_1868_ VGND VPWR net124 daisychain\[89\] _0568_ net64 sg13g2_a21oi_1
X_1799_ net198 VPWR _0513_ VGND daisychain\[76\] net41 sg13g2_o21ai_1
XFILLER_29_213 VPWR VGND sg13g2_decap_8
XFILLER_16_76 VPWR VGND sg13g2_decap_8
XFILLER_25_452 VPWR VGND sg13g2_fill_2
XFILLER_44_238 VPWR VGND sg13g2_decap_8
X_2453__278 VPWR VGND net277 sg13g2_tiehi
XFILLER_12_168 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_8_117 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_16_430 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_31_466 VPWR VGND sg13g2_decap_8
XFILLER_8_640 VPWR VGND sg13g2_fill_1
X_2547__416 VPWR VGND net415 sg13g2_tiehi
X_2840_ daisychain\[120\] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_194 VPWR VGND sg13g2_decap_8
X_1722_ _0451_ net172 _0450_ VPWR VGND sg13g2_nand2_1
X_1653_ VGND VPWR net117 daisychain\[46\] _0396_ net58 sg13g2_a21oi_1
X_1584_ net193 VPWR _0985_ VGND daisychain\[33\] net36 sg13g2_o21ai_1
XFILLER_39_500 VPWR VGND sg13g2_decap_4
X_2205_ VGND VPWR _0503_ _0792_ _0330_ net84 sg13g2_a21oi_1
XFILLER_34_271 VPWR VGND sg13g2_decap_8
XFILLER_35_772 VPWR VGND sg13g2_fill_1
X_2136_ _0758_ net115 state\[40\] VPWR VGND sg13g2_nand2_1
X_2067_ VGND VPWR _0871_ _0723_ _0261_ net67 sg13g2_a21oi_1
XFILLER_10_617 VPWR VGND sg13g2_fill_2
XFILLER_22_499 VPWR VGND sg13g2_fill_1
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_13_444 VPWR VGND sg13g2_decap_8
XFILLER_27_97 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_41_753 VPWR VGND sg13g2_decap_8
XFILLER_41_764 VPWR VGND sg13g2_fill_1
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_9_448 VPWR VGND sg13g2_decap_4
XFILLER_4_164 VPWR VGND sg13g2_decap_8
XFILLER_5_687 VPWR VGND sg13g2_fill_2
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_36_503 VPWR VGND sg13g2_fill_1
XFILLER_16_293 VPWR VGND sg13g2_decap_8
XFILLER_17_794 VPWR VGND sg13g2_fill_1
XFILLER_44_591 VPWR VGND sg13g2_fill_1
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_31_263 VPWR VGND sg13g2_decap_8
X_1705_ VGND VPWR _0435_ _0436_ _0185_ _0437_ sg13g2_a21oi_1
X_1636_ state\[44\] daisychain\[44\] net146 _1026_ VPWR VGND sg13g2_mux2_1
X_1567_ _0971_ net164 _0970_ VPWR VGND sg13g2_nand2_1
XFILLER_27_536 VPWR VGND sg13g2_fill_2
XFILLER_39_385 VPWR VGND sg13g2_decap_8
X_1498_ VGND VPWR net99 daisychain\[15\] _0916_ net49 sg13g2_a21oi_1
X_2119_ VGND VPWR _0975_ _0749_ _0287_ net74 sg13g2_a21oi_1
XFILLER_10_425 VPWR VGND sg13g2_fill_1
XFILLER_13_22 VPWR VGND sg13g2_fill_2
XFILLER_14_219 VPWR VGND sg13g2_decap_8
Xfanout23 net44 net23 VPWR VGND sg13g2_buf_1
Xfanout34 net44 net34 VPWR VGND sg13g2_buf_1
Xfanout89 _0847_ net89 VPWR VGND sg13g2_buf_1
Xfanout78 net79 net78 VPWR VGND sg13g2_buf_1
Xfanout67 net69 net67 VPWR VGND sg13g2_buf_1
Xfanout56 net66 net56 VPWR VGND sg13g2_buf_1
Xfanout45 net47 net45 VPWR VGND sg13g2_buf_1
X_2415__379 VPWR VGND net378 sg13g2_tiehi
XFILLER_13_55 VPWR VGND sg13g2_decap_8
XFILLER_6_429 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_fill_2
XFILLER_14_731 VPWR VGND sg13g2_decap_8
XFILLER_33_528 VPWR VGND sg13g2_fill_2
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_13_230 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_fill_1
XFILLER_9_245 VPWR VGND sg13g2_decap_8
XFILLER_5_440 VPWR VGND sg13g2_decap_8
X_1421_ state\[1\] daisychain\[1\] net133 _0854_ VPWR VGND sg13g2_mux2_1
X_2470_ net209 VGND VPWR _0286_ state\[30\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
X_1352_ VPWR _0084_ state\[60\] VGND sg13g2_inv_1
XFILLER_17_580 VPWR VGND sg13g2_fill_1
XFILLER_20_723 VPWR VGND sg13g2_fill_1
XFILLER_20_756 VPWR VGND sg13g2_fill_1
XFILLER_20_789 VPWR VGND sg13g2_fill_1
Xclkload9 clkload9/Y clknet_leaf_9_clk VPWR VGND sg13g2_inv_2
X_1619_ net192 VPWR _1013_ VGND daisychain\[40\] net35 sg13g2_o21ai_1
XFILLER_15_528 VPWR VGND sg13g2_fill_2
XFILLER_27_344 VPWR VGND sg13g2_decap_8
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_43_815 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_10_255 VPWR VGND sg13g2_decap_8
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_6_226 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_18_344 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_2_476 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_46_620 VPWR VGND sg13g2_fill_2
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_18_355 VPWR VGND sg13g2_fill_1
XFILLER_45_196 VPWR VGND sg13g2_decap_8
X_2318__317 VPWR VGND net316 sg13g2_tiehi
X_1970_ VGND VPWR _0647_ _0648_ _0238_ _0649_ sg13g2_a21oi_1
X_2522_ net443 VGND VPWR _0338_ state\[82\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1335_ VPWR _0102_ state\[77\] VGND sg13g2_inv_1
X_1404_ VPWR _0116_ state\[8\] VGND sg13g2_inv_1
X_2453_ net277 VGND VPWR _0269_ state\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2384_ net440 VGND VPWR _0200_ daisychain\[72\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_37_620 VPWR VGND sg13g2_fill_1
XFILLER_49_480 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_2369__215 VPWR VGND net214 sg13g2_tiehi
XFILLER_10_45 VPWR VGND sg13g2_fill_2
XFILLER_3_218 VPWR VGND sg13g2_decap_8
X_2449__294 VPWR VGND net293 sg13g2_tiehi
XFILLER_19_43 VPWR VGND sg13g2_fill_2
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_27_174 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_43_656 VPWR VGND sg13g2_fill_1
XFILLER_11_575 VPWR VGND sg13g2_decap_4
XFILLER_2_273 VPWR VGND sg13g2_decap_8
XFILLER_3_796 VPWR VGND sg13g2_fill_1
XFILLER_18_152 VPWR VGND sg13g2_decap_8
XFILLER_34_634 VPWR VGND sg13g2_decap_4
XFILLER_38_406 VPWR VGND sg13g2_fill_2
XFILLER_38_428 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_21_306 VPWR VGND sg13g2_decap_4
XFILLER_33_144 VPWR VGND sg13g2_decap_8
X_1953_ VGND VPWR net107 daisychain\[106\] _0636_ net53 sg13g2_a21oi_1
X_1884_ net189 VPWR _0581_ VGND daisychain\[93\] net32 sg13g2_o21ai_1
X_2505_ net323 VGND VPWR _0321_ state\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_29_439 VPWR VGND sg13g2_fill_1
X_1318_ VPWR _0121_ state\[94\] VGND sg13g2_inv_1
X_2436_ net336 VGND VPWR _0252_ daisychain\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2367_ net218 VGND VPWR _0183_ daisychain\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2298_ _0839_ net90 state\[121\] VPWR VGND sg13g2_nand2_1
XFILLER_24_155 VPWR VGND sg13g2_decap_8
XFILLER_20_372 VPWR VGND sg13g2_decap_4
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_40_659 VPWR VGND sg13g2_decap_8
XFILLER_0_755 VPWR VGND sg13g2_fill_1
XFILLER_21_66 VPWR VGND sg13g2_decap_8
XFILLER_15_100 VPWR VGND sg13g2_decap_8
XFILLER_16_623 VPWR VGND sg13g2_decap_4
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_48_748 VPWR VGND sg13g2_decap_4
XFILLER_15_177 VPWR VGND sg13g2_decap_8
XFILLER_16_645 VPWR VGND sg13g2_decap_8
XFILLER_30_158 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_8_822 VPWR VGND sg13g2_fill_1
XFILLER_7_376 VPWR VGND sg13g2_decap_8
XFILLER_7_68 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_4
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_3_582 VPWR VGND sg13g2_fill_2
X_2221_ VGND VPWR _0535_ _0800_ _0338_ net84 sg13g2_a21oi_1
X_2152_ _0766_ net122 state\[48\] VPWR VGND sg13g2_nand2_1
XFILLER_19_461 VPWR VGND sg13g2_decap_4
XFILLER_46_280 VPWR VGND sg13g2_decap_8
X_2083_ VGND VPWR _0903_ _0731_ _0269_ net68 sg13g2_a21oi_1
XFILLER_21_136 VPWR VGND sg13g2_decap_8
XFILLER_30_681 VPWR VGND sg13g2_fill_1
X_1936_ state\[104\] daisychain\[104\] net143 _0622_ VPWR VGND sg13g2_mux2_1
X_1867_ _0567_ net173 _0566_ VPWR VGND sg13g2_nand2_1
X_2524__428 VPWR VGND net427 sg13g2_tiehi
X_1798_ VGND VPWR net128 daisychain\[75\] _0512_ net62 sg13g2_a21oi_1
XFILLER_29_269 VPWR VGND sg13g2_decap_8
XFILLER_44_217 VPWR VGND sg13g2_decap_8
X_2419_ net370 VGND VPWR _0235_ daisychain\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_12_147 VPWR VGND sg13g2_decap_8
XFILLER_13_626 VPWR VGND sg13g2_fill_2
XFILLER_16_55 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_9_608 VPWR VGND sg13g2_decap_8
XFILLER_20_180 VPWR VGND sg13g2_decap_8
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_8
X_2425__359 VPWR VGND net358 sg13g2_tiehi
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_fill_1
XFILLER_16_497 VPWR VGND sg13g2_fill_2
XFILLER_43_294 VPWR VGND sg13g2_decap_8
X_1721_ state\[61\] daisychain\[61\] net149 _0450_ VPWR VGND sg13g2_mux2_1
XFILLER_7_173 VPWR VGND sg13g2_decap_8
X_1652_ _0395_ net170 _0394_ VPWR VGND sg13g2_nand2_1
X_1583_ VGND VPWR net105 daisychain\[32\] _0984_ net51 sg13g2_a21oi_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
X_2204_ _0792_ net125 state\[74\] VPWR VGND sg13g2_nand2_1
X_2135_ VGND VPWR _1007_ _0757_ _0295_ net80 sg13g2_a21oi_1
XFILLER_34_250 VPWR VGND sg13g2_decap_8
XFILLER_35_784 VPWR VGND sg13g2_decap_8
X_2066_ _0723_ net93 state\[5\] VPWR VGND sg13g2_nand2_1
X_1919_ net190 VPWR _0609_ VGND daisychain\[100\] net33 sg13g2_o21ai_1
XFILLER_2_817 VPWR VGND sg13g2_decap_4
XFILLER_17_239 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_4
XFILLER_27_76 VPWR VGND sg13g2_decap_8
XFILLER_45_559 VPWR VGND sg13g2_decap_4
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_41_776 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_decap_8
XFILLER_4_143 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_4
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_16_272 VPWR VGND sg13g2_decap_8
XFILLER_31_242 VPWR VGND sg13g2_decap_8
XFILLER_8_460 VPWR VGND sg13g2_decap_4
XFILLER_8_493 VPWR VGND sg13g2_decap_4
X_1704_ net194 VPWR _0437_ VGND daisychain\[57\] net37 sg13g2_o21ai_1
X_1497_ _0915_ net162 _0914_ VPWR VGND sg13g2_nand2_1
X_1635_ VGND VPWR _1023_ _1024_ _0171_ _1025_ sg13g2_a21oi_1
X_1566_ state\[30\] daisychain\[30\] net140 _0970_ VPWR VGND sg13g2_mux2_1
XFILLER_39_364 VPWR VGND sg13g2_decap_8
XFILLER_42_529 VPWR VGND sg13g2_fill_2
X_2378__453 VPWR VGND net452 sg13g2_tiehi
X_2118_ _0749_ net105 state\[31\] VPWR VGND sg13g2_nand2_1
X_2049_ net179 VPWR _0713_ VGND daisychain\[126\] net25 sg13g2_o21ai_1
XFILLER_22_264 VPWR VGND sg13g2_decap_8
XFILLER_6_408 VPWR VGND sg13g2_decap_8
Xfanout24 net44 net24 VPWR VGND sg13g2_buf_1
Xfanout79 net89 net79 VPWR VGND sg13g2_buf_1
Xfanout68 net69 net68 VPWR VGND sg13g2_buf_1
Xfanout57 net58 net57 VPWR VGND sg13g2_buf_1
Xfanout46 net47 net46 VPWR VGND sg13g2_buf_1
Xfanout35 net36 net35 VPWR VGND sg13g2_buf_1
XFILLER_2_625 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_13_286 VPWR VGND sg13g2_decap_8
XFILLER_14_776 VPWR VGND sg13g2_fill_1
XFILLER_14_787 VPWR VGND sg13g2_fill_2
XFILLER_41_584 VPWR VGND sg13g2_decap_8
XFILLER_9_224 VPWR VGND sg13g2_decap_8
X_1351_ VPWR _0085_ state\[61\] VGND sg13g2_inv_1
X_1420_ VGND VPWR _0849_ _0852_ _0128_ _0853_ sg13g2_a21oi_1
Xdigitalen.g\[1\].u.inv1 VPWR digitalen.g\[1\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_49_673 VPWR VGND sg13g2_decap_8
XFILLER_17_592 VPWR VGND sg13g2_fill_2
XFILLER_20_702 VPWR VGND sg13g2_fill_1
XFILLER_20_735 VPWR VGND sg13g2_fill_1
XFILLER_36_389 VPWR VGND sg13g2_fill_2
X_1618_ VGND VPWR net116 daisychain\[39\] _1012_ net57 sg13g2_a21oi_1
XFILLER_39_161 VPWR VGND sg13g2_decap_8
XFILLER_5_90 VPWR VGND sg13g2_decap_8
X_1549_ net184 VPWR _0957_ VGND daisychain\[26\] net27 sg13g2_o21ai_1
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_27_378 VPWR VGND sg13g2_decap_8
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_10_234 VPWR VGND sg13g2_decap_8
XFILLER_11_735 VPWR VGND sg13g2_fill_1
XFILLER_11_768 VPWR VGND sg13g2_decap_8
XFILLER_11_779 VPWR VGND sg13g2_fill_1
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_6_205 VPWR VGND sg13g2_decap_8
XFILLER_2_455 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_14_562 VPWR VGND sg13g2_decap_8
XFILLER_14_573 VPWR VGND sg13g2_decap_4
XFILLER_33_326 VPWR VGND sg13g2_fill_2
XFILLER_41_392 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
X_2521_ net451 VGND VPWR _0337_ state\[81\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_28_109 VPWR VGND sg13g2_decap_8
XFILLER_5_293 VPWR VGND sg13g2_decap_8
X_1334_ VPWR _0103_ state\[78\] VGND sg13g2_inv_1
X_1403_ VPWR _0127_ state\[9\] VGND sg13g2_inv_1
X_2452_ net281 VGND VPWR _0268_ state\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2383_ net442 VGND VPWR _0199_ daisychain\[71\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_37_676 VPWR VGND sg13g2_fill_1
XFILLER_37_698 VPWR VGND sg13g2_fill_1
XFILLER_40_808 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_20_576 VPWR VGND sg13g2_fill_1
XFILLER_32_370 VPWR VGND sg13g2_decap_8
X_2527__404 VPWR VGND net403 sg13g2_tiehi
XFILLER_19_99 VPWR VGND sg13g2_decap_8
XFILLER_27_153 VPWR VGND sg13g2_decap_8
X_2456__266 VPWR VGND net265 sg13g2_tiehi
XFILLER_15_337 VPWR VGND sg13g2_decap_8
XFILLER_31_808 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_43_635 VPWR VGND sg13g2_decap_4
XFILLER_43_668 VPWR VGND sg13g2_decap_8
XFILLER_2_252 VPWR VGND sg13g2_decap_8
XFILLER_18_131 VPWR VGND sg13g2_decap_8
XFILLER_19_665 VPWR VGND sg13g2_decap_4
XFILLER_33_123 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
X_2435__339 VPWR VGND net338 sg13g2_tiehi
XFILLER_21_318 VPWR VGND sg13g2_decap_4
X_1952_ _0635_ net165 _0634_ VPWR VGND sg13g2_nand2_1
X_1883_ VGND VPWR net110 daisychain\[92\] _0580_ net55 sg13g2_a21oi_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_2504_ net329 VGND VPWR _0320_ state\[64\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2435_ net338 VGND VPWR _0251_ daisychain\[123\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
X_1317_ VPWR _0122_ state\[95\] VGND sg13g2_inv_1
X_2366_ net220 VGND VPWR _0182_ daisychain\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2297_ VGND VPWR _0687_ _0838_ _0376_ net70 sg13g2_a21oi_1
XFILLER_12_329 VPWR VGND sg13g2_decap_8
XFILLER_40_605 VPWR VGND sg13g2_decap_8
XFILLER_40_649 VPWR VGND sg13g2_fill_1
XFILLER_21_45 VPWR VGND sg13g2_decap_8
XFILLER_4_506 VPWR VGND sg13g2_decap_4
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_28_473 VPWR VGND sg13g2_decap_4
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_15_156 VPWR VGND sg13g2_decap_8
XFILLER_30_137 VPWR VGND sg13g2_decap_8
XFILLER_31_605 VPWR VGND sg13g2_fill_1
XFILLER_43_476 VPWR VGND sg13g2_decap_4
XFILLER_11_395 VPWR VGND sg13g2_decap_8
XFILLER_7_355 VPWR VGND sg13g2_decap_8
XFILLER_38_259 VPWR VGND sg13g2_decap_8
X_2220_ _0800_ net126 state\[82\] VPWR VGND sg13g2_nand2_1
X_2151_ VGND VPWR _0395_ _0765_ _0303_ net83 sg13g2_a21oi_1
X_2082_ _0731_ net93 state\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_19_484 VPWR VGND sg13g2_decap_4
XFILLER_21_115 VPWR VGND sg13g2_decap_8
XFILLER_34_454 VPWR VGND sg13g2_decap_4
XFILLER_30_693 VPWR VGND sg13g2_fill_1
X_1935_ VGND VPWR _0619_ _0620_ _0231_ _0621_ sg13g2_a21oi_1
X_1866_ state\[90\] daisychain\[90\] net152 _0566_ VPWR VGND sg13g2_mux2_1
X_1797_ _0511_ net175 _0510_ VPWR VGND sg13g2_nand2_1
X_2418_ net372 VGND VPWR _0234_ daisychain\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_29_248 VPWR VGND sg13g2_decap_8
XFILLER_38_771 VPWR VGND sg13g2_fill_2
X_2349_ net254 VGND VPWR _0165_ daisychain\[37\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_12_126 VPWR VGND sg13g2_decap_8
XFILLER_25_454 VPWR VGND sg13g2_fill_1
XFILLER_32_11 VPWR VGND sg13g2_decap_8
XFILLER_40_468 VPWR VGND sg13g2_decap_8
X_2388__433 VPWR VGND net432 sg13g2_tiehi
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_5_815 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_0_575 VPWR VGND sg13g2_fill_1
XFILLER_0_586 VPWR VGND sg13g2_fill_2
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_28_270 VPWR VGND sg13g2_decap_8
XFILLER_28_281 VPWR VGND sg13g2_fill_1
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_11_192 VPWR VGND sg13g2_decap_8
XFILLER_7_152 VPWR VGND sg13g2_decap_8
X_1720_ VGND VPWR _0447_ _0448_ _0188_ _0449_ sg13g2_a21oi_1
X_1651_ state\[47\] daisychain\[47\] net147 _0394_ VPWR VGND sg13g2_mux2_1
X_1582_ _0983_ net170 _0982_ VPWR VGND sg13g2_nand2_1
XFILLER_19_281 VPWR VGND sg13g2_decap_8
XFILLER_26_218 VPWR VGND sg13g2_decap_8
X_2203_ VGND VPWR _0499_ _0791_ _0329_ net86 sg13g2_a21oi_1
X_2134_ _0757_ net116 state\[39\] VPWR VGND sg13g2_nand2_1
X_2065_ VGND VPWR _0867_ _0722_ _0260_ net67 sg13g2_a21oi_1
XFILLER_22_435 VPWR VGND sg13g2_fill_2
XFILLER_35_763 VPWR VGND sg13g2_decap_8
X_2487__398 VPWR VGND net397 sg13g2_tiehi
X_1918_ VGND VPWR net112 daisychain\[99\] _0608_ net54 sg13g2_a21oi_1
X_1849_ net196 VPWR _0553_ VGND daisychain\[86\] net39 sg13g2_o21ai_1
XFILLER_17_218 VPWR VGND sg13g2_decap_8
XFILLER_27_55 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_41_788 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_9_406 VPWR VGND sg13g2_decap_8
XFILLER_4_122 VPWR VGND sg13g2_decap_8
XFILLER_4_199 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_fill_2
XFILLER_5_645 VPWR VGND sg13g2_decap_4
XFILLER_5_689 VPWR VGND sg13g2_fill_1
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_49_822 VPWR VGND sg13g2_fill_1
XFILLER_16_251 VPWR VGND sg13g2_decap_8
XFILLER_31_221 VPWR VGND sg13g2_decap_8
XFILLER_31_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_1703_ VGND VPWR net119 daisychain\[56\] _0436_ net59 sg13g2_a21oi_1
X_1634_ net192 VPWR _1025_ VGND daisychain\[43\] net35 sg13g2_o21ai_1
XFILLER_39_343 VPWR VGND sg13g2_decap_8
X_1496_ state\[16\] daisychain\[16\] net137 _0914_ VPWR VGND sg13g2_mux2_1
X_1565_ VGND VPWR _0967_ _0968_ _0157_ _0969_ sg13g2_a21oi_1
X_2117_ VGND VPWR _0971_ _0748_ _0286_ net74 sg13g2_a21oi_1
X_2048_ VGND VPWR net91 daisychain\[125\] _0712_ net48 sg13g2_a21oi_1
XFILLER_10_416 VPWR VGND sg13g2_decap_8
XFILLER_13_24 VPWR VGND sg13g2_fill_1
XFILLER_13_35 VPWR VGND sg13g2_decap_8
XFILLER_22_221 VPWR VGND sg13g2_decap_8
Xfanout25 net44 net25 VPWR VGND sg13g2_buf_1
Xfanout69 net89 net69 VPWR VGND sg13g2_buf_1
Xfanout58 net65 net58 VPWR VGND sg13g2_buf_1
Xfanout47 net66 net47 VPWR VGND sg13g2_buf_1
Xfanout36 net43 net36 VPWR VGND sg13g2_buf_1
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_8_6 VPWR VGND sg13g2_fill_1
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_13_265 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[1\].u.inv2 VPWR digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_1_692 VPWR VGND sg13g2_fill_2
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_1350_ VPWR _0086_ state\[62\] VGND sg13g2_inv_1
XFILLER_24_508 VPWR VGND sg13g2_fill_2
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_2_1__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_20_714 VPWR VGND sg13g2_fill_2
XFILLER_20_769 VPWR VGND sg13g2_fill_1
X_2414__381 VPWR VGND net380 sg13g2_tiehi
XFILLER_9_792 VPWR VGND sg13g2_fill_2
X_1617_ _1011_ net169 _1010_ VPWR VGND sg13g2_nand2_1
XFILLER_39_140 VPWR VGND sg13g2_decap_8
X_1479_ net180 VPWR _0901_ VGND daisychain\[12\] net23 sg13g2_o21ai_1
X_1548_ VGND VPWR net100 daisychain\[25\] _0956_ net49 sg13g2_a21oi_1
XFILLER_15_519 VPWR VGND sg13g2_decap_4
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_10_213 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_19_803 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_46_633 VPWR VGND sg13g2_decap_4
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_decap_8
XFILLER_26_390 VPWR VGND sg13g2_fill_1
XFILLER_41_371 VPWR VGND sg13g2_decap_8
XFILLER_10_780 VPWR VGND sg13g2_fill_1
XFILLER_5_272 VPWR VGND sg13g2_decap_8
X_1402_ VPWR _0011_ state\[10\] VGND sg13g2_inv_1
X_2520_ net203 VGND VPWR _0336_ state\[80\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2451_ net285 VGND VPWR _0267_ state\[11\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1333_ VPWR _0104_ state\[79\] VGND sg13g2_inv_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_2382_ net444 VGND VPWR _0198_ daisychain\[70\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_24_349 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_decap_8
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_10_47 VPWR VGND sg13g2_fill_1
XFILLER_19_45 VPWR VGND sg13g2_fill_1
XFILLER_19_78 VPWR VGND sg13g2_decap_8
XFILLER_27_132 VPWR VGND sg13g2_decap_8
XFILLER_43_614 VPWR VGND sg13g2_decap_8
XFILLER_11_511 VPWR VGND sg13g2_decap_8
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_2_231 VPWR VGND sg13g2_decap_8
XFILLER_3_732 VPWR VGND sg13g2_fill_2
X_2463__238 VPWR VGND net237 sg13g2_tiehi
X_2398__413 VPWR VGND net412 sg13g2_tiehi
XFILLER_18_110 VPWR VGND sg13g2_decap_8
XFILLER_18_187 VPWR VGND sg13g2_decap_8
XFILLER_33_102 VPWR VGND sg13g2_decap_8
XFILLER_33_179 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
X_1951_ state\[107\] daisychain\[107\] net142 _0634_ VPWR VGND sg13g2_mux2_1
X_1882_ _0579_ net166 _0578_ VPWR VGND sg13g2_nand2_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_2503_ net333 VGND VPWR _0319_ state\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2434_ net340 VGND VPWR _0250_ daisychain\[122\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2365_ net222 VGND VPWR _0181_ daisychain\[53\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_1316_ VPWR _0123_ state\[96\] VGND sg13g2_inv_1
X_2296_ _0838_ net98 state\[120\] VPWR VGND sg13g2_nand2_1
XFILLER_12_308 VPWR VGND sg13g2_decap_8
XFILLER_24_113 VPWR VGND sg13g2_fill_2
XFILLER_33_680 VPWR VGND sg13g2_fill_2
XFILLER_33_691 VPWR VGND sg13g2_fill_2
XFILLER_0_713 VPWR VGND sg13g2_fill_2
XFILLER_15_135 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_11_374 VPWR VGND sg13g2_decap_8
XFILLER_30_116 VPWR VGND sg13g2_decap_8
XFILLER_31_639 VPWR VGND sg13g2_decap_8
XFILLER_43_499 VPWR VGND sg13g2_fill_2
XFILLER_7_15 VPWR VGND sg13g2_fill_1
XFILLER_7_26 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_decap_8
XFILLER_7_48 VPWR VGND sg13g2_fill_2
XFILLER_3_595 VPWR VGND sg13g2_decap_8
XFILLER_19_441 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
X_2150_ _0765_ net123 state\[47\] VPWR VGND sg13g2_nand2_1
X_2081_ VGND VPWR _0899_ _0730_ _0268_ net67 sg13g2_a21oi_1
XFILLER_19_496 VPWR VGND sg13g2_fill_2
X_1934_ net189 VPWR _0621_ VGND daisychain\[103\] net32 sg13g2_o21ai_1
XFILLER_30_672 VPWR VGND sg13g2_fill_1
X_2563__424 VPWR VGND net423 sg13g2_tiehi
X_1865_ VGND VPWR _0563_ _0564_ _0217_ _0565_ sg13g2_a21oi_1
X_1796_ state\[76\] daisychain\[76\] net153 _0510_ VPWR VGND sg13g2_mux2_1
XFILLER_29_227 VPWR VGND sg13g2_decap_8
X_2417_ net374 VGND VPWR _0233_ daisychain\[105\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2348_ net256 VGND VPWR _0164_ daisychain\[36\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_16_35 VPWR VGND sg13g2_fill_2
XFILLER_38_794 VPWR VGND sg13g2_fill_2
X_2279_ VGND VPWR _0651_ _0829_ _0367_ net79 sg13g2_a21oi_1
XFILLER_12_105 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_4_304 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_36_709 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_16_422 VPWR VGND sg13g2_fill_2
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_44_775 VPWR VGND sg13g2_decap_4
XFILLER_11_171 VPWR VGND sg13g2_decap_8
XFILLER_12_661 VPWR VGND sg13g2_fill_1
XFILLER_12_672 VPWR VGND sg13g2_fill_1
XFILLER_7_131 VPWR VGND sg13g2_decap_8
XFILLER_8_687 VPWR VGND sg13g2_fill_1
X_1650_ VGND VPWR _0391_ _0392_ _0174_ _0393_ sg13g2_a21oi_1
X_1581_ state\[33\] daisychain\[33\] net147 _0982_ VPWR VGND sg13g2_mux2_1
X_2202_ _0791_ net130 state\[73\] VPWR VGND sg13g2_nand2_1
XFILLER_14_2 VPWR VGND sg13g2_fill_1
XFILLER_19_260 VPWR VGND sg13g2_decap_8
XFILLER_35_753 VPWR VGND sg13g2_decap_4
XFILLER_39_536 VPWR VGND sg13g2_decap_8
XFILLER_39_547 VPWR VGND sg13g2_fill_2
X_2133_ VGND VPWR _1003_ _0756_ _0294_ net73 sg13g2_a21oi_1
X_2064_ _0722_ net93 state\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_22_403 VPWR VGND sg13g2_fill_1
XFILLER_22_469 VPWR VGND sg13g2_fill_1
XFILLER_34_285 VPWR VGND sg13g2_decap_8
X_1917_ _0607_ net167 _0606_ VPWR VGND sg13g2_nand2_1
XFILLER_1_329 VPWR VGND sg13g2_decap_8
X_2528__396 VPWR VGND net395 sg13g2_tiehi
X_2424__361 VPWR VGND net360 sg13g2_tiehi
X_1848_ VGND VPWR net124 daisychain\[85\] _0552_ net61 sg13g2_a21oi_1
X_1779_ net198 VPWR _0497_ VGND daisychain\[72\] net41 sg13g2_o21ai_1
XFILLER_13_414 VPWR VGND sg13g2_fill_1
XFILLER_25_263 VPWR VGND sg13g2_decap_4
XFILLER_25_285 VPWR VGND sg13g2_decap_8
XFILLER_38_580 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_4_101 VPWR VGND sg13g2_decap_8
XFILLER_4_178 VPWR VGND sg13g2_decap_8
XFILLER_16_230 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_31_200 VPWR VGND sg13g2_decap_8
XFILLER_31_277 VPWR VGND sg13g2_decap_8
X_1702_ _0435_ net171 _0434_ VPWR VGND sg13g2_nand2_1
X_1633_ VGND VPWR net115 daisychain\[42\] _1024_ net57 sg13g2_a21oi_1
X_1564_ net185 VPWR _0969_ VGND daisychain\[29\] net28 sg13g2_o21ai_1
XFILLER_39_322 VPWR VGND sg13g2_decap_8
X_1495_ VGND VPWR _0911_ _0912_ _0143_ _0913_ sg13g2_a21oi_1
XFILLER_22_200 VPWR VGND sg13g2_decap_8
XFILLER_39_399 VPWR VGND sg13g2_decap_8
Xfanout26 net29 net26 VPWR VGND sg13g2_buf_1
Xfanout37 net38 net37 VPWR VGND sg13g2_buf_1
X_2116_ _0748_ net105 state\[30\] VPWR VGND sg13g2_nand2_1
X_2047_ _0711_ net157 _0710_ VPWR VGND sg13g2_nand2_1
XFILLER_13_69 VPWR VGND sg13g2_decap_8
Xfanout59 net60 net59 VPWR VGND sg13g2_buf_1
Xfanout48 net66 net48 VPWR VGND sg13g2_buf_1
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_46_815 VPWR VGND sg13g2_decap_8
X_2459__254 VPWR VGND net253 sg13g2_tiehi
XFILLER_13_244 VPWR VGND sg13g2_decap_8
XFILLER_14_745 VPWR VGND sg13g2_decap_4
XFILLER_14_789 VPWR VGND sg13g2_fill_1
XFILLER_41_553 VPWR VGND sg13g2_decap_4
XFILLER_9_259 VPWR VGND sg13g2_decap_8
XFILLER_5_454 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_17_594 VPWR VGND sg13g2_fill_1
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_20_748 VPWR VGND sg13g2_fill_1
X_2564__360 VPWR VGND net359 sg13g2_tiehi
XFILLER_8_292 VPWR VGND sg13g2_decap_8
X_1547_ _0955_ net161 _0954_ VPWR VGND sg13g2_nand2_1
X_1616_ state\[40\] daisychain\[40\] net146 _1010_ VPWR VGND sg13g2_mux2_1
XFILLER_27_358 VPWR VGND sg13g2_decap_8
XFILLER_39_196 VPWR VGND sg13g2_decap_8
X_1478_ VGND VPWR net92 daisychain\[11\] _0900_ net45 sg13g2_a21oi_1
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_269 VPWR VGND sg13g2_decap_8
XFILLER_2_413 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_46_601 VPWR VGND sg13g2_fill_2
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_33_328 VPWR VGND sg13g2_fill_1
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
X_2544__208 VPWR VGND net207 sg13g2_tiehi
XFILLER_5_251 VPWR VGND sg13g2_decap_8
X_1401_ VPWR _0022_ state\[11\] VGND sg13g2_inv_1
X_2450_ net289 VGND VPWR _0266_ state\[10\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2381_ net446 VGND VPWR _0197_ daisychain\[69\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_37_634 VPWR VGND sg13g2_decap_8
XFILLER_49_494 VPWR VGND sg13g2_decap_8
X_1332_ VPWR _0106_ state\[80\] VGND sg13g2_inv_1
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_32_350 VPWR VGND sg13g2_fill_2
XFILLER_37_689 VPWR VGND sg13g2_decap_8
XFILLER_20_589 VPWR VGND sg13g2_fill_1
XFILLER_10_59 VPWR VGND sg13g2_decap_8
XFILLER_16_818 VPWR VGND sg13g2_decap_4
XFILLER_19_57 VPWR VGND sg13g2_decap_8
XFILLER_27_111 VPWR VGND sg13g2_decap_8
XFILLER_27_188 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_11_534 VPWR VGND sg13g2_fill_2
XFILLER_11_556 VPWR VGND sg13g2_fill_1
XFILLER_11_589 VPWR VGND sg13g2_fill_2
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_2_210 VPWR VGND sg13g2_decap_8
XFILLER_2_287 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_14_383 VPWR VGND sg13g2_decap_8
XFILLER_18_166 VPWR VGND sg13g2_decap_8
XFILLER_30_810 VPWR VGND sg13g2_fill_1
XFILLER_33_158 VPWR VGND sg13g2_decap_8
XFILLER_34_604 VPWR VGND sg13g2_fill_2
XFILLER_46_497 VPWR VGND sg13g2_decap_8
X_1950_ VGND VPWR _0631_ _0632_ _0234_ _0633_ sg13g2_a21oi_1
X_2502_ net337 VGND VPWR _0318_ state\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1881_ state\[93\] daisychain\[93\] net143 _0578_ VPWR VGND sg13g2_mux2_1
X_1315_ VPWR _0124_ state\[97\] VGND sg13g2_inv_1
X_2433_ net342 VGND VPWR _0249_ daisychain\[121\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2364_ net224 VGND VPWR _0180_ daisychain\[52\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_37_453 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
X_2295_ VGND VPWR _0683_ _0837_ _0375_ net69 sg13g2_a21oi_1
XFILLER_24_169 VPWR VGND sg13g2_decap_8
XFILLER_40_629 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_15_114 VPWR VGND sg13g2_decap_8
XFILLER_16_659 VPWR VGND sg13g2_fill_2
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
X_2434__341 VPWR VGND net340 sg13g2_tiehi
XFILLER_11_353 VPWR VGND sg13g2_decap_8
XFILLER_7_313 VPWR VGND sg13g2_decap_8
XFILLER_8_803 VPWR VGND sg13g2_fill_1
X_2510__284 VPWR VGND net283 sg13g2_tiehi
XFILLER_11_80 VPWR VGND sg13g2_decap_8
XFILLER_30_8 VPWR VGND sg13g2_fill_2
XFILLER_3_530 VPWR VGND sg13g2_fill_1
XFILLER_3_552 VPWR VGND sg13g2_fill_2
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
X_2080_ _0730_ net92 state\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_14_191 VPWR VGND sg13g2_decap_8
XFILLER_30_651 VPWR VGND sg13g2_fill_1
X_2335__283 VPWR VGND net282 sg13g2_tiehi
X_1933_ VGND VPWR net110 daisychain\[102\] _0620_ net55 sg13g2_a21oi_1
X_1864_ net196 VPWR _0565_ VGND daisychain\[89\] net39 sg13g2_o21ai_1
X_1795_ VGND VPWR _0507_ _0508_ _0203_ _0509_ sg13g2_a21oi_1
XFILLER_29_206 VPWR VGND sg13g2_decap_8
X_2416_ net376 VGND VPWR _0232_ daisychain\[104\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2347_ net258 VGND VPWR _0163_ daisychain\[35\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2278_ _0829_ net114 state\[111\] VPWR VGND sg13g2_nand2_1
XFILLER_16_69 VPWR VGND sg13g2_decap_8
XFILLER_25_478 VPWR VGND sg13g2_fill_2
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_38_762 VPWR VGND sg13g2_fill_1
XFILLER_20_194 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_fill_1
XFILLER_16_412 VPWR VGND sg13g2_decap_4
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_11_150 VPWR VGND sg13g2_decap_8
XFILLER_12_640 VPWR VGND sg13g2_fill_1
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_7_110 VPWR VGND sg13g2_decap_8
XFILLER_7_187 VPWR VGND sg13g2_decap_8
XFILLER_8_633 VPWR VGND sg13g2_decap_8
XFILLER_8_677 VPWR VGND sg13g2_decap_4
XFILLER_8_699 VPWR VGND sg13g2_decap_8
X_1580_ VGND VPWR _0979_ _0980_ _0160_ _0981_ sg13g2_a21oi_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_fill_2
XFILLER_39_515 VPWR VGND sg13g2_fill_1
XFILLER_3_393 VPWR VGND sg13g2_decap_8
X_2201_ VGND VPWR _0495_ _0790_ _0328_ net86 sg13g2_a21oi_1
X_2132_ _0756_ net103 state\[38\] VPWR VGND sg13g2_nand2_1
XFILLER_34_264 VPWR VGND sg13g2_decap_8
XFILLER_35_710 VPWR VGND sg13g2_decap_4
X_2452__282 VPWR VGND net281 sg13g2_tiehi
X_2063_ VGND VPWR _0863_ _0721_ _0259_ net67 sg13g2_a21oi_1
X_1916_ state\[100\] daisychain\[100\] net144 _0606_ VPWR VGND sg13g2_mux2_1
X_1847_ _0551_ net174 _0550_ VPWR VGND sg13g2_nand2_1
XFILLER_1_308 VPWR VGND sg13g2_decap_8
X_1778_ VGND VPWR net128 daisychain\[71\] _0496_ net63 sg13g2_a21oi_1
XFILLER_38_570 VPWR VGND sg13g2_fill_1
XFILLER_25_242 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_decap_4
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_4_157 VPWR VGND sg13g2_decap_8
XFILLER_5_636 VPWR VGND sg13g2_fill_1
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_fill_2
XFILLER_17_743 VPWR VGND sg13g2_fill_2
XFILLER_17_787 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_fill_2
XFILLER_44_584 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_16_286 VPWR VGND sg13g2_decap_8
XFILLER_31_256 VPWR VGND sg13g2_decap_8
X_1701_ state\[57\] daisychain\[57\] net148 _0434_ VPWR VGND sg13g2_mux2_1
XFILLER_3_190 VPWR VGND sg13g2_decap_8
X_1494_ net183 VPWR _0913_ VGND daisychain\[15\] net26 sg13g2_o21ai_1
X_1632_ _1023_ net169 _1022_ VPWR VGND sg13g2_nand2_1
X_1563_ VGND VPWR net100 daisychain\[28\] _0968_ net52 sg13g2_a21oi_1
XFILLER_27_507 VPWR VGND sg13g2_fill_2
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_39_378 VPWR VGND sg13g2_decap_8
X_2115_ VGND VPWR _0967_ _0747_ _0285_ net74 sg13g2_a21oi_1
Xfanout27 net29 net27 VPWR VGND sg13g2_buf_1
Xfanout49 net52 net49 VPWR VGND sg13g2_buf_1
Xfanout38 net43 net38 VPWR VGND sg13g2_buf_1
X_2046_ state\[126\] daisychain\[126\] net135 _0710_ VPWR VGND sg13g2_mux2_1
XFILLER_13_48 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_2_639 VPWR VGND sg13g2_fill_2
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_13_223 VPWR VGND sg13g2_decap_8
XFILLER_41_598 VPWR VGND sg13g2_fill_2
XFILLER_9_238 VPWR VGND sg13g2_decap_8
X_2466__226 VPWR VGND net225 sg13g2_tiehi
XFILLER_5_433 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_1_694 VPWR VGND sg13g2_fill_1
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_32_510 VPWR VGND sg13g2_decap_8
XFILLER_32_565 VPWR VGND sg13g2_decap_4
XFILLER_44_392 VPWR VGND sg13g2_decap_8
XFILLER_20_727 VPWR VGND sg13g2_fill_1
XFILLER_8_271 VPWR VGND sg13g2_decap_8
XFILLER_9_794 VPWR VGND sg13g2_fill_1
X_1477_ _0899_ net158 _0898_ VPWR VGND sg13g2_nand2_1
X_1546_ state\[26\] daisychain\[26\] net138 _0954_ VPWR VGND sg13g2_mux2_1
X_1615_ VGND VPWR _1007_ _1008_ _0167_ _1009_ sg13g2_a21oi_1
XFILLER_27_326 VPWR VGND sg13g2_decap_4
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_43_808 VPWR VGND sg13g2_decap_8
XFILLER_10_248 VPWR VGND sg13g2_decap_8
XFILLER_11_749 VPWR VGND sg13g2_decap_8
XFILLER_23_510 VPWR VGND sg13g2_fill_2
XFILLER_23_521 VPWR VGND sg13g2_fill_1
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_42_329 VPWR VGND sg13g2_decap_8
X_2029_ net179 VPWR _0697_ VGND daisychain\[122\] net25 sg13g2_o21ai_1
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_6_219 VPWR VGND sg13g2_decap_8
XFILLER_2_469 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
X_2513__260 VPWR VGND net259 sg13g2_tiehi
XFILLER_10_771 VPWR VGND sg13g2_decap_8
XFILLER_14_587 VPWR VGND sg13g2_fill_2
XFILLER_5_230 VPWR VGND sg13g2_decap_8
X_1331_ VPWR _0107_ state\[81\] VGND sg13g2_inv_1
X_1400_ VPWR _0031_ state\[12\] VGND sg13g2_inv_1
Xwires dac/Iout dac/VcascP[1] dac/VcascP[0] dac/VbiasP[1] dac/VbiasP[0] wires/VDDA[1]
+ wires/VDDA[0] i_in i_out analog_wires
X_2380_ net448 VGND VPWR _0196_ daisychain\[68\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_20_535 VPWR VGND sg13g2_fill_1
XFILLER_32_362 VPWR VGND sg13g2_fill_2
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_10_38 VPWR VGND sg13g2_decap_8
X_2345__263 VPWR VGND net262 sg13g2_tiehi
XFILLER_19_36 VPWR VGND sg13g2_fill_2
X_1529_ net185 VPWR _0941_ VGND daisychain\[22\] net28 sg13g2_o21ai_1
XFILLER_27_167 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_11_568 VPWR VGND sg13g2_decap_8
XFILLER_11_579 VPWR VGND sg13g2_fill_2
XFILLER_2_266 VPWR VGND sg13g2_decap_8
XFILLER_3_756 VPWR VGND sg13g2_decap_4
XFILLER_18_145 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_25_90 VPWR VGND sg13g2_fill_1
XFILLER_33_137 VPWR VGND sg13g2_decap_8
XFILLER_34_638 VPWR VGND sg13g2_fill_2
X_1880_ VGND VPWR _0575_ _0576_ _0220_ _0577_ sg13g2_a21oi_1
XFILLER_6_594 VPWR VGND sg13g2_decap_8
X_2501_ net341 VGND VPWR _0317_ state\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1314_ VPWR _0125_ state\[98\] VGND sg13g2_inv_1
X_2432_ net344 VGND VPWR _0248_ daisychain\[120\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2363_ net226 VGND VPWR _0179_ daisychain\[51\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2294_ _0837_ net97 state\[119\] VPWR VGND sg13g2_nand2_1
XFILLER_24_115 VPWR VGND sg13g2_fill_1
XFILLER_24_148 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_20_365 VPWR VGND sg13g2_decap_8
XFILLER_20_398 VPWR VGND sg13g2_decap_8
XFILLER_33_682 VPWR VGND sg13g2_fill_1
XFILLER_21_59 VPWR VGND sg13g2_decap_8
XFILLER_16_616 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
X_2497__358 VPWR VGND net357 sg13g2_tiehi
XFILLER_11_332 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_3_520 VPWR VGND sg13g2_fill_1
XFILLER_7_369 VPWR VGND sg13g2_decap_8
XFILLER_8_815 VPWR VGND sg13g2_decap_8
XFILLER_23_8 VPWR VGND sg13g2_fill_1
XFILLER_19_454 VPWR VGND sg13g2_decap_8
XFILLER_19_465 VPWR VGND sg13g2_fill_2
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_14_170 VPWR VGND sg13g2_decap_8
XFILLER_21_129 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_fill_2
XFILLER_30_685 VPWR VGND sg13g2_fill_1
X_1932_ _0619_ net166 _0618_ VPWR VGND sg13g2_nand2_1
X_1863_ VGND VPWR net111 daisychain\[88\] _0564_ net54 sg13g2_a21oi_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_6_380 VPWR VGND sg13g2_decap_8
X_2415_ net378 VGND VPWR _0231_ daisychain\[103\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1794_ net196 VPWR _0509_ VGND daisychain\[75\] net39 sg13g2_o21ai_1
X_2346_ net260 VGND VPWR _0162_ daisychain\[34\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2277_ VGND VPWR _0647_ _0828_ _0366_ net79 sg13g2_a21oi_1
XFILLER_13_619 VPWR VGND sg13g2_decap_8
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_20_173 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_fill_2
XFILLER_16_424 VPWR VGND sg13g2_fill_1
XFILLER_43_210 VPWR VGND sg13g2_decap_8
X_2551__352 VPWR VGND net351 sg13g2_tiehi
XFILLER_12_652 VPWR VGND sg13g2_fill_2
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_3_372 VPWR VGND sg13g2_decap_8
XFILLER_7_166 VPWR VGND sg13g2_decap_8
X_2200_ _0790_ net128 state\[72\] VPWR VGND sg13g2_nand2_1
X_2131_ VGND VPWR _0999_ _0755_ _0293_ net73 sg13g2_a21oi_1
X_2062_ _0721_ net92 state\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_19_295 VPWR VGND sg13g2_decap_8
XFILLER_34_243 VPWR VGND sg13g2_decap_8
XFILLER_30_493 VPWR VGND sg13g2_fill_1
XFILLER_8_82 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_2_0__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_1915_ VGND VPWR _0603_ _0604_ _0227_ _0605_ sg13g2_a21oi_1
X_1846_ state\[86\] daisychain\[86\] net152 _0550_ VPWR VGND sg13g2_mux2_1
X_1777_ _0495_ net175 _0494_ VPWR VGND sg13g2_nand2_1
XFILLER_25_221 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_27_69 VPWR VGND sg13g2_decap_8
X_2329_ net294 VGND VPWR _0145_ daisychain\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_41_769 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_4_136 VPWR VGND sg13g2_decap_8
X_2546__432 VPWR VGND net431 sg13g2_tiehi
X_2403__403 VPWR VGND net402 sg13g2_tiehi
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_1_821 VPWR VGND sg13g2_fill_2
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_16_265 VPWR VGND sg13g2_decap_8
XFILLER_17_777 VPWR VGND sg13g2_decap_4
XFILLER_31_235 VPWR VGND sg13g2_decap_8
XFILLER_8_453 VPWR VGND sg13g2_decap_8
XFILLER_8_464 VPWR VGND sg13g2_fill_2
X_1700_ VGND VPWR _0431_ _0432_ _0184_ _0433_ sg13g2_a21oi_1
X_1631_ state\[43\] daisychain\[43\] net146 _1022_ VPWR VGND sg13g2_mux2_1
X_1493_ VGND VPWR net94 daisychain\[14\] _0912_ net47 sg13g2_a21oi_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_1562_ _0967_ net163 _0966_ VPWR VGND sg13g2_nand2_1
XFILLER_39_357 VPWR VGND sg13g2_decap_8
X_2114_ _0747_ net105 state\[29\] VPWR VGND sg13g2_nand2_1
X_2045_ VGND VPWR _0707_ _0708_ _0253_ _0709_ sg13g2_a21oi_1
XFILLER_35_585 VPWR VGND sg13g2_fill_2
Xfanout28 net29 net28 VPWR VGND sg13g2_buf_1
Xfanout39 net40 net39 VPWR VGND sg13g2_buf_1
X_2385__439 VPWR VGND net438 sg13g2_tiehi
X_1829_ net197 VPWR _0537_ VGND daisychain\[82\] net40 sg13g2_o21ai_1
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_13_202 VPWR VGND sg13g2_decap_8
XFILLER_41_522 VPWR VGND sg13g2_decap_4
X_2355__243 VPWR VGND net242 sg13g2_tiehi
XFILLER_13_279 VPWR VGND sg13g2_decap_8
XFILLER_41_577 VPWR VGND sg13g2_decap_8
XFILLER_5_412 VPWR VGND sg13g2_decap_8
XFILLER_9_217 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_49_666 VPWR VGND sg13g2_decap_8
XFILLER_49_688 VPWR VGND sg13g2_decap_4
XFILLER_17_585 VPWR VGND sg13g2_decap_8
XFILLER_20_706 VPWR VGND sg13g2_fill_1
XFILLER_20_739 VPWR VGND sg13g2_fill_2
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_8_250 VPWR VGND sg13g2_decap_8
X_1614_ net192 VPWR _1009_ VGND daisychain\[39\] net35 sg13g2_o21ai_1
XFILLER_5_83 VPWR VGND sg13g2_decap_8
X_1476_ state\[12\] daisychain\[12\] net134 _0898_ VPWR VGND sg13g2_mux2_1
X_1545_ VGND VPWR _0951_ _0952_ _0153_ _0953_ sg13g2_a21oi_1
XFILLER_27_338 VPWR VGND sg13g2_fill_2
XFILLER_35_371 VPWR VGND sg13g2_fill_2
XFILLER_39_154 VPWR VGND sg13g2_decap_8
XFILLER_42_308 VPWR VGND sg13g2_decap_8
X_2028_ VGND VPWR net90 daisychain\[121\] _0696_ net48 sg13g2_a21oi_1
XFILLER_10_227 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_2_448 VPWR VGND sg13g2_decap_8
XFILLER_19_817 VPWR VGND sg13g2_fill_2
XFILLER_46_658 VPWR VGND sg13g2_decap_4
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_14_511 VPWR VGND sg13g2_decap_8
XFILLER_14_555 VPWR VGND sg13g2_decap_8
XFILLER_14_577 VPWR VGND sg13g2_fill_1
XFILLER_26_360 VPWR VGND sg13g2_fill_1
XFILLER_33_319 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_42_820 VPWR VGND sg13g2_fill_2
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_6_732 VPWR VGND sg13g2_fill_2
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_5_286 VPWR VGND sg13g2_decap_8
X_1330_ VPWR _0108_ state\[82\] VGND sg13g2_inv_1
XFILLER_33_820 VPWR VGND sg13g2_fill_2
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_37_647 VPWR VGND sg13g2_decap_4
XFILLER_49_452 VPWR VGND sg13g2_decap_8
X_2490__386 VPWR VGND net385 sg13g2_tiehi
XFILLER_32_330 VPWR VGND sg13g2_decap_4
X_2531__372 VPWR VGND net371 sg13g2_tiehi
X_1459_ net183 VPWR _0885_ VGND daisychain\[8\] net26 sg13g2_o21ai_1
X_1528_ VGND VPWR net104 daisychain\[21\] _0940_ net50 sg13g2_a21oi_1
XFILLER_23_363 VPWR VGND sg13g2_fill_2
XFILLER_27_146 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_43_628 VPWR VGND sg13g2_decap_8
XFILLER_43_639 VPWR VGND sg13g2_fill_2
XFILLER_11_536 VPWR VGND sg13g2_fill_1
XFILLER_11_547 VPWR VGND sg13g2_decap_4
XFILLER_3_713 VPWR VGND sg13g2_fill_1
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_18_124 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_decap_8
XFILLER_33_116 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_26_190 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
X_2411__387 VPWR VGND net386 sg13g2_tiehi
X_2500_ net345 VGND VPWR _0316_ state\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2431_ net346 VGND VPWR _0247_ daisychain\[119\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_2_790 VPWR VGND sg13g2_fill_2
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_1313_ VPWR _0126_ state\[99\] VGND sg13g2_inv_1
X_2362_ net228 VGND VPWR _0178_ daisychain\[50\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2293_ VGND VPWR _0679_ _0836_ _0374_ net69 sg13g2_a21oi_1
XFILLER_17_190 VPWR VGND sg13g2_decap_8
XFILLER_18_691 VPWR VGND sg13g2_fill_2
XFILLER_33_672 VPWR VGND sg13g2_fill_2
XFILLER_37_466 VPWR VGND sg13g2_decap_4
X_2455__270 VPWR VGND net269 sg13g2_tiehi
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_28_488 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_11_311 VPWR VGND sg13g2_decap_8
XFILLER_15_149 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_11_388 VPWR VGND sg13g2_decap_8
XFILLER_3_554 VPWR VGND sg13g2_fill_1
XFILLER_7_348 VPWR VGND sg13g2_decap_8
XFILLER_47_731 VPWR VGND sg13g2_fill_1
XFILLER_19_477 VPWR VGND sg13g2_decap_8
XFILLER_21_108 VPWR VGND sg13g2_decap_8
XFILLER_34_458 VPWR VGND sg13g2_fill_1
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_30_664 VPWR VGND sg13g2_fill_1
XFILLER_30_697 VPWR VGND sg13g2_fill_1
X_1931_ state\[103\] daisychain\[103\] net143 _0618_ VPWR VGND sg13g2_mux2_1
X_1862_ _0563_ net173 _0562_ VPWR VGND sg13g2_nand2_1
X_1793_ VGND VPWR net125 daisychain\[74\] _0508_ net61 sg13g2_a21oi_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
X_2414_ net380 VGND VPWR _0230_ daisychain\[102\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_37_252 VPWR VGND sg13g2_decap_8
X_2345_ net262 VGND VPWR _0161_ daisychain\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2276_ _0828_ net109 state\[110\] VPWR VGND sg13g2_nand2_1
XFILLER_12_119 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_4
X_2314__325 VPWR VGND net324 sg13g2_tiehi
XFILLER_20_152 VPWR VGND sg13g2_decap_8
XFILLER_4_318 VPWR VGND sg13g2_decap_8
XFILLER_5_808 VPWR VGND sg13g2_decap_8
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
X_2395__419 VPWR VGND net418 sg13g2_tiehi
XFILLER_28_263 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_11_185 VPWR VGND sg13g2_decap_8
XFILLER_12_631 VPWR VGND sg13g2_decap_8
XFILLER_31_428 VPWR VGND sg13g2_decap_4
XFILLER_7_145 VPWR VGND sg13g2_decap_8
XFILLER_8_613 VPWR VGND sg13g2_fill_1
X_2469__214 VPWR VGND net213 sg13g2_tiehi
X_2365__223 VPWR VGND net222 sg13g2_tiehi
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_3_351 VPWR VGND sg13g2_decap_8
XFILLER_19_274 VPWR VGND sg13g2_decap_8
X_2130_ _0755_ net103 state\[37\] VPWR VGND sg13g2_nand2_1
X_2061_ VGND VPWR _0859_ _0720_ _0258_ net67 sg13g2_a21oi_1
XFILLER_34_222 VPWR VGND sg13g2_decap_8
XFILLER_34_299 VPWR VGND sg13g2_decap_8
XFILLER_35_778 VPWR VGND sg13g2_fill_1
X_1914_ net190 VPWR _0605_ VGND daisychain\[99\] net33 sg13g2_o21ai_1
XFILLER_30_450 VPWR VGND sg13g2_fill_1
XFILLER_8_61 VPWR VGND sg13g2_decap_8
X_1845_ VGND VPWR _0547_ _0548_ _0213_ _0549_ sg13g2_a21oi_1
X_1776_ state\[72\] daisychain\[72\] net153 _0494_ VPWR VGND sg13g2_mux2_1
X_2328_ net296 VGND VPWR _0144_ daisychain\[16\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_25_200 VPWR VGND sg13g2_decap_8
XFILLER_25_233 VPWR VGND sg13g2_fill_1
XFILLER_27_48 VPWR VGND sg13g2_decap_8
XFILLER_38_594 VPWR VGND sg13g2_decap_8
XFILLER_41_715 VPWR VGND sg13g2_decap_4
XFILLER_43_14 VPWR VGND sg13g2_decap_8
X_2259_ VGND VPWR _0611_ _0819_ _0357_ net78 sg13g2_a21oi_1
XFILLER_25_299 VPWR VGND sg13g2_fill_2
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_fill_2
XFILLER_4_115 VPWR VGND sg13g2_decap_8
XFILLER_5_649 VPWR VGND sg13g2_fill_2
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_17_701 VPWR VGND sg13g2_fill_1
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_16_244 VPWR VGND sg13g2_decap_8
XFILLER_17_92 VPWR VGND sg13g2_decap_8
XFILLER_31_214 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_decap_8
XFILLER_44_553 VPWR VGND sg13g2_fill_1
XFILLER_8_432 VPWR VGND sg13g2_decap_8
X_1630_ VGND VPWR _1019_ _1020_ _0170_ _1021_ sg13g2_a21oi_1
X_1492_ _0911_ net161 _0910_ VPWR VGND sg13g2_nand2_1
X_1561_ state\[29\] daisychain\[29\] net140 _0966_ VPWR VGND sg13g2_mux2_1
XFILLER_39_336 VPWR VGND sg13g2_decap_8
X_2113_ VGND VPWR _0963_ _0746_ _0284_ net72 sg13g2_a21oi_1
X_2044_ net179 VPWR _0709_ VGND daisychain\[125\] net25 sg13g2_o21ai_1
XFILLER_10_409 VPWR VGND sg13g2_decap_8
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_30_291 VPWR VGND sg13g2_fill_2
Xfanout29 net44 net29 VPWR VGND sg13g2_buf_1
X_1828_ VGND VPWR net126 daisychain\[81\] _0536_ net61 sg13g2_a21oi_1
X_1759_ net198 VPWR _0481_ VGND daisychain\[68\] net41 sg13g2_o21ai_1
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_13_258 VPWR VGND sg13g2_decap_8
XFILLER_14_726 VPWR VGND sg13g2_fill_1
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_1_663 VPWR VGND sg13g2_fill_2
XFILLER_49_634 VPWR VGND sg13g2_fill_1
XFILLER_5_468 VPWR VGND sg13g2_fill_2
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_12_280 VPWR VGND sg13g2_decap_8
XFILLER_32_589 VPWR VGND sg13g2_fill_2
XFILLER_5_62 VPWR VGND sg13g2_decap_8
X_1544_ net184 VPWR _0953_ VGND daisychain\[25\] net27 sg13g2_o21ai_1
X_1613_ VGND VPWR net103 daisychain\[38\] _1008_ net50 sg13g2_a21oi_1
XFILLER_39_133 VPWR VGND sg13g2_decap_8
X_1475_ VGND VPWR _0895_ _0896_ _0139_ _0897_ sg13g2_a21oi_1
X_2421__367 VPWR VGND net366 sg13g2_tiehi
XFILLER_23_534 VPWR VGND sg13g2_decap_4
XFILLER_35_350 VPWR VGND sg13g2_decap_8
X_2027_ _0695_ net157 _0694_ VPWR VGND sg13g2_nand2_1
XFILLER_10_206 VPWR VGND sg13g2_decap_8
XFILLER_2_427 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_18_306 VPWR VGND sg13g2_fill_2
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_46_626 VPWR VGND sg13g2_decap_8
XFILLER_46_637 VPWR VGND sg13g2_fill_2
XFILLER_14_589 VPWR VGND sg13g2_fill_1
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_14_93 VPWR VGND sg13g2_decap_8
XFILLER_30_81 VPWR VGND sg13g2_decap_8
XFILLER_5_265 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_4
XFILLER_6_755 VPWR VGND sg13g2_decap_4
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_17_372 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_32_364 VPWR VGND sg13g2_fill_1
XFILLER_9_560 VPWR VGND sg13g2_decap_8
X_1527_ _0939_ net163 _0938_ VPWR VGND sg13g2_nand2_1
XFILLER_27_125 VPWR VGND sg13g2_decap_8
X_1389_ VPWR _0043_ state\[23\] VGND sg13g2_inv_1
X_1458_ VGND VPWR net101 daisychain\[7\] _0884_ net49 sg13g2_a21oi_1
XFILLER_11_504 VPWR VGND sg13g2_decap_8
XFILLER_3_725 VPWR VGND sg13g2_decap_8
X_2324__305 VPWR VGND net304 sg13g2_tiehi
XFILLER_19_615 VPWR VGND sg13g2_decap_4
XFILLER_2_224 VPWR VGND sg13g2_decap_8
XFILLER_14_331 VPWR VGND sg13g2_decap_8
XFILLER_15_821 VPWR VGND sg13g2_fill_2
XFILLER_18_103 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_14_397 VPWR VGND sg13g2_fill_1
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_552 VPWR VGND sg13g2_fill_1
XFILLER_6_574 VPWR VGND sg13g2_decap_4
X_2430_ net348 VGND VPWR _0246_ daisychain\[118\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2361_ net230 VGND VPWR _0177_ daisychain\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XFILLER_2_780 VPWR VGND sg13g2_decap_4
X_1312_ VPWR _0001_ state\[100\] VGND sg13g2_inv_1
X_2375__203 VPWR VGND net202 sg13g2_tiehi
X_2292_ _0836_ net95 state\[118\] VPWR VGND sg13g2_nand2_1
XFILLER_32_172 VPWR VGND sg13g2_decap_8
X_2462__242 VPWR VGND net241 sg13g2_tiehi
X_2559_ net375 VGND VPWR _0375_ state\[119\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_15_128 VPWR VGND sg13g2_decap_8
XFILLER_28_412 VPWR VGND sg13g2_decap_4
XFILLER_28_456 VPWR VGND sg13g2_decap_4
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_11_367 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_30_109 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_8
XFILLER_11_94 VPWR VGND sg13g2_decap_8
XFILLER_3_588 VPWR VGND sg13g2_decap_8
X_2441__326 VPWR VGND net325 sg13g2_tiehi
XFILLER_19_423 VPWR VGND sg13g2_decap_4
XFILLER_19_434 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_fill_1
XFILLER_15_662 VPWR VGND sg13g2_fill_2
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_42_470 VPWR VGND sg13g2_fill_1
X_1930_ VGND VPWR _0615_ _0616_ _0230_ _0617_ sg13g2_a21oi_1
XFILLER_30_643 VPWR VGND sg13g2_fill_1
XFILLER_30_676 VPWR VGND sg13g2_fill_2
X_1861_ state\[89\] daisychain\[89\] net143 _0562_ VPWR VGND sg13g2_mux2_1
X_1792_ _0507_ net173 _0506_ VPWR VGND sg13g2_nand2_1
X_2413_ net382 VGND VPWR _0229_ daisychain\[101\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2344_ net264 VGND VPWR _0160_ daisychain\[32\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_37_231 VPWR VGND sg13g2_decap_8
XFILLER_38_787 VPWR VGND sg13g2_fill_2
X_2275_ VGND VPWR _0643_ _0827_ _0365_ net76 sg13g2_a21oi_1
XFILLER_20_131 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_0_569 VPWR VGND sg13g2_fill_1
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_16_437 VPWR VGND sg13g2_fill_1
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_44_779 VPWR VGND sg13g2_fill_1
XFILLER_11_164 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_7_124 VPWR VGND sg13g2_decap_8
XFILLER_3_330 VPWR VGND sg13g2_decap_8
XFILLER_19_253 VPWR VGND sg13g2_decap_8
XFILLER_34_201 VPWR VGND sg13g2_decap_8
XFILLER_35_746 VPWR VGND sg13g2_decap_8
XFILLER_35_757 VPWR VGND sg13g2_fill_2
XFILLER_47_551 VPWR VGND sg13g2_decap_8
XFILLER_47_562 VPWR VGND sg13g2_fill_1
XFILLER_47_595 VPWR VGND sg13g2_decap_4
X_2060_ _0720_ net94 state\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_34_278 VPWR VGND sg13g2_decap_8
X_1913_ VGND VPWR net109 daisychain\[98\] _0604_ net54 sg13g2_a21oi_1
X_1844_ net196 VPWR _0549_ VGND daisychain\[85\] net39 sg13g2_o21ai_1
X_1775_ VGND VPWR _0491_ _0492_ _0199_ _0493_ sg13g2_a21oi_1
X_2327_ net298 VGND VPWR _0143_ daisychain\[15\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2258_ _0819_ net110 state\[101\] VPWR VGND sg13g2_nand2_1
XFILLER_25_256 VPWR VGND sg13g2_decap_8
XFILLER_25_267 VPWR VGND sg13g2_fill_2
XFILLER_25_278 VPWR VGND sg13g2_decap_8
X_2431__347 VPWR VGND net346 sg13g2_tiehi
X_2189_ VGND VPWR _0471_ _0784_ _0322_ net86 sg13g2_a21oi_1
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_16_223 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_12_462 VPWR VGND sg13g2_decap_8
XFILLER_17_71 VPWR VGND sg13g2_decap_8
XFILLER_8_411 VPWR VGND sg13g2_decap_8
X_2332__289 VPWR VGND net288 sg13g2_tiehi
XFILLER_33_81 VPWR VGND sg13g2_decap_8
X_1560_ VGND VPWR _0963_ _0964_ _0156_ _0965_ sg13g2_a21oi_1
XFILLER_39_315 VPWR VGND sg13g2_decap_8
X_1491_ state\[15\] daisychain\[15\] net137 _0910_ VPWR VGND sg13g2_mux2_1
X_2112_ _0746_ net102 state\[28\] VPWR VGND sg13g2_nand2_1
XFILLER_35_587 VPWR VGND sg13g2_fill_1
XFILLER_47_392 VPWR VGND sg13g2_decap_8
X_2493__374 VPWR VGND net373 sg13g2_tiehi
X_2043_ VGND VPWR net90 daisychain\[124\] _0708_ net48 sg13g2_a21oi_1
XFILLER_30_270 VPWR VGND sg13g2_decap_8
XFILLER_31_793 VPWR VGND sg13g2_decap_4
X_1827_ _0535_ net174 _0534_ VPWR VGND sg13g2_nand2_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
X_1758_ VGND VPWR net129 daisychain\[67\] _0480_ net62 sg13g2_a21oi_1
X_1689_ net194 VPWR _0425_ VGND daisychain\[54\] net37 sg13g2_o21ai_1
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_46_808 VPWR VGND sg13g2_decap_8
XFILLER_13_237 VPWR VGND sg13g2_decap_8
XFILLER_14_705 VPWR VGND sg13g2_decap_4
XFILLER_14_738 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_4
XFILLER_41_557 VPWR VGND sg13g2_fill_1
XFILLER_41_568 VPWR VGND sg13g2_decap_4
XFILLER_21_292 VPWR VGND sg13g2_decap_8
XFILLER_5_447 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_49_646 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_29_392 VPWR VGND sg13g2_fill_2
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_20_719 VPWR VGND sg13g2_fill_1
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_9_742 VPWR VGND sg13g2_decap_8
XFILLER_8_285 VPWR VGND sg13g2_decap_8
X_1474_ net180 VPWR _0897_ VGND daisychain\[11\] net23 sg13g2_o21ai_1
X_1543_ VGND VPWR net100 daisychain\[24\] _0952_ net50 sg13g2_a21oi_1
X_2384__441 VPWR VGND net440 sg13g2_tiehi
X_1612_ _1007_ net169 _1006_ VPWR VGND sg13g2_nand2_1
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_35_384 VPWR VGND sg13g2_fill_2
X_2026_ state\[122\] daisychain\[122\] net135 _0694_ VPWR VGND sg13g2_mux2_1
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_2_406 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_19_819 VPWR VGND sg13g2_fill_1
XFILLER_39_690 VPWR VGND sg13g2_decap_8
XFILLER_42_822 VPWR VGND sg13g2_fill_1
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_46_616 VPWR VGND sg13g2_decap_4
XFILLER_14_72 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_30_60 VPWR VGND sg13g2_decap_8
XFILLER_5_244 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_32_343 VPWR VGND sg13g2_decap_8
XFILLER_33_822 VPWR VGND sg13g2_fill_1
XFILLER_45_660 VPWR VGND sg13g2_decap_8
XFILLER_20_527 VPWR VGND sg13g2_fill_2
X_1457_ _0883_ net161 _0882_ VPWR VGND sg13g2_nand2_1
X_1526_ state\[22\] daisychain\[22\] net139 _0938_ VPWR VGND sg13g2_mux2_1
XFILLER_27_104 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
X_1388_ VPWR _0044_ state\[24\] VGND sg13g2_inv_1
X_2009_ net181 VPWR _0681_ VGND daisychain\[118\] net24 sg13g2_o21ai_1
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_14_310 VPWR VGND sg13g2_decap_8
XFILLER_18_159 VPWR VGND sg13g2_decap_8
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_42_641 VPWR VGND sg13g2_fill_2
XFILLER_10_593 VPWR VGND sg13g2_fill_2
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_531 VPWR VGND sg13g2_decap_8
X_1311_ VPWR _0002_ state\[101\] VGND sg13g2_inv_1
X_2360_ net232 VGND VPWR _0176_ daisychain\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2291_ VGND VPWR _0675_ _0835_ _0373_ net69 sg13g2_a21oi_1
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XFILLER_37_446 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_20_313 VPWR VGND sg13g2_decap_4
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_33_674 VPWR VGND sg13g2_fill_1
XFILLER_21_18 VPWR VGND sg13g2_decap_4
X_1509_ net183 VPWR _0925_ VGND daisychain\[18\] net26 sg13g2_o21ai_1
X_2558_ net407 VGND VPWR _0374_ state\[118\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2489_ net389 VGND VPWR _0305_ state\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_15_107 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_11_346 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_7_306 VPWR VGND sg13g2_decap_8
XFILLER_11_73 VPWR VGND sg13g2_decap_8
XFILLER_3_512 VPWR VGND sg13g2_fill_2
XFILLER_3_545 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_47_722 VPWR VGND sg13g2_decap_8
XFILLER_14_184 VPWR VGND sg13g2_decap_8
XFILLER_30_622 VPWR VGND sg13g2_fill_1
XFILLER_30_655 VPWR VGND sg13g2_fill_1
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
X_2489__390 VPWR VGND net389 sg13g2_tiehi
X_1860_ VGND VPWR _0559_ _0560_ _0216_ _0561_ sg13g2_a21oi_1
XFILLER_6_394 VPWR VGND sg13g2_decap_8
X_1791_ state\[75\] daisychain\[75\] net151 _0506_ VPWR VGND sg13g2_mux2_1
X_2412_ net384 VGND VPWR _0228_ daisychain\[100\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2343_ net266 VGND VPWR _0159_ daisychain\[31\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2342__269 VPWR VGND net268 sg13g2_tiehi
X_2274_ _0827_ net109 state\[109\] VPWR VGND sg13g2_nand2_1
XFILLER_37_210 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_38_755 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_2_1__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_20_110 VPWR VGND sg13g2_decap_8
XFILLER_20_187 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
X_1989_ net181 VPWR _0665_ VGND daisychain\[114\] net24 sg13g2_o21ai_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
X_2505__324 VPWR VGND net323 sg13g2_tiehi
XFILLER_16_405 VPWR VGND sg13g2_decap_8
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_44_703 VPWR VGND sg13g2_decap_8
XFILLER_16_416 VPWR VGND sg13g2_fill_2
XFILLER_28_298 VPWR VGND sg13g2_fill_2
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_11_143 VPWR VGND sg13g2_decap_8
XFILLER_7_103 VPWR VGND sg13g2_decap_8
XFILLER_3_386 VPWR VGND sg13g2_decap_8
XFILLER_19_232 VPWR VGND sg13g2_decap_8
XFILLER_34_257 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
X_2517__228 VPWR VGND net227 sg13g2_tiehi
X_1912_ _0603_ net167 _0602_ VPWR VGND sg13g2_nand2_1
X_1843_ VGND VPWR net124 daisychain\[84\] _0548_ net61 sg13g2_a21oi_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_6_191 VPWR VGND sg13g2_decap_8
XFILLER_8_96 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_6_clk clknet_2_3__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_1774_ net199 VPWR _0493_ VGND daisychain\[71\] net42 sg13g2_o21ai_1
X_2394__421 VPWR VGND net420 sg13g2_tiehi
X_2326_ net300 VGND VPWR _0142_ daisychain\[14\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2257_ VGND VPWR _0607_ _0818_ _0356_ net77 sg13g2_a21oi_1
XFILLER_13_408 VPWR VGND sg13g2_fill_2
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
X_2188_ _0784_ net129 state\[66\] VPWR VGND sg13g2_nand2_1
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_16_202 VPWR VGND sg13g2_decap_8
XFILLER_17_736 VPWR VGND sg13g2_decap_8
XFILLER_44_511 VPWR VGND sg13g2_decap_8
XFILLER_44_566 VPWR VGND sg13g2_decap_4
XFILLER_16_279 VPWR VGND sg13g2_decap_8
XFILLER_31_249 VPWR VGND sg13g2_decap_8
XFILLER_32_728 VPWR VGND sg13g2_fill_1
XFILLER_33_60 VPWR VGND sg13g2_decap_8
XFILLER_40_750 VPWR VGND sg13g2_decap_8
XFILLER_40_794 VPWR VGND sg13g2_fill_1
X_1490_ VGND VPWR _0907_ _0908_ _0142_ _0909_ sg13g2_a21oi_1
XFILLER_12_4 VPWR VGND sg13g2_decap_4
XFILLER_3_183 VPWR VGND sg13g2_decap_8
X_2111_ VGND VPWR _0959_ _0745_ _0283_ net72 sg13g2_a21oi_1
X_2042_ _0707_ net157 _0706_ VPWR VGND sg13g2_nand2_1
XFILLER_35_500 VPWR VGND sg13g2_fill_2
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_30_293 VPWR VGND sg13g2_fill_1
XFILLER_31_750 VPWR VGND sg13g2_decap_8
XFILLER_31_772 VPWR VGND sg13g2_decap_4
X_1826_ state\[82\] daisychain\[82\] net151 _0534_ VPWR VGND sg13g2_mux2_1
X_2502__338 VPWR VGND net337 sg13g2_tiehi
X_1757_ _0479_ net175 _0478_ VPWR VGND sg13g2_nand2_1
X_1688_ VGND VPWR net118 daisychain\[53\] _0424_ net59 sg13g2_a21oi_1
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
X_2309_ VGND VPWR _0711_ _0844_ _0382_ net70 sg13g2_a21oi_1
XFILLER_13_216 VPWR VGND sg13g2_decap_8
XFILLER_5_426 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_49_658 VPWR VGND sg13g2_decap_4
XFILLER_17_522 VPWR VGND sg13g2_decap_4
XFILLER_17_544 VPWR VGND sg13g2_decap_4
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_fill_2
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_13_794 VPWR VGND sg13g2_fill_2
XFILLER_8_264 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_4
X_1611_ state\[39\] daisychain\[39\] net146 _1006_ VPWR VGND sg13g2_mux2_1
XFILLER_4_492 VPWR VGND sg13g2_decap_8
XFILLER_5_97 VPWR VGND sg13g2_decap_8
X_1473_ VGND VPWR net92 daisychain\[10\] _0896_ net45 sg13g2_a21oi_1
X_1542_ _0951_ net161 _0950_ VPWR VGND sg13g2_nand2_1
XFILLER_39_168 VPWR VGND sg13g2_decap_8
X_2025_ VGND VPWR _0691_ _0692_ _0249_ _0693_ sg13g2_a21oi_1
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
X_2465__230 VPWR VGND net229 sg13g2_tiehi
X_1809_ net198 VPWR _0521_ VGND daisychain\[78\] net41 sg13g2_o21ai_1
X_2400__409 VPWR VGND net408 sg13g2_tiehi
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_5_223 VPWR VGND sg13g2_decap_8
X_2444__314 VPWR VGND net313 sg13g2_tiehi
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_32_377 VPWR VGND sg13g2_decap_4
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_9_551 VPWR VGND sg13g2_decap_4
X_1387_ VPWR _0045_ state\[25\] VGND sg13g2_inv_1
X_1456_ state\[8\] daisychain\[8\] net137 _0882_ VPWR VGND sg13g2_mux2_1
X_1525_ VGND VPWR _0935_ _0936_ _0149_ _0937_ sg13g2_a21oi_1
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
X_2352__249 VPWR VGND net248 sg13g2_tiehi
X_2008_ VGND VPWR net95 daisychain\[117\] _0680_ net47 sg13g2_a21oi_1
X_2508__300 VPWR VGND net299 sg13g2_tiehi
XFILLER_2_259 VPWR VGND sg13g2_decap_8
XFILLER_3_705 VPWR VGND sg13g2_fill_2
XFILLER_3_749 VPWR VGND sg13g2_decap_8
X_2543__224 VPWR VGND net223 sg13g2_tiehi
XFILLER_18_138 VPWR VGND sg13g2_decap_8
XFILLER_14_355 VPWR VGND sg13g2_fill_1
XFILLER_14_366 VPWR VGND sg13g2_decap_4
XFILLER_25_83 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_6_587 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
X_1310_ VPWR _0003_ state\[102\] VGND sg13g2_inv_1
Xheichips25_pudding VPWR VGND uio_oe[0] sg13g2_tiehi
X_2290_ _0835_ net95 state\[117\] VPWR VGND sg13g2_nand2_1
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_20_358 VPWR VGND sg13g2_decap_8
XFILLER_32_130 VPWR VGND sg13g2_decap_8
XFILLER_9_392 VPWR VGND sg13g2_decap_8
X_2557_ net439 VGND VPWR _0373_ state\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_46_49 VPWR VGND sg13g2_decap_8
X_1439_ net181 VPWR _0869_ VGND daisychain\[4\] net24 sg13g2_o21ai_1
X_1508_ VGND VPWR net99 daisychain\[17\] _0924_ net49 sg13g2_a21oi_1
X_2538__304 VPWR VGND net303 sg13g2_tiehi
X_2488_ net393 VGND VPWR _0304_ state\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_16_609 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_11_325 VPWR VGND sg13g2_decap_8
XFILLER_8_808 VPWR VGND sg13g2_decap_8
XFILLER_11_52 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_14_163 VPWR VGND sg13g2_decap_8
XFILLER_30_601 VPWR VGND sg13g2_fill_1
XFILLER_30_689 VPWR VGND sg13g2_fill_1
XFILLER_42_461 VPWR VGND sg13g2_decap_8
XFILLER_42_494 VPWR VGND sg13g2_decap_4
X_1790_ VGND VPWR _0503_ _0504_ _0202_ _0505_ sg13g2_a21oi_1
XFILLER_6_373 VPWR VGND sg13g2_decap_8
X_2411_ net386 VGND VPWR _0227_ daisychain\[99\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_38_712 VPWR VGND sg13g2_fill_1
X_2496__362 VPWR VGND net361 sg13g2_tiehi
X_2342_ net268 VGND VPWR _0158_ daisychain\[30\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2273_ VGND VPWR _0639_ _0826_ _0364_ net76 sg13g2_a21oi_1
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_38_767 VPWR VGND sg13g2_decap_4
XFILLER_38_789 VPWR VGND sg13g2_fill_1
XFILLER_20_166 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
X_1988_ VGND VPWR net95 daisychain\[113\] _0664_ net46 sg13g2_a21oi_1
XFILLER_28_200 VPWR VGND sg13g2_decap_8
XFILLER_28_277 VPWR VGND sg13g2_decap_4
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_44_737 VPWR VGND sg13g2_fill_2
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
X_2475__446 VPWR VGND net445 sg13g2_tiehi
XFILLER_11_122 VPWR VGND sg13g2_decap_8
XFILLER_12_645 VPWR VGND sg13g2_decap_8
XFILLER_11_199 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_7_159 VPWR VGND sg13g2_decap_8
X_2523__436 VPWR VGND net435 sg13g2_tiehi
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_19_211 VPWR VGND sg13g2_decap_8
XFILLER_3_365 VPWR VGND sg13g2_decap_8
Xfanout190 net191 net190 VPWR VGND sg13g2_buf_1
XFILLER_19_288 VPWR VGND sg13g2_decap_8
XFILLER_34_236 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_4
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_30_475 VPWR VGND sg13g2_decap_8
XFILLER_30_486 VPWR VGND sg13g2_decap_8
XFILLER_42_280 VPWR VGND sg13g2_decap_8
XFILLER_7_660 VPWR VGND sg13g2_decap_8
XFILLER_8_75 VPWR VGND sg13g2_decap_8
X_1911_ state\[99\] daisychain\[99\] net144 _0602_ VPWR VGND sg13g2_mux2_1
X_1842_ _0547_ net173 _0546_ VPWR VGND sg13g2_nand2_1
X_1773_ VGND VPWR net129 daisychain\[70\] _0492_ net63 sg13g2_a21oi_1
XFILLER_6_170 VPWR VGND sg13g2_decap_8
XFILLER_25_214 VPWR VGND sg13g2_decap_8
X_2325_ net302 VGND VPWR _0141_ daisychain\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2256_ _0818_ net112 state\[100\] VPWR VGND sg13g2_nand2_1
X_2187_ VGND VPWR _0467_ _0783_ _0321_ net87 sg13g2_a21oi_1
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_4_129 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_4
XFILLER_16_258 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_fill_1
XFILLER_31_228 VPWR VGND sg13g2_decap_8
XFILLER_8_446 VPWR VGND sg13g2_decap_8
XFILLER_3_162 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
X_2110_ _0745_ net100 state\[27\] VPWR VGND sg13g2_nand2_1
X_2041_ state\[125\] daisychain\[125\] net135 _0706_ VPWR VGND sg13g2_mux2_1
XFILLER_35_578 VPWR VGND sg13g2_decap_8
X_1825_ VGND VPWR _0531_ _0532_ _0209_ _0533_ sg13g2_a21oi_1
X_1756_ state\[68\] daisychain\[68\] net153 _0478_ VPWR VGND sg13g2_mux2_1
XFILLER_38_28 VPWR VGND sg13g2_decap_8
X_2308_ _0844_ net91 state\[126\] VPWR VGND sg13g2_nand2_1
X_1687_ _0423_ net171 _0422_ VPWR VGND sg13g2_nand2_1
XFILLER_38_350 VPWR VGND sg13g2_decap_8
X_2239_ VGND VPWR _0571_ _0809_ _0347_ net84 sg13g2_a21oi_1
XFILLER_21_261 VPWR VGND sg13g2_decap_8
X_2331__291 VPWR VGND net290 sg13g2_tiehi
XFILLER_5_405 VPWR VGND sg13g2_decap_8
X_2407__395 VPWR VGND net394 sg13g2_tiehi
X_2362__229 VPWR VGND net228 sg13g2_tiehi
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_17_501 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_13_740 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_12_294 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_8_243 VPWR VGND sg13g2_decap_8
X_1610_ VGND VPWR _1003_ _1004_ _0166_ _1005_ sg13g2_a21oi_1
XFILLER_5_76 VPWR VGND sg13g2_decap_8
X_1472_ _0895_ net158 _0894_ VPWR VGND sg13g2_nand2_1
X_1541_ state\[25\] daisychain\[25\] net138 _0950_ VPWR VGND sg13g2_mux2_1
XFILLER_35_364 VPWR VGND sg13g2_decap_8
XFILLER_39_147 VPWR VGND sg13g2_decap_8
X_2024_ net179 VPWR _0693_ VGND daisychain\[121\] net25 sg13g2_o21ai_1
XFILLER_31_592 VPWR VGND sg13g2_decap_4
X_1808_ VGND VPWR net128 daisychain\[77\] _0520_ net62 sg13g2_a21oi_1
X_1739_ net199 VPWR _0465_ VGND daisychain\[64\] net42 sg13g2_o21ai_1
X_2472__202 VPWR VGND net sg13g2_tiehi
XFILLER_14_548 VPWR VGND sg13g2_decap_8
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_42_813 VPWR VGND sg13g2_decap_8
XFILLER_10_710 VPWR VGND sg13g2_fill_1
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_5_202 VPWR VGND sg13g2_decap_8
XFILLER_6_725 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_30_95 VPWR VGND sg13g2_decap_8
XFILLER_5_279 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_fill_2
XFILLER_33_813 VPWR VGND sg13g2_decap_8
XFILLER_37_607 VPWR VGND sg13g2_fill_2
XFILLER_37_618 VPWR VGND sg13g2_fill_2
XFILLER_45_673 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_fill_1
XFILLER_32_334 VPWR VGND sg13g2_fill_1
XFILLER_44_161 VPWR VGND sg13g2_decap_8
XFILLER_9_574 VPWR VGND sg13g2_fill_2
X_1524_ net185 VPWR _0937_ VGND daisychain\[21\] net28 sg13g2_o21ai_1
XFILLER_4_290 VPWR VGND sg13g2_decap_8
X_1386_ VPWR _0046_ state\[26\] VGND sg13g2_inv_1
X_1455_ VGND VPWR _0879_ _0880_ _0135_ _0881_ sg13g2_a21oi_1
XFILLER_23_301 VPWR VGND sg13g2_fill_1
XFILLER_27_139 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
X_2007_ _0679_ net159 _0678_ VPWR VGND sg13g2_nand2_1
XFILLER_2_238 VPWR VGND sg13g2_decap_8
XFILLER_18_117 VPWR VGND sg13g2_decap_8
XFILLER_33_109 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_14_345 VPWR VGND sg13g2_decap_4
XFILLER_25_62 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_decap_8
XFILLER_26_183 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
X_2526__412 VPWR VGND net411 sg13g2_tiehi
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_17_183 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_decap_8
XFILLER_18_684 VPWR VGND sg13g2_decap_8
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_33_687 VPWR VGND sg13g2_decap_4
XFILLER_9_371 VPWR VGND sg13g2_decap_8
X_1507_ _0923_ net162 _0922_ VPWR VGND sg13g2_nand2_1
X_2556_ net215 VGND VPWR _0372_ state\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2487_ net397 VGND VPWR _0303_ state\[47\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_46_28 VPWR VGND sg13g2_decap_8
X_1369_ VPWR _0065_ state\[43\] VGND sg13g2_inv_1
X_1438_ VGND VPWR net95 daisychain\[3\] _0868_ net46 sg13g2_a21oi_1
XFILLER_11_304 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_36_492 VPWR VGND sg13g2_decap_8
XFILLER_3_514 VPWR VGND sg13g2_fill_1
XFILLER_2_4 VPWR VGND sg13g2_decap_4
Xdac dac/VbiasP[1] dac/Iout dac/VbiasP[0] dac/VcascP[1] dac/VcascP[0] state\[64\]
+ _0088_ state\[65\] _0089_ state\[66\] _0090_ state\[67\] _0091_ state\[68\] _0092_
+ state\[69\] _0093_ state\[70\] _0095_ state\[71\] _0096_ state\[72\] _0097_ digitalen.g\[2\].u.OUTP
+ digitalen.g\[2\].u.OUTN state\[73\] _0098_ state\[74\] _0099_ state\[75\] _0100_
+ state\[76\] _0101_ state\[77\] _0102_ state\[78\] _0103_ state\[79\] _0104_ state\[80\]
+ _0106_ state\[81\] _0107_ state\[82\] _0108_ state\[83\] _0109_ state\[84\] _0110_
+ state\[85\] _0111_ state\[86\] _0112_ state\[87\] _0113_ state\[88\] _0114_ state\[89\]
+ _0115_ state\[90\] _0117_ state\[91\] _0118_ state\[92\] _0119_ state\[93\] _0120_
+ state\[94\] _0121_ state\[95\] _0122_ state\[96\] _0123_ state\[97\] _0124_ state\[98\]
+ _0125_ state\[99\] _0126_ state\[100\] _0001_ state\[101\] _0002_ state\[102\] _0003_
+ state\[103\] _0004_ state\[104\] _0005_ state\[105\] _0006_ state\[106\] _0007_
+ state\[107\] _0008_ state\[108\] _0009_ state\[109\] _0010_ state\[110\] _0012_
+ state\[111\] _0013_ state\[112\] _0014_ state\[113\] _0015_ state\[114\] _0016_
+ state\[115\] _0017_ state\[116\] _0018_ state\[117\] _0019_ state\[118\] _0020_
+ state\[119\] _0021_ state\[120\] _0023_ state\[121\] _0024_ state\[122\] _0025_
+ digitalen.g\[3\].u.OUTP digitalen.g\[3\].u.OUTN state\[123\] _0026_ state\[124\]
+ _0027_ state\[125\] _0028_ state\[126\] _0029_ state\[127\] _0030_ state\[0\] _0000_
+ state\[1\] _0039_ state\[2\] _0050_ state\[3\] _0061_ state\[4\] _0072_ state\[5\]
+ _0083_ state\[6\] digitalen.g\[0\].u.OUTP digitalen.g\[0\].u.OUTN _0094_ state\[7\]
+ _0105_ state\[8\] _0116_ state\[9\] _0127_ state\[10\] _0011_ state\[11\] _0022_
+ state\[12\] _0031_ state\[13\] _0032_ state\[14\] _0033_ state\[15\] _0034_ state\[16\]
+ _0035_ state\[17\] _0036_ state\[18\] _0037_ state\[19\] _0038_ state\[20\] _0040_
+ state\[21\] _0041_ state\[22\] _0042_ state\[23\] _0043_ state\[24\] _0044_ state\[25\]
+ _0045_ state\[26\] _0046_ state\[27\] _0047_ state\[28\] _0048_ state\[29\] _0049_
+ state\[30\] _0051_ state\[31\] _0052_ state\[33\] _0054_ state\[32\] _0053_ state\[34\]
+ _0055_ state\[35\] _0056_ state\[36\] _0057_ state\[37\] _0058_ state\[38\] _0059_
+ state\[39\] _0060_ state\[40\] _0062_ state\[41\] _0063_ state\[42\] _0064_ state\[43\]
+ _0065_ state\[44\] _0066_ state\[45\] _0067_ state\[46\] _0068_ state\[47\] _0069_
+ state\[48\] _0070_ state\[49\] _0071_ state\[50\] _0073_ state\[51\] _0074_ state\[52\]
+ _0075_ state\[53\] _0076_ state\[54\] _0077_ state\[55\] _0078_ state\[56\] _0079_
+ state\[57\] _0080_ state\[58\] _0081_ state\[59\] _0082_ state\[60\] _0084_ state\[61\]
+ _0085_ state\[62\] _0086_ state\[63\] _0087_ digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN
+ VGND VPWR dac128module
XFILLER_15_610 VPWR VGND sg13g2_fill_1
XFILLER_19_448 VPWR VGND sg13g2_fill_2
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_14_142 VPWR VGND sg13g2_decap_8
XFILLER_30_635 VPWR VGND sg13g2_fill_1
XFILLER_30_668 VPWR VGND sg13g2_fill_1
XFILLER_10_381 VPWR VGND sg13g2_decap_8
XFILLER_6_352 VPWR VGND sg13g2_decap_8
X_2410_ net388 VGND VPWR _0226_ daisychain\[98\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2341_ net270 VGND VPWR _0157_ daisychain\[29\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_37_245 VPWR VGND sg13g2_decap_8
X_2272_ _0826_ net108 state\[108\] VPWR VGND sg13g2_nand2_1
XFILLER_18_492 VPWR VGND sg13g2_fill_1
XFILLER_20_145 VPWR VGND sg13g2_decap_8
X_1987_ _0663_ net165 _0662_ VPWR VGND sg13g2_nand2_1
XFILLER_0_539 VPWR VGND sg13g2_decap_8
X_2539_ net287 VGND VPWR _0355_ state\[99\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_256 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_11_101 VPWR VGND sg13g2_decap_8
XFILLER_11_178 VPWR VGND sg13g2_decap_8
XFILLER_12_624 VPWR VGND sg13g2_decap_8
XFILLER_7_138 VPWR VGND sg13g2_decap_8
X_2482__418 VPWR VGND net417 sg13g2_tiehi
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_3_344 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_decap_8
Xfanout180 net182 net180 VPWR VGND sg13g2_buf_1
Xfanout191 net201 net191 VPWR VGND sg13g2_buf_1
X_2372__209 VPWR VGND net208 sg13g2_tiehi
X_2341__271 VPWR VGND net270 sg13g2_tiehi
XFILLER_15_451 VPWR VGND sg13g2_decap_8
XFILLER_19_267 VPWR VGND sg13g2_decap_8
XFILLER_34_215 VPWR VGND sg13g2_decap_8
XFILLER_35_738 VPWR VGND sg13g2_decap_4
X_2417__375 VPWR VGND net374 sg13g2_tiehi
X_1910_ VGND VPWR _0599_ _0600_ _0226_ _0601_ sg13g2_a21oi_1
XFILLER_30_443 VPWR VGND sg13g2_decap_8
XFILLER_8_54 VPWR VGND sg13g2_decap_8
X_1841_ state\[85\] daisychain\[85\] net152 _0546_ VPWR VGND sg13g2_mux2_1
X_1772_ _0491_ net176 _0490_ VPWR VGND sg13g2_nand2_1
X_2324_ net304 VGND VPWR _0140_ daisychain\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_38_554 VPWR VGND sg13g2_decap_8
XFILLER_38_587 VPWR VGND sg13g2_decap_8
X_2255_ VGND VPWR _0603_ _0817_ _0355_ net77 sg13g2_a21oi_1
X_2186_ _0783_ net131 state\[65\] VPWR VGND sg13g2_nand2_1
XFILLER_33_270 VPWR VGND sg13g2_decap_8
XFILLER_41_719 VPWR VGND sg13g2_fill_1
XFILLER_4_108 VPWR VGND sg13g2_decap_8
X_2509__292 VPWR VGND net291 sg13g2_tiehi
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_16_237 VPWR VGND sg13g2_decap_8
XFILLER_17_716 VPWR VGND sg13g2_fill_2
XFILLER_17_85 VPWR VGND sg13g2_decap_8
XFILLER_31_207 VPWR VGND sg13g2_decap_8
XFILLER_12_443 VPWR VGND sg13g2_decap_4
XFILLER_33_95 VPWR VGND sg13g2_decap_8
XFILLER_8_425 VPWR VGND sg13g2_decap_8
X_2447__302 VPWR VGND net301 sg13g2_tiehi
XFILLER_3_141 VPWR VGND sg13g2_decap_8
XFILLER_39_329 VPWR VGND sg13g2_decap_8
X_2040_ VGND VPWR _0703_ _0704_ _0252_ _0705_ sg13g2_a21oi_1
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_30_284 VPWR VGND sg13g2_decap_8
X_1824_ net197 VPWR _0533_ VGND daisychain\[81\] net40 sg13g2_o21ai_1
X_1755_ VGND VPWR _0475_ _0476_ _0195_ _0477_ sg13g2_a21oi_1
X_1686_ state\[54\] daisychain\[54\] net148 _0422_ VPWR VGND sg13g2_mux2_1
X_2307_ VGND VPWR _0707_ _0843_ _0381_ net70 sg13g2_a21oi_1
X_2238_ _0809_ net126 state\[91\] VPWR VGND sg13g2_nand2_1
X_2169_ VGND VPWR _0431_ _0774_ _0312_ net81 sg13g2_a21oi_1
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_17_535 VPWR VGND sg13g2_decap_4
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_29_384 VPWR VGND sg13g2_fill_2
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_8
XFILLER_32_527 VPWR VGND sg13g2_fill_1
XFILLER_40_571 VPWR VGND sg13g2_fill_2
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_12_273 VPWR VGND sg13g2_decap_8
XFILLER_5_55 VPWR VGND sg13g2_decap_8
XFILLER_8_222 VPWR VGND sg13g2_decap_8
XFILLER_8_299 VPWR VGND sg13g2_decap_8
XFILLER_9_756 VPWR VGND sg13g2_decap_4
X_1540_ VGND VPWR _0947_ _0948_ _0152_ _0949_ sg13g2_a21oi_1
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_4_472 VPWR VGND sg13g2_decap_8
X_1471_ state\[11\] daisychain\[11\] net133 _0894_ VPWR VGND sg13g2_mux2_1
XFILLER_23_516 VPWR VGND sg13g2_fill_1
XFILLER_35_343 VPWR VGND sg13g2_decap_8
X_2023_ VGND VPWR net90 daisychain\[120\] _0692_ net48 sg13g2_a21oi_1
X_1807_ _0519_ net175 _0518_ VPWR VGND sg13g2_nand2_1
XFILLER_49_39 VPWR VGND sg13g2_decap_8
X_1738_ VGND VPWR net127 daisychain\[63\] _0464_ net63 sg13g2_a21oi_1
X_1669_ net194 VPWR _0409_ VGND daisychain\[50\] net37 sg13g2_o21ai_1
XFILLER_14_505 VPWR VGND sg13g2_fill_1
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_14_86 VPWR VGND sg13g2_decap_8
XFILLER_30_74 VPWR VGND sg13g2_decap_8
XFILLER_5_258 VPWR VGND sg13g2_decap_8
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_6_748 VPWR VGND sg13g2_decap_8
XFILLER_6_759 VPWR VGND sg13g2_fill_1
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
X_2520__204 VPWR VGND net203 sg13g2_tiehi
XFILLER_17_321 VPWR VGND sg13g2_fill_2
XFILLER_17_365 VPWR VGND sg13g2_decap_8
XFILLER_29_192 VPWR VGND sg13g2_decap_8
XFILLER_32_302 VPWR VGND sg13g2_fill_1
XFILLER_44_140 VPWR VGND sg13g2_decap_8
X_1454_ net183 VPWR _0881_ VGND daisychain\[7\] net26 sg13g2_o21ai_1
X_1523_ VGND VPWR net104 daisychain\[20\] _0936_ net50 sg13g2_a21oi_1
X_2499__350 VPWR VGND net349 sg13g2_tiehi
XFILLER_27_118 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
X_1385_ VPWR _0047_ state\[27\] VGND sg13g2_inv_1
XFILLER_35_140 VPWR VGND sg13g2_decap_8
X_2006_ state\[118\] daisychain\[118\] net136 _0678_ VPWR VGND sg13g2_mux2_1
XFILLER_31_390 VPWR VGND sg13g2_decap_8
XFILLER_3_707 VPWR VGND sg13g2_fill_1
X_2839_ state\[127\] net14 VPWR VGND sg13g2_buf_1
XFILLER_2_217 VPWR VGND sg13g2_decap_8
XFILLER_4_8 VPWR VGND sg13g2_fill_2
X_2478__434 VPWR VGND net433 sg13g2_tiehi
XFILLER_19_619 VPWR VGND sg13g2_fill_1
XFILLER_26_162 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_14_324 VPWR VGND sg13g2_decap_8
XFILLER_30_806 VPWR VGND sg13g2_fill_1
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_6_567 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_fill_1
X_2381__447 VPWR VGND net446 sg13g2_tiehi
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_fill_2
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_17_162 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_33_600 VPWR VGND sg13g2_fill_1
XFILLER_33_611 VPWR VGND sg13g2_fill_1
XFILLER_33_633 VPWR VGND sg13g2_fill_2
X_2351__251 VPWR VGND net250 sg13g2_tiehi
XFILLER_9_350 VPWR VGND sg13g2_decap_8
X_2427__355 VPWR VGND net354 sg13g2_tiehi
X_1437_ _0867_ net158 _0866_ VPWR VGND sg13g2_nand2_1
X_1506_ state\[18\] daisychain\[18\] net137 _0922_ VPWR VGND sg13g2_mux2_1
X_2555_ net247 VGND VPWR _0371_ state\[115\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2486_ net401 VGND VPWR _0302_ state\[46\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_28_405 VPWR VGND sg13g2_decap_8
XFILLER_28_416 VPWR VGND sg13g2_fill_1
XFILLER_28_449 VPWR VGND sg13g2_decap_8
X_1299_ VPWR _0015_ state\[113\] VGND sg13g2_inv_1
X_1368_ VPWR _0066_ state\[44\] VGND sg13g2_inv_1
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_11_87 VPWR VGND sg13g2_decap_8
XFILLER_3_526 VPWR VGND sg13g2_decap_4
X_2328__297 VPWR VGND net296 sg13g2_tiehi
XFILLER_19_427 VPWR VGND sg13g2_fill_2
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_14_121 VPWR VGND sg13g2_decap_8
XFILLER_15_644 VPWR VGND sg13g2_decap_8
XFILLER_30_614 VPWR VGND sg13g2_fill_1
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_10_360 VPWR VGND sg13g2_decap_8
XFILLER_14_198 VPWR VGND sg13g2_decap_8
XFILLER_30_647 VPWR VGND sg13g2_fill_1
XFILLER_6_331 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
X_2340_ net272 VGND VPWR _0156_ daisychain\[28\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2271_ VGND VPWR _0635_ _0825_ _0363_ net76 sg13g2_a21oi_1
XFILLER_18_471 VPWR VGND sg13g2_fill_2
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
XFILLER_20_124 VPWR VGND sg13g2_decap_8
X_1986_ state\[114\] daisychain\[114\] net142 _0662_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
X_2538_ net303 VGND VPWR _0354_ state\[98\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2469_ net213 VGND VPWR _0285_ state\[29\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_11_157 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_7_117 VPWR VGND sg13g2_decap_8
XFILLER_3_323 VPWR VGND sg13g2_decap_8
XFILLER_19_246 VPWR VGND sg13g2_decap_8
XFILLER_35_728 VPWR VGND sg13g2_fill_1
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_47_544 VPWR VGND sg13g2_decap_8
Xfanout170 net177 net170 VPWR VGND sg13g2_buf_1
Xfanout181 net182 net181 VPWR VGND sg13g2_buf_1
Xfanout192 net193 net192 VPWR VGND sg13g2_buf_1
X_1840_ VGND VPWR _0543_ _0544_ _0212_ _0545_ sg13g2_a21oi_1
XFILLER_7_651 VPWR VGND sg13g2_decap_4
X_1771_ state\[71\] daisychain\[71\] net154 _0490_ VPWR VGND sg13g2_mux2_1
X_2323_ net306 VGND VPWR _0139_ daisychain\[11\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2254_ _0817_ net112 state\[99\] VPWR VGND sg13g2_nand2_1
XFILLER_19_780 VPWR VGND sg13g2_decap_8
XFILLER_19_791 VPWR VGND sg13g2_fill_1
XFILLER_25_249 VPWR VGND sg13g2_decap_8
X_2185_ VGND VPWR _0463_ _0782_ _0320_ net87 sg13g2_a21oi_1
XFILLER_21_455 VPWR VGND sg13g2_fill_2
X_1969_ net188 VPWR _0649_ VGND daisychain\[110\] net31 sg13g2_o21ai_1
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_17_20 VPWR VGND sg13g2_fill_1
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_12_400 VPWR VGND sg13g2_decap_4
XFILLER_16_216 VPWR VGND sg13g2_decap_8
XFILLER_40_720 VPWR VGND sg13g2_decap_8
XFILLER_8_404 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_decap_8
XFILLER_3_120 VPWR VGND sg13g2_decap_8
XFILLER_4_643 VPWR VGND sg13g2_decap_4
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_3_197 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_15_282 VPWR VGND sg13g2_decap_8
XFILLER_30_263 VPWR VGND sg13g2_decap_8
XFILLER_31_764 VPWR VGND sg13g2_fill_2
X_1823_ VGND VPWR net126 daisychain\[80\] _0532_ net61 sg13g2_a21oi_1
XFILLER_7_481 VPWR VGND sg13g2_decap_4
X_1754_ net198 VPWR _0477_ VGND daisychain\[67\] net41 sg13g2_o21ai_1
X_1685_ VGND VPWR _0419_ _0420_ _0181_ _0421_ sg13g2_a21oi_1
X_2306_ _0843_ net91 state\[125\] VPWR VGND sg13g2_nand2_1
X_2237_ VGND VPWR _0567_ _0808_ _0346_ net85 sg13g2_a21oi_1
XFILLER_14_709 VPWR VGND sg13g2_fill_2
XFILLER_38_385 VPWR VGND sg13g2_decap_8
XFILLER_38_396 VPWR VGND sg13g2_fill_2
Xheichips25_pudding_460 VPWR VGND uio_oe[3] sg13g2_tiehi
X_2168_ _0774_ net119 state\[56\] VPWR VGND sg13g2_nand2_1
X_2099_ VGND VPWR _0935_ _0739_ _0277_ net73 sg13g2_a21oi_1
XFILLER_21_285 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_49_639 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_29_352 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_12_252 VPWR VGND sg13g2_decap_8
XFILLER_32_517 VPWR VGND sg13g2_fill_2
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_8_201 VPWR VGND sg13g2_decap_8
XFILLER_4_451 VPWR VGND sg13g2_decap_8
XFILLER_8_278 VPWR VGND sg13g2_decap_8
X_1470_ VGND VPWR _0891_ _0892_ _0138_ _0893_ sg13g2_a21oi_1
XFILLER_10_4 VPWR VGND sg13g2_fill_2
XFILLER_36_812 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_35_377 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
X_2391__427 VPWR VGND net426 sg13g2_tiehi
X_2022_ _0691_ net157 _0690_ VPWR VGND sg13g2_nand2_1
X_1806_ state\[78\] daisychain\[78\] net153 _0518_ VPWR VGND sg13g2_mux2_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
X_2361__231 VPWR VGND net230 sg13g2_tiehi
X_1737_ _0463_ net176 _0462_ VPWR VGND sg13g2_nand2_1
X_1668_ VGND VPWR net122 daisychain\[49\] _0408_ net60 sg13g2_a21oi_1
X_1599_ net192 VPWR _0997_ VGND daisychain\[36\] net35 sg13g2_o21ai_1
XFILLER_26_322 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
X_2437__335 VPWR VGND net334 sg13g2_tiehi
XFILLER_26_388 VPWR VGND sg13g2_fill_2
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_10_778 VPWR VGND sg13g2_fill_2
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_5_237 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_fill_2
XFILLER_29_171 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
X_2338__277 VPWR VGND net276 sg13g2_tiehi
XFILLER_5_771 VPWR VGND sg13g2_decap_8
XFILLER_5_782 VPWR VGND sg13g2_fill_2
XFILLER_5_793 VPWR VGND sg13g2_fill_2
X_1453_ VGND VPWR net101 daisychain\[6\] _0880_ net49 sg13g2_a21oi_1
X_1522_ _0935_ net163 _0934_ VPWR VGND sg13g2_nand2_1
X_1384_ VPWR _0048_ state\[28\] VGND sg13g2_inv_1
X_2005_ VGND VPWR _0675_ _0676_ _0245_ _0677_ sg13g2_a21oi_1
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_36_675 VPWR VGND sg13g2_fill_2
XFILLER_3_719 VPWR VGND sg13g2_fill_1
X_2838_ state\[126\] net13 VPWR VGND sg13g2_buf_1
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_14_303 VPWR VGND sg13g2_decap_8
XFILLER_26_141 VPWR VGND sg13g2_decap_8
XFILLER_39_480 VPWR VGND sg13g2_fill_1
XFILLER_42_634 VPWR VGND sg13g2_decap_8
XFILLER_10_542 VPWR VGND sg13g2_decap_4
XFILLER_10_586 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_6_524 VPWR VGND sg13g2_decap_8
X_2485__406 VPWR VGND net405 sg13g2_tiehi
XFILLER_2_730 VPWR VGND sg13g2_decap_4
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_2_13 VPWR VGND sg13g2_decap_4
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_37_439 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_17_141 VPWR VGND sg13g2_decap_8
XFILLER_20_306 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_fill_1
X_2554_ net279 VGND VPWR _0370_ state\[114\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1367_ VPWR _0067_ state\[45\] VGND sg13g2_inv_1
X_1436_ state\[4\] daisychain\[4\] net133 _0866_ VPWR VGND sg13g2_mux2_1
X_1505_ VGND VPWR _0919_ _0920_ _0145_ _0921_ sg13g2_a21oi_1
X_2485_ net405 VGND VPWR _0301_ state\[45\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_36_461 VPWR VGND sg13g2_fill_1
XFILLER_36_472 VPWR VGND sg13g2_decap_8
X_1298_ VPWR _0016_ state\[114\] VGND sg13g2_inv_1
XFILLER_11_339 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_11_66 VPWR VGND sg13g2_decap_8
XFILLER_3_505 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_14_100 VPWR VGND sg13g2_decap_8
XFILLER_14_177 VPWR VGND sg13g2_decap_8
XFILLER_15_634 VPWR VGND sg13g2_decap_4
XFILLER_30_626 VPWR VGND sg13g2_fill_1
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_42_420 VPWR VGND sg13g2_decap_8
XFILLER_42_442 VPWR VGND sg13g2_decap_8
XFILLER_30_659 VPWR VGND sg13g2_fill_2
XFILLER_6_310 VPWR VGND sg13g2_decap_8
XFILLER_6_387 VPWR VGND sg13g2_decap_8
XFILLER_2_560 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_2270_ _0825_ net107 state\[107\] VPWR VGND sg13g2_nand2_1
XFILLER_18_461 VPWR VGND sg13g2_fill_2
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_38_748 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_46_792 VPWR VGND sg13g2_decap_4
XFILLER_20_103 VPWR VGND sg13g2_decap_8
XFILLER_33_431 VPWR VGND sg13g2_fill_1
XFILLER_33_475 VPWR VGND sg13g2_fill_1
X_1985_ VGND VPWR _0659_ _0660_ _0241_ _0661_ sg13g2_a21oi_1
X_2537_ net319 VGND VPWR _0353_ state\[97\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_28_214 VPWR VGND sg13g2_decap_8
X_1419_ net180 VPWR _0853_ VGND daisychain\[0\] net23 sg13g2_o21ai_1
X_2468_ net217 VGND VPWR _0284_ state\[28\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2399_ net410 VGND VPWR _0215_ daisychain\[87\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_11_136 VPWR VGND sg13g2_decap_8
XFILLER_12_659 VPWR VGND sg13g2_fill_2
XFILLER_20_681 VPWR VGND sg13g2_fill_1
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_3_302 VPWR VGND sg13g2_decap_8
XFILLER_3_379 VPWR VGND sg13g2_decap_8
XFILLER_19_225 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
Xfanout160 net178 net160 VPWR VGND sg13g2_buf_1
Xfanout171 net172 net171 VPWR VGND sg13g2_buf_1
Xfanout182 net201 net182 VPWR VGND sg13g2_buf_1
Xfanout193 net200 net193 VPWR VGND sg13g2_buf_1
XFILLER_30_434 VPWR VGND sg13g2_decap_4
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_8_34 VPWR VGND sg13g2_fill_1
X_1770_ VGND VPWR _0487_ _0488_ _0198_ _0489_ sg13g2_a21oi_1
XFILLER_6_184 VPWR VGND sg13g2_decap_8
XFILLER_7_674 VPWR VGND sg13g2_fill_2
XFILLER_8_89 VPWR VGND sg13g2_decap_8
X_2322_ net308 VGND VPWR _0138_ daisychain\[10\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2320__313 VPWR VGND net312 sg13g2_tiehi
X_2253_ VGND VPWR _0599_ _0816_ _0354_ net76 sg13g2_a21oi_1
X_2184_ _0782_ net127 state\[64\] VPWR VGND sg13g2_nand2_1
Xdigitalen.g\[0\].u.inv1 VPWR digitalen.g\[0\].u.OUTN net6 VGND sg13g2_inv_1
X_1968_ VGND VPWR net109 daisychain\[109\] _0648_ net56 sg13g2_a21oi_1
X_1899_ net190 VPWR _0593_ VGND daisychain\[96\] net33 sg13g2_o21ai_1
XFILLER_1_817 VPWR VGND sg13g2_decap_4
X_2371__211 VPWR VGND net210 sg13g2_tiehi
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_40_787 VPWR VGND sg13g2_decap_8
XFILLER_44_559 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_1
XFILLER_3_176 VPWR VGND sg13g2_decap_8
XFILLER_48_821 VPWR VGND sg13g2_fill_2
XFILLER_15_261 VPWR VGND sg13g2_decap_8
XFILLER_16_740 VPWR VGND sg13g2_fill_2
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_30_242 VPWR VGND sg13g2_decap_8
XFILLER_31_743 VPWR VGND sg13g2_decap_8
XFILLER_31_776 VPWR VGND sg13g2_fill_2
XFILLER_7_460 VPWR VGND sg13g2_decap_8
X_2348__257 VPWR VGND net256 sg13g2_tiehi
X_1822_ _0531_ net174 _0530_ VPWR VGND sg13g2_nand2_1
X_1753_ VGND VPWR net129 daisychain\[66\] _0476_ net62 sg13g2_a21oi_1
X_1684_ net194 VPWR _0421_ VGND daisychain\[53\] net37 sg13g2_o21ai_1
XFILLER_38_364 VPWR VGND sg13g2_decap_8
X_2305_ VGND VPWR _0703_ _0842_ _0380_ net70 sg13g2_a21oi_1
X_2236_ _0808_ net124 state\[90\] VPWR VGND sg13g2_nand2_1
X_2167_ VGND VPWR _0427_ _0773_ _0311_ net81 sg13g2_a21oi_1
XFILLER_13_209 VPWR VGND sg13g2_decap_8
XFILLER_21_220 VPWR VGND sg13g2_decap_8
XFILLER_34_592 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_461 VPWR VGND uio_oe[4] sg13g2_tiehi
X_2098_ _0739_ net103 state\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_21_275 VPWR VGND sg13g2_fill_2
XFILLER_5_419 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_13_710 VPWR VGND sg13g2_fill_1
XFILLER_17_515 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_29_386 VPWR VGND sg13g2_fill_1
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
XFILLER_12_231 VPWR VGND sg13g2_decap_8
XFILLER_13_765 VPWR VGND sg13g2_decap_4
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_8_257 VPWR VGND sg13g2_decap_8
XFILLER_9_736 VPWR VGND sg13g2_fill_1
XFILLER_4_430 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
X_2501__342 VPWR VGND net341 sg13g2_tiehi
X_2021_ state\[121\] daisychain\[121\] net135 _0690_ VPWR VGND sg13g2_mux2_1
X_1805_ VGND VPWR _0515_ _0516_ _0205_ _0517_ sg13g2_a21oi_1
X_1736_ state\[64\] daisychain\[64\] net154 _0462_ VPWR VGND sg13g2_mux2_1
X_1667_ _0407_ net171 _0406_ VPWR VGND sg13g2_nand2_1
X_1598_ VGND VPWR net116 daisychain\[35\] _0996_ net57 sg13g2_a21oi_1
XFILLER_14_518 VPWR VGND sg13g2_decap_4
XFILLER_26_356 VPWR VGND sg13g2_decap_4
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
X_2219_ VGND VPWR _0531_ _0799_ _0337_ net84 sg13g2_a21oi_1
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_5_216 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_29_150 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_45_654 VPWR VGND sg13g2_fill_2
XFILLER_40_392 VPWR VGND sg13g2_decap_8
X_1383_ VPWR _0049_ state\[29\] VGND sg13g2_inv_1
X_1452_ _0879_ net161 _0878_ VPWR VGND sg13g2_nand2_1
X_1521_ state\[21\] daisychain\[21\] net139 _0934_ VPWR VGND sg13g2_mux2_1
XFILLER_36_632 VPWR VGND sg13g2_decap_4
X_2004_ net181 VPWR _0677_ VGND daisychain\[117\] net24 sg13g2_o21ai_1
XFILLER_35_175 VPWR VGND sg13g2_decap_8
X_2837_ state\[125\] net12 VPWR VGND sg13g2_buf_1
X_1719_ net195 VPWR _0449_ VGND daisychain\[60\] net38 sg13g2_o21ai_1
XFILLER_39_470 VPWR VGND sg13g2_fill_2
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_25_76 VPWR VGND sg13g2_decap_8
XFILLER_26_120 VPWR VGND sg13g2_decap_8
XFILLER_26_197 VPWR VGND sg13g2_decap_8
XFILLER_39_492 VPWR VGND sg13g2_decap_4
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_22_381 VPWR VGND sg13g2_decap_8
XFILLER_22_392 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_17_120 VPWR VGND sg13g2_decap_8
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_13_370 VPWR VGND sg13g2_fill_2
XFILLER_13_392 VPWR VGND sg13g2_fill_2
XFILLER_17_197 VPWR VGND sg13g2_decap_8
XFILLER_32_123 VPWR VGND sg13g2_decap_8
XFILLER_45_495 VPWR VGND sg13g2_decap_4
XFILLER_9_385 VPWR VGND sg13g2_decap_8
X_1504_ net183 VPWR _0921_ VGND daisychain\[17\] net26 sg13g2_o21ai_1
X_2553_ net311 VGND VPWR _0369_ state\[113\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1366_ VPWR _0068_ state\[46\] VGND sg13g2_inv_1
X_1435_ VGND VPWR _0863_ _0864_ _0131_ _0865_ sg13g2_a21oi_1
X_2484_ net409 VGND VPWR _0300_ state\[44\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_23_101 VPWR VGND sg13g2_fill_2
XFILLER_23_123 VPWR VGND sg13g2_decap_8
X_1297_ VPWR _0017_ state\[115\] VGND sg13g2_inv_1
XFILLER_11_318 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_14_156 VPWR VGND sg13g2_decap_8
XFILLER_30_605 VPWR VGND sg13g2_fill_1
XFILLER_42_454 VPWR VGND sg13g2_decap_8
XFILLER_10_395 VPWR VGND sg13g2_decap_8
XFILLER_6_366 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_38_727 VPWR VGND sg13g2_fill_2
XFILLER_33_421 VPWR VGND sg13g2_fill_1
XFILLER_33_443 VPWR VGND sg13g2_decap_4
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_20_159 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_8
X_1984_ net187 VPWR _0661_ VGND daisychain\[113\] net30 sg13g2_o21ai_1
X_2536_ net331 VGND VPWR _0352_ state\[96\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2467_ net221 VGND VPWR _0283_ state\[27\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1349_ VPWR _0087_ state\[63\] VGND sg13g2_inv_1
X_1418_ VGND VPWR net98 net2 _0852_ net48 sg13g2_a21oi_1
X_2398_ net412 VGND VPWR _0214_ daisychain\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2358__237 VPWR VGND net236 sg13g2_tiehi
XFILLER_11_115 VPWR VGND sg13g2_decap_8
XFILLER_12_638 VPWR VGND sg13g2_fill_2
XFILLER_24_410 VPWR VGND sg13g2_fill_2
XFILLER_20_660 VPWR VGND sg13g2_fill_1
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_19_204 VPWR VGND sg13g2_decap_8
XFILLER_3_358 VPWR VGND sg13g2_decap_8
X_2556__216 VPWR VGND net215 sg13g2_tiehi
Xfanout150 net155 net150 VPWR VGND sg13g2_buf_1
Xfanout161 net162 net161 VPWR VGND sg13g2_buf_1
Xfanout172 net177 net172 VPWR VGND sg13g2_buf_1
Xfanout183 net186 net183 VPWR VGND sg13g2_buf_1
XFILLER_34_229 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
Xfanout194 net195 net194 VPWR VGND sg13g2_buf_1
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_7_631 VPWR VGND sg13g2_fill_2
XFILLER_8_68 VPWR VGND sg13g2_decap_8
XFILLER_10_192 VPWR VGND sg13g2_decap_8
XFILLER_6_163 VPWR VGND sg13g2_decap_8
X_2321_ net310 VGND VPWR _0137_ daisychain\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2474__450 VPWR VGND net449 sg13g2_tiehi
X_2252_ _0816_ net109 state\[98\] VPWR VGND sg13g2_nand2_1
X_2183_ VGND VPWR _0459_ _0781_ _0319_ net83 sg13g2_a21oi_1
XFILLER_18_292 VPWR VGND sg13g2_decap_8
XFILLER_21_446 VPWR VGND sg13g2_fill_1
XFILLER_25_207 VPWR VGND sg13g2_decap_8
XFILLER_33_284 VPWR VGND sg13g2_decap_8
XFILLER_34_752 VPWR VGND sg13g2_fill_2
XFILLER_46_590 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[0\].u.inv2 VPWR digitalen.g\[0\].u.OUTP digitalen.g\[0\].u.OUTN VGND
+ sg13g2_inv_1
X_1967_ _0647_ net168 _0646_ VPWR VGND sg13g2_nand2_1
X_1898_ VGND VPWR net111 daisychain\[95\] _0592_ net55 sg13g2_a21oi_1
X_2519_ net211 VGND VPWR _0335_ state\[79\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_17_99 VPWR VGND sg13g2_decap_8
XFILLER_44_549 VPWR VGND sg13g2_decap_4
XFILLER_33_32 VPWR VGND sg13g2_decap_8
XFILLER_40_799 VPWR VGND sg13g2_fill_1
XFILLER_8_439 VPWR VGND sg13g2_decap_8
XFILLER_3_155 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_15_240 VPWR VGND sg13g2_decap_8
XFILLER_30_221 VPWR VGND sg13g2_decap_8
XFILLER_31_711 VPWR VGND sg13g2_decap_8
XFILLER_43_593 VPWR VGND sg13g2_decap_8
XFILLER_11_490 VPWR VGND sg13g2_decap_8
XFILLER_30_298 VPWR VGND sg13g2_decap_8
XFILLER_31_766 VPWR VGND sg13g2_fill_1
XFILLER_31_788 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_10_clk clknet_2_0__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_1821_ state\[81\] daisychain\[81\] net151 _0530_ VPWR VGND sg13g2_mux2_1
X_1752_ _0475_ net175 _0474_ VPWR VGND sg13g2_nand2_1
X_1683_ VGND VPWR net118 daisychain\[52\] _0420_ net59 sg13g2_a21oi_1
X_2304_ _0842_ net91 state\[124\] VPWR VGND sg13g2_nand2_1
XFILLER_38_343 VPWR VGND sg13g2_decap_8
X_2539__288 VPWR VGND net287 sg13g2_tiehi
X_2235_ VGND VPWR _0563_ _0807_ _0345_ net77 sg13g2_a21oi_1
X_2166_ _0773_ net119 state\[55\] VPWR VGND sg13g2_nand2_1
X_2097_ VGND VPWR _0931_ _0738_ _0276_ net73 sg13g2_a21oi_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_21_254 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_462 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_321 VPWR VGND sg13g2_fill_2
XFILLER_12_210 VPWR VGND sg13g2_decap_8
XFILLER_32_519 VPWR VGND sg13g2_fill_1
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_12_287 VPWR VGND sg13g2_decap_8
XFILLER_8_236 VPWR VGND sg13g2_decap_8
XFILLER_9_704 VPWR VGND sg13g2_fill_1
XFILLER_4_486 VPWR VGND sg13g2_fill_1
XFILLER_5_69 VPWR VGND sg13g2_decap_8
XFILLER_10_6 VPWR VGND sg13g2_fill_1
XFILLER_47_140 VPWR VGND sg13g2_decap_8
X_2020_ VGND VPWR _0687_ _0688_ _0248_ _0689_ sg13g2_a21oi_1
XFILLER_31_552 VPWR VGND sg13g2_decap_8
XFILLER_31_563 VPWR VGND sg13g2_fill_2
XFILLER_31_596 VPWR VGND sg13g2_fill_2
XFILLER_35_357 VPWR VGND sg13g2_decap_8
X_1804_ net198 VPWR _0517_ VGND daisychain\[77\] net41 sg13g2_o21ai_1
X_1735_ VGND VPWR _0459_ _0460_ _0191_ _0461_ sg13g2_a21oi_1
X_1666_ state\[50\] daisychain\[50\] net148 _0406_ VPWR VGND sg13g2_mux2_1
X_1597_ _0995_ net169 _0994_ VPWR VGND sg13g2_nand2_1
XFILLER_26_302 VPWR VGND sg13g2_fill_2
XFILLER_38_140 VPWR VGND sg13g2_decap_8
XFILLER_39_685 VPWR VGND sg13g2_fill_1
X_2218_ _0799_ net126 state\[81\] VPWR VGND sg13g2_nand2_1
X_2149_ VGND VPWR _0391_ _0764_ _0302_ net83 sg13g2_a21oi_1
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_30_88 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_17_302 VPWR VGND sg13g2_decap_8
XFILLER_18_814 VPWR VGND sg13g2_decap_8
XFILLER_45_600 VPWR VGND sg13g2_fill_2
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_17_379 VPWR VGND sg13g2_fill_2
XFILLER_33_806 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_44_154 VPWR VGND sg13g2_decap_8
XFILLER_9_567 VPWR VGND sg13g2_decap_8
X_1520_ VGND VPWR _0931_ _0932_ _0148_ _0933_ sg13g2_a21oi_1
XFILLER_4_283 VPWR VGND sg13g2_decap_8
X_1382_ VPWR _0051_ state\[30\] VGND sg13g2_inv_1
X_1451_ state\[7\] daisychain\[7\] net137 _0878_ VPWR VGND sg13g2_mux2_1
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_36_600 VPWR VGND sg13g2_fill_2
XFILLER_36_677 VPWR VGND sg13g2_fill_1
X_2317__319 VPWR VGND net318 sg13g2_tiehi
X_2003_ VGND VPWR net95 daisychain\[116\] _0676_ net46 sg13g2_a21oi_1
X_2836_ state\[124\] net11 VPWR VGND sg13g2_buf_1
X_1718_ VGND VPWR net119 daisychain\[59\] _0448_ net60 sg13g2_a21oi_1
X_1649_ net193 VPWR _0393_ VGND daisychain\[46\] net36 sg13g2_o21ai_1
XFILLER_10_511 VPWR VGND sg13g2_decap_8
XFILLER_14_338 VPWR VGND sg13g2_decap_8
XFILLER_14_349 VPWR VGND sg13g2_fill_2
XFILLER_22_360 VPWR VGND sg13g2_decap_8
XFILLER_22_371 VPWR VGND sg13g2_fill_2
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_25_55 VPWR VGND sg13g2_decap_8
XFILLER_26_176 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
X_2530__380 VPWR VGND net379 sg13g2_tiehi
XFILLER_10_522 VPWR VGND sg13g2_fill_2
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_6_548 VPWR VGND sg13g2_decap_4
X_2368__217 VPWR VGND net216 sg13g2_tiehi
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_17_176 VPWR VGND sg13g2_decap_8
XFILLER_18_677 VPWR VGND sg13g2_fill_2
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_9_364 VPWR VGND sg13g2_decap_8
X_1503_ VGND VPWR net99 daisychain\[16\] _0920_ net49 sg13g2_a21oi_1
X_2542__240 VPWR VGND net239 sg13g2_tiehi
X_2552_ net335 VGND VPWR _0368_ state\[112\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2483_ net413 VGND VPWR _0299_ state\[43\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1296_ VPWR _0018_ state\[116\] VGND sg13g2_inv_1
X_1365_ VPWR _0069_ state\[47\] VGND sg13g2_inv_1
X_1434_ net181 VPWR _0865_ VGND daisychain\[3\] net24 sg13g2_o21ai_1
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_11_35 VPWR VGND sg13g2_decap_4
XFILLER_2_8 VPWR VGND sg13g2_fill_1
XFILLER_15_603 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_14_135 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_fill_1
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_10_374 VPWR VGND sg13g2_decap_8
XFILLER_6_345 VPWR VGND sg13g2_decap_8
XFILLER_37_238 VPWR VGND sg13g2_decap_8
X_2537__320 VPWR VGND net319 sg13g2_tiehi
XFILLER_46_783 VPWR VGND sg13g2_decap_4
XFILLER_14_691 VPWR VGND sg13g2_fill_2
XFILLER_20_138 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
X_1983_ VGND VPWR net95 daisychain\[112\] _0660_ net53 sg13g2_a21oi_1
X_1417_ VGND VPWR _0851_ net3 net160 sg13g2_or2_1
X_2535_ net339 VGND VPWR _0351_ state\[95\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2466_ net225 VGND VPWR _0282_ state\[26\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_28_249 VPWR VGND sg13g2_decap_8
X_1348_ VPWR _0088_ state\[64\] VGND sg13g2_inv_1
X_2397_ net414 VGND VPWR _0213_ daisychain\[85\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_12_617 VPWR VGND sg13g2_decap_8
XFILLER_20_694 VPWR VGND sg13g2_fill_1
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_3_337 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
Xfanout140 net141 net140 VPWR VGND sg13g2_buf_1
Xfanout151 net155 net151 VPWR VGND sg13g2_buf_1
Xfanout162 net164 net162 VPWR VGND sg13g2_buf_1
Xfanout173 net174 net173 VPWR VGND sg13g2_buf_1
Xfanout184 net186 net184 VPWR VGND sg13g2_buf_1
Xfanout195 net200 net195 VPWR VGND sg13g2_buf_1
XFILLER_15_444 VPWR VGND sg13g2_decap_8
XFILLER_34_208 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_43_720 VPWR VGND sg13g2_fill_1
XFILLER_47_558 VPWR VGND sg13g2_decap_4
XFILLER_10_171 VPWR VGND sg13g2_decap_8
XFILLER_43_797 VPWR VGND sg13g2_fill_1
XFILLER_6_142 VPWR VGND sg13g2_decap_8
XFILLER_7_676 VPWR VGND sg13g2_fill_1
XFILLER_8_47 VPWR VGND sg13g2_decap_8
XFILLER_2_392 VPWR VGND sg13g2_decap_8
XFILLER_7_687 VPWR VGND sg13g2_fill_1
X_2504__330 VPWR VGND net329 sg13g2_tiehi
X_2320_ net312 VGND VPWR _0136_ daisychain\[8\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2251_ VGND VPWR _0595_ _0815_ _0353_ net77 sg13g2_a21oi_1
XFILLER_19_761 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ _0781_ net123 state\[63\] VPWR VGND sg13g2_nand2_1
XFILLER_18_271 VPWR VGND sg13g2_decap_8
XFILLER_33_263 VPWR VGND sg13g2_decap_8
X_1966_ state\[110\] daisychain\[110\] net145 _0646_ VPWR VGND sg13g2_mux2_1
X_2481__422 VPWR VGND net421 sg13g2_tiehi
X_1897_ _0591_ net167 _0590_ VPWR VGND sg13g2_nand2_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_503 VPWR VGND sg13g2_decap_4
X_2518_ net219 VGND VPWR _0334_ state\[78\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2449_ net293 VGND VPWR _0265_ state\[9\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_17_78 VPWR VGND sg13g2_decap_8
XFILLER_12_436 VPWR VGND sg13g2_decap_8
XFILLER_12_469 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_decap_8
XFILLER_8_418 VPWR VGND sg13g2_decap_8
X_2562__232 VPWR VGND net231 sg13g2_tiehi
XFILLER_3_134 VPWR VGND sg13g2_decap_8
XFILLER_4_602 VPWR VGND sg13g2_decap_4
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_4_624 VPWR VGND sg13g2_fill_2
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_15_296 VPWR VGND sg13g2_fill_2
XFILLER_16_731 VPWR VGND sg13g2_fill_1
XFILLER_30_200 VPWR VGND sg13g2_decap_8
XFILLER_43_572 VPWR VGND sg13g2_fill_2
XFILLER_47_399 VPWR VGND sg13g2_decap_8
X_1820_ VGND VPWR _0527_ _0528_ _0208_ _0529_ sg13g2_a21oi_1
XFILLER_30_277 VPWR VGND sg13g2_decap_8
XFILLER_7_495 VPWR VGND sg13g2_decap_8
X_1751_ state\[67\] daisychain\[67\] net153 _0474_ VPWR VGND sg13g2_mux2_1
X_1682_ _0419_ net171 _0418_ VPWR VGND sg13g2_nand2_1
XFILLER_38_322 VPWR VGND sg13g2_decap_8
X_2303_ VGND VPWR _0699_ _0841_ _0379_ net70 sg13g2_a21oi_1
X_2234_ _0807_ net111 state\[89\] VPWR VGND sg13g2_nand2_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_19_580 VPWR VGND sg13g2_decap_8
X_2165_ VGND VPWR _0423_ _0772_ _0310_ net81 sg13g2_a21oi_1
X_2096_ _0738_ net104 state\[20\] VPWR VGND sg13g2_nand2_1
XFILLER_21_299 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_463 VPWR VGND uio_oe[6] sg13g2_tiehi
X_1949_ net187 VPWR _0633_ VGND daisychain\[106\] net30 sg13g2_o21ai_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
X_2377__455 VPWR VGND net454 sg13g2_tiehi
XFILLER_17_539 VPWR VGND sg13g2_fill_1
XFILLER_40_542 VPWR VGND sg13g2_fill_2
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_12_266 VPWR VGND sg13g2_decap_8
XFILLER_8_215 VPWR VGND sg13g2_decap_8
XFILLER_9_749 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_4_465 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_16_572 VPWR VGND sg13g2_decap_4
XFILLER_31_531 VPWR VGND sg13g2_decap_4
X_1803_ VGND VPWR net128 daisychain\[76\] _0516_ net62 sg13g2_a21oi_1
XFILLER_7_292 VPWR VGND sg13g2_decap_8
XFILLER_8_793 VPWR VGND sg13g2_fill_1
X_1734_ net200 VPWR _0461_ VGND daisychain\[63\] net43 sg13g2_o21ai_1
X_1665_ VGND VPWR _0403_ _0404_ _0177_ _0405_ sg13g2_a21oi_1
X_1596_ state\[36\] daisychain\[36\] net146 _0994_ VPWR VGND sg13g2_mux2_1
X_2217_ VGND VPWR _0527_ _0798_ _0336_ net84 sg13g2_a21oi_1
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_39_697 VPWR VGND sg13g2_decap_8
X_2148_ _0764_ net117 state\[46\] VPWR VGND sg13g2_nand2_1
X_2079_ VGND VPWR _0895_ _0729_ _0267_ net68 sg13g2_a21oi_1
XFILLER_14_79 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_30_67 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_29_185 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_45_667 VPWR VGND sg13g2_fill_2
XFILLER_25_380 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_4_262 VPWR VGND sg13g2_decap_8
XFILLER_5_752 VPWR VGND sg13g2_decap_8
X_1450_ VGND VPWR _0875_ _0876_ _0134_ _0877_ sg13g2_a21oi_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
X_1381_ VPWR _0052_ state\[31\] VGND sg13g2_inv_1
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
X_2002_ _0675_ net159 _0674_ VPWR VGND sg13g2_nand2_1
X_2835_ state\[123\] net10 VPWR VGND sg13g2_buf_1
X_1717_ _0447_ net172 _0446_ VPWR VGND sg13g2_nand2_1
X_1648_ VGND VPWR net117 daisychain\[45\] _0392_ net58 sg13g2_a21oi_1
X_1579_ net186 VPWR _0981_ VGND daisychain\[32\] net29 sg13g2_o21ai_1
XFILLER_26_155 VPWR VGND sg13g2_decap_8
XFILLER_39_472 VPWR VGND sg13g2_fill_1
XFILLER_14_317 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_10_556 VPWR VGND sg13g2_fill_2
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_17_155 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_13_372 VPWR VGND sg13g2_fill_1
XFILLER_32_158 VPWR VGND sg13g2_decap_8
XFILLER_9_343 VPWR VGND sg13g2_decap_8
X_1433_ VGND VPWR net92 daisychain\[2\] _0864_ net45 sg13g2_a21oi_1
X_1502_ _0919_ net162 _0918_ VPWR VGND sg13g2_nand2_1
X_2551_ net351 VGND VPWR _0367_ state\[111\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2482_ net417 VGND VPWR _0298_ state\[42\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_49_792 VPWR VGND sg13g2_fill_2
X_1295_ VPWR _0019_ state\[117\] VGND sg13g2_inv_1
X_1364_ VPWR _0070_ state\[48\] VGND sg13g2_inv_1
XFILLER_20_821 VPWR VGND sg13g2_fill_2
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_36_486 VPWR VGND sg13g2_fill_2
XFILLER_47_729 VPWR VGND sg13g2_fill_2
XFILLER_14_114 VPWR VGND sg13g2_decap_8
XFILLER_15_615 VPWR VGND sg13g2_fill_1
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_42_434 VPWR VGND sg13g2_decap_4
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_10_353 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_fill_1
XFILLER_6_324 VPWR VGND sg13g2_decap_8
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_38_729 VPWR VGND sg13g2_fill_1
XFILLER_20_117 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_decap_8
X_1982_ _0659_ net165 _0658_ VPWR VGND sg13g2_nand2_1
XFILLER_9_140 VPWR VGND sg13g2_decap_8
X_2534_ net347 VGND VPWR _0350_ state\[94\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_3_92 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_1347_ VPWR _0089_ state\[65\] VGND sg13g2_inv_1
X_1416_ net160 net3 _0850_ VPWR VGND sg13g2_nor2_1
X_2465_ net229 VGND VPWR _0281_ state\[25\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2396_ net416 VGND VPWR _0212_ daisychain\[84\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_37_751 VPWR VGND sg13g2_decap_8
XFILLER_37_795 VPWR VGND sg13g2_fill_1
XFILLER_20_673 VPWR VGND sg13g2_fill_1
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_3_316 VPWR VGND sg13g2_decap_8
XFILLER_19_239 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
Xfanout130 net131 net130 VPWR VGND sg13g2_buf_1
Xfanout141 net156 net141 VPWR VGND sg13g2_buf_1
Xfanout152 net155 net152 VPWR VGND sg13g2_buf_1
Xfanout163 net164 net163 VPWR VGND sg13g2_buf_1
Xfanout174 net177 net174 VPWR VGND sg13g2_buf_1
Xfanout185 net186 net185 VPWR VGND sg13g2_buf_1
Xfanout196 net197 net196 VPWR VGND sg13g2_buf_1
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_43_732 VPWR VGND sg13g2_decap_8
XFILLER_10_150 VPWR VGND sg13g2_decap_8
XFILLER_11_684 VPWR VGND sg13g2_decap_4
XFILLER_6_121 VPWR VGND sg13g2_decap_8
XFILLER_7_644 VPWR VGND sg13g2_decap_8
XFILLER_7_655 VPWR VGND sg13g2_fill_1
X_2387__435 VPWR VGND net434 sg13g2_tiehi
XFILLER_2_371 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_6_198 VPWR VGND sg13g2_decap_8
X_2250_ _0815_ net112 state\[97\] VPWR VGND sg13g2_nand2_1
XFILLER_18_250 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_fill_1
XFILLER_19_740 VPWR VGND sg13g2_decap_8
XFILLER_34_710 VPWR VGND sg13g2_fill_2
X_2181_ VGND VPWR _0455_ _0780_ _0318_ net82 sg13g2_a21oi_1
XFILLER_33_242 VPWR VGND sg13g2_decap_8
X_1965_ VGND VPWR _0643_ _0644_ _0237_ _0645_ sg13g2_a21oi_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_2517_ net227 VGND VPWR _0333_ state\[77\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1896_ state\[96\] daisychain\[96\] net144 _0590_ VPWR VGND sg13g2_mux2_1
X_2448_ net297 VGND VPWR _0264_ state\[8\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2379_ net450 VGND VPWR _0195_ daisychain\[67\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_16_209 VPWR VGND sg13g2_decap_8
XFILLER_40_713 VPWR VGND sg13g2_decap_8
XFILLER_44_518 VPWR VGND sg13g2_fill_1
XFILLER_44_529 VPWR VGND sg13g2_decap_4
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_40_757 VPWR VGND sg13g2_fill_2
XFILLER_3_113 VPWR VGND sg13g2_decap_8
XFILLER_4_636 VPWR VGND sg13g2_decap_8
XFILLER_4_647 VPWR VGND sg13g2_fill_1
XFILLER_35_529 VPWR VGND sg13g2_fill_2
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_15_275 VPWR VGND sg13g2_decap_8
XFILLER_30_256 VPWR VGND sg13g2_decap_8
XFILLER_31_757 VPWR VGND sg13g2_decap_8
X_1750_ VGND VPWR _0471_ _0472_ _0194_ _0473_ sg13g2_a21oi_1
XFILLER_7_474 VPWR VGND sg13g2_decap_8
X_1681_ state\[53\] daisychain\[53\] net148 _0418_ VPWR VGND sg13g2_mux2_1
XFILLER_38_301 VPWR VGND sg13g2_decap_8
XFILLER_3_691 VPWR VGND sg13g2_decap_8
X_2302_ _0841_ net90 state\[123\] VPWR VGND sg13g2_nand2_1
X_2233_ VGND VPWR _0559_ _0806_ _0344_ net77 sg13g2_a21oi_1
X_2164_ _0772_ net118 state\[54\] VPWR VGND sg13g2_nand2_1
XFILLER_34_540 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_464 VPWR VGND uio_oe[7] sg13g2_tiehi
X_2095_ VGND VPWR _0927_ _0737_ _0275_ net71 sg13g2_a21oi_1
XFILLER_21_234 VPWR VGND sg13g2_fill_1
XFILLER_9_91 VPWR VGND sg13g2_decap_8
X_1948_ VGND VPWR net108 daisychain\[105\] _0632_ net53 sg13g2_a21oi_1
X_1879_ net197 VPWR _0577_ VGND daisychain\[92\] net40 sg13g2_o21ai_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_29_323 VPWR VGND sg13g2_fill_1
XFILLER_29_345 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_12_245 VPWR VGND sg13g2_decap_8
XFILLER_25_540 VPWR VGND sg13g2_decap_4
XFILLER_40_510 VPWR VGND sg13g2_fill_1
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_fill_2
XFILLER_4_499 VPWR VGND sg13g2_decap_8
XFILLER_16_551 VPWR VGND sg13g2_decap_8
XFILLER_31_510 VPWR VGND sg13g2_decap_4
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_36_805 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_8_772 VPWR VGND sg13g2_decap_8
X_1802_ _0515_ net175 _0514_ VPWR VGND sg13g2_nand2_1
X_1733_ VGND VPWR net122 daisychain\[62\] _0460_ net65 sg13g2_a21oi_1
XFILLER_7_271 VPWR VGND sg13g2_decap_8
X_1664_ net195 VPWR _0405_ VGND daisychain\[49\] net38 sg13g2_o21ai_1
X_1595_ VGND VPWR _0991_ _0992_ _0163_ _0993_ sg13g2_a21oi_1
XFILLER_26_315 VPWR VGND sg13g2_decap_8
XFILLER_38_175 VPWR VGND sg13g2_decap_8
X_2216_ _0798_ net126 state\[80\] VPWR VGND sg13g2_nand2_1
X_2147_ VGND VPWR _0387_ _0763_ _0301_ net83 sg13g2_a21oi_1
XFILLER_41_329 VPWR VGND sg13g2_decap_8
X_2413__383 VPWR VGND net382 sg13g2_tiehi
X_2078_ _0729_ net92 state\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_30_46 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_29_164 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_45_613 VPWR VGND sg13g2_decap_4
XFILLER_4_241 VPWR VGND sg13g2_decap_8
XFILLER_5_720 VPWR VGND sg13g2_decap_8
X_1380_ VPWR _0053_ state\[32\] VGND sg13g2_inv_1
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
X_2001_ state\[117\] daisychain\[117\] net136 _0674_ VPWR VGND sg13g2_mux2_1
XFILLER_23_329 VPWR VGND sg13g2_fill_2
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_31_384 VPWR VGND sg13g2_fill_2
XFILLER_8_580 VPWR VGND sg13g2_decap_4
X_2834_ state\[122\] net9 VPWR VGND sg13g2_buf_1
X_1716_ state\[60\] daisychain\[60\] net149 _0446_ VPWR VGND sg13g2_mux2_1
X_1647_ _0391_ net170 _0390_ VPWR VGND sg13g2_nand2_1
X_1578_ VGND VPWR net105 daisychain\[31\] _0980_ net51 sg13g2_a21oi_1
XFILLER_26_134 VPWR VGND sg13g2_decap_8
XFILLER_10_535 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_2_701 VPWR VGND sg13g2_fill_2
XFILLER_2_723 VPWR VGND sg13g2_decap_8
XFILLER_2_734 VPWR VGND sg13g2_fill_2
X_2448__298 VPWR VGND net297 sg13g2_tiehi
XFILLER_18_602 VPWR VGND sg13g2_fill_2
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_17 VPWR VGND sg13g2_fill_1
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_17_134 VPWR VGND sg13g2_decap_8
XFILLER_18_679 VPWR VGND sg13g2_fill_1
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_decap_8
X_2316__321 VPWR VGND net320 sg13g2_tiehi
XFILLER_9_322 VPWR VGND sg13g2_decap_8
XFILLER_9_399 VPWR VGND sg13g2_decap_8
X_2550_ net367 VGND VPWR _0366_ state\[110\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_49_4 VPWR VGND sg13g2_decap_8
X_1363_ VPWR _0071_ state\[49\] VGND sg13g2_inv_1
X_1432_ _0863_ net158 _0862_ VPWR VGND sg13g2_nand2_1
X_1501_ state\[17\] daisychain\[17\] net137 _0918_ VPWR VGND sg13g2_mux2_1
X_2481_ net421 VGND VPWR _0297_ state\[41\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2397__415 VPWR VGND net414 sg13g2_tiehi
X_1294_ VPWR _0020_ state\[118\] VGND sg13g2_inv_1
XFILLER_20_800 VPWR VGND sg13g2_fill_1
XFILLER_20_811 VPWR VGND sg13g2_fill_1
XFILLER_23_137 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[3\].u.inv1 VPWR digitalen.g\[3\].u.OUTN net6 VGND sg13g2_inv_1
X_2484__410 VPWR VGND net409 sg13g2_tiehi
XFILLER_11_59 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_15_638 VPWR VGND sg13g2_fill_1
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_42_468 VPWR VGND sg13g2_fill_2
XFILLER_10_332 VPWR VGND sg13g2_decap_8
XFILLER_6_303 VPWR VGND sg13g2_decap_8
X_2565__264 VPWR VGND net263 sg13g2_tiehi
XFILLER_2_553 VPWR VGND sg13g2_fill_2
XFILLER_18_454 VPWR VGND sg13g2_decap_8
XFILLER_38_708 VPWR VGND sg13g2_decap_4
XFILLER_13_181 VPWR VGND sg13g2_decap_8
XFILLER_14_671 VPWR VGND sg13g2_fill_2
XFILLER_14_693 VPWR VGND sg13g2_fill_1
XFILLER_33_413 VPWR VGND sg13g2_fill_2
XFILLER_45_273 VPWR VGND sg13g2_decap_8
X_1981_ state\[113\] daisychain\[113\] net134 _0658_ VPWR VGND sg13g2_mux2_1
XFILLER_5_391 VPWR VGND sg13g2_decap_8
XFILLER_9_196 VPWR VGND sg13g2_decap_8
X_2533_ net355 VGND VPWR _0349_ state\[93\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_28_207 VPWR VGND sg13g2_decap_8
XFILLER_3_71 VPWR VGND sg13g2_decap_8
X_1346_ VPWR _0090_ state\[66\] VGND sg13g2_inv_1
X_1415_ _0849_ net158 _0848_ VPWR VGND sg13g2_nand2_1
X_2464_ net233 VGND VPWR _0280_ state\[24\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2395_ net418 VGND VPWR _0211_ daisychain\[83\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_24_435 VPWR VGND sg13g2_fill_2
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_11_129 VPWR VGND sg13g2_decap_8
XFILLER_20_652 VPWR VGND sg13g2_fill_1
XFILLER_20_685 VPWR VGND sg13g2_fill_1
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xfanout120 net121 net120 VPWR VGND sg13g2_buf_1
Xfanout131 net132 net131 VPWR VGND sg13g2_buf_1
XFILLER_19_218 VPWR VGND sg13g2_decap_8
XFILLER_27_251 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
Xfanout142 net145 net142 VPWR VGND sg13g2_buf_1
Xfanout153 net154 net153 VPWR VGND sg13g2_buf_1
Xfanout164 net178 net164 VPWR VGND sg13g2_buf_1
Xfanout175 net176 net175 VPWR VGND sg13g2_buf_1
Xfanout186 net201 net186 VPWR VGND sg13g2_buf_1
Xfanout197 net200 net197 VPWR VGND sg13g2_buf_1
XFILLER_30_427 VPWR VGND sg13g2_decap_8
XFILLER_30_438 VPWR VGND sg13g2_fill_1
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_12_91 VPWR VGND sg13g2_decap_8
XFILLER_6_100 VPWR VGND sg13g2_decap_8
XFILLER_6_177 VPWR VGND sg13g2_decap_8
XFILLER_7_667 VPWR VGND sg13g2_decap_8
XFILLER_2_350 VPWR VGND sg13g2_decap_8
X_2180_ _0780_ net122 state\[62\] VPWR VGND sg13g2_nand2_1
XFILLER_19_796 VPWR VGND sg13g2_decap_8
XFILLER_33_221 VPWR VGND sg13g2_decap_8
XFILLER_46_571 VPWR VGND sg13g2_fill_1
XFILLER_14_490 VPWR VGND sg13g2_fill_1
XFILLER_21_416 VPWR VGND sg13g2_fill_2
XFILLER_33_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_1964_ net188 VPWR _0645_ VGND daisychain\[109\] net31 sg13g2_o21ai_1
X_1895_ VGND VPWR _0587_ _0588_ _0223_ _0589_ sg13g2_a21oi_1
X_2516_ net235 VGND VPWR _0332_ state\[76\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2447_ net301 VGND VPWR _0263_ state\[7\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_17_36 VPWR VGND sg13g2_fill_2
X_1329_ VPWR _0109_ state\[83\] VGND sg13g2_inv_1
X_2516__236 VPWR VGND net235 sg13g2_tiehi
X_2378_ net452 VGND VPWR _0194_ daisychain\[66\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_33_46 VPWR VGND sg13g2_decap_8
X_2566__392 VPWR VGND net391 sg13g2_tiehi
XFILLER_3_169 VPWR VGND sg13g2_decap_8
XFILLER_48_814 VPWR VGND sg13g2_decap_8
X_2423__363 VPWR VGND net362 sg13g2_tiehi
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_15_254 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_fill_2
XFILLER_16_799 VPWR VGND sg13g2_fill_1
XFILLER_23_90 VPWR VGND sg13g2_decap_8
XFILLER_30_235 VPWR VGND sg13g2_decap_8
XFILLER_31_725 VPWR VGND sg13g2_decap_4
XFILLER_43_574 VPWR VGND sg13g2_fill_1
XFILLER_7_453 VPWR VGND sg13g2_decap_8
X_2301_ VGND VPWR _0695_ _0840_ _0378_ net70 sg13g2_a21oi_1
X_1680_ VGND VPWR _0415_ _0416_ _0180_ _0417_ sg13g2_a21oi_1
XFILLER_31_4 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2232_ _0806_ net111 state\[88\] VPWR VGND sg13g2_nand2_1
X_2163_ VGND VPWR _0419_ _0771_ _0309_ net81 sg13g2_a21oi_1
XFILLER_21_213 VPWR VGND sg13g2_decap_8
XFILLER_34_585 VPWR VGND sg13g2_decap_8
X_2094_ _0737_ net102 state\[19\] VPWR VGND sg13g2_nand2_1
XFILLER_21_268 VPWR VGND sg13g2_decap_8
XFILLER_30_780 VPWR VGND sg13g2_fill_1
XFILLER_9_70 VPWR VGND sg13g2_decap_8
X_1947_ _0631_ net165 _0630_ VPWR VGND sg13g2_nand2_1
X_1878_ VGND VPWR net110 daisychain\[91\] _0576_ net61 sg13g2_a21oi_1
XFILLER_17_508 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_12_224 VPWR VGND sg13g2_decap_8
XFILLER_13_703 VPWR VGND sg13g2_decap_8
XFILLER_13_747 VPWR VGND sg13g2_decap_8
XFILLER_13_758 VPWR VGND sg13g2_decap_8
XFILLER_13_769 VPWR VGND sg13g2_fill_2
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_4
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_11_290 VPWR VGND sg13g2_decap_8
XFILLER_7_250 VPWR VGND sg13g2_decap_8
XFILLER_8_751 VPWR VGND sg13g2_decap_8
X_2326__301 VPWR VGND net300 sg13g2_tiehi
X_1801_ state\[77\] daisychain\[77\] net153 _0514_ VPWR VGND sg13g2_mux2_1
X_1732_ _0459_ net177 _0458_ VPWR VGND sg13g2_nand2_1
X_1663_ VGND VPWR net122 daisychain\[48\] _0404_ net60 sg13g2_a21oi_1
X_1594_ net192 VPWR _0993_ VGND daisychain\[35\] net35 sg13g2_o21ai_1
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_39_644 VPWR VGND sg13g2_decap_4
X_2215_ VGND VPWR _0523_ _0797_ _0335_ net87 sg13g2_a21oi_1
X_2146_ _0763_ net117 state\[45\] VPWR VGND sg13g2_nand2_1
X_2077_ VGND VPWR _0891_ _0728_ _0266_ net68 sg13g2_a21oi_1
XFILLER_10_728 VPWR VGND sg13g2_fill_2
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_30_25 VPWR VGND sg13g2_decap_8
XFILLER_5_209 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_29_143 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_710 VPWR VGND sg13g2_fill_1
XFILLER_4_220 VPWR VGND sg13g2_decap_8
XFILLER_4_297 VPWR VGND sg13g2_decap_8
XFILLER_36_636 VPWR VGND sg13g2_fill_2
XFILLER_48_441 VPWR VGND sg13g2_decap_8
X_2000_ VGND VPWR _0671_ _0672_ _0244_ _0673_ sg13g2_a21oi_1
XFILLER_31_352 VPWR VGND sg13g2_decap_4
XFILLER_35_168 VPWR VGND sg13g2_decap_8
X_2833_ state\[121\] net8 VPWR VGND sg13g2_buf_1
XFILLER_6_93 VPWR VGND sg13g2_decap_8
X_1715_ VGND VPWR _0443_ _0444_ _0187_ _0445_ sg13g2_a21oi_1
X_1646_ state\[46\] daisychain\[46\] net147 _0390_ VPWR VGND sg13g2_mux2_1
XFILLER_39_430 VPWR VGND sg13g2_decap_4
X_1577_ _0979_ net164 _0978_ VPWR VGND sg13g2_nand2_1
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_25_69 VPWR VGND sg13g2_decap_8
XFILLER_26_113 VPWR VGND sg13g2_decap_8
XFILLER_39_463 VPWR VGND sg13g2_decap_8
XFILLER_39_485 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
X_2129_ VGND VPWR _0995_ _0754_ _0292_ net80 sg13g2_a21oi_1
XFILLER_10_558 VPWR VGND sg13g2_fill_1
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_fill_1
XFILLER_17_113 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_13_363 VPWR VGND sg13g2_decap_8
XFILLER_32_116 VPWR VGND sg13g2_decap_8
XFILLER_45_488 VPWR VGND sg13g2_decap_8
XFILLER_9_301 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_5_562 VPWR VGND sg13g2_decap_8
XFILLER_9_378 VPWR VGND sg13g2_decap_8
X_1500_ VGND VPWR _0915_ _0916_ _0144_ _0917_ sg13g2_a21oi_1
X_2480_ net425 VGND VPWR _0296_ state\[40\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1293_ VPWR _0021_ state\[119\] VGND sg13g2_inv_1
X_1362_ VPWR _0073_ state\[50\] VGND sg13g2_inv_1
X_1431_ state\[3\] daisychain\[3\] net133 _0862_ VPWR VGND sg13g2_mux2_1
XFILLER_36_499 VPWR VGND sg13g2_decap_4
XFILLER_49_783 VPWR VGND sg13g2_fill_1
XFILLER_31_193 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[3\].u.inv2 VPWR digitalen.g\[3\].u.OUTP digitalen.g\[3\].u.OUTN VGND
+ sg13g2_inv_1
X_1629_ net192 VPWR _1021_ VGND daisychain\[42\] net35 sg13g2_o21ai_1
XFILLER_27_433 VPWR VGND sg13g2_fill_2
XFILLER_36_35 VPWR VGND sg13g2_decap_8
X_2519__212 VPWR VGND net211 sg13g2_tiehi
XFILLER_11_812 VPWR VGND sg13g2_decap_8
XFILLER_14_149 VPWR VGND sg13g2_decap_8
XFILLER_27_499 VPWR VGND sg13g2_fill_2
XFILLER_30_609 VPWR VGND sg13g2_fill_2
XFILLER_10_311 VPWR VGND sg13g2_decap_8
XFILLER_10_388 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_359 VPWR VGND sg13g2_decap_8
XFILLER_2_532 VPWR VGND sg13g2_decap_8
XFILLER_33_436 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_46_731 VPWR VGND sg13g2_decap_8
X_2433__343 VPWR VGND net342 sg13g2_tiehi
XFILLER_13_160 VPWR VGND sg13g2_decap_8
XFILLER_33_447 VPWR VGND sg13g2_fill_1
XFILLER_9_175 VPWR VGND sg13g2_decap_8
X_1980_ VGND VPWR _0655_ _0656_ _0240_ _0657_ sg13g2_a21oi_1
XFILLER_5_370 VPWR VGND sg13g2_decap_8
X_2532_ net363 VGND VPWR _0348_ state\[92\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2463_ net237 VGND VPWR _0279_ state\[23\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_3_50 VPWR VGND sg13g2_decap_8
X_1345_ VPWR _0091_ state\[67\] VGND sg13g2_inv_1
X_1414_ state\[0\] daisychain\[0\] net133 _0848_ VPWR VGND sg13g2_mux2_1
X_2394_ net420 VGND VPWR _0210_ daisychain\[82\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_11_108 VPWR VGND sg13g2_decap_8
XFILLER_24_425 VPWR VGND sg13g2_fill_1
XFILLER_36_252 VPWR VGND sg13g2_decap_8
X_2334__285 VPWR VGND net284 sg13g2_tiehi
XFILLER_20_664 VPWR VGND sg13g2_fill_1
Xfanout110 net113 net110 VPWR VGND sg13g2_buf_1
Xfanout121 net123 net121 VPWR VGND sg13g2_buf_1
Xfanout132 _0846_ net132 VPWR VGND sg13g2_buf_1
Xfanout143 net145 net143 VPWR VGND sg13g2_buf_1
Xfanout154 net155 net154 VPWR VGND sg13g2_buf_1
Xfanout165 net168 net165 VPWR VGND sg13g2_buf_1
XFILLER_27_230 VPWR VGND sg13g2_decap_8
XFILLER_27_296 VPWR VGND sg13g2_fill_2
XFILLER_47_539 VPWR VGND sg13g2_fill_1
XFILLER_47_56 VPWR VGND sg13g2_decap_8
Xfanout176 net177 net176 VPWR VGND sg13g2_buf_1
Xfanout187 net191 net187 VPWR VGND sg13g2_buf_1
Xfanout198 net199 net198 VPWR VGND sg13g2_buf_1
XFILLER_15_458 VPWR VGND sg13g2_decap_8
XFILLER_42_266 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_43_778 VPWR VGND sg13g2_decap_4
XFILLER_7_624 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_4
XFILLER_10_185 VPWR VGND sg13g2_decap_8
XFILLER_12_70 VPWR VGND sg13g2_decap_8
XFILLER_6_156 VPWR VGND sg13g2_decap_8
XFILLER_18_285 VPWR VGND sg13g2_decap_8
XFILLER_19_775 VPWR VGND sg13g2_fill_1
XFILLER_33_200 VPWR VGND sg13g2_decap_8
XFILLER_33_277 VPWR VGND sg13g2_decap_8
XFILLER_34_712 VPWR VGND sg13g2_fill_1
X_1963_ VGND VPWR net107 daisychain\[108\] _0644_ net53 sg13g2_a21oi_1
X_1894_ net189 VPWR _0589_ VGND daisychain\[95\] net32 sg13g2_o21ai_1
XFILLER_6_690 VPWR VGND sg13g2_fill_2
X_2515_ net243 VGND VPWR _0331_ state\[75\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2522__444 VPWR VGND net443 sg13g2_tiehi
X_2446_ net305 VGND VPWR _0262_ state\[6\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_24_211 VPWR VGND sg13g2_decap_8
X_1328_ VPWR _0110_ state\[84\] VGND sg13g2_inv_1
X_2377_ net454 VGND VPWR _0193_ daisychain\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_33_25 VPWR VGND sg13g2_decap_8
XFILLER_40_704 VPWR VGND sg13g2_decap_4
XFILLER_40_759 VPWR VGND sg13g2_fill_1
XFILLER_3_148 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_15_233 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_decap_8
X_2534__348 VPWR VGND net347 sg13g2_tiehi
XFILLER_30_214 VPWR VGND sg13g2_decap_8
XFILLER_7_432 VPWR VGND sg13g2_decap_8
X_2300_ _0840_ net90 state\[122\] VPWR VGND sg13g2_nand2_1
X_2231_ VGND VPWR _0555_ _0805_ _0343_ net77 sg13g2_a21oi_1
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_38_336 VPWR VGND sg13g2_decap_8
X_2162_ _0771_ net118 state\[53\] VPWR VGND sg13g2_nand2_1
X_2093_ VGND VPWR _0923_ _0736_ _0274_ net71 sg13g2_a21oi_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_21_247 VPWR VGND sg13g2_decap_8
XFILLER_34_597 VPWR VGND sg13g2_fill_2
X_1946_ state\[106\] daisychain\[106\] net142 _0630_ VPWR VGND sg13g2_mux2_1
X_1877_ _0575_ net174 _0574_ VPWR VGND sg13g2_nand2_1
XFILLER_28_25 VPWR VGND sg13g2_decap_8
X_2429_ net350 VGND VPWR _0245_ daisychain\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_12_203 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_8_229 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_4
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_4_479 VPWR VGND sg13g2_decap_8
XFILLER_0_641 VPWR VGND sg13g2_fill_1
XFILLER_0_652 VPWR VGND sg13g2_decap_4
XFILLER_0_674 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_31_545 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
X_1800_ VGND VPWR _0511_ _0512_ _0204_ _0513_ sg13g2_a21oi_1
X_1731_ state\[63\] daisychain\[63\] net150 _0458_ VPWR VGND sg13g2_mux2_1
X_1662_ _0403_ net172 _0402_ VPWR VGND sg13g2_nand2_1
X_2214_ _0797_ net127 state\[79\] VPWR VGND sg13g2_nand2_1
X_1593_ VGND VPWR net103 daisychain\[34\] _0992_ net57 sg13g2_a21oi_1
XFILLER_38_133 VPWR VGND sg13g2_decap_8
X_2145_ VGND VPWR _1027_ _0762_ _0300_ net80 sg13g2_a21oi_1
X_2076_ _0728_ net93 state\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_14_38 VPWR VGND sg13g2_fill_2
X_1929_ net189 VPWR _0617_ VGND daisychain\[102\] net32 sg13g2_o21ai_1
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_17_317 VPWR VGND sg13g2_decap_4
XFILLER_29_122 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_13_545 VPWR VGND sg13g2_fill_1
XFILLER_25_361 VPWR VGND sg13g2_fill_2
XFILLER_29_199 VPWR VGND sg13g2_decap_8
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_766 VPWR VGND sg13g2_fill_1
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_4_276 VPWR VGND sg13g2_decap_8
XFILLER_5_799 VPWR VGND sg13g2_fill_1
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_31_397 VPWR VGND sg13g2_decap_4
X_2832_ state\[120\] net7 VPWR VGND sg13g2_buf_1
XFILLER_6_72 VPWR VGND sg13g2_decap_8
X_1714_ net195 VPWR _0445_ VGND daisychain\[59\] net38 sg13g2_o21ai_1
X_1645_ VGND VPWR _0387_ _0388_ _0173_ _0389_ sg13g2_a21oi_1
X_1576_ state\[32\] daisychain\[32\] net140 _0978_ VPWR VGND sg13g2_mux2_1
XFILLER_25_48 VPWR VGND sg13g2_decap_8
XFILLER_26_169 VPWR VGND sg13g2_decap_8
XFILLER_34_180 VPWR VGND sg13g2_decap_8
XFILLER_35_670 VPWR VGND sg13g2_fill_2
XFILLER_35_681 VPWR VGND sg13g2_fill_2
X_2128_ _0754_ net116 state\[36\] VPWR VGND sg13g2_nand2_1
X_2059_ VGND VPWR _0855_ _0719_ _0257_ net67 sg13g2_a21oi_1
XFILLER_22_353 VPWR VGND sg13g2_fill_2
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
X_2344__265 VPWR VGND net264 sg13g2_tiehi
XFILLER_17_169 VPWR VGND sg13g2_decap_8
XFILLER_18_615 VPWR VGND sg13g2_decap_4
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_13_342 VPWR VGND sg13g2_decap_8
XFILLER_14_810 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_fill_2
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_357 VPWR VGND sg13g2_decap_8
X_1430_ VGND VPWR _0859_ _0860_ _0130_ _0861_ sg13g2_a21oi_1
X_1292_ VPWR _0023_ state\[120\] VGND sg13g2_inv_1
X_1361_ VPWR _0074_ state\[51\] VGND sg13g2_inv_1
XFILLER_23_117 VPWR VGND sg13g2_fill_2
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_31_172 VPWR VGND sg13g2_decap_8
XFILLER_8_390 VPWR VGND sg13g2_decap_8
X_2525__420 VPWR VGND net419 sg13g2_tiehi
X_2560__344 VPWR VGND net343 sg13g2_tiehi
X_1628_ VGND VPWR net115 daisychain\[41\] _1020_ net57 sg13g2_a21oi_1
X_1559_ net184 VPWR _0965_ VGND daisychain\[28\] net27 sg13g2_o21ai_1
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_14_128 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_10_367 VPWR VGND sg13g2_decap_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
XFILLER_6_338 VPWR VGND sg13g2_decap_8
XFILLER_2_555 VPWR VGND sg13g2_fill_1
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_46_710 VPWR VGND sg13g2_decap_4
XFILLER_18_434 VPWR VGND sg13g2_decap_4
XFILLER_18_467 VPWR VGND sg13g2_decap_4
XFILLER_18_478 VPWR VGND sg13g2_decap_4
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_46_776 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_decap_8
XFILLER_9_154 VPWR VGND sg13g2_decap_8
X_1413_ VPWR _0847_ net182 VGND sg13g2_inv_1
X_2531_ net371 VGND VPWR _0347_ state\[91\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2462_ net241 VGND VPWR _0278_ state\[22\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2393_ net422 VGND VPWR _0209_ daisychain\[81\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_36_231 VPWR VGND sg13g2_decap_8
X_1344_ VPWR _0092_ state\[68\] VGND sg13g2_inv_1
XFILLER_20_610 VPWR VGND sg13g2_fill_1
XFILLER_24_437 VPWR VGND sg13g2_fill_1
XFILLER_20_698 VPWR VGND sg13g2_fill_1
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
Xfanout100 net102 net100 VPWR VGND sg13g2_buf_1
Xfanout111 net112 net111 VPWR VGND sg13g2_buf_1
Xfanout122 net123 net122 VPWR VGND sg13g2_buf_1
Xfanout133 net134 net133 VPWR VGND sg13g2_buf_1
Xfanout144 net145 net144 VPWR VGND sg13g2_buf_1
Xfanout155 net156 net155 VPWR VGND sg13g2_buf_1
Xfanout166 net168 net166 VPWR VGND sg13g2_buf_1
Xfanout177 net178 net177 VPWR VGND sg13g2_buf_1
Xfanout188 net191 net188 VPWR VGND sg13g2_buf_1
Xfanout199 net200 net199 VPWR VGND sg13g2_buf_1
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_43_702 VPWR VGND sg13g2_decap_8
XFILLER_10_164 VPWR VGND sg13g2_decap_8
XFILLER_23_492 VPWR VGND sg13g2_decap_4
XFILLER_30_407 VPWR VGND sg13g2_decap_4
XFILLER_6_135 VPWR VGND sg13g2_decap_8
XFILLER_19_754 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_decap_8
XFILLER_14_481 VPWR VGND sg13g2_decap_8
XFILLER_18_264 VPWR VGND sg13g2_decap_8
XFILLER_19_787 VPWR VGND sg13g2_decap_4
XFILLER_21_418 VPWR VGND sg13g2_fill_1
XFILLER_33_256 VPWR VGND sg13g2_decap_8
XFILLER_46_562 VPWR VGND sg13g2_decap_8
X_1962_ _0643_ net168 _0642_ VPWR VGND sg13g2_nand2_1
X_1893_ VGND VPWR net111 daisychain\[94\] _0588_ net54 sg13g2_a21oi_1
XFILLER_29_507 VPWR VGND sg13g2_fill_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2514_ net251 VGND VPWR _0330_ state\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2445_ net309 VGND VPWR _0261_ state\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2376_ net456 VGND VPWR _0192_ daisychain\[64\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_17_38 VPWR VGND sg13g2_fill_1
X_1327_ VPWR _0111_ state\[85\] VGND sg13g2_inv_1
XFILLER_40_727 VPWR VGND sg13g2_fill_1
XFILLER_20_495 VPWR VGND sg13g2_decap_4
XFILLER_3_127 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_fill_2
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_15_212 VPWR VGND sg13g2_decap_8
XFILLER_15_289 VPWR VGND sg13g2_decap_8
XFILLER_11_462 VPWR VGND sg13g2_decap_8
XFILLER_7_411 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_decap_8
X_2402__405 VPWR VGND net404 sg13g2_tiehi
X_2230_ _0805_ net125 state\[87\] VPWR VGND sg13g2_nand2_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_19_573 VPWR VGND sg13g2_decap_8
XFILLER_34_510 VPWR VGND sg13g2_decap_4
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
X_2161_ VGND VPWR _0415_ _0770_ _0308_ net81 sg13g2_a21oi_1
X_2092_ _0736_ net99 state\[18\] VPWR VGND sg13g2_nand2_1
XFILLER_30_760 VPWR VGND sg13g2_fill_1
XFILLER_30_793 VPWR VGND sg13g2_fill_1
XFILLER_34_554 VPWR VGND sg13g2_decap_4
X_1945_ VGND VPWR _0627_ _0628_ _0233_ _0629_ sg13g2_a21oi_1
X_1876_ state\[92\] daisychain\[92\] net151 _0574_ VPWR VGND sg13g2_mux2_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_337 VPWR VGND sg13g2_decap_4
XFILLER_29_359 VPWR VGND sg13g2_decap_8
X_2428_ net352 VGND VPWR _0244_ daisychain\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2359_ net234 VGND VPWR _0175_ daisychain\[47\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_37_392 VPWR VGND sg13g2_fill_1
XFILLER_40_535 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_12_259 VPWR VGND sg13g2_decap_8
XFILLER_20_292 VPWR VGND sg13g2_decap_8
XFILLER_8_208 VPWR VGND sg13g2_decap_8
XFILLER_4_458 VPWR VGND sg13g2_decap_8
XFILLER_28_392 VPWR VGND sg13g2_decap_4
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_36_819 VPWR VGND sg13g2_decap_4
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
X_2458__258 VPWR VGND net257 sg13g2_tiehi
X_2354__245 VPWR VGND net244 sg13g2_tiehi
XFILLER_16_565 VPWR VGND sg13g2_fill_2
XFILLER_16_576 VPWR VGND sg13g2_fill_1
XFILLER_16_587 VPWR VGND sg13g2_decap_8
XFILLER_31_535 VPWR VGND sg13g2_fill_1
XFILLER_7_285 VPWR VGND sg13g2_decap_8
X_1730_ VGND VPWR _0455_ _0456_ _0190_ _0457_ sg13g2_a21oi_1
X_1661_ state\[49\] daisychain\[49\] net149 _0402_ VPWR VGND sg13g2_mux2_1
X_1592_ _0991_ net169 _0990_ VPWR VGND sg13g2_nand2_1
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_3_491 VPWR VGND sg13g2_decap_8
X_2213_ VGND VPWR _0519_ _0796_ _0334_ net87 sg13g2_a21oi_1
X_2144_ _0762_ net117 state\[44\] VPWR VGND sg13g2_nand2_1
XFILLER_34_395 VPWR VGND sg13g2_fill_1
XFILLER_38_189 VPWR VGND sg13g2_decap_8
X_2075_ VGND VPWR _0887_ _0727_ _0265_ net67 sg13g2_a21oi_1
XFILLER_10_708 VPWR VGND sg13g2_fill_2
X_1928_ VGND VPWR net110 daisychain\[101\] _0616_ net55 sg13g2_a21oi_1
X_1859_ net189 VPWR _0561_ VGND daisychain\[88\] net32 sg13g2_o21ai_1
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_29_101 VPWR VGND sg13g2_decap_8
XFILLER_29_178 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_25_340 VPWR VGND sg13g2_fill_1
XFILLER_25_373 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_4_255 VPWR VGND sg13g2_decap_8
XFILLER_5_701 VPWR VGND sg13g2_decap_8
XFILLER_5_734 VPWR VGND sg13g2_decap_4
XFILLER_5_778 VPWR VGND sg13g2_decap_4
XFILLER_5_789 VPWR VGND sg13g2_decap_4
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_20_82 VPWR VGND sg13g2_decap_8
XFILLER_29_80 VPWR VGND sg13g2_decap_8
XFILLER_16_340 VPWR VGND sg13g2_fill_2
XFILLER_16_362 VPWR VGND sg13g2_decap_8
XFILLER_16_373 VPWR VGND sg13g2_fill_1
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
X_1713_ VGND VPWR net119 daisychain\[58\] _0444_ net60 sg13g2_a21oi_1
X_1644_ net193 VPWR _0389_ VGND daisychain\[45\] net36 sg13g2_o21ai_1
X_1575_ VGND VPWR _0975_ _0976_ _0159_ _0977_ sg13g2_a21oi_1
XFILLER_39_421 VPWR VGND sg13g2_decap_4
X_2127_ VGND VPWR _0991_ _0753_ _0291_ net80 sg13g2_a21oi_1
XFILLER_26_148 VPWR VGND sg13g2_decap_8
X_2058_ _0719_ net94 state\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_17_148 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_13_321 VPWR VGND sg13g2_decap_8
XFILLER_15_93 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_9_336 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_decap_8
XFILLER_5_520 VPWR VGND sg13g2_decap_8
X_1360_ VPWR _0075_ state\[52\] VGND sg13g2_inv_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_36_402 VPWR VGND sg13g2_fill_2
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_49_752 VPWR VGND sg13g2_decap_8
X_1291_ VPWR _0024_ state\[121\] VGND sg13g2_inv_1
XFILLER_16_181 VPWR VGND sg13g2_decap_8
XFILLER_17_693 VPWR VGND sg13g2_fill_1
XFILLER_31_151 VPWR VGND sg13g2_decap_8
XFILLER_36_479 VPWR VGND sg13g2_decap_8
X_2410__389 VPWR VGND net388 sg13g2_tiehi
X_1489_ net180 VPWR _0909_ VGND daisychain\[14\] net23 sg13g2_o21ai_1
X_1558_ VGND VPWR net100 daisychain\[27\] _0964_ net52 sg13g2_a21oi_1
X_1627_ _1019_ net169 _1018_ VPWR VGND sg13g2_nand2_1
XFILLER_14_107 VPWR VGND sg13g2_decap_8
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_42_427 VPWR VGND sg13g2_decap_8
XFILLER_10_346 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_42_449 VPWR VGND sg13g2_fill_1
XFILLER_6_317 VPWR VGND sg13g2_decap_8
XFILLER_2_567 VPWR VGND sg13g2_fill_2
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_26_92 VPWR VGND sg13g2_decap_8
XFILLER_33_427 VPWR VGND sg13g2_decap_4
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_13_195 VPWR VGND sg13g2_decap_8
XFILLER_42_91 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_8
X_2530_ net379 VGND VPWR _0346_ state\[90\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1343_ VPWR _0093_ state\[69\] VGND sg13g2_inv_1
X_1412_ VPWR _0000_ state\[0\] VGND sg13g2_inv_1
X_2461_ net245 VGND VPWR _0277_ state\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2392_ net424 VGND VPWR _0208_ daisychain\[80\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_37_744 VPWR VGND sg13g2_decap_8
XFILLER_3_85 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_49_582 VPWR VGND sg13g2_fill_2
XFILLER_20_622 VPWR VGND sg13g2_fill_1
XFILLER_22_39 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_2_0__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_20_677 VPWR VGND sg13g2_fill_1
XFILLER_3_309 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
Xfanout101 net102 net101 VPWR VGND sg13g2_buf_1
Xfanout112 net113 net112 VPWR VGND sg13g2_buf_1
Xfanout123 net132 net123 VPWR VGND sg13g2_buf_1
Xfanout134 net136 net134 VPWR VGND sg13g2_buf_1
Xfanout145 net156 net145 VPWR VGND sg13g2_buf_1
Xfanout156 net5 net156 VPWR VGND sg13g2_buf_1
Xfanout167 net168 net167 VPWR VGND sg13g2_buf_1
Xfanout178 net4 net178 VPWR VGND sg13g2_buf_1
Xfanout189 net191 net189 VPWR VGND sg13g2_buf_1
XFILLER_27_298 VPWR VGND sg13g2_fill_1
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_43_725 VPWR VGND sg13g2_decap_8
X_2313__327 VPWR VGND net326 sg13g2_tiehi
XFILLER_10_143 VPWR VGND sg13g2_decap_8
XFILLER_11_677 VPWR VGND sg13g2_decap_8
XFILLER_11_688 VPWR VGND sg13g2_fill_2
XFILLER_23_460 VPWR VGND sg13g2_decap_8
XFILLER_6_114 VPWR VGND sg13g2_decap_8
XFILLER_7_615 VPWR VGND sg13g2_decap_4
XFILLER_7_637 VPWR VGND sg13g2_decap_8
XFILLER_2_364 VPWR VGND sg13g2_decap_8
XFILLER_18_243 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_33_235 VPWR VGND sg13g2_decap_8
X_1961_ state\[109\] daisychain\[109\] net142 _0642_ VPWR VGND sg13g2_mux2_1
X_1892_ _0587_ net166 _0586_ VPWR VGND sg13g2_nand2_1
XFILLER_6_692 VPWR VGND sg13g2_fill_1
X_2513_ net259 VGND VPWR _0329_ state\[73\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2409__391 VPWR VGND net390 sg13g2_tiehi
X_2364__225 VPWR VGND net224 sg13g2_tiehi
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_1326_ VPWR _0112_ state\[86\] VGND sg13g2_inv_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2444_ net313 VGND VPWR _0260_ state\[4\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2375_ net202 VGND VPWR _0191_ daisychain\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2451__286 VPWR VGND net285 sg13g2_tiehi
XFILLER_3_106 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_15_268 VPWR VGND sg13g2_decap_8
XFILLER_16_736 VPWR VGND sg13g2_decap_4
XFILLER_23_290 VPWR VGND sg13g2_fill_2
XFILLER_30_249 VPWR VGND sg13g2_decap_8
XFILLER_7_467 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
X_2160_ _0770_ net121 state\[52\] VPWR VGND sg13g2_nand2_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
X_2091_ VGND VPWR _0919_ _0735_ _0273_ net71 sg13g2_a21oi_1
XFILLER_21_227 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_fill_1
XFILLER_34_599 VPWR VGND sg13g2_fill_1
XFILLER_9_84 VPWR VGND sg13g2_decap_8
X_1944_ net187 VPWR _0629_ VGND daisychain\[105\] net30 sg13g2_o21ai_1
X_1875_ VGND VPWR _0571_ _0572_ _0219_ _0573_ sg13g2_a21oi_1
X_2427_ net354 VGND VPWR _0243_ daisychain\[115\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_44_308 VPWR VGND sg13g2_decap_8
X_1309_ VPWR _0004_ state\[103\] VGND sg13g2_inv_1
X_2358_ net236 VGND VPWR _0174_ daisychain\[46\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2289_ VGND VPWR _0671_ _0834_ _0372_ net69 sg13g2_a21oi_1
XFILLER_12_238 VPWR VGND sg13g2_decap_8
XFILLER_25_533 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_20_271 VPWR VGND sg13g2_decap_8
XFILLER_4_437 VPWR VGND sg13g2_decap_8
XFILLER_48_625 VPWR VGND sg13g2_decap_4
XFILLER_16_533 VPWR VGND sg13g2_fill_1
XFILLER_16_544 VPWR VGND sg13g2_decap_8
XFILLER_18_82 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_31_503 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_8_765 VPWR VGND sg13g2_decap_8
XFILLER_3_470 VPWR VGND sg13g2_decap_8
XFILLER_7_264 VPWR VGND sg13g2_decap_8
XFILLER_8_798 VPWR VGND sg13g2_fill_1
X_1660_ VGND VPWR _0399_ _0400_ _0176_ _0401_ sg13g2_a21oi_1
X_1591_ state\[35\] daisychain\[35\] net146 _0990_ VPWR VGND sg13g2_mux2_1
XFILLER_26_308 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_decap_8
X_2212_ _0796_ net127 state\[78\] VPWR VGND sg13g2_nand2_1
X_2143_ VGND VPWR _1023_ _0761_ _0299_ net80 sg13g2_a21oi_1
XFILLER_47_680 VPWR VGND sg13g2_decap_4
XFILLER_47_691 VPWR VGND sg13g2_fill_2
X_2074_ _0727_ net101 state\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_30_39 VPWR VGND sg13g2_decap_8
X_1927_ _0615_ net166 _0614_ VPWR VGND sg13g2_nand2_1
X_1858_ VGND VPWR net111 daisychain\[87\] _0560_ net54 sg13g2_a21oi_1
X_2420__369 VPWR VGND net368 sg13g2_tiehi
X_1789_ net196 VPWR _0505_ VGND daisychain\[74\] net39 sg13g2_o21ai_1
XFILLER_25_352 VPWR VGND sg13g2_decap_4
XFILLER_29_157 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_45_606 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_4
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_4_234 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_31_333 VPWR VGND sg13g2_fill_1
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_8_562 VPWR VGND sg13g2_fill_2
XFILLER_8_573 VPWR VGND sg13g2_decap_8
XFILLER_8_584 VPWR VGND sg13g2_fill_2
X_1712_ _0443_ net172 _0442_ VPWR VGND sg13g2_nand2_1
X_1643_ VGND VPWR net116 daisychain\[44\] _0388_ net58 sg13g2_a21oi_1
X_1574_ net186 VPWR _0977_ VGND daisychain\[31\] net29 sg13g2_o21ai_1
XFILLER_19_190 VPWR VGND sg13g2_decap_8
XFILLER_26_127 VPWR VGND sg13g2_decap_8
XFILLER_35_650 VPWR VGND sg13g2_decap_8
X_2126_ _0753_ net116 state\[35\] VPWR VGND sg13g2_nand2_1
X_2057_ VGND VPWR _0849_ _0718_ _0256_ net67 sg13g2_a21oi_1
XFILLER_10_528 VPWR VGND sg13g2_decap_8
XFILLER_22_344 VPWR VGND sg13g2_decap_4
XFILLER_22_355 VPWR VGND sg13g2_fill_1
XFILLER_22_399 VPWR VGND sg13g2_decap_4
XFILLER_25_39 VPWR VGND sg13g2_fill_2
XFILLER_35_694 VPWR VGND sg13g2_fill_1
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_13_300 VPWR VGND sg13g2_decap_8
XFILLER_17_127 VPWR VGND sg13g2_decap_8
XFILLER_25_193 VPWR VGND sg13g2_decap_8
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_13_388 VPWR VGND sg13g2_decap_4
XFILLER_15_72 VPWR VGND sg13g2_decap_8
XFILLER_31_60 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_41_675 VPWR VGND sg13g2_fill_2
XFILLER_9_315 VPWR VGND sg13g2_decap_8
X_2323__307 VPWR VGND net306 sg13g2_tiehi
XFILLER_48_252 VPWR VGND sg13g2_decap_8
X_1290_ VPWR _0025_ state\[122\] VGND sg13g2_inv_1
XFILLER_16_160 VPWR VGND sg13g2_decap_8
XFILLER_20_804 VPWR VGND sg13g2_fill_1
XFILLER_31_130 VPWR VGND sg13g2_decap_8
XFILLER_32_620 VPWR VGND sg13g2_fill_1
X_1626_ state\[42\] daisychain\[42\] net146 _1018_ VPWR VGND sg13g2_mux2_1
XFILLER_39_252 VPWR VGND sg13g2_decap_8
X_1488_ VGND VPWR net93 daisychain\[13\] _0908_ net45 sg13g2_a21oi_1
X_1557_ _0963_ net162 _0962_ VPWR VGND sg13g2_nand2_1
X_2374__205 VPWR VGND net204 sg13g2_tiehi
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
X_2419__371 VPWR VGND net370 sg13g2_tiehi
X_2109_ VGND VPWR _0955_ _0744_ _0282_ net72 sg13g2_a21oi_1
XFILLER_10_325 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_2_546 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_decap_8
XFILLER_18_447 VPWR VGND sg13g2_decap_8
XFILLER_13_174 VPWR VGND sg13g2_decap_8
XFILLER_14_642 VPWR VGND sg13g2_decap_4
XFILLER_26_71 VPWR VGND sg13g2_decap_8
XFILLER_41_472 VPWR VGND sg13g2_fill_1
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
X_2548__400 VPWR VGND net399 sg13g2_tiehi
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_decap_8
X_2460_ net249 VGND VPWR _0276_ state\[20\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_3_64 VPWR VGND sg13g2_decap_8
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_5_384 VPWR VGND sg13g2_decap_8
X_1342_ VPWR _0095_ state\[70\] VGND sg13g2_inv_1
X_1411_ VPWR _0039_ state\[1\] VGND sg13g2_inv_1
X_2391_ net426 VGND VPWR _0207_ daisychain\[79\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_20_656 VPWR VGND sg13g2_fill_1
XFILLER_20_689 VPWR VGND sg13g2_fill_2
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_9_690 VPWR VGND sg13g2_decap_8
Xfanout102 net106 net102 VPWR VGND sg13g2_buf_1
Xfanout113 net114 net113 VPWR VGND sg13g2_buf_1
X_1609_ net185 VPWR _1005_ VGND daisychain\[38\] net28 sg13g2_o21ai_1
XFILLER_27_244 VPWR VGND sg13g2_decap_8
Xfanout124 net125 net124 VPWR VGND sg13g2_buf_1
Xfanout135 net156 net135 VPWR VGND sg13g2_buf_1
Xfanout146 net150 net146 VPWR VGND sg13g2_buf_1
Xfanout157 net160 net157 VPWR VGND sg13g2_buf_1
Xfanout168 net178 net168 VPWR VGND sg13g2_buf_1
Xfanout179 net182 net179 VPWR VGND sg13g2_buf_1
XFILLER_15_428 VPWR VGND sg13g2_fill_2
XFILLER_15_439 VPWR VGND sg13g2_fill_1
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_10_122 VPWR VGND sg13g2_decap_8
XFILLER_10_199 VPWR VGND sg13g2_decap_8
XFILLER_12_84 VPWR VGND sg13g2_decap_8
XFILLER_2_343 VPWR VGND sg13g2_decap_8
XFILLER_18_222 VPWR VGND sg13g2_decap_8
XFILLER_18_299 VPWR VGND sg13g2_decap_8
XFILLER_33_214 VPWR VGND sg13g2_decap_8
XFILLER_34_748 VPWR VGND sg13g2_decap_4
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_46_597 VPWR VGND sg13g2_decap_4
XFILLER_21_409 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
X_1960_ VGND VPWR _0639_ _0640_ _0236_ _0641_ sg13g2_a21oi_1
X_1891_ state\[95\] daisychain\[95\] net144 _0586_ VPWR VGND sg13g2_mux2_1
XFILLER_5_181 VPWR VGND sg13g2_decap_8
X_2512_ net267 VGND VPWR _0328_ state\[72\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2443_ net317 VGND VPWR _0259_ state\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1325_ VPWR _0113_ state\[87\] VGND sg13g2_inv_1
X_2374_ net204 VGND VPWR _0190_ daisychain\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_33_39 VPWR VGND sg13g2_decap_8
XFILLER_33_781 VPWR VGND sg13g2_decap_8
XFILLER_33_792 VPWR VGND sg13g2_fill_2
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_16_704 VPWR VGND sg13g2_fill_2
XFILLER_43_501 VPWR VGND sg13g2_fill_1
XFILLER_15_247 VPWR VGND sg13g2_decap_8
XFILLER_30_228 VPWR VGND sg13g2_decap_8
XFILLER_31_718 VPWR VGND sg13g2_decap_8
XFILLER_31_729 VPWR VGND sg13g2_fill_1
X_2430__349 VPWR VGND net348 sg13g2_tiehi
XFILLER_11_497 VPWR VGND sg13g2_decap_8
XFILLER_23_83 VPWR VGND sg13g2_decap_8
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_7_446 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
X_2090_ _0735_ net99 state\[17\] VPWR VGND sg13g2_nand2_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_21_206 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_458 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_30_751 VPWR VGND sg13g2_fill_1
XFILLER_30_784 VPWR VGND sg13g2_fill_2
X_1943_ VGND VPWR net107 daisychain\[104\] _0628_ net53 sg13g2_a21oi_1
X_1874_ net197 VPWR _0573_ VGND daisychain\[91\] net40 sg13g2_o21ai_1
XFILLER_6_490 VPWR VGND sg13g2_decap_4
X_2426_ net356 VGND VPWR _0242_ daisychain\[114\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_25_501 VPWR VGND sg13g2_decap_4
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
X_1308_ VPWR _0005_ state\[104\] VGND sg13g2_inv_1
X_2357_ net238 VGND VPWR _0173_ daisychain\[45\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2288_ _0834_ net96 state\[116\] VPWR VGND sg13g2_nand2_1
XFILLER_12_217 VPWR VGND sg13g2_decap_8
XFILLER_20_250 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_4_416 VPWR VGND sg13g2_decap_8
XFILLER_18_61 VPWR VGND sg13g2_decap_8
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_11_283 VPWR VGND sg13g2_decap_8
XFILLER_31_559 VPWR VGND sg13g2_decap_4
XFILLER_34_82 VPWR VGND sg13g2_decap_8
XFILLER_7_243 VPWR VGND sg13g2_decap_8
XFILLER_8_744 VPWR VGND sg13g2_fill_2
X_1590_ VGND VPWR _0987_ _0988_ _0162_ _0989_ sg13g2_a21oi_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_decap_8
XFILLER_39_648 VPWR VGND sg13g2_fill_2
X_2211_ VGND VPWR _0515_ _0795_ _0333_ net86 sg13g2_a21oi_1
X_2142_ _0761_ net115 state\[43\] VPWR VGND sg13g2_nand2_1
X_2073_ VGND VPWR _0883_ _0726_ _0264_ net71 sg13g2_a21oi_1
XFILLER_34_320 VPWR VGND sg13g2_decap_8
XFILLER_34_353 VPWR VGND sg13g2_decap_8
XFILLER_30_18 VPWR VGND sg13g2_decap_8
X_2383__443 VPWR VGND net442 sg13g2_tiehi
X_1926_ state\[102\] daisychain\[102\] net143 _0614_ VPWR VGND sg13g2_mux2_1
X_1857_ _0559_ net166 _0558_ VPWR VGND sg13g2_nand2_1
X_1788_ VGND VPWR net125 daisychain\[73\] _0504_ net62 sg13g2_a21oi_1
XFILLER_29_136 VPWR VGND sg13g2_decap_8
XFILLER_39_49 VPWR VGND sg13g2_decap_8
X_2409_ net390 VGND VPWR _0225_ daisychain\[97\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_17_309 VPWR VGND sg13g2_decap_4
XFILLER_38_670 VPWR VGND sg13g2_fill_1
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_40_378 VPWR VGND sg13g2_decap_8
X_2429__351 VPWR VGND net350 sg13g2_tiehi
XFILLER_4_213 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_16_342 VPWR VGND sg13g2_fill_1
XFILLER_31_312 VPWR VGND sg13g2_decap_8
XFILLER_31_356 VPWR VGND sg13g2_fill_1
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
X_1711_ state\[59\] daisychain\[59\] net149 _0442_ VPWR VGND sg13g2_mux2_1
X_1642_ _0387_ net170 _0386_ VPWR VGND sg13g2_nand2_1
XFILLER_6_86 VPWR VGND sg13g2_decap_8
X_1573_ VGND VPWR net105 daisychain\[30\] _0976_ net51 sg13g2_a21oi_1
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_26_106 VPWR VGND sg13g2_decap_8
XFILLER_39_478 VPWR VGND sg13g2_fill_2
X_2125_ VGND VPWR _0987_ _0752_ _0290_ net73 sg13g2_a21oi_1
X_2056_ _0718_ net94 state\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_10_518 VPWR VGND sg13g2_decap_4
XFILLER_22_367 VPWR VGND sg13g2_decap_4
XFILLER_34_194 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
X_1909_ net188 VPWR _0601_ VGND daisychain\[98\] net31 sg13g2_o21ai_1
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_17_106 VPWR VGND sg13g2_decap_8
XFILLER_13_356 VPWR VGND sg13g2_decap_8
XFILLER_25_172 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_41_621 VPWR VGND sg13g2_fill_1
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_555 VPWR VGND sg13g2_decap_8
XFILLER_36_459 VPWR VGND sg13g2_fill_2
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_31_186 VPWR VGND sg13g2_decap_8
XFILLER_32_687 VPWR VGND sg13g2_decap_4
X_1556_ state\[28\] daisychain\[28\] net138 _0962_ VPWR VGND sg13g2_mux2_1
X_1625_ VGND VPWR _1015_ _1016_ _0169_ _1017_ sg13g2_a21oi_1
XFILLER_27_415 VPWR VGND sg13g2_decap_8
XFILLER_27_426 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_39_231 VPWR VGND sg13g2_decap_8
X_1487_ _0907_ net159 _0906_ VPWR VGND sg13g2_nand2_1
XFILLER_11_805 VPWR VGND sg13g2_decap_8
X_2454__274 VPWR VGND net273 sg13g2_tiehi
X_2108_ _0744_ net100 state\[26\] VPWR VGND sg13g2_nand2_1
X_2039_ net179 VPWR _0705_ VGND daisychain\[124\] net25 sg13g2_o21ai_1
XFILLER_10_304 VPWR VGND sg13g2_decap_8
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_2_525 VPWR VGND sg13g2_decap_8
XFILLER_18_415 VPWR VGND sg13g2_decap_8
XFILLER_26_50 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_46_724 VPWR VGND sg13g2_decap_8
XFILLER_13_153 VPWR VGND sg13g2_decap_8
XFILLER_14_698 VPWR VGND sg13g2_decap_8
XFILLER_26_481 VPWR VGND sg13g2_decap_8
XFILLER_5_363 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
X_1410_ VPWR _0050_ state\[2\] VGND sg13g2_inv_1
X_2440__329 VPWR VGND net328 sg13g2_tiehi
X_1341_ VPWR _0096_ state\[71\] VGND sg13g2_inv_1
X_2390_ net428 VGND VPWR _0206_ daisychain\[78\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_37_735 VPWR VGND sg13g2_fill_1
XFILLER_49_595 VPWR VGND sg13g2_decap_4
XFILLER_20_668 VPWR VGND sg13g2_fill_2
X_1539_ net185 VPWR _0949_ VGND daisychain\[24\] net28 sg13g2_o21ai_1
Xfanout103 net104 net103 VPWR VGND sg13g2_buf_1
Xfanout114 net132 net114 VPWR VGND sg13g2_buf_1
Xfanout125 net126 net125 VPWR VGND sg13g2_buf_1
Xfanout136 net156 net136 VPWR VGND sg13g2_buf_1
Xfanout147 net150 net147 VPWR VGND sg13g2_buf_1
X_1608_ VGND VPWR net103 daisychain\[37\] _1004_ net50 sg13g2_a21oi_1
XFILLER_27_223 VPWR VGND sg13g2_decap_8
XFILLER_43_716 VPWR VGND sg13g2_decap_4
XFILLER_47_49 VPWR VGND sg13g2_decap_8
Xfanout158 net159 net158 VPWR VGND sg13g2_buf_1
Xfanout169 net170 net169 VPWR VGND sg13g2_buf_1
XFILLER_10_101 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_10_178 VPWR VGND sg13g2_decap_8
XFILLER_2_322 VPWR VGND sg13g2_decap_8
XFILLER_6_149 VPWR VGND sg13g2_decap_8
XFILLER_18_201 VPWR VGND sg13g2_decap_8
XFILLER_19_713 VPWR VGND sg13g2_decap_4
XFILLER_2_399 VPWR VGND sg13g2_decap_8
XFILLER_18_278 VPWR VGND sg13g2_decap_8
XFILLER_19_768 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_fill_2
X_2550__368 VPWR VGND net367 sg13g2_tiehi
X_2468__218 VPWR VGND net217 sg13g2_tiehi
X_1890_ VGND VPWR _0583_ _0584_ _0222_ _0585_ sg13g2_a21oi_1
XFILLER_5_160 VPWR VGND sg13g2_decap_8
XFILLER_6_683 VPWR VGND sg13g2_fill_2
X_2511_ net275 VGND VPWR _0327_ state\[71\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2442_ net321 VGND VPWR _0258_ state\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2373_ net206 VGND VPWR _0189_ daisychain\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1324_ VPWR _0114_ state\[88\] VGND sg13g2_inv_1
XFILLER_24_204 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_33_760 VPWR VGND sg13g2_decap_4
XFILLER_40_708 VPWR VGND sg13g2_fill_1
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_15_226 VPWR VGND sg13g2_decap_8
XFILLER_16_727 VPWR VGND sg13g2_decap_4
X_2393__423 VPWR VGND net422 sg13g2_tiehi
XFILLER_23_62 VPWR VGND sg13g2_decap_8
XFILLER_30_207 VPWR VGND sg13g2_decap_8
XFILLER_43_579 VPWR VGND sg13g2_decap_8
XFILLER_7_425 VPWR VGND sg13g2_decap_8
X_2545__448 VPWR VGND net447 sg13g2_tiehi
XFILLER_3_642 VPWR VGND sg13g2_decap_8
XFILLER_3_675 VPWR VGND sg13g2_decap_8
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
X_2439__331 VPWR VGND net330 sg13g2_tiehi
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_15_793 VPWR VGND sg13g2_fill_1
XFILLER_19_587 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_459 VPWR VGND uio_oe[2] sg13g2_tiehi
X_1942_ _0627_ net165 _0626_ VPWR VGND sg13g2_nand2_1
XFILLER_6_480 VPWR VGND sg13g2_decap_4
X_1873_ VGND VPWR net124 daisychain\[90\] _0572_ net64 sg13g2_a21oi_1
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_2425_ net358 VGND VPWR _0241_ daisychain\[113\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2356_ net240 VGND VPWR _0172_ daisychain\[44\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_25_513 VPWR VGND sg13g2_fill_2
XFILLER_44_28 VPWR VGND sg13g2_decap_8
X_1307_ VPWR _0006_ state\[105\] VGND sg13g2_inv_1
X_2287_ VGND VPWR _0667_ _0833_ _0371_ net69 sg13g2_a21oi_1
XFILLER_33_590 VPWR VGND sg13g2_fill_2
XFILLER_0_601 VPWR VGND sg13g2_fill_2
XFILLER_0_634 VPWR VGND sg13g2_fill_2
XFILLER_18_40 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_28_362 VPWR VGND sg13g2_fill_2
XFILLER_34_61 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_11_262 VPWR VGND sg13g2_decap_8
XFILLER_7_222 VPWR VGND sg13g2_decap_8
XFILLER_7_299 VPWR VGND sg13g2_decap_8
XFILLER_8_789 VPWR VGND sg13g2_decap_4
X_2210_ _0795_ net128 state\[77\] VPWR VGND sg13g2_nand2_1
XFILLER_15_4 VPWR VGND sg13g2_fill_1
XFILLER_19_340 VPWR VGND sg13g2_fill_1
XFILLER_19_351 VPWR VGND sg13g2_decap_4
XFILLER_19_362 VPWR VGND sg13g2_fill_1
XFILLER_38_126 VPWR VGND sg13g2_decap_8
X_2141_ VGND VPWR _1019_ _0760_ _0298_ net80 sg13g2_a21oi_1
X_2072_ _0726_ net101 state\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_22_505 VPWR VGND sg13g2_fill_2
XFILLER_30_571 VPWR VGND sg13g2_fill_2
X_1925_ VGND VPWR _0611_ _0612_ _0229_ _0613_ sg13g2_a21oi_1
XFILLER_30_593 VPWR VGND sg13g2_fill_1
X_1856_ state\[88\] daisychain\[88\] net143 _0558_ VPWR VGND sg13g2_mux2_1
X_1787_ _0503_ net173 _0502_ VPWR VGND sg13g2_nand2_1
XFILLER_29_115 VPWR VGND sg13g2_decap_8
XFILLER_39_28 VPWR VGND sg13g2_decap_8
X_2408_ net392 VGND VPWR _0224_ daisychain\[96\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2339_ net274 VGND VPWR _0155_ daisychain\[27\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_25_310 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_20_96 VPWR VGND sg13g2_decap_8
XFILLER_4_269 VPWR VGND sg13g2_decap_8
XFILLER_5_759 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_16_321 VPWR VGND sg13g2_decap_8
XFILLER_17_822 VPWR VGND sg13g2_fill_1
XFILLER_29_94 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_12_571 VPWR VGND sg13g2_decap_8
XFILLER_16_354 VPWR VGND sg13g2_fill_2
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_4_770 VPWR VGND sg13g2_decap_4
XFILLER_8_542 VPWR VGND sg13g2_fill_1
XFILLER_8_553 VPWR VGND sg13g2_decap_4
XFILLER_8_564 VPWR VGND sg13g2_fill_1
X_1710_ VGND VPWR _0439_ _0440_ _0186_ _0441_ sg13g2_a21oi_1
X_1641_ state\[45\] daisychain\[45\] net147 _0386_ VPWR VGND sg13g2_mux2_1
X_1572_ _0975_ net164 _0974_ VPWR VGND sg13g2_nand2_1
XFILLER_39_413 VPWR VGND sg13g2_decap_4
X_2124_ _0752_ net116 state\[34\] VPWR VGND sg13g2_nand2_1
XFILLER_34_173 VPWR VGND sg13g2_decap_8
XFILLER_35_663 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
X_2055_ VGND VPWR _0715_ _0716_ _0255_ _0717_ sg13g2_a21oi_1
X_1908_ VGND VPWR net109 daisychain\[97\] _0600_ net54 sg13g2_a21oi_1
X_1839_ net197 VPWR _0545_ VGND daisychain\[84\] net40 sg13g2_o21ai_1
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_18_608 VPWR VGND sg13g2_decap_8
XFILLER_18_619 VPWR VGND sg13g2_fill_1
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_13_335 VPWR VGND sg13g2_decap_8
XFILLER_14_803 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_41_677 VPWR VGND sg13g2_fill_1
XFILLER_31_95 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_fill_2
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_4
XFILLER_16_195 VPWR VGND sg13g2_decap_8
XFILLER_31_165 VPWR VGND sg13g2_decap_8
XFILLER_8_383 VPWR VGND sg13g2_decap_8
X_1555_ VGND VPWR _0959_ _0960_ _0155_ _0961_ sg13g2_a21oi_1
X_1624_ net192 VPWR _1017_ VGND daisychain\[41\] net35 sg13g2_o21ai_1
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
X_1486_ state\[14\] daisychain\[14\] net134 _0906_ VPWR VGND sg13g2_mux2_1
X_2107_ VGND VPWR _0951_ _0743_ _0281_ net72 sg13g2_a21oi_1
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_35_493 VPWR VGND sg13g2_decap_8
X_2038_ VGND VPWR net90 daisychain\[123\] _0704_ net48 sg13g2_a21oi_1
XFILLER_2_504 VPWR VGND sg13g2_decap_8
X_2461__246 VPWR VGND net245 sg13g2_tiehi
XFILLER_18_427 VPWR VGND sg13g2_decap_8
XFILLER_33_419 VPWR VGND sg13g2_fill_2
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_46_703 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_fill_1
XFILLER_46_747 VPWR VGND sg13g2_decap_4
XFILLER_46_769 VPWR VGND sg13g2_decap_8
XFILLER_13_132 VPWR VGND sg13g2_decap_8
XFILLER_14_677 VPWR VGND sg13g2_decap_8
XFILLER_9_147 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_342 VPWR VGND sg13g2_decap_8
X_1340_ VPWR _0097_ state\[72\] VGND sg13g2_inv_1
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_3_99 VPWR VGND sg13g2_decap_8
XFILLER_20_614 VPWR VGND sg13g2_fill_1
XFILLER_8_180 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_8_clk clknet_2_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
X_1469_ net180 VPWR _0893_ VGND daisychain\[10\] net23 sg13g2_o21ai_1
X_1538_ VGND VPWR net104 daisychain\[23\] _0948_ net50 sg13g2_a21oi_1
Xfanout104 net106 net104 VPWR VGND sg13g2_buf_1
Xfanout115 net116 net115 VPWR VGND sg13g2_buf_1
Xfanout126 net131 net126 VPWR VGND sg13g2_buf_1
Xfanout137 net141 net137 VPWR VGND sg13g2_buf_1
Xfanout148 net149 net148 VPWR VGND sg13g2_buf_1
Xfanout159 net160 net159 VPWR VGND sg13g2_buf_1
X_1607_ _1003_ net163 _1002_ VPWR VGND sg13g2_nand2_1
XFILLER_27_202 VPWR VGND sg13g2_decap_8
XFILLER_36_791 VPWR VGND sg13g2_fill_1
XFILLER_10_157 VPWR VGND sg13g2_decap_8
XFILLER_23_474 VPWR VGND sg13g2_decap_4
XFILLER_23_485 VPWR VGND sg13g2_fill_2
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_2_301 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_6_128 VPWR VGND sg13g2_decap_8
XFILLER_19_747 VPWR VGND sg13g2_fill_2
XFILLER_2_378 VPWR VGND sg13g2_decap_8
XFILLER_14_474 VPWR VGND sg13g2_decap_8
XFILLER_18_257 VPWR VGND sg13g2_decap_8
XFILLER_33_249 VPWR VGND sg13g2_decap_8
X_2510_ net283 VGND VPWR _0326_ state\[70\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_1323_ VPWR _0115_ state\[89\] VGND sg13g2_inv_1
X_2441_ net325 VGND VPWR _0257_ state\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2372_ net208 VGND VPWR _0188_ daisychain\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_37_577 VPWR VGND sg13g2_fill_2
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_20_477 VPWR VGND sg13g2_fill_2
XFILLER_20_488 VPWR VGND sg13g2_decap_8
XFILLER_20_499 VPWR VGND sg13g2_fill_1
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_15_205 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_fill_1
XFILLER_16_717 VPWR VGND sg13g2_fill_2
XFILLER_43_525 VPWR VGND sg13g2_decap_4
XFILLER_11_422 VPWR VGND sg13g2_fill_2
XFILLER_11_444 VPWR VGND sg13g2_decap_8
XFILLER_11_455 VPWR VGND sg13g2_fill_2
XFILLER_23_271 VPWR VGND sg13g2_fill_1
XFILLER_23_41 VPWR VGND sg13g2_decap_8
XFILLER_7_404 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_3_698 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_544 VPWR VGND sg13g2_fill_2
XFILLER_34_514 VPWR VGND sg13g2_fill_1
XFILLER_34_525 VPWR VGND sg13g2_fill_1
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
X_2554__280 VPWR VGND net279 sg13g2_tiehi
XFILLER_14_282 VPWR VGND sg13g2_decap_8
XFILLER_15_761 VPWR VGND sg13g2_decap_4
XFILLER_30_731 VPWR VGND sg13g2_fill_1
XFILLER_30_764 VPWR VGND sg13g2_fill_1
XFILLER_34_547 VPWR VGND sg13g2_fill_2
X_1941_ state\[105\] daisychain\[105\] net142 _0626_ VPWR VGND sg13g2_mux2_1
X_1872_ _0571_ net174 _0570_ VPWR VGND sg13g2_nand2_1
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_38_820 VPWR VGND sg13g2_fill_2
X_1306_ VPWR _0007_ state\[106\] VGND sg13g2_inv_1
X_2424_ net360 VGND VPWR _0240_ daisychain\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2355_ net242 VGND VPWR _0171_ daisychain\[43\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2286_ _0833_ net96 state\[115\] VPWR VGND sg13g2_nand2_1
XFILLER_37_385 VPWR VGND sg13g2_decap_8
X_2492__378 VPWR VGND net377 sg13g2_tiehi
XFILLER_20_285 VPWR VGND sg13g2_decap_8
XFILLER_16_503 VPWR VGND sg13g2_fill_2
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_11_241 VPWR VGND sg13g2_decap_8
XFILLER_16_558 VPWR VGND sg13g2_fill_2
XFILLER_18_96 VPWR VGND sg13g2_decap_8
XFILLER_34_40 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_8_713 VPWR VGND sg13g2_fill_1
XFILLER_7_201 VPWR VGND sg13g2_decap_8
XFILLER_7_278 VPWR VGND sg13g2_decap_8
XFILLER_8_746 VPWR VGND sg13g2_fill_1
X_2330__293 VPWR VGND net292 sg13g2_tiehi
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_3_484 VPWR VGND sg13g2_decap_8
X_2406__397 VPWR VGND net396 sg13g2_tiehi
X_2140_ _0760_ net115 state\[42\] VPWR VGND sg13g2_nand2_1
XFILLER_19_396 VPWR VGND sg13g2_decap_4
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
X_2071_ VGND VPWR _0879_ _0725_ _0263_ net71 sg13g2_a21oi_1
XFILLER_15_591 VPWR VGND sg13g2_decap_4
X_1924_ net189 VPWR _0613_ VGND daisychain\[101\] net32 sg13g2_o21ai_1
X_1855_ VGND VPWR _0555_ _0556_ _0215_ _0557_ sg13g2_a21oi_1
X_1786_ state\[74\] daisychain\[74\] net151 _0502_ VPWR VGND sg13g2_mux2_1
XFILLER_38_661 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
X_2457__262 VPWR VGND net261 sg13g2_tiehi
X_2407_ net394 VGND VPWR _0223_ daisychain\[95\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2338_ net276 VGND VPWR _0154_ daisychain\[26\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2269_ VGND VPWR _0631_ _0824_ _0362_ net76 sg13g2_a21oi_1
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_4_248 VPWR VGND sg13g2_decap_8
XFILLER_5_727 VPWR VGND sg13g2_decap_8
XFILLER_5_738 VPWR VGND sg13g2_fill_1
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_20_75 VPWR VGND sg13g2_decap_8
XFILLER_16_300 VPWR VGND sg13g2_decap_8
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_29_73 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_44_631 VPWR VGND sg13g2_fill_2
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_8_532 VPWR VGND sg13g2_fill_2
XFILLER_3_281 VPWR VGND sg13g2_decap_8
XFILLER_6_33 VPWR VGND sg13g2_fill_2
X_1640_ VGND VPWR _1027_ _0384_ _0172_ _0385_ sg13g2_a21oi_1
X_1571_ state\[31\] daisychain\[31\] net140 _0974_ VPWR VGND sg13g2_mux2_1
XFILLER_39_447 VPWR VGND sg13g2_fill_2
X_2123_ VGND VPWR _0983_ _0751_ _0289_ net74 sg13g2_a21oi_1
XFILLER_22_303 VPWR VGND sg13g2_fill_1
XFILLER_22_336 VPWR VGND sg13g2_decap_4
XFILLER_34_152 VPWR VGND sg13g2_decap_8
XFILLER_35_620 VPWR VGND sg13g2_fill_2
X_2054_ net179 VPWR _0717_ VGND daisychain\[127\] net25 sg13g2_o21ai_1
X_1907_ _0599_ net165 _0598_ VPWR VGND sg13g2_nand2_1
X_1838_ VGND VPWR net124 daisychain\[83\] _0544_ net61 sg13g2_a21oi_1
X_1769_ net199 VPWR _0489_ VGND daisychain\[70\] net42 sg13g2_o21ai_1
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_13_314 VPWR VGND sg13g2_decap_8
XFILLER_15_86 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_9_329 VPWR VGND sg13g2_decap_8
XFILLER_31_74 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_36_417 VPWR VGND sg13g2_fill_2
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_decap_8
X_2553__312 VPWR VGND net311 sg13g2_tiehi
XFILLER_16_174 VPWR VGND sg13g2_decap_8
XFILLER_31_144 VPWR VGND sg13g2_decap_8
XFILLER_8_362 VPWR VGND sg13g2_decap_8
X_1485_ VGND VPWR _0903_ _0904_ _0141_ _0905_ sg13g2_a21oi_1
X_1554_ net184 VPWR _0961_ VGND daisychain\[27\] net27 sg13g2_o21ai_1
X_1623_ VGND VPWR net115 daisychain\[40\] _1016_ net57 sg13g2_a21oi_1
.ends

