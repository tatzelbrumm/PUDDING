VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO heichips25_pudding
  CLASS BLOCK ;
  FOREIGN heichips25_pudding ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 21.580 3.150 23.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 81.580 3.150 83.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 141.580 3.150 143.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 201.580 3.150 203.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 261.580 3.150 263.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 321.580 3.150 323.780 193.410 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 381.580 3.150 383.780 193.410 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 15.380 3.560 17.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 75.380 3.560 77.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 135.380 3.560 137.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 195.380 3.560 197.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 255.380 3.560 257.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 315.380 3.560 317.580 193.000 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 375.380 3.560 377.580 193.000 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.340 0.400 183.740 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.140 0.400 179.540 ;
    END
  END ena
  PIN i_in
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13075.336914 ;
    ANTENNADIFFAREA 13852.298828 ;
    PORT
      LAYER Metal3 ;
        RECT 438.885 107.930 500.000 108.630 ;
    END
  END i_in
  PIN i_out
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13075.336914 ;
    ANTENNADIFFAREA 13852.298828 ;
    PORT
      LAYER Metal3 ;
        RECT 400.000 99.745 500.000 100.445 ;
    END
  END i_out
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.540 0.400 187.940 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.940 0.400 112.340 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.140 0.400 116.540 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.340 0.400 120.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.540 0.400 124.940 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.740 0.400 129.140 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.940 0.400 133.340 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.140 0.400 137.540 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.340 0.400 141.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.540 0.400 145.940 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.740 0.400 150.140 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.940 0.400 154.340 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.140 0.400 158.540 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.340 0.400 162.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.540 0.400 166.940 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.740 0.400 171.140 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.940 0.400 175.340 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.340 0.400 78.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.540 0.400 82.940 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.400 87.140 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.940 0.400 91.340 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.140 0.400 95.540 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.340 0.400 99.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.540 0.400 103.940 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.740 0.400 108.140 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.740 0.400 45.140 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.140 0.400 53.540 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.540 0.400 61.940 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.740 0.400 66.140 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.940 0.400 70.340 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.140 0.400 74.540 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.140 0.400 11.540 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.540 0.400 19.940 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.940 0.400 28.340 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.340 0.400 36.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 421.405 192.930 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 421.945 196.060 ;
      LAYER Metal2 ;
        RECT 2.295 3.635 421.945 196.060 ;
      LAYER Metal3 ;
        RECT 0.400 188.150 438.885 192.880 ;
        RECT 0.610 187.330 438.885 188.150 ;
        RECT 0.400 183.950 438.885 187.330 ;
        RECT 0.610 183.130 438.885 183.950 ;
        RECT 0.400 179.750 438.885 183.130 ;
        RECT 0.610 178.930 438.885 179.750 ;
        RECT 0.400 175.550 438.885 178.930 ;
        RECT 0.610 174.730 438.885 175.550 ;
        RECT 0.400 171.350 438.885 174.730 ;
        RECT 0.610 170.530 438.885 171.350 ;
        RECT 0.400 167.150 438.885 170.530 ;
        RECT 0.610 166.330 438.885 167.150 ;
        RECT 0.400 162.950 438.885 166.330 ;
        RECT 0.610 162.130 438.885 162.950 ;
        RECT 0.400 158.750 438.885 162.130 ;
        RECT 0.610 157.930 438.885 158.750 ;
        RECT 0.400 154.550 438.885 157.930 ;
        RECT 0.610 153.730 438.885 154.550 ;
        RECT 0.400 150.350 438.885 153.730 ;
        RECT 0.610 149.530 438.885 150.350 ;
        RECT 0.400 146.150 438.885 149.530 ;
        RECT 0.610 145.330 438.885 146.150 ;
        RECT 0.400 141.950 438.885 145.330 ;
        RECT 0.610 141.130 438.885 141.950 ;
        RECT 0.400 137.750 438.885 141.130 ;
        RECT 0.610 136.930 438.885 137.750 ;
        RECT 0.400 133.550 438.885 136.930 ;
        RECT 0.610 132.730 438.885 133.550 ;
        RECT 0.400 129.350 438.885 132.730 ;
        RECT 0.610 128.530 438.885 129.350 ;
        RECT 0.400 125.150 438.885 128.530 ;
        RECT 0.610 124.330 438.885 125.150 ;
        RECT 0.400 120.950 438.885 124.330 ;
        RECT 0.610 120.130 438.885 120.950 ;
        RECT 0.400 116.750 438.885 120.130 ;
        RECT 0.610 115.930 438.885 116.750 ;
        RECT 0.400 112.550 438.885 115.930 ;
        RECT 0.610 111.730 438.885 112.550 ;
        RECT 0.400 108.840 438.885 111.730 ;
        RECT 0.400 108.350 438.675 108.840 ;
        RECT 0.610 107.720 438.675 108.350 ;
        RECT 0.610 107.530 438.885 107.720 ;
        RECT 0.400 104.150 438.885 107.530 ;
        RECT 0.610 103.330 438.885 104.150 ;
        RECT 0.400 100.655 438.885 103.330 ;
        RECT 0.400 99.950 399.790 100.655 ;
        RECT 0.610 99.535 399.790 99.950 ;
        RECT 0.610 99.130 438.885 99.535 ;
        RECT 0.400 95.750 438.885 99.130 ;
        RECT 0.610 94.930 438.885 95.750 ;
        RECT 0.400 91.550 438.885 94.930 ;
        RECT 0.610 90.730 438.885 91.550 ;
        RECT 0.400 87.350 438.885 90.730 ;
        RECT 0.610 86.530 438.885 87.350 ;
        RECT 0.400 83.150 438.885 86.530 ;
        RECT 0.610 82.330 438.885 83.150 ;
        RECT 0.400 78.950 438.885 82.330 ;
        RECT 0.610 78.130 438.885 78.950 ;
        RECT 0.400 74.750 438.885 78.130 ;
        RECT 0.610 73.930 438.885 74.750 ;
        RECT 0.400 70.550 438.885 73.930 ;
        RECT 0.610 69.730 438.885 70.550 ;
        RECT 0.400 66.350 438.885 69.730 ;
        RECT 0.610 65.530 438.885 66.350 ;
        RECT 0.400 62.150 438.885 65.530 ;
        RECT 0.610 61.330 438.885 62.150 ;
        RECT 0.400 57.950 438.885 61.330 ;
        RECT 0.610 57.130 438.885 57.950 ;
        RECT 0.400 53.750 438.885 57.130 ;
        RECT 0.610 52.930 438.885 53.750 ;
        RECT 0.400 49.550 438.885 52.930 ;
        RECT 0.610 48.730 438.885 49.550 ;
        RECT 0.400 45.350 438.885 48.730 ;
        RECT 0.610 44.530 438.885 45.350 ;
        RECT 0.400 41.150 438.885 44.530 ;
        RECT 0.610 40.330 438.885 41.150 ;
        RECT 0.400 36.950 438.885 40.330 ;
        RECT 0.610 36.130 438.885 36.950 ;
        RECT 0.400 32.750 438.885 36.130 ;
        RECT 0.610 31.930 438.885 32.750 ;
        RECT 0.400 28.550 438.885 31.930 ;
        RECT 0.610 27.730 438.885 28.550 ;
        RECT 0.400 24.350 438.885 27.730 ;
        RECT 0.610 23.530 438.885 24.350 ;
        RECT 0.400 20.150 438.885 23.530 ;
        RECT 0.610 19.330 438.885 20.150 ;
        RECT 0.400 15.950 438.885 19.330 ;
        RECT 0.610 15.130 438.885 15.950 ;
        RECT 0.400 11.750 438.885 15.130 ;
        RECT 0.610 10.930 438.885 11.750 ;
        RECT 0.400 3.680 438.885 10.930 ;
      LAYER Metal4 ;
        RECT 15.560 3.635 400.000 192.925 ;
      LAYER Metal5 ;
        RECT 15.515 3.470 400.000 193.090 ;
      LAYER TopMetal1 ;
        RECT 358.780 80.240 373.740 119.680 ;
        RECT 379.220 80.240 379.940 119.680 ;
        RECT 385.420 80.240 394.620 119.680 ;
  END
END heichips25_pudding
END LIBRARY

