* NGSPICE file created from heichips25_pudding.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for analog_wires abstract view
.subckt analog_wires Iout VcascP[1] VcascP[0] VbiasP[1] VbiasP[0] VDDA[1] VDDA[0]
+ i_in i_out
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for dac128module abstract view
.subckt dac128module VbiasP[1] Iout VbiasP[0] VcascP[1] VcascP[0] ON[64] ONB[64] ON[65]
+ ONB[65] ON[66] ONB[66] ON[67] ONB[67] ON[68] ONB[68] ON[69] ONB[69] ON[70] ONB[70]
+ ON[71] ONB[71] ON[72] ONB[72] EN[2] ENB[2] ON[73] ONB[73] ON[74] ONB[74] ON[75]
+ ONB[75] ON[76] ONB[76] ON[77] ONB[77] ON[78] ONB[78] ON[79] ONB[79] ON[80] ONB[80]
+ ON[81] ONB[81] ON[82] ONB[82] ON[83] ONB[83] ON[84] ONB[84] ON[85] ONB[85] ON[86]
+ ONB[86] ON[87] ONB[87] ON[88] ONB[88] ON[89] ONB[89] ON[90] ONB[90] ON[91] ONB[91]
+ ON[92] ONB[92] ON[93] ONB[93] ON[94] ONB[94] ON[95] ONB[95] ON[96] ONB[96] ON[97]
+ ONB[97] ON[98] ONB[98] ON[99] ONB[99] ON[100] ONB[100] ON[101] ONB[101] ON[102]
+ ONB[102] ON[103] ONB[103] ON[104] ONB[104] ON[105] ONB[105] ON[106] ONB[106] ON[107]
+ ONB[107] ON[108] ONB[108] ON[109] ONB[109] ON[110] ONB[110] ON[111] ONB[111] ON[112]
+ ONB[112] ON[113] ONB[113] ON[114] ONB[114] ON[115] ONB[115] ON[116] ONB[116] ON[117]
+ ONB[117] ON[118] ONB[118] ON[119] ONB[119] ON[120] ONB[120] ON[121] ONB[121] ON[122]
+ ONB[122] EN[3] ENB[3] ON[123] ONB[123] ON[124] ONB[124] ON[125] ONB[125] ON[126]
+ ONB[126] ON[127] ONB[127] ON[0] ONB[0] ON[1] ONB[1] ON[2] ONB[2] ON[3] ONB[3] ON[4]
+ ONB[4] ON[5] ONB[5] ON[6] EN[0] ENB[0] ONB[6] ON[7] ONB[7] ON[8] ONB[8] ON[9] ONB[9]
+ ON[10] ONB[10] ON[11] ONB[11] ON[12] ONB[12] ON[13] ONB[13] ON[14] ONB[14] ON[15]
+ ONB[15] ON[16] ONB[16] ON[17] ONB[17] ON[18] ONB[18] ON[19] ONB[19] ON[20] ONB[20]
+ ON[21] ONB[21] ON[22] ONB[22] ON[23] ONB[23] ON[24] ONB[24] ON[25] ONB[25] ON[26]
+ ONB[26] ON[27] ONB[27] ON[28] ONB[28] ON[29] ONB[29] ON[30] ONB[30] ON[31] ONB[31]
+ ON[33] ONB[33] ON[32] ONB[32] ON[34] ONB[34] ON[35] ONB[35] ON[36] ONB[36] ON[37]
+ ONB[37] ON[38] ONB[38] ON[39] ONB[39] ON[40] ONB[40] ON[41] ONB[41] ON[42] ONB[42]
+ ON[43] ONB[43] ON[44] ONB[44] ON[45] ONB[45] ON[46] ONB[46] ON[47] ONB[47] ON[48]
+ ONB[48] ON[49] ONB[49] ON[50] ONB[50] ON[51] ONB[51] ON[52] ONB[52] ON[53] ONB[53]
+ ON[54] ONB[54] ON[55] ONB[55] ON[56] ONB[56] ON[57] ONB[57] ON[58] ONB[58] ON[59]
+ ONB[59] ON[60] ONB[60] ON[61] ONB[61] ON[62] ONB[62] ON[63] ONB[63] EN[1] ENB[1]
+ VSS VDD
.ends

.subckt heichips25_pudding VGND VPWR clk ena i_in i_out rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_266 VPWR VGND sg13g2_decap_8
X_2037_ net198 VGND VPWR _0369_ state\[113\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_166 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_46_726 VPWR VGND sg13g2_decap_8
XFILLER_14_612 VPWR VGND sg13g2_fill_1
XFILLER_26_483 VPWR VGND sg13g2_fill_1
XFILLER_26_494 VPWR VGND sg13g2_decap_8
XFILLER_41_420 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_14_689 VPWR VGND sg13g2_fill_1
XFILLER_41_497 VPWR VGND sg13g2_decap_8
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
X_1270_ VGND VPWR net72 daisychain\[27\] _0397_ net34 sg13g2_a21oi_1
XFILLER_44_280 VPWR VGND sg13g2_decap_8
X_1606_ VGND VPWR net75 daisychain\[111\] _0649_ net37 sg13g2_a21oi_1
X_0985_ VPWR _0103_ state\[78\] VGND sg13g2_inv_1
Xfanout105 net106 net105 VPWR VGND sg13g2_buf_1
Xfanout116 net135 net116 VPWR VGND sg13g2_buf_1
Xfanout127 net134 net127 VPWR VGND sg13g2_buf_1
Xfanout138 net141 net138 VPWR VGND sg13g2_buf_1
Xfanout149 net157 net149 VPWR VGND sg13g2_buf_1
X_1537_ _0796_ net109 _0596_ _0597_ VPWR VGND sg13g2_a21o_1
X_1468_ net175 VPWR _0545_ VGND net128 state\[78\] sg13g2_o21ai_1
X_1399_ _0188_ _0492_ _0493_ net52 _0761_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_214 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_11_615 VPWR VGND sg13g2_decap_4
XFILLER_12_76 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
XFILLER_33_228 VPWR VGND sg13g2_decap_8
XFILLER_34_729 VPWR VGND sg13g2_fill_2
XFILLER_41_294 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_6_663 VPWR VGND sg13g2_fill_2
X_1322_ VGND VPWR net79 daisychain\[40\] _0436_ net46 sg13g2_a21oi_1
X_1253_ _0725_ net102 _0897_ _0384_ VPWR VGND sg13g2_a21o_1
XFILLER_49_361 VPWR VGND sg13g2_decap_8
X_1184_ net139 VPWR _0846_ VGND net92 state\[7\] sg13g2_o21ai_1
X_0968_ VPWR _0085_ state\[61\] VGND sg13g2_inv_1
X_0899_ VPWR _0696_ net138 VGND sg13g2_inv_1
XFILLER_23_20 VPWR VGND sg13g2_decap_8
XFILLER_23_261 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_fill_2
XFILLER_43_537 VPWR VGND sg13g2_fill_1
XFILLER_3_611 VPWR VGND sg13g2_decap_4
XFILLER_7_427 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_501 VPWR VGND sg13g2_fill_2
XFILLER_19_523 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_14_272 VPWR VGND sg13g2_decap_8
XFILLER_15_784 VPWR VGND sg13g2_decap_4
XFILLER_15_795 VPWR VGND sg13g2_fill_2
XFILLER_30_754 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
X_1940_ net189 VGND VPWR _0272_ state\[16\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1871_ net220 VGND VPWR _0203_ daisychain\[75\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_9_88 VPWR VGND sg13g2_decap_8
X_1305_ _0738_ net115 _0422_ _0423_ VPWR VGND sg13g2_a21o_1
X_1236_ net147 VPWR _0885_ VGND net101 state\[20\] sg13g2_o21ai_1
XFILLER_12_209 VPWR VGND sg13g2_decap_8
XFILLER_37_364 VPWR VGND sg13g2_decap_8
X_1167_ _0130_ _0832_ _0833_ net38 _0703_ VPWR VGND sg13g2_a22oi_1
X_1098_ VPWR _0767_ daisychain\[66\] VGND sg13g2_inv_1
XFILLER_20_231 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_28_331 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_44_813 VPWR VGND sg13g2_decap_8
XFILLER_11_242 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_decap_8
X_2070_ daisychain\[122\] net17 VPWR VGND sg13g2_buf_1
XFILLER_34_301 VPWR VGND sg13g2_decap_8
XFILLER_34_378 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
X_1021_ VPWR _0016_ state\[114\] VGND sg13g2_inv_1
X_1923_ net184 VGND VPWR _0255_ daisychain\[127\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1854_ net209 VGND VPWR _0186_ daisychain\[58\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1785_ _0663_ VPWR _0373_ VGND net140 _0019_ sg13g2_o21ai_1
XFILLER_29_139 VPWR VGND sg13g2_decap_8
XFILLER_37_161 VPWR VGND sg13g2_decap_8
X_1219_ _0143_ _0871_ _0872_ net31 _0716_ VPWR VGND sg13g2_a22oi_1
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_29_41 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_16_356 VPWR VGND sg13g2_decap_8
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_12_595 VPWR VGND sg13g2_decap_4
XANTENNA_5 VPWR VGND state\[56\] sg13g2_antennanp
XFILLER_6_67 VPWR VGND sg13g2_decap_8
X_1570_ VGND VPWR net77 daisychain\[102\] _0622_ net40 sg13g2_a21oi_1
XFILLER_20_4 VPWR VGND sg13g2_decap_4
XFILLER_39_448 VPWR VGND sg13g2_decap_8
XFILLER_34_175 VPWR VGND sg13g2_decap_8
X_1004_ VPWR _0124_ state\[97\] VGND sg13g2_inv_1
X_1906_ net197 VGND VPWR _0238_ daisychain\[110\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1837_ net204 VGND VPWR _0169_ daisychain\[41\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1768_ _0612_ VPWR _0356_ VGND net171 _0001_ sg13g2_o21ai_1
X_1699_ _0405_ VPWR _0287_ VGND net158 _0052_ sg13g2_o21ai_1
XFILLER_25_131 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_15_76 VPWR VGND sg13g2_decap_8
XFILLER_31_20 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_41_646 VPWR VGND sg13g2_fill_1
XFILLER_9_319 VPWR VGND sg13g2_decap_8
XFILLER_31_97 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_fill_1
XFILLER_5_547 VPWR VGND sg13g2_fill_2
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_decap_8
XFILLER_16_153 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_fill_1
XFILLER_31_167 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_8
XFILLER_12_370 VPWR VGND sg13g2_decap_8
XFILLER_8_396 VPWR VGND sg13g2_decap_8
X_1622_ VGND VPWR net68 daisychain\[115\] _0661_ net27 sg13g2_a21oi_1
X_1553_ _0800_ net108 _0608_ _0609_ VPWR VGND sg13g2_a21o_1
X_1484_ net170 VPWR _0557_ VGND net127 state\[82\] sg13g2_o21ai_1
XFILLER_27_429 VPWR VGND sg13g2_fill_2
XFILLER_39_245 VPWR VGND sg13g2_decap_8
X_2036_ net196 VGND VPWR _0368_ state\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_145 VPWR VGND sg13g2_decap_8
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_14_635 VPWR VGND sg13g2_decap_4
XFILLER_14_646 VPWR VGND sg13g2_fill_1
XFILLER_26_473 VPWR VGND sg13g2_decap_4
XFILLER_41_476 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_5_333 VPWR VGND sg13g2_decap_8
XFILLER_6_812 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_37_705 VPWR VGND sg13g2_fill_1
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_20_616 VPWR VGND sg13g2_fill_2
XFILLER_32_454 VPWR VGND sg13g2_fill_2
XFILLER_32_498 VPWR VGND sg13g2_decap_8
X_0984_ VPWR _0102_ state\[77\] VGND sg13g2_inv_1
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_1605_ _0813_ net104 _0647_ _0648_ VPWR VGND sg13g2_a21o_1
X_1536_ net154 VPWR _0596_ VGND net108 state\[95\] sg13g2_o21ai_1
XFILLER_9_672 VPWR VGND sg13g2_decap_4
Xfanout106 net111 net106 VPWR VGND sg13g2_buf_1
Xfanout117 net118 net117 VPWR VGND sg13g2_buf_1
Xfanout128 net134 net128 VPWR VGND sg13g2_buf_1
Xfanout139 net140 net139 VPWR VGND sg13g2_buf_1
X_1467_ _0205_ _0543_ _0544_ net61 _0778_ VPWR VGND sg13g2_a22oi_1
X_1398_ VGND VPWR net82 daisychain\[59\] _0493_ net52 sg13g2_a21oi_1
X_2019_ net202 VGND VPWR _0351_ state\[95\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_12_55 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_19_716 VPWR VGND sg13g2_fill_1
XFILLER_33_207 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_6_642 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
X_1321_ _0742_ net114 _0434_ _0435_ VPWR VGND sg13g2_a21o_1
X_1252_ net148 VPWR _0897_ VGND net102 state\[24\] sg13g2_o21ai_1
XFILLER_33_774 VPWR VGND sg13g2_fill_2
XFILLER_37_579 VPWR VGND sg13g2_fill_2
X_1183_ _0134_ _0844_ _0845_ net25 _0707_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_424 VPWR VGND sg13g2_decap_8
XFILLER_32_284 VPWR VGND sg13g2_decap_8
X_0967_ VPWR _0084_ state\[60\] VGND sg13g2_inv_1
XFILLER_9_491 VPWR VGND sg13g2_fill_1
X_1519_ _0218_ _0582_ _0583_ net43 _0791_ VPWR VGND sg13g2_a22oi_1
X_0898_ VPWR _0695_ daisychain\[123\] VGND sg13g2_inv_1
XFILLER_11_424 VPWR VGND sg13g2_decap_8
XFILLER_11_435 VPWR VGND sg13g2_fill_2
XFILLER_23_240 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_3_623 VPWR VGND sg13g2_fill_1
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_14_251 VPWR VGND sg13g2_decap_8
X_1870_ net220 VGND VPWR _0202_ daisychain\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_6_494 VPWR VGND sg13g2_decap_8
XFILLER_37_343 VPWR VGND sg13g2_decap_8
X_1304_ net161 VPWR _0422_ VGND net115 state\[37\] sg13g2_o21ai_1
X_1235_ _0147_ _0883_ _0884_ net34 _0720_ VPWR VGND sg13g2_a22oi_1
X_1166_ VGND VPWR net75 daisychain\[1\] _0833_ net38 sg13g2_a21oi_1
XFILLER_20_210 VPWR VGND sg13g2_decap_8
X_1097_ VPWR _0766_ daisychain\[65\] VGND sg13g2_inv_1
X_1999_ net221 VGND VPWR _0331_ state\[75\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_16_516 VPWR VGND sg13g2_fill_1
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_11_221 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_fill_1
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_3_420 VPWR VGND sg13g2_decap_8
XFILLER_3_497 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
X_1020_ VPWR _0015_ state\[113\] VGND sg13g2_inv_1
XFILLER_15_593 VPWR VGND sg13g2_fill_1
XFILLER_19_398 VPWR VGND sg13g2_decap_8
XFILLER_34_357 VPWR VGND sg13g2_decap_8
X_1922_ net183 VGND VPWR _0254_ daisychain\[126\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1853_ net209 VGND VPWR _0185_ daisychain\[57\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1784_ _0660_ VPWR _0372_ VGND net151 _0018_ sg13g2_o21ai_1
XFILLER_29_118 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_38_663 VPWR VGND sg13g2_decap_4
X_1218_ VGND VPWR net74 daisychain\[14\] _0872_ net31 sg13g2_a21oi_1
X_1149_ VPWR _0818_ daisychain\[117\] VGND sg13g2_inv_1
XFILLER_20_55 VPWR VGND sg13g2_decap_4
XFILLER_4_228 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_29_20 VPWR VGND sg13g2_decap_8
XFILLER_29_97 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_16_335 VPWR VGND sg13g2_decap_8
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_31_349 VPWR VGND sg13g2_decap_8
XFILLER_32_806 VPWR VGND sg13g2_fill_1
XFILLER_32_817 VPWR VGND sg13g2_decap_4
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XANTENNA_6 VPWR VGND state\[83\] sg13g2_antennanp
XFILLER_12_563 VPWR VGND sg13g2_fill_1
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_8_512 VPWR VGND sg13g2_fill_2
XFILLER_3_294 VPWR VGND sg13g2_decap_8
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_19_195 VPWR VGND sg13g2_decap_8
XFILLER_35_622 VPWR VGND sg13g2_fill_2
XFILLER_39_427 VPWR VGND sg13g2_decap_8
X_1003_ VPWR _0123_ state\[96\] VGND sg13g2_inv_1
XFILLER_34_154 VPWR VGND sg13g2_decap_8
X_1905_ net199 VGND VPWR _0237_ daisychain\[109\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_30_393 VPWR VGND sg13g2_fill_2
X_1836_ net205 VGND VPWR _0168_ daisychain\[40\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1767_ _0609_ VPWR _0355_ VGND net156 _0126_ sg13g2_o21ai_1
X_1698_ _0402_ VPWR _0286_ VGND net158 _0051_ sg13g2_o21ai_1
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_55 VPWR VGND sg13g2_decap_8
XFILLER_25_187 VPWR VGND sg13g2_decap_8
XFILLER_38_460 VPWR VGND sg13g2_decap_4
XFILLER_41_625 VPWR VGND sg13g2_fill_1
XFILLER_31_76 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_5_515 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_16_132 VPWR VGND sg13g2_decap_8
XFILLER_29_471 VPWR VGND sg13g2_fill_1
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_31_146 VPWR VGND sg13g2_decap_8
XFILLER_8_375 VPWR VGND sg13g2_decap_8
X_1621_ _0817_ net94 _0659_ _0660_ VPWR VGND sg13g2_a21o_1
X_1552_ net155 VPWR _0608_ VGND net110 state\[99\] sg13g2_o21ai_1
XFILLER_39_224 VPWR VGND sg13g2_decap_8
X_1483_ _0209_ _0555_ _0556_ net56 _0782_ VPWR VGND sg13g2_a22oi_1
X_2035_ net197 VGND VPWR _0367_ state\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_31_680 VPWR VGND sg13g2_decap_8
XFILLER_2_529 VPWR VGND sg13g2_decap_8
X_1819_ net193 VGND VPWR _0151_ daisychain\[23\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_26_452 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_4
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_17_485 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_45_750 VPWR VGND sg13g2_fill_2
XFILLER_32_466 VPWR VGND sg13g2_fill_2
XFILLER_8_172 VPWR VGND sg13g2_decap_8
X_0983_ VPWR _0101_ state\[76\] VGND sg13g2_inv_1
XFILLER_9_640 VPWR VGND sg13g2_fill_1
Xfanout107 net110 net107 VPWR VGND sg13g2_buf_1
Xfanout118 net122 net118 VPWR VGND sg13g2_buf_1
Xfanout129 net134 net129 VPWR VGND sg13g2_buf_1
X_1604_ net150 VPWR _0647_ VGND net104 state\[112\] sg13g2_o21ai_1
X_1535_ _0222_ _0594_ _0595_ net41 _0795_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_249 VPWR VGND sg13g2_decap_8
X_1466_ VGND VPWR net87 daisychain\[76\] _0544_ net61 sg13g2_a21oi_1
X_1397_ _0761_ net122 _0491_ _0492_ VPWR VGND sg13g2_a21o_1
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_36_750 VPWR VGND sg13g2_fill_1
X_2018_ net201 VGND VPWR _0350_ state\[94\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_12_34 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_42_775 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
X_1320_ net159 VPWR _0434_ VGND net114 state\[41\] sg13g2_o21ai_1
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
X_1251_ _0151_ _0895_ _0896_ net35 _0724_ VPWR VGND sg13g2_a22oi_1
X_1182_ VGND VPWR net71 daisychain\[5\] _0845_ net30 sg13g2_a21oi_1
XFILLER_17_293 VPWR VGND sg13g2_decap_8
XFILLER_18_783 VPWR VGND sg13g2_fill_1
XFILLER_24_219 VPWR VGND sg13g2_decap_8
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_20_469 VPWR VGND sg13g2_fill_2
X_0966_ VPWR _0082_ state\[59\] VGND sg13g2_inv_1
X_1518_ VGND VPWR net76 daisychain\[89\] _0583_ net41 sg13g2_a21oi_1
X_1449_ _0774_ net130 _0530_ _0531_ VPWR VGND sg13g2_a21o_1
XFILLER_43_506 VPWR VGND sg13g2_fill_1
XFILLER_11_403 VPWR VGND sg13g2_decap_8
XFILLER_11_469 VPWR VGND sg13g2_fill_2
XFILLER_23_296 VPWR VGND sg13g2_decap_8
XFILLER_23_66 VPWR VGND sg13g2_fill_2
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_19_503 VPWR VGND sg13g2_fill_1
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_14_230 VPWR VGND sg13g2_decap_8
XFILLER_19_569 VPWR VGND sg13g2_fill_1
XFILLER_30_712 VPWR VGND sg13g2_fill_1
XFILLER_42_561 VPWR VGND sg13g2_fill_1
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_30_734 VPWR VGND sg13g2_fill_1
XFILLER_30_778 VPWR VGND sg13g2_fill_2
XFILLER_42_594 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_6_473 VPWR VGND sg13g2_decap_8
X_1303_ _0164_ _0420_ _0421_ net48 _0737_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_37_399 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
X_1234_ VGND VPWR net72 daisychain\[18\] _0884_ net34 sg13g2_a21oi_1
X_1165_ _0703_ net101 _0831_ _0832_ VPWR VGND sg13g2_a21o_1
X_1096_ VPWR _0765_ daisychain\[64\] VGND sg13g2_inv_1
XFILLER_20_266 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_fill_1
X_1998_ net221 VGND VPWR _0330_ state\[74\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_0949_ VPWR _0064_ state\[42\] VGND sg13g2_inv_1
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_28_344 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_11_200 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_476 VPWR VGND sg13g2_decap_8
XFILLER_15_8 VPWR VGND sg13g2_fill_1
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_30_553 VPWR VGND sg13g2_fill_1
XFILLER_34_336 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_decap_8
X_1921_ net183 VGND VPWR _0253_ daisychain\[125\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1852_ net211 VGND VPWR _0184_ daisychain\[56\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_30_575 VPWR VGND sg13g2_fill_1
XFILLER_6_270 VPWR VGND sg13g2_decap_8
X_1783_ _0657_ VPWR _0371_ VGND net150 _0017_ sg13g2_o21ai_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_25_325 VPWR VGND sg13g2_fill_1
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_38_642 VPWR VGND sg13g2_decap_8
X_1217_ _0716_ net97 _0870_ _0871_ VPWR VGND sg13g2_a21o_1
X_1148_ VPWR _0817_ daisychain\[116\] VGND sg13g2_inv_1
X_1079_ VPWR _0748_ daisychain\[47\] VGND sg13g2_inv_1
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_20_34 VPWR VGND sg13g2_decap_8
XFILLER_20_89 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
XFILLER_16_314 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_29_76 VPWR VGND sg13g2_decap_8
XFILLER_44_601 VPWR VGND sg13g2_fill_1
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_12_520 VPWR VGND sg13g2_fill_2
XFILLER_12_531 VPWR VGND sg13g2_fill_1
XFILLER_31_328 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_44_634 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_3_273 VPWR VGND sg13g2_decap_8
XFILLER_19_174 VPWR VGND sg13g2_decap_8
XFILLER_22_306 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
XFILLER_35_601 VPWR VGND sg13g2_decap_4
XFILLER_35_689 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
X_2051_ net184 VGND VPWR _0383_ state\[127\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1002_ VPWR _0122_ state\[95\] VGND sg13g2_inv_1
XFILLER_15_391 VPWR VGND sg13g2_decap_8
XFILLER_30_361 VPWR VGND sg13g2_decap_8
X_1904_ net197 VGND VPWR _0236_ daisychain\[108\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1835_ net204 VGND VPWR _0167_ daisychain\[39\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1766_ _0606_ VPWR _0354_ VGND net154 _0125_ sg13g2_o21ai_1
X_1697_ _0399_ VPWR _0285_ VGND net149 _0049_ sg13g2_o21ai_1
XFILLER_15_34 VPWR VGND sg13g2_decap_8
XFILLER_25_166 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_31_11 VPWR VGND sg13g2_fill_1
XFILLER_31_55 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
Xoutput9 net9 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_16_111 VPWR VGND sg13g2_decap_8
XFILLER_17_656 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_16_188 VPWR VGND sg13g2_decap_8
XFILLER_31_125 VPWR VGND sg13g2_decap_8
XFILLER_44_497 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
X_1620_ net150 VPWR _0659_ VGND net94 state\[116\] sg13g2_o21ai_1
X_1551_ _0226_ _0606_ _0607_ net42 _0799_ VPWR VGND sg13g2_a22oi_1
X_1482_ VGND VPWR net85 daisychain\[80\] _0556_ net56 sg13g2_a21oi_1
XFILLER_39_203 VPWR VGND sg13g2_decap_8
XFILLER_35_475 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
X_2034_ net199 VGND VPWR _0366_ state\[110\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1818_ net193 VGND VPWR _0150_ daisychain\[22\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_2_508 VPWR VGND sg13g2_decap_8
X_1749_ _0555_ VPWR _0337_ VGND net174 _0107_ sg13g2_o21ai_1
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_442 VPWR VGND sg13g2_decap_4
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_10_821 VPWR VGND sg13g2_fill_2
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_21_180 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_49_578 VPWR VGND sg13g2_decap_8
XFILLER_17_442 VPWR VGND sg13g2_decap_8
XFILLER_32_423 VPWR VGND sg13g2_decap_4
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_45_784 VPWR VGND sg13g2_decap_8
XFILLER_20_618 VPWR VGND sg13g2_fill_1
XFILLER_32_478 VPWR VGND sg13g2_decap_8
XFILLER_32_489 VPWR VGND sg13g2_fill_2
XFILLER_8_151 VPWR VGND sg13g2_decap_8
X_0982_ VPWR _0100_ state\[75\] VGND sg13g2_inv_1
Xfanout108 net109 net108 VPWR VGND sg13g2_buf_1
Xfanout119 net122 net119 VPWR VGND sg13g2_buf_1
X_1603_ _0239_ _0645_ _0646_ net39 _0812_ VPWR VGND sg13g2_a22oi_1
X_1534_ VGND VPWR net76 daisychain\[93\] _0595_ net41 sg13g2_a21oi_1
X_1465_ _0778_ net128 _0542_ _0543_ VPWR VGND sg13g2_a21o_1
XFILLER_27_228 VPWR VGND sg13g2_decap_8
XFILLER_36_740 VPWR VGND sg13g2_fill_1
X_2017_ net216 VGND VPWR _0349_ state\[93\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_1396_ net165 VPWR _0491_ VGND net118 state\[60\] sg13g2_o21ai_1
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_12_13 VPWR VGND sg13g2_decap_8
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_14_412 VPWR VGND sg13g2_decap_8
XFILLER_18_228 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_42_754 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_6_688 VPWR VGND sg13g2_decap_8
XFILLER_18_762 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
X_1250_ VGND VPWR net73 daisychain\[22\] _0896_ net35 sg13g2_a21oi_1
X_1181_ _0707_ net96 _0843_ _0844_ VPWR VGND sg13g2_a21o_1
XFILLER_17_272 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_33_776 VPWR VGND sg13g2_fill_1
X_0965_ VPWR _0081_ state\[58\] VGND sg13g2_inv_1
X_1517_ _0791_ net126 _0581_ _0582_ VPWR VGND sg13g2_a21o_1
X_1448_ net177 VPWR _0530_ VGND net130 state\[73\] sg13g2_o21ai_1
XFILLER_15_209 VPWR VGND sg13g2_decap_8
XFILLER_36_570 VPWR VGND sg13g2_decap_8
X_1379_ _0183_ _0477_ _0478_ net50 _0756_ VPWR VGND sg13g2_a22oi_1
XFILLER_23_275 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_19_537 VPWR VGND sg13g2_fill_1
XFILLER_34_507 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_14_286 VPWR VGND sg13g2_decap_8
XFILLER_30_746 VPWR VGND sg13g2_fill_1
XFILLER_42_573 VPWR VGND sg13g2_fill_2
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_30_768 VPWR VGND sg13g2_decap_4
XFILLER_6_452 VPWR VGND sg13g2_decap_8
Xfanout90 net136 net90 VPWR VGND sg13g2_buf_1
X_1302_ VGND VPWR net80 daisychain\[35\] _0421_ net48 sg13g2_a21oi_1
X_1233_ _0720_ net99 _0882_ _0883_ VPWR VGND sg13g2_a21o_1
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
X_1164_ net147 VPWR _0831_ VGND net101 state\[2\] sg13g2_o21ai_1
X_1095_ VPWR _0764_ daisychain\[63\] VGND sg13g2_inv_1
XFILLER_20_245 VPWR VGND sg13g2_decap_8
XFILLER_33_573 VPWR VGND sg13g2_fill_2
X_1997_ net222 VGND VPWR _0329_ state\[73\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_0948_ VPWR _0063_ state\[41\] VGND sg13g2_inv_1
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_28_312 VPWR VGND sg13g2_decap_4
XFILLER_12_735 VPWR VGND sg13g2_decap_4
XFILLER_28_389 VPWR VGND sg13g2_decap_8
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
XFILLER_12_779 VPWR VGND sg13g2_decap_8
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_3_455 VPWR VGND sg13g2_decap_8
XFILLER_34_315 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_47_632 VPWR VGND sg13g2_decap_4
Xheichips25_pudding_228 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_15_562 VPWR VGND sg13g2_decap_4
XFILLER_30_598 VPWR VGND sg13g2_decap_8
XFILLER_42_392 VPWR VGND sg13g2_decap_8
X_1920_ net183 VGND VPWR _0252_ daisychain\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1851_ net211 VGND VPWR _0183_ daisychain\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_7_783 VPWR VGND sg13g2_decap_8
X_1782_ _0654_ VPWR _0370_ VGND net152 _0016_ sg13g2_o21ai_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
X_1216_ net143 VPWR _0870_ VGND net97 state\[15\] sg13g2_o21ai_1
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_38_687 VPWR VGND sg13g2_fill_1
XFILLER_40_329 VPWR VGND sg13g2_decap_8
X_1147_ VPWR _0816_ daisychain\[115\] VGND sg13g2_inv_1
X_1078_ VPWR _0747_ daisychain\[46\] VGND sg13g2_inv_1
XFILLER_20_13 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_20_68 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_29_55 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv1 VPWR digitalen.g\[2\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_24_370 VPWR VGND sg13g2_fill_1
XFILLER_31_307 VPWR VGND sg13g2_decap_8
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_8_514 VPWR VGND sg13g2_fill_1
XFILLER_3_252 VPWR VGND sg13g2_decap_8
X_2050_ net184 VGND VPWR _0382_ state\[126\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_15_370 VPWR VGND sg13g2_decap_8
XFILLER_19_153 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_34_189 VPWR VGND sg13g2_decap_8
XFILLER_35_624 VPWR VGND sg13g2_fill_1
XFILLER_47_462 VPWR VGND sg13g2_decap_8
X_1001_ VPWR _0121_ state\[94\] VGND sg13g2_inv_1
XFILLER_30_340 VPWR VGND sg13g2_decap_8
XFILLER_30_395 VPWR VGND sg13g2_fill_1
X_1903_ net197 VGND VPWR _0235_ daisychain\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1834_ net204 VGND VPWR _0166_ daisychain\[38\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1765_ _0603_ VPWR _0353_ VGND net154 _0124_ sg13g2_o21ai_1
X_1696_ _0396_ VPWR _0284_ VGND net149 _0048_ sg13g2_o21ai_1
XFILLER_15_13 VPWR VGND sg13g2_decap_8
XFILLER_25_145 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_31_34 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_1_778 VPWR VGND sg13g2_fill_1
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_49_749 VPWR VGND sg13g2_decap_8
XFILLER_16_167 VPWR VGND sg13g2_decap_8
XFILLER_31_104 VPWR VGND sg13g2_decap_8
XFILLER_44_476 VPWR VGND sg13g2_decap_8
XFILLER_12_384 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_4
X_1550_ VGND VPWR net76 daisychain\[97\] _0607_ net42 sg13g2_a21oi_1
X_1481_ _0782_ net123 _0554_ _0555_ VPWR VGND sg13g2_a21o_1
XFILLER_35_410 VPWR VGND sg13g2_fill_2
XFILLER_35_421 VPWR VGND sg13g2_decap_8
XFILLER_39_259 VPWR VGND sg13g2_decap_8
X_2033_ net199 VGND VPWR _0365_ state\[109\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_22_159 VPWR VGND sg13g2_decap_8
XFILLER_35_465 VPWR VGND sg13g2_decap_4
XFILLER_7_91 VPWR VGND sg13g2_decap_8
X_1817_ net193 VGND VPWR _0149_ daisychain\[21\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1748_ _0552_ VPWR _0336_ VGND net170 _0106_ sg13g2_o21ai_1
X_1679_ _0859_ VPWR _0267_ VGND net140 _0022_ sg13g2_o21ai_1
XFILLER_14_605 VPWR VGND sg13g2_fill_2
XFILLER_26_487 VPWR VGND sg13g2_decap_8
XFILLER_41_413 VPWR VGND sg13g2_decap_8
XFILLER_46_719 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_32_402 VPWR VGND sg13g2_fill_1
XFILLER_44_273 VPWR VGND sg13g2_decap_8
X_0981_ VPWR _0099_ state\[74\] VGND sg13g2_inv_1
XFILLER_12_181 VPWR VGND sg13g2_decap_8
XFILLER_40_490 VPWR VGND sg13g2_decap_8
XFILLER_8_130 VPWR VGND sg13g2_decap_8
X_1602_ VGND VPWR net75 daisychain\[110\] _0646_ net39 sg13g2_a21oi_1
Xfanout109 net110 net109 VPWR VGND sg13g2_buf_1
X_1533_ _0795_ net108 _0593_ _0594_ VPWR VGND sg13g2_a21o_1
X_1464_ net175 VPWR _0542_ VGND net128 state\[77\] sg13g2_o21ai_1
X_1395_ _0187_ _0489_ _0490_ net52 _0760_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_207 VPWR VGND sg13g2_decap_8
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_36_763 VPWR VGND sg13g2_decap_4
X_2016_ net217 VGND VPWR _0348_ state\[92\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_12_69 VPWR VGND sg13g2_decap_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_39_590 VPWR VGND sg13g2_fill_1
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_10_674 VPWR VGND sg13g2_decap_4
XFILLER_22_490 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_6_656 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_17_251 VPWR VGND sg13g2_decap_8
XFILLER_37_505 VPWR VGND sg13g2_fill_2
XFILLER_45_560 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
X_1180_ net142 VPWR _0843_ VGND net96 state\[6\] sg13g2_o21ai_1
XFILLER_20_438 VPWR VGND sg13g2_fill_1
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_8
XFILLER_33_755 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_0964_ VPWR _0080_ state\[57\] VGND sg13g2_inv_1
X_1516_ net171 VPWR _0581_ VGND net124 state\[90\] sg13g2_o21ai_1
XFILLER_4_81 VPWR VGND sg13g2_decap_8
X_1447_ _0200_ _0528_ _0529_ net63 _0773_ VPWR VGND sg13g2_a22oi_1
X_1378_ VGND VPWR net81 daisychain\[54\] _0478_ net50 sg13g2_a21oi_1
XFILLER_23_254 VPWR VGND sg13g2_decap_8
XFILLER_23_13 VPWR VGND sg13g2_decap_8
XFILLER_23_68 VPWR VGND sg13g2_fill_1
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_3_604 VPWR VGND sg13g2_decap_8
XFILLER_3_615 VPWR VGND sg13g2_fill_1
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_19_516 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_14_265 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_15_788 VPWR VGND sg13g2_fill_1
Xfanout91 net136 net91 VPWR VGND sg13g2_buf_1
Xfanout80 net88 net80 VPWR VGND sg13g2_buf_1
XFILLER_10_471 VPWR VGND sg13g2_decap_8
XFILLER_10_493 VPWR VGND sg13g2_decap_4
XFILLER_6_431 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_2_692 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_1_clk clknet_2_1__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_1301_ _0737_ net115 _0419_ _0420_ VPWR VGND sg13g2_a21o_1
X_1232_ net146 VPWR _0882_ VGND net99 state\[19\] sg13g2_o21ai_1
XFILLER_18_593 VPWR VGND sg13g2_decap_8
XFILLER_37_357 VPWR VGND sg13g2_decap_8
X_1163_ _0129_ _0829_ _0830_ net38 _0702_ VPWR VGND sg13g2_a22oi_1
X_1094_ VPWR _0763_ daisychain\[62\] VGND sg13g2_inv_1
XFILLER_20_224 VPWR VGND sg13g2_decap_8
X_1996_ net222 VGND VPWR _0328_ state\[72\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_0947_ VPWR _0062_ state\[40\] VGND sg13g2_inv_1
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_11_235 VPWR VGND sg13g2_decap_8
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_7_217 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_2_1__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_19_302 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_229 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_30_500 VPWR VGND sg13g2_fill_1
XFILLER_30_511 VPWR VGND sg13g2_fill_1
XFILLER_42_371 VPWR VGND sg13g2_decap_8
X_1850_ net211 VGND VPWR _0182_ daisychain\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1781_ _0651_ VPWR _0369_ VGND net150 _0015_ sg13g2_o21ai_1
XFILLER_37_154 VPWR VGND sg13g2_decap_8
X_1215_ _0142_ _0868_ _0869_ net30 _0715_ VPWR VGND sg13g2_a22oi_1
X_1146_ VPWR _0815_ daisychain\[114\] VGND sg13g2_inv_1
XFILLER_25_349 VPWR VGND sg13g2_decap_4
XFILLER_40_308 VPWR VGND sg13g2_decap_8
X_1077_ VPWR _0746_ daisychain\[45\] VGND sg13g2_inv_1
X_1979_ net209 VGND VPWR _0311_ state\[55\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_34 VPWR VGND sg13g2_decap_8
XFILLER_16_349 VPWR VGND sg13g2_decap_8
XFILLER_28_165 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[2\].u.inv2 VPWR digitalen.g\[2\].u.OUTP digitalen.g\[2\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_12_588 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_decap_8
XFILLER_4_732 VPWR VGND sg13g2_fill_1
XFILLER_19_132 VPWR VGND sg13g2_decap_8
XFILLER_20_8 VPWR VGND sg13g2_fill_1
XFILLER_47_441 VPWR VGND sg13g2_decap_8
X_1000_ VPWR _0120_ state\[93\] VGND sg13g2_inv_1
XFILLER_34_168 VPWR VGND sg13g2_decap_8
XFILLER_35_636 VPWR VGND sg13g2_decap_8
X_1902_ net203 VGND VPWR _0234_ daisychain\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1833_ net207 VGND VPWR _0165_ daisychain\[37\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1764_ _0600_ VPWR _0352_ VGND net154 _0123_ sg13g2_o21ai_1
X_1695_ _0393_ VPWR _0283_ VGND net146 _0047_ sg13g2_o21ai_1
XFILLER_25_124 VPWR VGND sg13g2_decap_8
XFILLER_38_496 VPWR VGND sg13g2_fill_1
X_1129_ VPWR _0798_ daisychain\[97\] VGND sg13g2_inv_1
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_69 VPWR VGND sg13g2_decap_8
XFILLER_21_363 VPWR VGND sg13g2_fill_1
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_41_639 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_16_146 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_12_363 VPWR VGND sg13g2_decap_8
XFILLER_40_650 VPWR VGND sg13g2_fill_2
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_8_389 VPWR VGND sg13g2_decap_8
X_1480_ net170 VPWR _0554_ VGND net123 state\[81\] sg13g2_o21ai_1
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_39_238 VPWR VGND sg13g2_decap_8
X_2032_ net197 VGND VPWR _0364_ state\[108\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_138 VPWR VGND sg13g2_decap_8
XFILLER_30_193 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
X_1816_ net188 VGND VPWR _0148_ daisychain\[20\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1747_ _0549_ VPWR _0335_ VGND net175 _0104_ sg13g2_o21ai_1
X_1678_ _0856_ VPWR _0266_ VGND net140 _0011_ sg13g2_o21ai_1
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_fill_2
XFILLER_26_466 VPWR VGND sg13g2_decap_8
XFILLER_26_477 VPWR VGND sg13g2_fill_2
XFILLER_26_68 VPWR VGND sg13g2_fill_2
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_17_433 VPWR VGND sg13g2_fill_2
XFILLER_29_293 VPWR VGND sg13g2_decap_8
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_12_160 VPWR VGND sg13g2_decap_8
XFILLER_16_90 VPWR VGND sg13g2_decap_8
XFILLER_32_414 VPWR VGND sg13g2_fill_2
XFILLER_44_252 VPWR VGND sg13g2_decap_8
X_0980_ VPWR _0098_ state\[73\] VGND sg13g2_inv_1
XFILLER_8_186 VPWR VGND sg13g2_decap_8
X_1601_ _0812_ net106 _0644_ _0645_ VPWR VGND sg13g2_a21o_1
X_1532_ net154 VPWR _0593_ VGND net108 state\[94\] sg13g2_o21ai_1
XFILLER_9_698 VPWR VGND sg13g2_fill_2
XFILLER_9_676 VPWR VGND sg13g2_fill_2
X_1463_ _0204_ _0540_ _0541_ net63 _0777_ VPWR VGND sg13g2_a22oi_1
X_1394_ VGND VPWR net82 daisychain\[58\] _0490_ net52 sg13g2_a21oi_1
XFILLER_35_252 VPWR VGND sg13g2_decap_8
X_2015_ net218 VGND VPWR _0347_ state\[91\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_12_48 VPWR VGND sg13g2_decap_8
XFILLER_19_709 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_26_263 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_42_712 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_6_635 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_17_230 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_4
XFILLER_18_797 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_45_594 VPWR VGND sg13g2_decap_8
XFILLER_20_417 VPWR VGND sg13g2_decap_4
XFILLER_32_277 VPWR VGND sg13g2_decap_8
XFILLER_33_767 VPWR VGND sg13g2_decap_8
X_0963_ VPWR _0079_ state\[56\] VGND sg13g2_inv_1
XFILLER_4_60 VPWR VGND sg13g2_decap_8
X_1515_ _0217_ _0579_ _0580_ net41 _0790_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_506 VPWR VGND sg13g2_fill_1
X_1446_ VGND VPWR net86 daisychain\[71\] _0529_ net63 sg13g2_a21oi_1
X_1377_ _0756_ net119 _0476_ _0477_ VPWR VGND sg13g2_a21o_1
XFILLER_11_417 VPWR VGND sg13g2_decap_8
XFILLER_23_233 VPWR VGND sg13g2_decap_8
XFILLER_36_550 VPWR VGND sg13g2_decap_8
XFILLER_23_58 VPWR VGND sg13g2_decap_4
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_15_712 VPWR VGND sg13g2_decap_4
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_14_244 VPWR VGND sg13g2_decap_8
XFILLER_6_410 VPWR VGND sg13g2_decap_8
Xfanout92 net93 net92 VPWR VGND sg13g2_buf_1
Xfanout81 net83 net81 VPWR VGND sg13g2_buf_1
Xfanout70 net89 net70 VPWR VGND sg13g2_buf_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_6_487 VPWR VGND sg13g2_decap_8
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
X_1300_ net161 VPWR _0419_ VGND net115 state\[36\] sg13g2_o21ai_1
X_1231_ _0146_ _0880_ _0881_ net32 _0719_ VPWR VGND sg13g2_a22oi_1
X_1162_ VGND VPWR net75 daisychain\[0\] _0830_ net37 sg13g2_a21oi_1
XFILLER_20_203 VPWR VGND sg13g2_decap_8
X_1093_ VPWR _0762_ daisychain\[61\] VGND sg13g2_inv_1
X_1995_ net222 VGND VPWR _0327_ state\[71\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_0946_ VPWR _0060_ state\[39\] VGND sg13g2_inv_1
XFILLER_9_270 VPWR VGND sg13g2_decap_8
X_1429_ _0769_ net131 _0515_ _0516_ VPWR VGND sg13g2_a21o_1
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_28_358 VPWR VGND sg13g2_decap_4
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_2_3__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_20_792 VPWR VGND sg13g2_decap_8
XFILLER_3_413 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_15_586 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_decap_8
X_1780_ _0648_ VPWR _0368_ VGND net150 _0014_ sg13g2_o21ai_1
XFILLER_6_284 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_38_656 VPWR VGND sg13g2_decap_8
XFILLER_38_667 VPWR VGND sg13g2_fill_1
X_1214_ VGND VPWR net74 daisychain\[13\] _0869_ net30 sg13g2_a21oi_1
X_1145_ VPWR _0814_ daisychain\[113\] VGND sg13g2_inv_1
XFILLER_33_361 VPWR VGND sg13g2_decap_8
X_1076_ VPWR _0745_ daisychain\[44\] VGND sg13g2_inv_1
XFILLER_20_48 VPWR VGND sg13g2_decap_8
X_1978_ net210 VGND VPWR _0310_ state\[54\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_0929_ VPWR _0042_ state\[22\] VGND sg13g2_inv_1
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_13 VPWR VGND sg13g2_decap_8
XFILLER_16_328 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_44_648 VPWR VGND sg13g2_fill_2
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_8_505 VPWR VGND sg13g2_decap_8
XFILLER_8_527 VPWR VGND sg13g2_decap_4
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_3_210 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_8
XFILLER_19_111 VPWR VGND sg13g2_decap_8
XFILLER_19_188 VPWR VGND sg13g2_decap_8
XFILLER_19_90 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_34_147 VPWR VGND sg13g2_decap_8
XFILLER_43_670 VPWR VGND sg13g2_decap_8
X_1901_ net199 VGND VPWR _0233_ daisychain\[105\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1832_ net207 VGND VPWR _0164_ daisychain\[36\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1763_ _0597_ VPWR _0351_ VGND net155 _0122_ sg13g2_o21ai_1
X_1694_ _0390_ VPWR _0282_ VGND net149 _0046_ sg13g2_o21ai_1
XFILLER_15_48 VPWR VGND sg13g2_decap_8
XFILLER_38_453 VPWR VGND sg13g2_decap_8
XFILLER_38_464 VPWR VGND sg13g2_fill_2
X_1128_ VPWR _0797_ daisychain\[96\] VGND sg13g2_inv_1
X_1059_ VPWR _0728_ daisychain\[27\] VGND sg13g2_inv_1
XFILLER_5_508 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_31_69 VPWR VGND sg13g2_decap_8
Xoutput14 net14 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_17_604 VPWR VGND sg13g2_decap_4
XFILLER_29_464 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_12_342 VPWR VGND sg13g2_decap_8
XFILLER_16_125 VPWR VGND sg13g2_decap_8
XFILLER_17_648 VPWR VGND sg13g2_fill_2
XFILLER_24_191 VPWR VGND sg13g2_decap_8
XFILLER_31_139 VPWR VGND sg13g2_decap_8
XFILLER_40_662 VPWR VGND sg13g2_decap_8
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
X_2031_ net199 VGND VPWR _0363_ state\[107\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_30_172 VPWR VGND sg13g2_decap_8
XFILLER_31_640 VPWR VGND sg13g2_decap_8
X_1815_ net191 VGND VPWR _0147_ daisychain\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1746_ _0546_ VPWR _0334_ VGND net175 _0103_ sg13g2_o21ai_1
X_1677_ _0853_ VPWR _0265_ VGND net139 _0127_ sg13g2_o21ai_1
XFILLER_26_401 VPWR VGND sg13g2_decap_8
XFILLER_14_629 VPWR VGND sg13g2_fill_2
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_21_194 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_1_599 VPWR VGND sg13g2_fill_2
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_17_456 VPWR VGND sg13g2_decap_4
XFILLER_29_272 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
X_1600_ net151 VPWR _0644_ VGND net105 state\[111\] sg13g2_o21ai_1
X_1531_ _0221_ _0591_ _0592_ net57 _0794_ VPWR VGND sg13g2_a22oi_1
X_1462_ VGND VPWR net86 daisychain\[75\] _0541_ net63 sg13g2_a21oi_1
XFILLER_48_581 VPWR VGND sg13g2_fill_1
X_1393_ _0760_ net118 _0488_ _0489_ VPWR VGND sg13g2_a21o_1
XFILLER_35_231 VPWR VGND sg13g2_decap_8
X_2014_ net218 VGND VPWR _0346_ state\[90\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_12_27 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_2_319 VPWR VGND sg13g2_decap_8
X_1729_ _0495_ VPWR _0317_ VGND net168 _0085_ sg13g2_o21ai_1
XFILLER_26_242 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_10_643 VPWR VGND sg13g2_decap_4
XFILLER_10_654 VPWR VGND sg13g2_fill_1
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_42_768 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_17_286 VPWR VGND sg13g2_decap_8
XFILLER_18_776 VPWR VGND sg13g2_fill_1
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_33_746 VPWR VGND sg13g2_decap_4
XFILLER_13_492 VPWR VGND sg13g2_decap_8
X_0962_ VPWR _0078_ state\[55\] VGND sg13g2_inv_1
XFILLER_9_463 VPWR VGND sg13g2_fill_1
XFILLER_9_452 VPWR VGND sg13g2_decap_8
X_1514_ VGND VPWR net76 daisychain\[88\] _0580_ net41 sg13g2_a21oi_1
X_1445_ _0773_ net130 _0527_ _0528_ VPWR VGND sg13g2_a21o_1
X_1376_ net164 VPWR _0476_ VGND net117 state\[55\] sg13g2_o21ai_1
XFILLER_23_212 VPWR VGND sg13g2_decap_8
XFILLER_23_289 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_14_223 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_30_727 VPWR VGND sg13g2_decap_8
XFILLER_42_587 VPWR VGND sg13g2_decap_8
Xfanout93 net95 net93 VPWR VGND sg13g2_buf_1
Xfanout82 net83 net82 VPWR VGND sg13g2_buf_1
Xfanout71 net74 net71 VPWR VGND sg13g2_buf_1
Xfanout60 net66 net60 VPWR VGND sg13g2_buf_1
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_4
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
X_1230_ VGND VPWR net71 daisychain\[17\] _0881_ net32 sg13g2_a21oi_1
X_1161_ _0702_ net97 _0828_ _0829_ VPWR VGND sg13g2_a21o_1
X_1092_ VPWR _0761_ daisychain\[60\] VGND sg13g2_inv_1
XFILLER_33_532 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
X_1994_ net222 VGND VPWR _0326_ state\[70\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_20_259 VPWR VGND sg13g2_decap_8
X_0945_ VPWR _0059_ state\[38\] VGND sg13g2_inv_1
XFILLER_0_609 VPWR VGND sg13g2_decap_4
X_1428_ net178 VPWR _0515_ VGND net131 state\[68\] sg13g2_o21ai_1
XFILLER_28_326 VPWR VGND sg13g2_fill_1
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
X_1359_ _0178_ _0462_ _0463_ net54 _0751_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_760 VPWR VGND sg13g2_decap_4
Xclkload2 clknet_leaf_9_clk clkload2/Y VPWR VGND sg13g2_inv_4
XFILLER_3_469 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_15_510 VPWR VGND sg13g2_fill_1
XFILLER_34_329 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_30_579 VPWR VGND sg13g2_fill_1
XFILLER_6_263 VPWR VGND sg13g2_decap_8
XFILLER_2_480 VPWR VGND sg13g2_decap_8
X_1213_ _0715_ net97 _0867_ _0868_ VPWR VGND sg13g2_a21o_1
XFILLER_18_392 VPWR VGND sg13g2_fill_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_25_307 VPWR VGND sg13g2_fill_2
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_38_679 VPWR VGND sg13g2_fill_1
X_1144_ VPWR _0813_ daisychain\[112\] VGND sg13g2_inv_1
X_1075_ VPWR _0744_ daisychain\[43\] VGND sg13g2_inv_1
XFILLER_33_340 VPWR VGND sg13g2_decap_8
X_1977_ net210 VGND VPWR _0309_ state\[53\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_20_27 VPWR VGND sg13g2_decap_8
X_0928_ VPWR _0041_ state\[21\] VGND sg13g2_inv_1
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_29_69 VPWR VGND sg13g2_decap_8
XFILLER_16_307 VPWR VGND sg13g2_decap_8
XFILLER_24_395 VPWR VGND sg13g2_fill_1
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_3_266 VPWR VGND sg13g2_decap_8
XFILLER_4_778 VPWR VGND sg13g2_decap_4
XFILLER_19_167 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_decap_8
XFILLER_35_605 VPWR VGND sg13g2_fill_1
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_15_384 VPWR VGND sg13g2_decap_8
XFILLER_30_354 VPWR VGND sg13g2_decap_8
XFILLER_31_822 VPWR VGND sg13g2_fill_1
X_1900_ net199 VGND VPWR _0232_ daisychain\[104\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1831_ net194 VGND VPWR _0163_ daisychain\[35\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1762_ _0594_ VPWR _0350_ VGND net155 _0121_ sg13g2_o21ai_1
X_1693_ _0387_ VPWR _0281_ VGND net148 _0045_ sg13g2_o21ai_1
XFILLER_25_0 VPWR VGND sg13g2_fill_1
XFILLER_38_432 VPWR VGND sg13g2_decap_8
XFILLER_15_27 VPWR VGND sg13g2_decap_8
XFILLER_21_321 VPWR VGND sg13g2_decap_8
XFILLER_25_159 VPWR VGND sg13g2_decap_8
XFILLER_34_693 VPWR VGND sg13g2_decap_8
X_1127_ VPWR _0796_ daisychain\[95\] VGND sg13g2_inv_1
X_1058_ VPWR _0727_ daisychain\[26\] VGND sg13g2_inv_1
XFILLER_21_398 VPWR VGND sg13g2_fill_2
XFILLER_31_48 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_16_104 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_12_321 VPWR VGND sg13g2_decap_8
XFILLER_13_822 VPWR VGND sg13g2_fill_1
XFILLER_24_170 VPWR VGND sg13g2_decap_8
XFILLER_31_118 VPWR VGND sg13g2_decap_8
XFILLER_12_398 VPWR VGND sg13g2_decap_8
XFILLER_4_586 VPWR VGND sg13g2_fill_1
XFILLER_8_347 VPWR VGND sg13g2_decap_8
X_2030_ net203 VGND VPWR _0362_ state\[106\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_35_435 VPWR VGND sg13g2_fill_1
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_15_181 VPWR VGND sg13g2_decap_8
XFILLER_30_151 VPWR VGND sg13g2_decap_8
XFILLER_31_696 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
X_1814_ net190 VGND VPWR _0146_ daisychain\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1745_ _0543_ VPWR _0333_ VGND net175 _0102_ sg13g2_o21ai_1
X_1676_ _0850_ VPWR _0264_ VGND net139 _0116_ sg13g2_o21ai_1
XFILLER_26_446 VPWR VGND sg13g2_fill_2
XFILLER_38_273 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_21_173 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_402 VPWR VGND sg13g2_fill_1
XFILLER_17_424 VPWR VGND sg13g2_fill_2
XFILLER_29_251 VPWR VGND sg13g2_decap_8
XFILLER_32_427 VPWR VGND sg13g2_fill_1
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_12_195 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
XFILLER_4_361 VPWR VGND sg13g2_decap_8
X_1530_ VGND VPWR net84 daisychain\[92\] _0592_ net57 sg13g2_a21oi_1
X_1461_ _0777_ net130 _0539_ _0540_ VPWR VGND sg13g2_a21o_1
X_1392_ net165 VPWR _0488_ VGND net118 state\[59\] sg13g2_o21ai_1
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_36_722 VPWR VGND sg13g2_decap_4
XFILLER_48_560 VPWR VGND sg13g2_decap_8
X_2013_ net202 VGND VPWR _0345_ state\[89\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_35_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_2_0__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_1728_ _0492_ VPWR _0316_ VGND net165 _0084_ sg13g2_o21ai_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
X_1659_ _0253_ _0687_ _0688_ net24 _0697_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_405 VPWR VGND sg13g2_decap_8
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_fill_2
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_10_600 VPWR VGND sg13g2_fill_2
XFILLER_2_821 VPWR VGND sg13g2_fill_2
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_18_700 VPWR VGND sg13g2_decap_4
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_17_265 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
X_0961_ VPWR _0077_ state\[54\] VGND sg13g2_inv_1
XFILLER_9_431 VPWR VGND sg13g2_decap_8
XFILLER_4_95 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_4_clk clknet_2_3__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_1513_ _0790_ net108 _0578_ _0579_ VPWR VGND sg13g2_a21o_1
X_1444_ net179 VPWR _0527_ VGND net132 state\[72\] sg13g2_o21ai_1
X_1375_ _0182_ _0474_ _0475_ net50 _0755_ VPWR VGND sg13g2_a22oi_1
XFILLER_23_268 VPWR VGND sg13g2_decap_8
XFILLER_23_27 VPWR VGND sg13g2_fill_2
XFILLER_3_629 VPWR VGND sg13g2_fill_2
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_14_202 VPWR VGND sg13g2_decap_8
XFILLER_14_279 VPWR VGND sg13g2_decap_8
XFILLER_15_747 VPWR VGND sg13g2_fill_2
XFILLER_42_511 VPWR VGND sg13g2_fill_1
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_4
XFILLER_10_485 VPWR VGND sg13g2_fill_2
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_6_445 VPWR VGND sg13g2_decap_8
Xfanout94 net95 net94 VPWR VGND sg13g2_buf_1
Xfanout83 net88 net83 VPWR VGND sg13g2_buf_1
Xfanout72 net73 net72 VPWR VGND sg13g2_buf_1
Xfanout61 net66 net61 VPWR VGND sg13g2_buf_1
Xfanout50 net53 net50 VPWR VGND sg13g2_buf_1
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_2_651 VPWR VGND sg13g2_fill_1
XFILLER_2_662 VPWR VGND sg13g2_fill_2
XFILLER_18_563 VPWR VGND sg13g2_decap_4
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
X_1160_ net143 VPWR _0828_ VGND net97 state\[1\] sg13g2_o21ai_1
X_1091_ VPWR _0760_ daisychain\[59\] VGND sg13g2_inv_1
XFILLER_20_238 VPWR VGND sg13g2_decap_8
X_1993_ net222 VGND VPWR _0325_ state\[69\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_0944_ VPWR _0058_ state\[37\] VGND sg13g2_inv_1
XFILLER_28_305 VPWR VGND sg13g2_decap_8
XFILLER_28_316 VPWR VGND sg13g2_fill_1
XFILLER_28_338 VPWR VGND sg13g2_fill_2
X_1427_ _0195_ _0513_ _0514_ net64 _0768_ VPWR VGND sg13g2_a22oi_1
X_1358_ VGND VPWR net83 daisychain\[49\] _0463_ net54 sg13g2_a21oi_1
XFILLER_12_728 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_43_308 VPWR VGND sg13g2_decap_8
X_1289_ _0734_ net112 _0410_ _0411_ VPWR VGND sg13g2_a21o_1
XFILLER_11_249 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_fill_1
Xclkload3 clkload3/Y clknet_leaf_10_clk VPWR VGND sg13g2_inv_2
XFILLER_3_448 VPWR VGND sg13g2_decap_8
XFILLER_19_316 VPWR VGND sg13g2_decap_8
XFILLER_34_308 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_15_555 VPWR VGND sg13g2_decap_8
XFILLER_15_566 VPWR VGND sg13g2_fill_2
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_30_569 VPWR VGND sg13g2_fill_2
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_11_772 VPWR VGND sg13g2_decap_4
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_38_625 VPWR VGND sg13g2_fill_1
X_1212_ net143 VPWR _0867_ VGND net97 state\[14\] sg13g2_o21ai_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
X_1143_ VPWR _0812_ daisychain\[111\] VGND sg13g2_inv_1
X_1074_ VPWR _0743_ daisychain\[42\] VGND sg13g2_inv_1
X_1976_ net210 VGND VPWR _0308_ state\[52\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_0927_ VPWR _0040_ state\[20\] VGND sg13g2_inv_1
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_29_48 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_8
XFILLER_15_363 VPWR VGND sg13g2_decap_8
XFILLER_19_146 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_30_333 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
X_1830_ net192 VGND VPWR _0162_ daisychain\[34\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1761_ _0591_ VPWR _0349_ VGND net171 _0120_ sg13g2_o21ai_1
XFILLER_3_790 VPWR VGND sg13g2_fill_2
XFILLER_7_562 VPWR VGND sg13g2_decap_4
X_1692_ _0384_ VPWR _0280_ VGND net148 _0044_ sg13g2_o21ai_1
X_1126_ VPWR _0795_ daisychain\[94\] VGND sg13g2_inv_1
XFILLER_25_138 VPWR VGND sg13g2_decap_8
XFILLER_33_193 VPWR VGND sg13g2_decap_8
XFILLER_34_672 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
X_1057_ VPWR _0726_ daisychain\[25\] VGND sg13g2_inv_1
XFILLER_31_27 VPWR VGND sg13g2_decap_8
X_1959_ net194 VGND VPWR _0291_ state\[35\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_29_455 VPWR VGND sg13g2_decap_4
XFILLER_44_469 VPWR VGND sg13g2_decap_8
XFILLER_12_300 VPWR VGND sg13g2_decap_8
XFILLER_12_377 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_4_543 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_48_753 VPWR VGND sg13g2_fill_2
XFILLER_15_160 VPWR VGND sg13g2_decap_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
XFILLER_35_458 VPWR VGND sg13g2_decap_8
XFILLER_35_469 VPWR VGND sg13g2_fill_2
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_7_392 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
X_1813_ net190 VGND VPWR _0145_ daisychain\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1744_ _0540_ VPWR _0332_ VGND net177 _0101_ sg13g2_o21ai_1
X_1675_ _0847_ VPWR _0263_ VGND net139 _0105_ sg13g2_o21ai_1
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_41_406 VPWR VGND sg13g2_decap_8
X_1109_ VPWR _0778_ daisychain\[77\] VGND sg13g2_inv_1
XFILLER_21_152 VPWR VGND sg13g2_decap_8
XFILLER_6_819 VPWR VGND sg13g2_decap_4
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_29_230 VPWR VGND sg13g2_decap_8
XFILLER_45_701 VPWR VGND sg13g2_fill_2
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_12_174 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
X_1460_ net177 VPWR _0539_ VGND net130 state\[76\] sg13g2_o21ai_1
X_1391_ _0186_ _0486_ _0487_ net52 _0759_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_756 VPWR VGND sg13g2_decap_4
XFILLER_36_767 VPWR VGND sg13g2_fill_2
X_2012_ net216 VGND VPWR _0344_ state\[88\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_35_266 VPWR VGND sg13g2_decap_8
X_1727_ _0489_ VPWR _0315_ VGND net165 _0082_ sg13g2_o21ai_1
X_1658_ VGND VPWR net70 daisychain\[124\] _0688_ net23 sg13g2_a21oi_1
X_1589_ _0809_ net105 _0635_ _0636_ VPWR VGND sg13g2_a21o_1
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_39_583 VPWR VGND sg13g2_decap_8
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_10_667 VPWR VGND sg13g2_decap_8
XFILLER_10_678 VPWR VGND sg13g2_fill_2
XFILLER_22_472 VPWR VGND sg13g2_fill_2
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_6_627 VPWR VGND sg13g2_fill_1
XFILLER_6_649 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_17_244 VPWR VGND sg13g2_decap_8
XFILLER_45_553 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_18_789 VPWR VGND sg13g2_fill_2
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_33_726 VPWR VGND sg13g2_fill_2
XFILLER_33_737 VPWR VGND sg13g2_decap_4
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
X_0960_ VPWR _0076_ state\[53\] VGND sg13g2_inv_1
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_5_660 VPWR VGND sg13g2_fill_1
X_1512_ net154 VPWR _0578_ VGND net108 state\[89\] sg13g2_o21ai_1
XFILLER_4_74 VPWR VGND sg13g2_decap_8
X_1443_ _0199_ _0525_ _0526_ net65 _0772_ VPWR VGND sg13g2_a22oi_1
X_1374_ VGND VPWR net81 daisychain\[53\] _0475_ net51 sg13g2_a21oi_1
XFILLER_23_247 VPWR VGND sg13g2_decap_8
XFILLER_36_564 VPWR VGND sg13g2_fill_2
XFILLER_32_792 VPWR VGND sg13g2_fill_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_19_509 VPWR VGND sg13g2_fill_2
XFILLER_14_258 VPWR VGND sg13g2_decap_8
XFILLER_30_718 VPWR VGND sg13g2_decap_4
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_1
Xfanout62 net66 net62 VPWR VGND sg13g2_buf_1
Xfanout51 net53 net51 VPWR VGND sg13g2_buf_1
Xfanout40 net43 net40 VPWR VGND sg13g2_buf_1
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_6_424 VPWR VGND sg13g2_decap_8
Xfanout95 net136 net95 VPWR VGND sg13g2_buf_1
Xfanout84 net85 net84 VPWR VGND sg13g2_buf_1
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_29_8 VPWR VGND sg13g2_fill_1
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_18_553 VPWR VGND sg13g2_fill_2
XFILLER_18_586 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
X_1090_ VPWR _0759_ daisychain\[58\] VGND sg13g2_inv_1
XFILLER_13_291 VPWR VGND sg13g2_decap_8
XFILLER_20_217 VPWR VGND sg13g2_decap_8
X_1992_ net221 VGND VPWR _0324_ state\[68\] clknet_leaf_6_clk sg13g2_dfrbpq_1
Xclkload10 VPWR clkload10/Y clknet_leaf_12_clk VGND sg13g2_inv_1
X_0943_ VPWR _0057_ state\[36\] VGND sg13g2_inv_1
XFILLER_9_284 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
X_1426_ VGND VPWR net86 daisychain\[66\] _0514_ net64 sg13g2_a21oi_1
X_1357_ _0751_ net120 _0461_ _0462_ VPWR VGND sg13g2_a21o_1
X_1288_ net158 VPWR _0410_ VGND net112 state\[33\] sg13g2_o21ai_1
XFILLER_11_228 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_20_751 VPWR VGND sg13g2_decap_4
XFILLER_3_427 VPWR VGND sg13g2_decap_8
Xclkload4 clkload4/Y clknet_leaf_15_clk VPWR VGND sg13g2_inv_2
XFILLER_43_810 VPWR VGND sg13g2_decap_8
XFILLER_43_821 VPWR VGND sg13g2_fill_2
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_30_504 VPWR VGND sg13g2_decap_8
XFILLER_30_559 VPWR VGND sg13g2_decap_8
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_7_700 VPWR VGND sg13g2_fill_1
XFILLER_7_733 VPWR VGND sg13g2_decap_4
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_7_744 VPWR VGND sg13g2_fill_2
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
X_1211_ _0141_ _0865_ _0866_ net30 _0714_ VPWR VGND sg13g2_a22oi_1
X_1142_ VPWR _0811_ daisychain\[110\] VGND sg13g2_inv_1
XFILLER_33_375 VPWR VGND sg13g2_fill_2
XFILLER_34_821 VPWR VGND sg13g2_fill_2
XFILLER_46_681 VPWR VGND sg13g2_decap_4
X_1073_ VPWR _0742_ daisychain\[41\] VGND sg13g2_inv_1
X_1975_ net213 VGND VPWR _0307_ state\[51\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0926_ VPWR _0038_ state\[19\] VGND sg13g2_inv_1
XFILLER_29_27 VPWR VGND sg13g2_decap_8
X_1409_ _0764_ net121 _0500_ _0501_ VPWR VGND sg13g2_a21o_1
XFILLER_28_158 VPWR VGND sg13g2_decap_8
XFILLER_12_559 VPWR VGND sg13g2_decap_4
XFILLER_24_342 VPWR VGND sg13g2_fill_1
XFILLER_20_592 VPWR VGND sg13g2_decap_4
XFILLER_3_224 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_19_125 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_15_342 VPWR VGND sg13g2_decap_8
XFILLER_30_312 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_43_684 VPWR VGND sg13g2_decap_4
X_1760_ _0588_ VPWR _0348_ VGND net171 _0119_ sg13g2_o21ai_1
X_1691_ _0895_ VPWR _0279_ VGND net148 _0043_ sg13g2_o21ai_1
XFILLER_25_117 VPWR VGND sg13g2_decap_8
X_1125_ VPWR _0794_ daisychain\[93\] VGND sg13g2_inv_1
XFILLER_33_172 VPWR VGND sg13g2_decap_8
XFILLER_34_640 VPWR VGND sg13g2_decap_8
X_1056_ VPWR _0725_ daisychain\[24\] VGND sg13g2_inv_1
Xoutput17 net17 uo_out[2] VPWR VGND sg13g2_buf_1
X_1958_ net207 VGND VPWR _0290_ state\[34\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1889_ net201 VGND VPWR _0221_ daisychain\[93\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0909_ VPWR _0050_ state\[2\] VGND sg13g2_inv_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_16_139 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_12_356 VPWR VGND sg13g2_decap_8
XFILLER_40_676 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_21_94 VPWR VGND sg13g2_fill_1
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_0_783 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_31_610 VPWR VGND sg13g2_fill_2
XFILLER_31_687 VPWR VGND sg13g2_decap_4
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_30_186 VPWR VGND sg13g2_decap_8
XFILLER_7_371 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
X_1812_ net190 VGND VPWR _0144_ daisychain\[16\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1743_ _0537_ VPWR _0331_ VGND net177 _0100_ sg13g2_o21ai_1
X_1674_ _0844_ VPWR _0262_ VGND net144 _0094_ sg13g2_o21ai_1
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
XFILLER_34_470 VPWR VGND sg13g2_decap_8
XFILLER_38_231 VPWR VGND sg13g2_decap_8
X_1108_ VPWR _0777_ daisychain\[76\] VGND sg13g2_inv_1
X_1039_ VPWR _0708_ daisychain\[7\] VGND sg13g2_inv_1
XFILLER_21_131 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_17_426 VPWR VGND sg13g2_fill_1
XFILLER_29_286 VPWR VGND sg13g2_decap_8
XFILLER_45_746 VPWR VGND sg13g2_decap_4
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_12_153 VPWR VGND sg13g2_decap_8
XFILLER_16_83 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_9_636 VPWR VGND sg13g2_decap_4
XFILLER_4_396 VPWR VGND sg13g2_decap_8
X_1390_ VGND VPWR net82 daisychain\[57\] _0487_ net52 sg13g2_a21oi_1
XFILLER_35_245 VPWR VGND sg13g2_decap_8
X_2011_ net217 VGND VPWR _0343_ state\[87\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1726_ _0486_ VPWR _0314_ VGND net164 _0081_ sg13g2_o21ai_1
X_1657_ net91 _0697_ _0686_ _0687_ VPWR VGND sg13g2_a21o_1
X_1588_ net151 VPWR _0635_ VGND net105 state\[108\] sg13g2_o21ai_1
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_10_602 VPWR VGND sg13g2_fill_1
XFILLER_26_256 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_42_705 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_17_223 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_18_757 VPWR VGND sg13g2_fill_1
XFILLER_33_716 VPWR VGND sg13g2_fill_1
XFILLER_45_532 VPWR VGND sg13g2_decap_8
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
X_1511_ _0216_ _0576_ _0577_ net57 _0789_ VPWR VGND sg13g2_a22oi_1
X_1442_ VGND VPWR net87 daisychain\[70\] _0526_ net65 sg13g2_a21oi_1
XFILLER_4_53 VPWR VGND sg13g2_decap_8
X_1373_ _0755_ net117 _0473_ _0474_ VPWR VGND sg13g2_a21o_1
XFILLER_23_226 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
X_1709_ _0435_ VPWR _0297_ VGND net159 _0063_ sg13g2_o21ai_1
XFILLER_15_705 VPWR VGND sg13g2_decap_8
XFILLER_15_716 VPWR VGND sg13g2_fill_1
XFILLER_27_543 VPWR VGND sg13g2_fill_1
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_4
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_14_237 VPWR VGND sg13g2_decap_8
XFILLER_15_749 VPWR VGND sg13g2_fill_1
XFILLER_22_292 VPWR VGND sg13g2_decap_8
Xfanout30 net32 net30 VPWR VGND sg13g2_buf_1
Xfanout96 net98 net96 VPWR VGND sg13g2_buf_1
Xfanout85 net88 net85 VPWR VGND sg13g2_buf_1
Xfanout74 net78 net74 VPWR VGND sg13g2_buf_1
Xfanout63 net65 net63 VPWR VGND sg13g2_buf_1
Xfanout52 net53 net52 VPWR VGND sg13g2_buf_1
Xfanout41 net42 net41 VPWR VGND sg13g2_buf_1
XFILLER_10_487 VPWR VGND sg13g2_fill_1
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_6_403 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_2_675 VPWR VGND sg13g2_fill_1
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_13_270 VPWR VGND sg13g2_decap_8
XFILLER_14_771 VPWR VGND sg13g2_decap_8
X_1991_ net221 VGND VPWR _0323_ state\[67\] clknet_leaf_6_clk sg13g2_dfrbpq_1
Xclkload11 VPWR clkload11/Y clknet_leaf_14_clk VGND sg13g2_inv_1
X_0942_ VPWR _0056_ state\[35\] VGND sg13g2_inv_1
XFILLER_9_263 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
X_1425_ _0768_ net131 _0512_ _0513_ VPWR VGND sg13g2_a21o_1
XFILLER_18_18 VPWR VGND sg13g2_decap_8
X_1356_ net167 VPWR _0461_ VGND net120 state\[50\] sg13g2_o21ai_1
X_1287_ _0160_ _0408_ _0409_ net45 _0733_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_207 VPWR VGND sg13g2_decap_8
XFILLER_34_28 VPWR VGND sg13g2_decap_8
Xclkload5 clknet_leaf_16_clk clkload5/X VPWR VGND sg13g2_buf_8
XFILLER_3_406 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
Xfanout220 net223 net220 VPWR VGND sg13g2_buf_1
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_24_50 VPWR VGND sg13g2_fill_2
XFILLER_30_549 VPWR VGND sg13g2_decap_4
XFILLER_6_200 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_6_277 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_8
XFILLER_18_351 VPWR VGND sg13g2_fill_1
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_38_649 VPWR VGND sg13g2_decap_8
X_1210_ VGND VPWR net71 daisychain\[12\] _0866_ net30 sg13g2_a21oi_1
X_1141_ VPWR _0810_ daisychain\[109\] VGND sg13g2_inv_1
X_1072_ VPWR _0741_ daisychain\[40\] VGND sg13g2_inv_1
XFILLER_33_354 VPWR VGND sg13g2_decap_8
X_1974_ net212 VGND VPWR _0306_ state\[50\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0925_ VPWR _0037_ state\[18\] VGND sg13g2_inv_1
X_1408_ net168 VPWR _0500_ VGND net121 state\[63\] sg13g2_o21ai_1
XFILLER_24_310 VPWR VGND sg13g2_fill_2
XFILLER_24_321 VPWR VGND sg13g2_fill_1
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_37_671 VPWR VGND sg13g2_fill_2
XFILLER_37_693 VPWR VGND sg13g2_fill_2
XFILLER_45_49 VPWR VGND sg13g2_decap_8
X_1339_ _0173_ _0447_ _0448_ net51 _0746_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_582 VPWR VGND sg13g2_fill_1
XFILLER_24_387 VPWR VGND sg13g2_fill_2
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_fill_1
XFILLER_16_800 VPWR VGND sg13g2_fill_1
XFILLER_19_104 VPWR VGND sg13g2_decap_8
XFILLER_19_83 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_15_321 VPWR VGND sg13g2_decap_8
XFILLER_15_398 VPWR VGND sg13g2_decap_8
XFILLER_16_811 VPWR VGND sg13g2_decap_8
XFILLER_16_822 VPWR VGND sg13g2_fill_1
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_43_641 VPWR VGND sg13g2_decap_8
XFILLER_11_582 VPWR VGND sg13g2_decap_4
XFILLER_30_368 VPWR VGND sg13g2_fill_2
X_1690_ _0892_ VPWR _0278_ VGND net148 _0042_ sg13g2_o21ai_1
XFILLER_2_291 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_38_413 VPWR VGND sg13g2_fill_1
XFILLER_19_660 VPWR VGND sg13g2_decap_8
XFILLER_19_682 VPWR VGND sg13g2_decap_8
XFILLER_38_446 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
X_1124_ VPWR _0793_ daisychain\[92\] VGND sg13g2_inv_1
X_1055_ VPWR _0724_ daisychain\[23\] VGND sg13g2_inv_1
XFILLER_33_151 VPWR VGND sg13g2_decap_8
XFILLER_34_663 VPWR VGND sg13g2_fill_1
X_1957_ net206 VGND VPWR _0289_ state\[33\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[3] VPWR VGND sg13g2_buf_1
X_1888_ net216 VGND VPWR _0220_ daisychain\[92\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0908_ VPWR _0039_ state\[1\] VGND sg13g2_inv_1
XFILLER_17_608 VPWR VGND sg13g2_fill_2
XFILLER_12_335 VPWR VGND sg13g2_decap_8
XFILLER_16_118 VPWR VGND sg13g2_decap_8
XFILLER_24_184 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_fill_2
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_21_51 VPWR VGND sg13g2_decap_4
XFILLER_40_688 VPWR VGND sg13g2_decap_4
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_16_652 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_15_195 VPWR VGND sg13g2_decap_8
XFILLER_30_165 VPWR VGND sg13g2_decap_8
X_1811_ net188 VGND VPWR _0143_ daisychain\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
X_1742_ _0534_ VPWR _0330_ VGND net177 _0099_ sg13g2_o21ai_1
X_1673_ _0841_ VPWR _0261_ VGND net142 _0083_ sg13g2_o21ai_1
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_21_110 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_4
XFILLER_38_287 VPWR VGND sg13g2_decap_8
X_1107_ VPWR _0776_ daisychain\[75\] VGND sg13g2_inv_1
X_1038_ VPWR _0707_ daisychain\[6\] VGND sg13g2_inv_1
XFILLER_21_187 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_17_449 VPWR VGND sg13g2_decap_8
XFILLER_29_265 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_12_132 VPWR VGND sg13g2_decap_8
XFILLER_13_666 VPWR VGND sg13g2_fill_2
XFILLER_16_62 VPWR VGND sg13g2_decap_8
XFILLER_25_493 VPWR VGND sg13g2_decap_4
XFILLER_40_441 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_5_821 VPWR VGND sg13g2_fill_2
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
X_2010_ net223 VGND VPWR _0342_ state\[86\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_16_493 VPWR VGND sg13g2_decap_8
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_8_681 VPWR VGND sg13g2_fill_1
X_1725_ _0483_ VPWR _0313_ VGND net164 _0080_ sg13g2_o21ai_1
Xclkbuf_leaf_7_clk clknet_2_3__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_1656_ net137 VPWR _0686_ VGND state\[125\] net91 sg13g2_o21ai_1
X_1587_ _0235_ _0633_ _0634_ net38 _0808_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_235 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_10_614 VPWR VGND sg13g2_fill_2
XFILLER_14_419 VPWR VGND sg13g2_decap_4
XFILLER_35_780 VPWR VGND sg13g2_fill_2
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_10_647 VPWR VGND sg13g2_fill_1
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_17_202 VPWR VGND sg13g2_decap_8
XFILLER_17_279 VPWR VGND sg13g2_decap_8
XFILLER_18_769 VPWR VGND sg13g2_decap_8
XFILLER_27_72 VPWR VGND sg13g2_fill_2
XFILLER_45_511 VPWR VGND sg13g2_decap_8
XFILLER_13_485 VPWR VGND sg13g2_decap_8
XFILLER_32_249 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_5_651 VPWR VGND sg13g2_decap_8
XFILLER_5_673 VPWR VGND sg13g2_fill_1
X_1510_ VGND VPWR net84 daisychain\[87\] _0577_ net57 sg13g2_a21oi_1
X_1441_ _0772_ net132 _0524_ _0525_ VPWR VGND sg13g2_a21o_1
XFILLER_36_500 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
X_1372_ net164 VPWR _0473_ VGND net117 state\[54\] sg13g2_o21ai_1
XFILLER_17_780 VPWR VGND sg13g2_fill_2
XFILLER_23_205 VPWR VGND sg13g2_decap_8
XFILLER_36_566 VPWR VGND sg13g2_fill_1
XFILLER_36_577 VPWR VGND sg13g2_fill_1
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_31_293 VPWR VGND sg13g2_decap_8
X_1708_ _0432_ VPWR _0296_ VGND net159 _0062_ sg13g2_o21ai_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_1639_ _0248_ _0672_ _0673_ net27 _0821_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_216 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_22_271 VPWR VGND sg13g2_decap_8
Xfanout31 net32 net31 VPWR VGND sg13g2_buf_1
Xfanout97 net98 net97 VPWR VGND sg13g2_buf_1
Xfanout86 net87 net86 VPWR VGND sg13g2_buf_1
Xfanout75 net78 net75 VPWR VGND sg13g2_buf_1
Xfanout64 net65 net64 VPWR VGND sg13g2_buf_1
Xfanout53 net55 net53 VPWR VGND sg13g2_buf_1
Xfanout42 net43 net42 VPWR VGND sg13g2_buf_1
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_18_500 VPWR VGND sg13g2_fill_1
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
XFILLER_33_558 VPWR VGND sg13g2_fill_2
XFILLER_33_569 VPWR VGND sg13g2_decap_4
XFILLER_45_385 VPWR VGND sg13g2_decap_8
X_1990_ net224 VGND VPWR _0322_ state\[66\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_0941_ VPWR _0055_ state\[34\] VGND sg13g2_inv_1
Xclkload12 VPWR clkload12/Y clknet_leaf_6_clk VGND sg13g2_inv_1
XFILLER_9_242 VPWR VGND sg13g2_decap_8
X_1424_ net178 VPWR _0512_ VGND net131 state\[67\] sg13g2_o21ai_1
X_1355_ _0177_ _0459_ _0460_ net54 _0750_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_385 VPWR VGND sg13g2_decap_8
X_1286_ VGND VPWR net79 daisychain\[31\] _0409_ net45 sg13g2_a21oi_1
XFILLER_12_709 VPWR VGND sg13g2_fill_2
XFILLER_20_764 VPWR VGND sg13g2_fill_1
XFILLER_20_775 VPWR VGND sg13g2_fill_2
XFILLER_32_591 VPWR VGND sg13g2_fill_1
Xclkload6 clknet_leaf_0_clk clkload6/Y VPWR VGND sg13g2_inv_4
XFILLER_46_105 VPWR VGND sg13g2_decap_8
Xfanout210 net214 net210 VPWR VGND sg13g2_buf_1
Xfanout221 net223 net221 VPWR VGND sg13g2_buf_1
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_11_731 VPWR VGND sg13g2_decap_8
XFILLER_11_742 VPWR VGND sg13g2_fill_1
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_6_256 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_18_385 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
X_1140_ VPWR _0809_ daisychain\[108\] VGND sg13g2_inv_1
X_1071_ VPWR _0740_ daisychain\[39\] VGND sg13g2_inv_1
XFILLER_14_591 VPWR VGND sg13g2_decap_8
XFILLER_33_333 VPWR VGND sg13g2_decap_8
XFILLER_33_377 VPWR VGND sg13g2_fill_1
XFILLER_45_182 VPWR VGND sg13g2_decap_8
X_1973_ net212 VGND VPWR _0305_ state\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0924_ VPWR _0036_ state\[17\] VGND sg13g2_inv_1
XFILLER_28_116 VPWR VGND sg13g2_decap_8
X_1407_ _0190_ _0498_ _0499_ net55 _0763_ VPWR VGND sg13g2_a22oi_1
X_1338_ VGND VPWR net81 daisychain\[44\] _0448_ net50 sg13g2_a21oi_1
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
X_1269_ _0729_ net100 _0395_ _0396_ VPWR VGND sg13g2_a21o_1
XFILLER_20_572 VPWR VGND sg13g2_fill_2
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_3_259 VPWR VGND sg13g2_decap_8
XFILLER_15_300 VPWR VGND sg13g2_decap_8
XFILLER_19_62 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_43_620 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_15_377 VPWR VGND sg13g2_decap_8
XFILLER_27_193 VPWR VGND sg13g2_decap_8
XFILLER_30_347 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_7_532 VPWR VGND sg13g2_decap_4
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_38_425 VPWR VGND sg13g2_decap_8
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_33_130 VPWR VGND sg13g2_decap_8
XFILLER_34_686 VPWR VGND sg13g2_decap_8
X_1123_ VPWR _0792_ daisychain\[91\] VGND sg13g2_inv_1
X_1054_ VPWR _0723_ daisychain\[22\] VGND sg13g2_inv_1
X_1956_ net206 VGND VPWR _0288_ state\[32\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1887_ net216 VGND VPWR _0219_ daisychain\[91\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0907_ VPWR _0000_ state\[0\] VGND sg13g2_inv_1
Xoutput19 net19 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_44_406 VPWR VGND sg13g2_decap_8
XFILLER_12_314 VPWR VGND sg13g2_decap_8
XFILLER_13_815 VPWR VGND sg13g2_decap_8
XFILLER_24_163 VPWR VGND sg13g2_decap_8
XFILLER_40_612 VPWR VGND sg13g2_decap_8
XFILLER_21_30 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_decap_4
XFILLER_35_428 VPWR VGND sg13g2_decap_4
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_48_789 VPWR VGND sg13g2_fill_1
XFILLER_15_174 VPWR VGND sg13g2_decap_8
XFILLER_30_144 VPWR VGND sg13g2_decap_8
XFILLER_31_612 VPWR VGND sg13g2_fill_1
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
X_1810_ net188 VGND VPWR _0142_ daisychain\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1741_ _0531_ VPWR _0329_ VGND net180 _0098_ sg13g2_o21ai_1
XFILLER_7_98 VPWR VGND sg13g2_decap_8
X_1672_ _0838_ VPWR _0260_ VGND net144 _0072_ sg13g2_o21ai_1
XFILLER_38_266 VPWR VGND sg13g2_decap_8
X_1106_ VPWR _0775_ daisychain\[74\] VGND sg13g2_inv_1
XFILLER_21_100 VPWR VGND sg13g2_fill_1
X_1037_ VPWR _0706_ daisychain\[5\] VGND sg13g2_inv_1
XFILLER_21_166 VPWR VGND sg13g2_decap_8
X_1939_ net188 VGND VPWR _0271_ state\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_16_41 VPWR VGND sg13g2_decap_8
XFILLER_29_244 VPWR VGND sg13g2_decap_8
XFILLER_44_203 VPWR VGND sg13g2_decap_8
XFILLER_12_111 VPWR VGND sg13g2_decap_8
XFILLER_12_188 VPWR VGND sg13g2_decap_8
XFILLER_13_634 VPWR VGND sg13g2_fill_2
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_40_497 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_36_715 VPWR VGND sg13g2_decap_8
XFILLER_36_726 VPWR VGND sg13g2_fill_1
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
X_1724_ _0480_ VPWR _0312_ VGND net163 _0079_ sg13g2_o21ai_1
X_1655_ _0252_ _0684_ _0685_ net24 _0698_ VPWR VGND sg13g2_a22oi_1
X_1586_ VGND VPWR net78 daisychain\[106\] _0634_ net39 sg13g2_a21oi_1
XFILLER_26_214 VPWR VGND sg13g2_decap_8
X_2069_ daisychain\[121\] net16 VPWR VGND sg13g2_buf_1
XFILLER_22_486 VPWR VGND sg13g2_fill_1
XFILLER_22_497 VPWR VGND sg13g2_fill_2
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_2_814 VPWR VGND sg13g2_decap_8
XFILLER_18_704 VPWR VGND sg13g2_fill_2
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_13_431 VPWR VGND sg13g2_decap_4
XFILLER_17_258 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
X_1440_ net179 VPWR _0524_ VGND net132 state\[71\] sg13g2_o21ai_1
X_1371_ _0181_ _0471_ _0472_ net51 _0754_ VPWR VGND sg13g2_a22oi_1
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_31_272 VPWR VGND sg13g2_decap_8
XFILLER_32_740 VPWR VGND sg13g2_fill_2
X_1707_ _0429_ VPWR _0295_ VGND net159 _0060_ sg13g2_o21ai_1
X_1638_ VGND VPWR net69 daisychain\[119\] _0673_ net27 sg13g2_a21oi_1
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_1569_ _0804_ net110 _0620_ _0621_ VPWR VGND sg13g2_a21o_1
XFILLER_42_504 VPWR VGND sg13g2_decap_8
XFILLER_42_559 VPWR VGND sg13g2_fill_2
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_10_478 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_22_250 VPWR VGND sg13g2_decap_8
XFILLER_6_438 VPWR VGND sg13g2_decap_8
Xfanout32 net44 net32 VPWR VGND sg13g2_buf_1
Xfanout98 net111 net98 VPWR VGND sg13g2_buf_1
Xfanout87 net88 net87 VPWR VGND sg13g2_buf_1
Xfanout76 net77 net76 VPWR VGND sg13g2_buf_1
Xfanout65 net66 net65 VPWR VGND sg13g2_buf_1
Xfanout54 net55 net54 VPWR VGND sg13g2_buf_1
Xfanout43 net44 net43 VPWR VGND sg13g2_buf_1
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_2_699 VPWR VGND sg13g2_decap_4
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_decap_8
X_0940_ VPWR _0054_ state\[33\] VGND sg13g2_inv_1
XFILLER_9_221 VPWR VGND sg13g2_decap_8
XFILLER_9_298 VPWR VGND sg13g2_decap_8
X_1423_ _0194_ _0510_ _0511_ net62 _0767_ VPWR VGND sg13g2_a22oi_1
X_1354_ VGND VPWR net83 daisychain\[48\] _0460_ net54 sg13g2_a21oi_1
X_1285_ _0733_ net112 _0407_ _0408_ VPWR VGND sg13g2_a21o_1
XFILLER_24_515 VPWR VGND sg13g2_fill_2
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_20_743 VPWR VGND sg13g2_fill_2
Xclkload7 clkload7/Y clknet_leaf_1_clk VPWR VGND sg13g2_inv_8
Xfanout200 net203 net200 VPWR VGND sg13g2_buf_1
Xfanout211 net214 net211 VPWR VGND sg13g2_buf_1
Xfanout222 net223 net222 VPWR VGND sg13g2_buf_1
XFILLER_19_309 VPWR VGND sg13g2_decap_8
XFILLER_24_52 VPWR VGND sg13g2_fill_1
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_11_765 VPWR VGND sg13g2_decap_8
XFILLER_11_776 VPWR VGND sg13g2_fill_2
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_38_618 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_33_312 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
X_1070_ VPWR _0739_ daisychain\[38\] VGND sg13g2_inv_1
X_1972_ net208 VGND VPWR _0304_ state\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0923_ VPWR _0035_ state\[16\] VGND sg13g2_inv_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_1406_ VGND VPWR net83 daisychain\[61\] _0499_ net54 sg13g2_a21oi_1
X_1337_ _0746_ net119 _0446_ _0447_ VPWR VGND sg13g2_a21o_1
X_1268_ net146 VPWR _0395_ VGND net100 state\[28\] sg13g2_o21ai_1
XFILLER_24_312 VPWR VGND sg13g2_fill_1
XFILLER_24_389 VPWR VGND sg13g2_fill_1
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_40_816 VPWR VGND sg13g2_decap_8
X_1199_ _0138_ _0856_ _0857_ net25 _0711_ VPWR VGND sg13g2_a22oi_1
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_238 VPWR VGND sg13g2_decap_8
XFILLER_19_139 VPWR VGND sg13g2_decap_8
XFILLER_19_41 VPWR VGND sg13g2_decap_8
XFILLER_27_172 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_15_356 VPWR VGND sg13g2_decap_8
XFILLER_30_326 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_decap_8
XFILLER_3_761 VPWR VGND sg13g2_fill_2
XFILLER_7_555 VPWR VGND sg13g2_decap_8
XFILLER_7_566 VPWR VGND sg13g2_fill_1
XFILLER_7_599 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_3_783 VPWR VGND sg13g2_decap_8
X_1122_ VPWR _0791_ daisychain\[90\] VGND sg13g2_inv_1
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_19_695 VPWR VGND sg13g2_fill_1
XFILLER_33_186 VPWR VGND sg13g2_decap_8
XFILLER_34_654 VPWR VGND sg13g2_fill_2
X_1053_ VPWR _0722_ daisychain\[21\] VGND sg13g2_inv_1
X_1955_ net204 VGND VPWR _0287_ state\[31\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1886_ net216 VGND VPWR _0218_ daisychain\[90\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0906_ VPWR _0700_ daisychain\[127\] VGND sg13g2_inv_1
XFILLER_29_448 VPWR VGND sg13g2_fill_2
XFILLER_29_459 VPWR VGND sg13g2_fill_2
XFILLER_37_492 VPWR VGND sg13g2_fill_1
XFILLER_24_142 VPWR VGND sg13g2_decap_8
XFILLER_40_646 VPWR VGND sg13g2_decap_4
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_15_153 VPWR VGND sg13g2_decap_8
XFILLER_16_632 VPWR VGND sg13g2_fill_2
XFILLER_28_492 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_30_123 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
X_1740_ _0528_ VPWR _0328_ VGND net180 _0097_ sg13g2_o21ai_1
X_1671_ _0835_ VPWR _0259_ VGND net147 _0061_ sg13g2_o21ai_1
XFILLER_39_702 VPWR VGND sg13g2_fill_1
XFILLER_7_385 VPWR VGND sg13g2_decap_8
XFILLER_38_245 VPWR VGND sg13g2_decap_8
X_1105_ VPWR _0774_ daisychain\[73\] VGND sg13g2_inv_1
XFILLER_21_145 VPWR VGND sg13g2_decap_8
X_1036_ VPWR _0705_ daisychain\[4\] VGND sg13g2_inv_1
X_1938_ net188 VGND VPWR _0270_ state\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1869_ net220 VGND VPWR _0201_ daisychain\[73\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_29_223 VPWR VGND sg13g2_decap_8
XFILLER_16_20 VPWR VGND sg13g2_decap_8
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_12_167 VPWR VGND sg13g2_decap_8
XFILLER_16_97 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_40_476 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_36_738 VPWR VGND sg13g2_fill_2
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_16_451 VPWR VGND sg13g2_fill_1
XFILLER_16_484 VPWR VGND sg13g2_decap_4
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_fill_1
XFILLER_7_182 VPWR VGND sg13g2_decap_8
XFILLER_8_650 VPWR VGND sg13g2_decap_8
X_1723_ _0477_ VPWR _0311_ VGND net163 _0078_ sg13g2_o21ai_1
X_1654_ VGND VPWR daisychain\[123\] net70 _0685_ net23 sg13g2_a21oi_1
X_1585_ _0808_ net105 _0632_ _0633_ VPWR VGND sg13g2_a21o_1
XFILLER_42_719 VPWR VGND sg13g2_fill_1
X_2068_ daisychain\[120\] net15 VPWR VGND sg13g2_buf_1
X_1019_ VPWR _0014_ state\[112\] VGND sg13g2_inv_1
XFILLER_22_465 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_17_237 VPWR VGND sg13g2_decap_8
XFILLER_45_546 VPWR VGND sg13g2_decap_8
XFILLER_13_410 VPWR VGND sg13g2_decap_8
XFILLER_13_465 VPWR VGND sg13g2_decap_4
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
X_1370_ VGND VPWR net81 daisychain\[52\] _0472_ net51 sg13g2_a21oi_1
XFILLER_36_557 VPWR VGND sg13g2_decap_8
XFILLER_31_251 VPWR VGND sg13g2_decap_8
XFILLER_8_480 VPWR VGND sg13g2_fill_1
XFILLER_8_491 VPWR VGND sg13g2_fill_1
X_1706_ _0426_ VPWR _0294_ VGND net161 _0059_ sg13g2_o21ai_1
X_1637_ _0821_ net94 _0671_ _0672_ VPWR VGND sg13g2_a21o_1
XFILLER_27_524 VPWR VGND sg13g2_fill_2
X_1568_ net153 VPWR _0620_ VGND net110 state\[103\] sg13g2_o21ai_1
X_1499_ _0213_ _0567_ _0568_ net58 _0786_ VPWR VGND sg13g2_a22oi_1
XFILLER_42_516 VPWR VGND sg13g2_fill_2
Xfanout33 net34 net33 VPWR VGND sg13g2_buf_1
Xfanout55 net67 net55 VPWR VGND sg13g2_buf_1
Xfanout44 net67 net44 VPWR VGND sg13g2_buf_1
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_6_417 VPWR VGND sg13g2_decap_8
Xfanout99 net103 net99 VPWR VGND sg13g2_buf_1
Xfanout88 net89 net88 VPWR VGND sg13g2_buf_1
Xfanout77 net78 net77 VPWR VGND sg13g2_buf_1
Xfanout66 net67 net66 VPWR VGND sg13g2_buf_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_601 VPWR VGND sg13g2_fill_1
XFILLER_2_634 VPWR VGND sg13g2_fill_2
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_18_579 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_fill_1
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_14_785 VPWR VGND sg13g2_decap_4
XFILLER_41_560 VPWR VGND sg13g2_fill_1
XFILLER_9_277 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
XFILLER_5_494 VPWR VGND sg13g2_decap_8
X_1422_ VGND VPWR net87 daisychain\[65\] _0511_ net62 sg13g2_a21oi_1
XFILLER_37_822 VPWR VGND sg13g2_fill_1
X_1353_ _0750_ net120 _0458_ _0459_ VPWR VGND sg13g2_a21o_1
X_1284_ net158 VPWR _0407_ VGND net112 state\[32\] sg13g2_o21ai_1
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_20_755 VPWR VGND sg13g2_fill_2
XFILLER_20_777 VPWR VGND sg13g2_fill_1
XFILLER_20_799 VPWR VGND sg13g2_decap_4
XFILLER_32_571 VPWR VGND sg13g2_decap_8
Xclkload8 clkload8/Y clknet_leaf_17_clk VPWR VGND sg13g2_inv_8
X_0999_ VPWR _0119_ state\[92\] VGND sg13g2_inv_1
Xfanout201 net202 net201 VPWR VGND sg13g2_buf_1
Xfanout212 net214 net212 VPWR VGND sg13g2_buf_1
Xfanout223 net224 net223 VPWR VGND sg13g2_buf_1
XFILLER_15_516 VPWR VGND sg13g2_decap_4
XFILLER_27_376 VPWR VGND sg13g2_fill_2
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_7_737 VPWR VGND sg13g2_fill_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_33_368 VPWR VGND sg13g2_decap_8
XFILLER_34_814 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
X_1971_ net208 VGND VPWR _0303_ state\[47\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_0922_ VPWR _0034_ state\[15\] VGND sg13g2_inv_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_5_291 VPWR VGND sg13g2_decap_8
X_1405_ _0763_ net121 _0497_ _0498_ VPWR VGND sg13g2_a21o_1
XFILLER_36_140 VPWR VGND sg13g2_decap_8
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
X_1336_ net163 VPWR _0446_ VGND net119 state\[45\] sg13g2_o21ai_1
X_1267_ _0155_ _0393_ _0394_ net34 _0728_ VPWR VGND sg13g2_a22oi_1
X_1198_ VGND VPWR net68 daisychain\[9\] _0857_ net25 sg13g2_a21oi_1
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_20_574 VPWR VGND sg13g2_fill_1
XFILLER_20_596 VPWR VGND sg13g2_fill_2
XFILLER_3_217 VPWR VGND sg13g2_decap_8
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_19_118 VPWR VGND sg13g2_decap_8
XFILLER_19_20 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_15_335 VPWR VGND sg13g2_decap_8
XFILLER_19_97 VPWR VGND sg13g2_decap_8
XFILLER_27_151 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_decap_8
XFILLER_43_677 VPWR VGND sg13g2_decap_8
XFILLER_30_305 VPWR VGND sg13g2_decap_8
XFILLER_43_688 VPWR VGND sg13g2_fill_1
XFILLER_18_151 VPWR VGND sg13g2_decap_8
X_1121_ VPWR _0790_ daisychain\[89\] VGND sg13g2_inv_1
X_1052_ VPWR _0721_ daisychain\[20\] VGND sg13g2_inv_1
XFILLER_33_165 VPWR VGND sg13g2_decap_8
X_1954_ net204 VGND VPWR _0286_ state\[30\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1885_ net201 VGND VPWR _0217_ daisychain\[89\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0905_ VPWR _0030_ state\[127\] VGND sg13g2_inv_1
XFILLER_40_603 VPWR VGND sg13g2_fill_1
X_1319_ _0168_ _0432_ _0433_ net46 _0741_ VPWR VGND sg13g2_a22oi_1
XFILLER_12_349 VPWR VGND sg13g2_decap_8
XFILLER_24_198 VPWR VGND sg13g2_decap_8
XFILLER_40_669 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_15_132 VPWR VGND sg13g2_decap_8
XFILLER_16_611 VPWR VGND sg13g2_decap_8
XFILLER_16_666 VPWR VGND sg13g2_decap_8
XFILLER_16_699 VPWR VGND sg13g2_decap_4
XFILLER_30_102 VPWR VGND sg13g2_decap_8
XFILLER_31_647 VPWR VGND sg13g2_fill_1
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_11_382 VPWR VGND sg13g2_decap_8
XFILLER_30_179 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_1670_ _0832_ VPWR _0258_ VGND net147 _0050_ sg13g2_o21ai_1
XFILLER_30_4 VPWR VGND sg13g2_decap_4
XFILLER_38_224 VPWR VGND sg13g2_decap_8
X_1104_ VPWR _0773_ daisychain\[72\] VGND sg13g2_inv_1
X_1035_ VPWR _0704_ daisychain\[3\] VGND sg13g2_inv_1
XFILLER_21_124 VPWR VGND sg13g2_decap_8
XFILLER_34_463 VPWR VGND sg13g2_decap_8
X_1937_ net189 VGND VPWR _0269_ state\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
X_1868_ net220 VGND VPWR _0200_ daisychain\[72\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1799_ net188 VGND VPWR _0131_ daisychain\[3\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_29_202 VPWR VGND sg13g2_decap_8
XFILLER_29_279 VPWR VGND sg13g2_decap_8
XFILLER_45_706 VPWR VGND sg13g2_decap_8
XFILLER_16_76 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_12_146 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_40_455 VPWR VGND sg13g2_decap_8
XFILLER_4_312 VPWR VGND sg13g2_decap_8
XFILLER_9_629 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_7_161 VPWR VGND sg13g2_decap_8
X_1722_ _0474_ VPWR _0310_ VGND net165 _0077_ sg13g2_o21ai_1
X_1653_ _0698_ net90 _0683_ _0684_ VPWR VGND sg13g2_a21o_1
X_1584_ net151 VPWR _0632_ VGND net105 state\[107\] sg13g2_o21ai_1
XFILLER_39_500 VPWR VGND sg13g2_decap_8
XFILLER_26_249 VPWR VGND sg13g2_decap_8
X_2067_ state\[127\] net14 VPWR VGND sg13g2_buf_1
X_1018_ VPWR _0013_ state\[111\] VGND sg13g2_inv_1
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_17_216 VPWR VGND sg13g2_decap_8
XFILLER_18_739 VPWR VGND sg13g2_fill_2
XFILLER_33_709 VPWR VGND sg13g2_fill_1
XFILLER_45_525 VPWR VGND sg13g2_decap_8
XFILLER_13_499 VPWR VGND sg13g2_decap_8
XFILLER_25_271 VPWR VGND sg13g2_fill_2
XFILLER_25_293 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_41_786 VPWR VGND sg13g2_fill_2
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_4
XFILLER_5_632 VPWR VGND sg13g2_fill_1
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_16_293 VPWR VGND sg13g2_decap_8
XFILLER_23_219 VPWR VGND sg13g2_decap_8
XFILLER_32_731 VPWR VGND sg13g2_fill_2
XFILLER_32_742 VPWR VGND sg13g2_fill_1
XFILLER_44_580 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_31_230 VPWR VGND sg13g2_decap_8
X_1705_ _0423_ VPWR _0293_ VGND net161 _0058_ sg13g2_o21ai_1
X_1636_ net140 VPWR _0671_ VGND net94 state\[120\] sg13g2_o21ai_1
X_1567_ _0230_ _0618_ _0619_ net56 _0803_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_536 VPWR VGND sg13g2_fill_1
XFILLER_39_385 VPWR VGND sg13g2_decap_8
X_1498_ VGND VPWR net84 daisychain\[84\] _0568_ net58 sg13g2_a21oi_1
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_22_285 VPWR VGND sg13g2_decap_8
Xfanout23 net24 net23 VPWR VGND sg13g2_buf_1
Xfanout34 net36 net34 VPWR VGND sg13g2_buf_1
Xfanout89 _0696_ net89 VPWR VGND sg13g2_buf_1
Xfanout78 net89 net78 VPWR VGND sg13g2_buf_1
Xfanout67 _0826_ net67 VPWR VGND sg13g2_buf_1
Xfanout56 net60 net56 VPWR VGND sg13g2_buf_1
Xfanout45 net47 net45 VPWR VGND sg13g2_buf_1
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_14_764 VPWR VGND sg13g2_decap_8
XFILLER_9_256 VPWR VGND sg13g2_decap_8
XFILLER_5_473 VPWR VGND sg13g2_decap_8
X_1421_ _0767_ net129 _0509_ _0510_ VPWR VGND sg13g2_a21o_1
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_49_650 VPWR VGND sg13g2_decap_8
XFILLER_49_694 VPWR VGND sg13g2_fill_2
X_1352_ net167 VPWR _0458_ VGND net120 state\[49\] sg13g2_o21ai_1
X_1283_ _0159_ _0405_ _0406_ net45 _0732_ VPWR VGND sg13g2_a22oi_1
XFILLER_17_591 VPWR VGND sg13g2_decap_8
XFILLER_36_399 VPWR VGND sg13g2_decap_8
Xclkload9 clkload9/Y clknet_leaf_8_clk VPWR VGND sg13g2_inv_2
X_0998_ VPWR _0118_ state\[91\] VGND sg13g2_inv_1
Xfanout202 net203 net202 VPWR VGND sg13g2_buf_1
Xfanout213 net214 net213 VPWR VGND sg13g2_buf_1
Xfanout224 net225 net224 VPWR VGND sg13g2_buf_1
X_1619_ _0243_ _0657_ _0658_ net38 _0816_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_24_43 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_46_653 VPWR VGND sg13g2_decap_4
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_33_347 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
X_1970_ net212 VGND VPWR _0302_ state\[46\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0921_ VPWR _0033_ state\[14\] VGND sg13g2_inv_1
XFILLER_6_760 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_8
XFILLER_6_793 VPWR VGND sg13g2_fill_1
X_1404_ net167 VPWR _0497_ VGND net121 state\[62\] sg13g2_o21ai_1
X_1335_ _0172_ _0444_ _0445_ net50 _0745_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_303 VPWR VGND sg13g2_decap_8
XFILLER_24_325 VPWR VGND sg13g2_decap_4
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_49_480 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_1266_ VGND VPWR net72 daisychain\[26\] _0394_ net34 sg13g2_a21oi_1
X_1197_ _0711_ net92 _0855_ _0856_ VPWR VGND sg13g2_a21o_1
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_19_76 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_15_314 VPWR VGND sg13g2_decap_8
XFILLER_31_818 VPWR VGND sg13g2_decap_4
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_43_634 VPWR VGND sg13g2_fill_2
XFILLER_11_586 VPWR VGND sg13g2_fill_2
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_3_763 VPWR VGND sg13g2_fill_1
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_19_653 VPWR VGND sg13g2_decap_8
XFILLER_19_675 VPWR VGND sg13g2_decap_8
XFILLER_34_601 VPWR VGND sg13g2_fill_1
XFILLER_38_406 VPWR VGND sg13g2_decap_8
XFILLER_38_439 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
X_1120_ VPWR _0789_ daisychain\[88\] VGND sg13g2_inv_1
X_1051_ VPWR _0720_ daisychain\[19\] VGND sg13g2_inv_1
XFILLER_14_391 VPWR VGND sg13g2_decap_8
XFILLER_21_328 VPWR VGND sg13g2_fill_1
XFILLER_33_144 VPWR VGND sg13g2_decap_8
XFILLER_34_656 VPWR VGND sg13g2_fill_1
X_1953_ net192 VGND VPWR _0285_ state\[29\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1884_ net201 VGND VPWR _0216_ daisychain\[88\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0904_ VPWR _0699_ daisychain\[126\] VGND sg13g2_inv_1
X_1318_ VGND VPWR net79 daisychain\[39\] _0433_ net46 sg13g2_a21oi_1
XFILLER_24_177 VPWR VGND sg13g2_decap_8
XFILLER_37_461 VPWR VGND sg13g2_decap_8
XFILLER_40_626 VPWR VGND sg13g2_fill_1
X_1249_ _0724_ net102 _0894_ _0895_ VPWR VGND sg13g2_a21o_1
XFILLER_12_328 VPWR VGND sg13g2_decap_8
XFILLER_20_383 VPWR VGND sg13g2_fill_2
XFILLER_21_44 VPWR VGND sg13g2_decap_8
XFILLER_21_55 VPWR VGND sg13g2_fill_1
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_15_111 VPWR VGND sg13g2_decap_8
XFILLER_15_188 VPWR VGND sg13g2_decap_8
XFILLER_30_158 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_fill_1
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_3_560 VPWR VGND sg13g2_decap_8
XFILLER_19_494 VPWR VGND sg13g2_decap_8
XFILLER_34_431 VPWR VGND sg13g2_fill_1
XFILLER_46_280 VPWR VGND sg13g2_decap_8
X_1103_ VPWR _0772_ daisychain\[71\] VGND sg13g2_inv_1
X_1034_ VPWR _0703_ daisychain\[2\] VGND sg13g2_inv_1
X_1936_ net189 VGND VPWR _0268_ state\[12\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1867_ net220 VGND VPWR _0199_ daisychain\[71\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1798_ net197 VGND VPWR _0130_ daisychain\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_29_258 VPWR VGND sg13g2_decap_8
XFILLER_44_217 VPWR VGND sg13g2_decap_8
XFILLER_12_125 VPWR VGND sg13g2_decap_8
XFILLER_13_659 VPWR VGND sg13g2_decap_8
XFILLER_16_55 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_5_814 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_28_291 VPWR VGND sg13g2_decap_8
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_36_707 VPWR VGND sg13g2_decap_4
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
X_1721_ _0471_ VPWR _0309_ VGND net166 _0076_ sg13g2_o21ai_1
X_1652_ net138 VPWR _0683_ VGND net90 state\[124\] sg13g2_o21ai_1
X_1583_ _0234_ _0630_ _0631_ net39 _0807_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_228 VPWR VGND sg13g2_decap_8
XFILLER_22_401 VPWR VGND sg13g2_decap_4
XFILLER_34_294 VPWR VGND sg13g2_decap_8
XFILLER_35_773 VPWR VGND sg13g2_decap_8
X_2066_ state\[126\] net13 VPWR VGND sg13g2_buf_1
X_1017_ VPWR _0012_ state\[110\] VGND sg13g2_inv_1
X_1919_ net183 VGND VPWR _0251_ daisychain\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_25_250 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_45_504 VPWR VGND sg13g2_decap_8
XFILLER_13_478 VPWR VGND sg13g2_decap_8
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_41_721 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_5_622 VPWR VGND sg13g2_fill_1
XFILLER_5_644 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_16_272 VPWR VGND sg13g2_decap_8
XFILLER_44_592 VPWR VGND sg13g2_decap_8
XFILLER_31_286 VPWR VGND sg13g2_decap_8
XFILLER_32_798 VPWR VGND sg13g2_fill_1
X_1704_ _0420_ VPWR _0292_ VGND net161 _0057_ sg13g2_o21ai_1
X_1635_ _0247_ _0669_ _0670_ net27 _0820_ VPWR VGND sg13g2_a22oi_1
X_1566_ VGND VPWR net85 daisychain\[101\] _0619_ net56 sg13g2_a21oi_1
X_1497_ _0786_ net125 _0566_ _0567_ VPWR VGND sg13g2_a21o_1
XFILLER_14_209 VPWR VGND sg13g2_decap_8
XFILLER_39_364 VPWR VGND sg13g2_decap_8
XFILLER_42_518 VPWR VGND sg13g2_fill_1
X_2049_ net184 VGND VPWR _0381_ state\[125\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_22_264 VPWR VGND sg13g2_decap_8
XFILLER_35_581 VPWR VGND sg13g2_decap_8
Xfanout24 net29 net24 VPWR VGND sg13g2_buf_1
Xfanout79 net80 net79 VPWR VGND sg13g2_buf_1
Xfanout68 net89 net68 VPWR VGND sg13g2_buf_1
Xfanout57 net59 net57 VPWR VGND sg13g2_buf_1
Xfanout46 net47 net46 VPWR VGND sg13g2_buf_1
Xfanout35 net36 net35 VPWR VGND sg13g2_buf_1
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_14_732 VPWR VGND sg13g2_decap_8
XFILLER_33_518 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[1\].u.inv1 VPWR digitalen.g\[1\].u.OUTN net6 VGND sg13g2_inv_1
X_1420_ net176 VPWR _0509_ VGND net129 state\[66\] sg13g2_o21ai_1
X_1351_ _0176_ _0456_ _0457_ net49 _0749_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
X_1282_ VGND VPWR net79 daisychain\[30\] _0406_ net45 sg13g2_a21oi_1
XFILLER_20_768 VPWR VGND sg13g2_decap_8
XFILLER_32_540 VPWR VGND sg13g2_decap_8
XFILLER_32_551 VPWR VGND sg13g2_fill_1
X_1618_ VGND VPWR net75 daisychain\[114\] _0658_ net38 sg13g2_a21oi_1
X_0997_ VPWR _0117_ state\[90\] VGND sg13g2_inv_1
XFILLER_39_161 VPWR VGND sg13g2_decap_8
Xfanout203 net226 net203 VPWR VGND sg13g2_buf_1
Xfanout214 net226 net214 VPWR VGND sg13g2_buf_1
Xfanout225 net226 net225 VPWR VGND sg13g2_buf_1
X_1549_ _0799_ net108 _0605_ _0606_ VPWR VGND sg13g2_a21o_1
XFILLER_24_22 VPWR VGND sg13g2_fill_2
XFILLER_24_33 VPWR VGND sg13g2_fill_1
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_14_584 VPWR VGND sg13g2_decap_8
XFILLER_33_326 VPWR VGND sg13g2_decap_8
XFILLER_41_392 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
X_0920_ VPWR _0032_ state\[13\] VGND sg13g2_inv_1
XFILLER_6_772 VPWR VGND sg13g2_decap_8
XFILLER_28_109 VPWR VGND sg13g2_decap_8
X_1403_ _0189_ _0495_ _0496_ net54 _0762_ VPWR VGND sg13g2_a22oi_1
X_1334_ VGND VPWR net81 daisychain\[43\] _0445_ net50 sg13g2_a21oi_1
X_1265_ _0728_ net99 _0392_ _0393_ VPWR VGND sg13g2_a21o_1
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_37_698 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
X_1196_ net139 VPWR _0855_ VGND net92 state\[10\] sg13g2_o21ai_1
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_19_55 VPWR VGND sg13g2_decap_8
XFILLER_27_186 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_7_525 VPWR VGND sg13g2_decap_8
XFILLER_7_536 VPWR VGND sg13g2_fill_2
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_38_418 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_33_123 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
X_1050_ VPWR _0719_ daisychain\[18\] VGND sg13g2_inv_1
XFILLER_14_370 VPWR VGND sg13g2_decap_8
XFILLER_34_679 VPWR VGND sg13g2_decap_8
X_1952_ net192 VGND VPWR _0284_ state\[28\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1883_ net216 VGND VPWR _0215_ daisychain\[87\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0903_ VPWR _0029_ state\[126\] VGND sg13g2_inv_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_1317_ _0741_ net113 _0431_ _0432_ VPWR VGND sg13g2_a21o_1
X_1248_ net148 VPWR _0894_ VGND net102 state\[23\] sg13g2_o21ai_1
XFILLER_12_307 VPWR VGND sg13g2_decap_8
XFILLER_13_808 VPWR VGND sg13g2_decap_8
XFILLER_24_112 VPWR VGND sg13g2_decap_8
XFILLER_24_156 VPWR VGND sg13g2_decap_8
X_1179_ _0133_ _0841_ _0842_ net30 _0706_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_340 VPWR VGND sg13g2_fill_1
XFILLER_20_351 VPWR VGND sg13g2_decap_8
XFILLER_20_362 VPWR VGND sg13g2_fill_1
XFILLER_21_23 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_decap_8
XFILLER_15_167 VPWR VGND sg13g2_decap_8
XFILLER_30_137 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_399 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_4
XFILLER_38_259 VPWR VGND sg13g2_decap_8
X_1102_ VPWR _0771_ daisychain\[70\] VGND sg13g2_inv_1
X_1033_ VPWR _0702_ daisychain\[1\] VGND sg13g2_inv_1
XFILLER_21_159 VPWR VGND sg13g2_decap_8
XFILLER_30_671 VPWR VGND sg13g2_fill_1
X_1935_ net187 VGND VPWR _0267_ state\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1866_ net221 VGND VPWR _0198_ daisychain\[70\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_1797_ net197 VGND VPWR _0129_ daisychain\[1\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_16_34 VPWR VGND sg13g2_decap_8
XFILLER_25_410 VPWR VGND sg13g2_fill_1
XFILLER_29_237 VPWR VGND sg13g2_decap_8
XFILLER_12_104 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_decap_8
XFILLER_40_413 VPWR VGND sg13g2_decap_8
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_4_347 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_28_270 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
X_1720_ _0468_ VPWR _0308_ VGND net163 _0075_ sg13g2_o21ai_1
X_1651_ _0251_ _0681_ _0682_ net23 _0695_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_196 VPWR VGND sg13g2_decap_8
X_1582_ VGND VPWR net76 daisychain\[105\] _0631_ net42 sg13g2_a21oi_1
XFILLER_26_207 VPWR VGND sg13g2_decap_8
X_2065_ state\[125\] net12 VPWR VGND sg13g2_buf_1
XFILLER_22_479 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_35_752 VPWR VGND sg13g2_decap_8
X_1016_ VPWR _0010_ state\[109\] VGND sg13g2_inv_1
XFILLER_2_807 VPWR VGND sg13g2_decap_8
X_1918_ net183 VGND VPWR _0250_ daisychain\[122\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1849_ net211 VGND VPWR _0181_ daisychain\[53\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_13_424 VPWR VGND sg13g2_decap_8
XFILLER_18_719 VPWR VGND sg13g2_decap_4
XFILLER_25_273 VPWR VGND sg13g2_fill_1
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_41_700 VPWR VGND sg13g2_decap_4
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_13_435 VPWR VGND sg13g2_fill_1
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_16_251 VPWR VGND sg13g2_decap_8
XFILLER_31_265 VPWR VGND sg13g2_decap_8
XFILLER_32_711 VPWR VGND sg13g2_fill_1
XFILLER_32_755 VPWR VGND sg13g2_fill_1
XFILLER_32_788 VPWR VGND sg13g2_decap_4
XFILLER_44_571 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_1703_ _0417_ VPWR _0291_ VGND net148 _0056_ sg13g2_o21ai_1
X_1634_ VGND VPWR net69 daisychain\[118\] _0670_ net27 sg13g2_a21oi_1
XFILLER_39_343 VPWR VGND sg13g2_decap_8
X_1565_ _0803_ net123 _0617_ _0618_ VPWR VGND sg13g2_a21o_1
X_1496_ net177 VPWR _0566_ VGND net130 state\[85\] sg13g2_o21ai_1
X_2048_ net184 VGND VPWR _0380_ state\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_22_243 VPWR VGND sg13g2_decap_8
Xfanout25 net29 net25 VPWR VGND sg13g2_buf_1
Xfanout69 net70 net69 VPWR VGND sg13g2_buf_1
Xfanout58 net59 net58 VPWR VGND sg13g2_buf_1
Xfanout47 net49 net47 VPWR VGND sg13g2_buf_1
Xfanout36 net44 net36 VPWR VGND sg13g2_buf_1
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
XFILLER_5_431 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[1\].u.inv2 VPWR digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_1350_ VGND VPWR net80 daisychain\[47\] _0457_ net49 sg13g2_a21oi_1
X_1281_ _0732_ net112 _0404_ _0405_ VPWR VGND sg13g2_a21o_1
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_2_1__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_20_736 VPWR VGND sg13g2_decap_4
X_0996_ VPWR _0115_ state\[89\] VGND sg13g2_inv_1
XFILLER_8_291 VPWR VGND sg13g2_decap_8
Xfanout204 net206 net204 VPWR VGND sg13g2_buf_1
X_1617_ _0816_ net105 _0656_ _0657_ VPWR VGND sg13g2_a21o_1
XFILLER_27_302 VPWR VGND sg13g2_fill_1
XFILLER_39_140 VPWR VGND sg13g2_decap_8
Xfanout215 net225 net215 VPWR VGND sg13g2_buf_1
Xfanout226 net227 net226 VPWR VGND sg13g2_buf_1
X_1548_ net155 VPWR _0605_ VGND net108 state\[98\] sg13g2_o21ai_1
X_1479_ _0208_ _0552_ _0553_ net56 _0781_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_508 VPWR VGND sg13g2_fill_2
XFILLER_43_817 VPWR VGND sg13g2_decap_4
XFILLER_10_235 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_decap_8
X_1402_ VGND VPWR net82 daisychain\[60\] _0496_ net53 sg13g2_a21oi_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_1333_ _0745_ net119 _0443_ _0444_ VPWR VGND sg13g2_a21o_1
X_1264_ net146 VPWR _0392_ VGND net99 state\[27\] sg13g2_o21ai_1
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_37_677 VPWR VGND sg13g2_fill_2
XFILLER_40_809 VPWR VGND sg13g2_decap_8
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
X_1195_ _0137_ _0853_ _0854_ net25 _0710_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_382 VPWR VGND sg13g2_decap_4
X_0979_ VPWR _0097_ state\[72\] VGND sg13g2_inv_1
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_16_806 VPWR VGND sg13g2_fill_2
XFILLER_19_34 VPWR VGND sg13g2_decap_8
XFILLER_27_165 VPWR VGND sg13g2_decap_8
XFILLER_15_349 VPWR VGND sg13g2_decap_8
XFILLER_23_371 VPWR VGND sg13g2_fill_2
XFILLER_30_319 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_43_636 VPWR VGND sg13g2_fill_1
XFILLER_43_658 VPWR VGND sg13g2_fill_2
XFILLER_7_504 VPWR VGND sg13g2_decap_8
XFILLER_11_577 VPWR VGND sg13g2_fill_1
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_3_776 VPWR VGND sg13g2_decap_8
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_19_699 VPWR VGND sg13g2_fill_2
XFILLER_33_102 VPWR VGND sg13g2_decap_8
XFILLER_33_179 VPWR VGND sg13g2_decap_8
XFILLER_34_647 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
X_1951_ net191 VGND VPWR _0283_ state\[27\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1882_ net217 VGND VPWR _0214_ daisychain\[86\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0902_ VPWR _0698_ daisychain\[124\] VGND sg13g2_inv_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_6_581 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
X_1316_ net159 VPWR _0431_ VGND net113 state\[40\] sg13g2_o21ai_1
X_1247_ _0150_ _0892_ _0893_ net35 _0723_ VPWR VGND sg13g2_a22oi_1
X_1178_ VGND VPWR net71 daisychain\[4\] _0842_ net30 sg13g2_a21oi_1
XFILLER_24_135 VPWR VGND sg13g2_decap_8
XFILLER_40_639 VPWR VGND sg13g2_decap_8
XFILLER_20_374 VPWR VGND sg13g2_fill_2
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_15_146 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_11_396 VPWR VGND sg13g2_decap_8
XFILLER_30_116 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_decap_8
XFILLER_7_378 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
X_1101_ VPWR _0770_ daisychain\[69\] VGND sg13g2_inv_1
X_1032_ VPWR _0701_ daisychain\[0\] VGND sg13g2_inv_1
XFILLER_15_691 VPWR VGND sg13g2_decap_8
XFILLER_21_138 VPWR VGND sg13g2_decap_8
XFILLER_30_650 VPWR VGND sg13g2_fill_1
XFILLER_34_422 VPWR VGND sg13g2_decap_8
XFILLER_34_477 VPWR VGND sg13g2_decap_8
X_1934_ net187 VGND VPWR _0266_ state\[10\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1865_ net221 VGND VPWR _0197_ daisychain\[69\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_1796_ net196 VGND VPWR _0128_ daisychain\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_29_216 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_fill_1
XFILLER_16_13 VPWR VGND sg13g2_decap_8
XFILLER_20_182 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_16_488 VPWR VGND sg13g2_fill_2
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_11_193 VPWR VGND sg13g2_decap_8
XFILLER_12_672 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_8_621 VPWR VGND sg13g2_decap_8
XFILLER_8_632 VPWR VGND sg13g2_fill_2
XFILLER_8_643 VPWR VGND sg13g2_decap_8
X_1650_ VGND VPWR net70 daisychain\[122\] _0682_ net23 sg13g2_a21oi_1
X_1581_ _0807_ net106 _0629_ _0630_ VPWR VGND sg13g2_a21o_1
XFILLER_39_514 VPWR VGND sg13g2_fill_2
XFILLER_3_392 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
X_2064_ state\[124\] net11 VPWR VGND sg13g2_buf_1
X_1015_ VPWR _0009_ state\[108\] VGND sg13g2_inv_1
XFILLER_30_491 VPWR VGND sg13g2_decap_4
X_1917_ net183 VGND VPWR _0249_ daisychain\[121\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_1_329 VPWR VGND sg13g2_decap_8
X_1848_ net211 VGND VPWR _0180_ daisychain\[52\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1779_ _0645_ VPWR _0367_ VGND net152 _0013_ sg13g2_o21ai_1
XFILLER_13_403 VPWR VGND sg13g2_decap_8
XFILLER_13_458 VPWR VGND sg13g2_decap_8
XFILLER_45_539 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_16_230 VPWR VGND sg13g2_decap_8
XFILLER_17_731 VPWR VGND sg13g2_fill_1
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_31_244 VPWR VGND sg13g2_decap_8
XFILLER_8_473 VPWR VGND sg13g2_decap_8
XFILLER_8_484 VPWR VGND sg13g2_decap_8
X_1702_ _0414_ VPWR _0290_ VGND net161 _0055_ sg13g2_o21ai_1
X_1633_ _0820_ net95 _0668_ _0669_ VPWR VGND sg13g2_a21o_1
X_1564_ net170 VPWR _0617_ VGND net123 state\[102\] sg13g2_o21ai_1
XFILLER_39_322 VPWR VGND sg13g2_decap_8
XFILLER_4_690 VPWR VGND sg13g2_decap_8
X_1495_ _0212_ _0564_ _0565_ net58 _0785_ VPWR VGND sg13g2_a22oi_1
XFILLER_22_222 VPWR VGND sg13g2_decap_8
XFILLER_39_399 VPWR VGND sg13g2_decap_8
X_2047_ net183 VGND VPWR _0379_ state\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
Xfanout26 net29 net26 VPWR VGND sg13g2_buf_1
Xfanout37 net38 net37 VPWR VGND sg13g2_buf_1
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_22_299 VPWR VGND sg13g2_decap_8
Xfanout59 net60 net59 VPWR VGND sg13g2_buf_1
Xfanout48 net49 net48 VPWR VGND sg13g2_buf_1
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_46_815 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_14_778 VPWR VGND sg13g2_decap_8
XFILLER_14_789 VPWR VGND sg13g2_fill_1
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_37_815 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_49_664 VPWR VGND sg13g2_fill_1
X_1280_ net158 VPWR _0404_ VGND net112 state\[31\] sg13g2_o21ai_1
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_32_564 VPWR VGND sg13g2_decap_8
XFILLER_32_597 VPWR VGND sg13g2_decap_4
XFILLER_8_270 VPWR VGND sg13g2_decap_8
X_0995_ VPWR _0114_ state\[88\] VGND sg13g2_inv_1
XFILLER_5_81 VPWR VGND sg13g2_decap_8
Xfanout205 net206 net205 VPWR VGND sg13g2_buf_1
Xfanout216 net218 net216 VPWR VGND sg13g2_buf_1
Xfanout227 net1 net227 VPWR VGND sg13g2_buf_1
X_1616_ net152 VPWR _0656_ VGND net105 state\[115\] sg13g2_o21ai_1
X_1547_ _0225_ _0603_ _0604_ net42 _0798_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_196 VPWR VGND sg13g2_decap_8
X_1478_ VGND VPWR net85 daisychain\[79\] _0553_ net56 sg13g2_a21oi_1
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_24_57 VPWR VGND sg13g2_fill_2
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_18_347 VPWR VGND sg13g2_decap_4
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_14_542 VPWR VGND sg13g2_decap_8
XFILLER_14_90 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_5_284 VPWR VGND sg13g2_decap_8
XFILLER_6_752 VPWR VGND sg13g2_fill_1
X_1401_ _0762_ net120 _0494_ _0495_ VPWR VGND sg13g2_a21o_1
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_49_494 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
X_1332_ net163 VPWR _0443_ VGND net119 state\[44\] sg13g2_o21ai_1
X_1263_ _0154_ _0390_ _0391_ net33 _0727_ VPWR VGND sg13g2_a22oi_1
X_1194_ VGND VPWR net68 daisychain\[8\] _0854_ net25 sg13g2_a21oi_1
XFILLER_24_317 VPWR VGND sg13g2_decap_4
XFILLER_32_361 VPWR VGND sg13g2_decap_8
X_0978_ VPWR _0096_ state\[71\] VGND sg13g2_inv_1
XFILLER_19_13 VPWR VGND sg13g2_decap_8
XFILLER_15_328 VPWR VGND sg13g2_decap_8
XFILLER_16_818 VPWR VGND sg13g2_decap_4
XFILLER_27_144 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_43_648 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_19_667 VPWR VGND sg13g2_decap_4
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_19_689 VPWR VGND sg13g2_fill_1
XFILLER_33_158 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
X_1950_ net192 VGND VPWR _0282_ state\[26\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1881_ net217 VGND VPWR _0213_ daisychain\[85\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0901_ VPWR _0697_ daisychain\[125\] VGND sg13g2_inv_1
X_1315_ _0167_ _0429_ _0430_ net47 _0740_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_37_475 VPWR VGND sg13g2_decap_4
XFILLER_49_291 VPWR VGND sg13g2_decap_8
X_1246_ VGND VPWR net73 daisychain\[21\] _0893_ net35 sg13g2_a21oi_1
X_1177_ _0706_ net96 _0840_ _0841_ VPWR VGND sg13g2_a21o_1
XFILLER_33_681 VPWR VGND sg13g2_fill_1
XFILLER_4_508 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_15_125 VPWR VGND sg13g2_decap_8
XFILLER_16_659 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_decap_8
XFILLER_23_191 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_30_8 VPWR VGND sg13g2_fill_2
XFILLER_3_574 VPWR VGND sg13g2_fill_2
XFILLER_19_464 VPWR VGND sg13g2_fill_2
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
X_1100_ VPWR _0769_ daisychain\[68\] VGND sg13g2_inv_1
X_1031_ VPWR _0027_ state\[124\] VGND sg13g2_inv_1
XFILLER_21_117 VPWR VGND sg13g2_decap_8
X_1933_ net185 VGND VPWR _0265_ state\[9\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1864_ net221 VGND VPWR _0196_ daisychain\[68\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_1795_ _0693_ VPWR _0383_ VGND net137 _0030_ sg13g2_o21ai_1
XFILLER_16_69 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
X_1229_ _0719_ net98 _0879_ _0880_ VPWR VGND sg13g2_a21o_1
XFILLER_12_139 VPWR VGND sg13g2_decap_8
XFILLER_20_161 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_40_448 VPWR VGND sg13g2_decap_8
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_44_721 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_fill_2
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
X_1580_ net152 VPWR _0629_ VGND net106 state\[106\] sg13g2_o21ai_1
XFILLER_39_548 VPWR VGND sg13g2_decap_4
XFILLER_3_371 VPWR VGND sg13g2_decap_8
XFILLER_19_272 VPWR VGND sg13g2_decap_4
XFILLER_34_231 VPWR VGND sg13g2_decap_8
X_2063_ state\[123\] net10 VPWR VGND sg13g2_buf_1
X_1014_ VPWR _0008_ state\[107\] VGND sg13g2_inv_1
XFILLER_8_81 VPWR VGND sg13g2_decap_8
X_1916_ net186 VGND VPWR _0248_ daisychain\[120\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1847_ net212 VGND VPWR _0179_ daisychain\[51\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_1_308 VPWR VGND sg13g2_decap_8
X_1778_ _0642_ VPWR _0366_ VGND net153 _0012_ sg13g2_o21ai_1
XFILLER_17_209 VPWR VGND sg13g2_decap_8
XFILLER_45_518 VPWR VGND sg13g2_decap_8
XFILLER_25_264 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_fill_2
XFILLER_41_779 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_5_658 VPWR VGND sg13g2_fill_2
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_17_776 VPWR VGND sg13g2_decap_4
XFILLER_17_90 VPWR VGND sg13g2_decap_8
XFILLER_36_507 VPWR VGND sg13g2_decap_4
XFILLER_44_540 VPWR VGND sg13g2_fill_1
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_16_286 VPWR VGND sg13g2_decap_8
XFILLER_31_223 VPWR VGND sg13g2_decap_8
XFILLER_8_452 VPWR VGND sg13g2_decap_8
X_1701_ _0411_ VPWR _0289_ VGND net160 _0054_ sg13g2_o21ai_1
X_1632_ net140 VPWR _0668_ VGND net95 state\[119\] sg13g2_o21ai_1
X_1563_ _0229_ _0615_ _0616_ net56 _0802_ VPWR VGND sg13g2_a22oi_1
X_1494_ VGND VPWR net84 daisychain\[83\] _0565_ net58 sg13g2_a21oi_1
XFILLER_27_529 VPWR VGND sg13g2_fill_1
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_39_378 VPWR VGND sg13g2_decap_8
XFILLER_22_201 VPWR VGND sg13g2_decap_8
X_2046_ net183 VGND VPWR _0378_ state\[122\] clknet_leaf_17_clk sg13g2_dfrbpq_1
Xfanout27 net28 net27 VPWR VGND sg13g2_buf_1
Xfanout49 net67 net49 VPWR VGND sg13g2_buf_1
Xfanout38 net39 net38 VPWR VGND sg13g2_buf_1
XFILLER_22_278 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_49_610 VPWR VGND sg13g2_decap_8
XFILLER_49_643 VPWR VGND sg13g2_decap_8
XFILLER_17_584 VPWR VGND sg13g2_decap_8
XFILLER_44_392 VPWR VGND sg13g2_decap_8
X_0994_ VPWR _0113_ state\[87\] VGND sg13g2_inv_1
XFILLER_5_60 VPWR VGND sg13g2_decap_8
Xfanout206 net208 net206 VPWR VGND sg13g2_buf_1
Xfanout217 net218 net217 VPWR VGND sg13g2_buf_1
X_1615_ _0242_ _0654_ _0655_ net37 _0815_ VPWR VGND sg13g2_a22oi_1
X_1546_ VGND VPWR net76 daisychain\[96\] _0604_ net42 sg13g2_a21oi_1
X_1477_ _0781_ net123 _0551_ _0552_ VPWR VGND sg13g2_a21o_1
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_11_738 VPWR VGND sg13g2_decap_4
XFILLER_23_543 VPWR VGND sg13g2_fill_1
XFILLER_35_392 VPWR VGND sg13g2_decap_8
XFILLER_42_329 VPWR VGND sg13g2_decap_8
X_2029_ net199 VGND VPWR _0361_ state\[105\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_19_816 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_26_381 VPWR VGND sg13g2_fill_2
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_46_646 VPWR VGND sg13g2_decap_8
XFILLER_46_657 VPWR VGND sg13g2_fill_1
XFILLER_14_598 VPWR VGND sg13g2_decap_8
XFILLER_6_742 VPWR VGND sg13g2_decap_4
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_6_786 VPWR VGND sg13g2_decap_8
Xwires dac/Iout dac/VcascP[1] dac/VcascP[0] dac/VbiasP[1] dac/VbiasP[0] wires/VDDA[1]
+ wires/VDDA[0] i_in i_out analog_wires
X_1400_ net167 VPWR _0494_ VGND net120 state\[61\] sg13g2_o21ai_1
X_1331_ _0171_ _0441_ _0442_ net46 _0744_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_37_602 VPWR VGND sg13g2_decap_4
XFILLER_49_473 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
X_1262_ VGND VPWR net72 daisychain\[25\] _0391_ net33 sg13g2_a21oi_1
X_1193_ _0710_ net92 _0852_ _0853_ VPWR VGND sg13g2_a21o_1
XFILLER_17_370 VPWR VGND sg13g2_decap_4
XFILLER_20_535 VPWR VGND sg13g2_fill_2
XFILLER_24_329 VPWR VGND sg13g2_fill_2
XFILLER_32_340 VPWR VGND sg13g2_decap_8
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_45_690 VPWR VGND sg13g2_decap_8
X_0977_ VPWR _0095_ state\[70\] VGND sg13g2_inv_1
XFILLER_9_580 VPWR VGND sg13g2_decap_8
XFILLER_19_69 VPWR VGND sg13g2_decap_8
XFILLER_27_101 VPWR VGND sg13g2_decap_8
X_1529_ _0794_ net124 _0590_ _0591_ VPWR VGND sg13g2_a21o_1
XFILLER_15_307 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_fill_1
XFILLER_43_627 VPWR VGND sg13g2_decap_8
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_3_756 VPWR VGND sg13g2_fill_2
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_19_624 VPWR VGND sg13g2_decap_4
XFILLER_19_646 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_14_384 VPWR VGND sg13g2_decap_8
XFILLER_30_800 VPWR VGND sg13g2_decap_8
XFILLER_30_811 VPWR VGND sg13g2_fill_2
XFILLER_33_137 VPWR VGND sg13g2_decap_8
X_1880_ net217 VGND VPWR _0212_ daisychain\[84\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_0900_ VPWR _0028_ state\[125\] VGND sg13g2_inv_1
X_1314_ VGND VPWR net79 daisychain\[38\] _0430_ net45 sg13g2_a21oi_1
XFILLER_37_454 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_8
X_1245_ _0723_ net101 _0891_ _0892_ VPWR VGND sg13g2_a21o_1
X_1176_ net142 VPWR _0840_ VGND net96 state\[5\] sg13g2_o21ai_1
XFILLER_21_15 VPWR VGND sg13g2_decap_4
XFILLER_21_37 VPWR VGND sg13g2_decap_8
XFILLER_40_619 VPWR VGND sg13g2_decap_8
XFILLER_28_421 VPWR VGND sg13g2_decap_4
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_15_104 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_39_708 VPWR VGND sg13g2_decap_4
XFILLER_3_553 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_47_774 VPWR VGND sg13g2_decap_4
X_1030_ VPWR _0026_ state\[123\] VGND sg13g2_inv_1
XFILLER_14_181 VPWR VGND sg13g2_decap_8
XFILLER_42_490 VPWR VGND sg13g2_decap_8
X_1932_ net185 VGND VPWR _0264_ state\[8\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1863_ net221 VGND VPWR _0195_ daisychain\[67\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_1794_ _0690_ VPWR _0382_ VGND net137 _0029_ sg13g2_o21ai_1
XFILLER_38_774 VPWR VGND sg13g2_decap_4
X_1228_ net145 VPWR _0879_ VGND net98 state\[18\] sg13g2_o21ai_1
XFILLER_12_118 VPWR VGND sg13g2_decap_8
XFILLER_16_48 VPWR VGND sg13g2_decap_8
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_decap_8
X_1159_ _0128_ _0827_ _0825_ net37 _0701_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_140 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_5_807 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_24_490 VPWR VGND sg13g2_fill_1
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_3_350 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_4
X_2062_ state\[122\] net9 VPWR VGND sg13g2_buf_1
XFILLER_19_251 VPWR VGND sg13g2_decap_8
XFILLER_19_295 VPWR VGND sg13g2_decap_8
XFILLER_22_405 VPWR VGND sg13g2_fill_2
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_8
XFILLER_35_733 VPWR VGND sg13g2_fill_1
XFILLER_35_766 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
X_1013_ VPWR _0007_ state\[106\] VGND sg13g2_inv_1
XFILLER_8_60 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_1915_ net186 VGND VPWR _0247_ daisychain\[119\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1846_ net212 VGND VPWR _0178_ daisychain\[50\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1777_ _0639_ VPWR _0365_ VGND net153 _0010_ sg13g2_o21ai_1
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_38_582 VPWR VGND sg13g2_fill_1
XFILLER_25_243 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_41_714 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_16_265 VPWR VGND sg13g2_decap_8
XFILLER_31_202 VPWR VGND sg13g2_decap_8
XFILLER_31_279 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_decap_8
X_1700_ _0408_ VPWR _0288_ VGND net158 _0053_ sg13g2_o21ai_1
X_1631_ _0246_ _0666_ _0667_ net28 _0819_ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_1562_ VGND VPWR net85 daisychain\[100\] _0616_ net56 sg13g2_a21oi_1
X_1493_ _0785_ net125 _0563_ _0564_ VPWR VGND sg13g2_a21o_1
XFILLER_39_357 VPWR VGND sg13g2_decap_8
X_2045_ net184 VGND VPWR _0377_ state\[121\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_22_257 VPWR VGND sg13g2_decap_8
XFILLER_35_574 VPWR VGND sg13g2_decap_8
Xfanout28 net29 net28 VPWR VGND sg13g2_buf_1
Xfanout39 net44 net39 VPWR VGND sg13g2_buf_1
X_1829_ net192 VGND VPWR _0161_ daisychain\[33\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_14_725 VPWR VGND sg13g2_decap_8
XFILLER_41_511 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_41_588 VPWR VGND sg13g2_fill_1
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_20_717 VPWR VGND sg13g2_fill_1
XFILLER_44_371 VPWR VGND sg13g2_decap_8
X_0993_ VPWR _0112_ state\[86\] VGND sg13g2_inv_1
X_1614_ VGND VPWR net75 daisychain\[113\] _0655_ net37 sg13g2_a21oi_1
XFILLER_9_784 VPWR VGND sg13g2_decap_4
Xfanout207 net208 net207 VPWR VGND sg13g2_buf_1
Xfanout218 net225 net218 VPWR VGND sg13g2_buf_1
X_1545_ _0798_ net109 _0602_ _0603_ VPWR VGND sg13g2_a21o_1
X_1476_ net170 VPWR _0551_ VGND net123 state\[80\] sg13g2_o21ai_1
XFILLER_23_522 VPWR VGND sg13g2_fill_2
XFILLER_35_371 VPWR VGND sg13g2_decap_8
XFILLER_39_154 VPWR VGND sg13g2_decap_8
XFILLER_42_308 VPWR VGND sg13g2_decap_8
X_2028_ net200 VGND VPWR _0360_ state\[104\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_33_319 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_10_772 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_6_721 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
X_1330_ VGND VPWR net79 daisychain\[42\] _0442_ net46 sg13g2_a21oi_1
X_1261_ _0727_ net99 _0389_ _0390_ VPWR VGND sg13g2_a21o_1
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_8
X_1192_ net139 VPWR _0852_ VGND net92 state\[9\] sg13g2_o21ai_1
X_0976_ VPWR _0093_ state\[69\] VGND sg13g2_inv_1
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_19_48 VPWR VGND sg13g2_decap_8
X_1528_ net171 VPWR _0590_ VGND net124 state\[93\] sg13g2_o21ai_1
X_1459_ _0203_ _0537_ _0538_ net63 _0776_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_179 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_7_518 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_3_746 VPWR VGND sg13g2_fill_2
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_decap_8
XFILLER_33_116 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_14_363 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
XFILLER_6_595 VPWR VGND sg13g2_fill_2
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_37_433 VPWR VGND sg13g2_decap_4
X_1313_ _0740_ net113 _0428_ _0429_ VPWR VGND sg13g2_a21o_1
X_1244_ net147 VPWR _0891_ VGND net102 state\[22\] sg13g2_o21ai_1
XFILLER_18_680 VPWR VGND sg13g2_decap_8
XFILLER_18_691 VPWR VGND sg13g2_fill_2
XFILLER_24_149 VPWR VGND sg13g2_decap_8
X_1175_ _0132_ _0838_ _0839_ net31 _0705_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_333 VPWR VGND sg13g2_fill_2
XFILLER_20_344 VPWR VGND sg13g2_decap_8
XFILLER_32_193 VPWR VGND sg13g2_decap_8
X_0959_ VPWR _0075_ state\[52\] VGND sg13g2_inv_1
XFILLER_0_716 VPWR VGND sg13g2_fill_1
XFILLER_16_628 VPWR VGND sg13g2_decap_4
XFILLER_28_499 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_11_333 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_8_816 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_532 VPWR VGND sg13g2_decap_8
XFILLER_16_8 VPWR VGND sg13g2_fill_1
XFILLER_3_576 VPWR VGND sg13g2_fill_1
XFILLER_19_466 VPWR VGND sg13g2_fill_1
XFILLER_34_403 VPWR VGND sg13g2_fill_1
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_14_160 VPWR VGND sg13g2_decap_8
X_1931_ net185 VGND VPWR _0263_ state\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1862_ net219 VGND VPWR _0194_ daisychain\[66\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1793_ _0687_ VPWR _0381_ VGND net137 _0028_ sg13g2_o21ai_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_37_252 VPWR VGND sg13g2_decap_8
X_1227_ _0145_ _0877_ _0878_ net32 _0718_ VPWR VGND sg13g2_a22oi_1
X_1158_ VGND VPWR net68 net2 _0827_ net27 sg13g2_a21oi_1
XFILLER_16_27 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_8
X_1089_ VPWR _0758_ daisychain\[57\] VGND sg13g2_inv_1
XFILLER_20_196 VPWR VGND sg13g2_decap_8
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_28_263 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_12_664 VPWR VGND sg13g2_fill_1
XFILLER_12_686 VPWR VGND sg13g2_decap_4
XFILLER_12_697 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_8_657 VPWR VGND sg13g2_fill_2
XFILLER_8_668 VPWR VGND sg13g2_fill_1
XFILLER_8_679 VPWR VGND sg13g2_fill_2
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_19_230 VPWR VGND sg13g2_decap_8
X_2061_ state\[121\] net8 VPWR VGND sg13g2_buf_1
X_1012_ VPWR _0006_ state\[105\] VGND sg13g2_inv_1
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_35_745 VPWR VGND sg13g2_decap_8
X_1914_ net186 VGND VPWR _0246_ daisychain\[118\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_30_472 VPWR VGND sg13g2_decap_8
X_1845_ net212 VGND VPWR _0177_ daisychain\[49\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1776_ _0636_ VPWR _0364_ VGND net151 _0009_ sg13g2_o21ai_1
XFILLER_25_222 VPWR VGND sg13g2_decap_8
XFILLER_27_37 VPWR VGND sg13g2_fill_2
XFILLER_41_704 VPWR VGND sg13g2_fill_2
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_13_417 VPWR VGND sg13g2_decap_8
XFILLER_21_450 VPWR VGND sg13g2_fill_2
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_41_737 VPWR VGND sg13g2_fill_1
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_16_244 VPWR VGND sg13g2_decap_8
XFILLER_31_258 VPWR VGND sg13g2_decap_8
XFILLER_32_748 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_8_498 VPWR VGND sg13g2_decap_8
X_1630_ VGND VPWR net69 daisychain\[117\] _0667_ net28 sg13g2_a21oi_1
X_1561_ _0802_ net123 _0614_ _0615_ VPWR VGND sg13g2_a21o_1
X_1492_ net177 VPWR _0563_ VGND net125 state\[84\] sg13g2_o21ai_1
XFILLER_39_336 VPWR VGND sg13g2_decap_8
X_2044_ net186 VGND VPWR _0376_ state\[120\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_22_236 VPWR VGND sg13g2_decap_8
XFILLER_30_291 VPWR VGND sg13g2_decap_8
XFILLER_35_597 VPWR VGND sg13g2_fill_1
Xfanout29 _0826_ net29 VPWR VGND sg13g2_buf_1
X_1828_ net204 VGND VPWR _0160_ daisychain\[32\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1759_ _0585_ VPWR _0347_ VGND net173 _0118_ sg13g2_o21ai_1
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_26_531 VPWR VGND sg13g2_decap_4
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_32_578 VPWR VGND sg13g2_decap_4
XFILLER_32_589 VPWR VGND sg13g2_fill_2
X_0992_ VPWR _0111_ state\[85\] VGND sg13g2_inv_1
XFILLER_8_284 VPWR VGND sg13g2_decap_8
X_1613_ _0815_ net104 _0653_ _0654_ VPWR VGND sg13g2_a21o_1
X_1544_ net154 VPWR _0602_ VGND net109 state\[97\] sg13g2_o21ai_1
XFILLER_39_133 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
Xfanout208 net226 net208 VPWR VGND sg13g2_buf_1
Xfanout219 net224 net219 VPWR VGND sg13g2_buf_1
X_1475_ _0207_ _0549_ _0550_ net61 _0780_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_350 VPWR VGND sg13g2_decap_8
X_2027_ net200 VGND VPWR _0359_ state\[103\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_26_394 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_10_762 VPWR VGND sg13g2_fill_2
XFILLER_30_81 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
X_1260_ net146 VPWR _0389_ VGND net99 state\[26\] sg13g2_o21ai_1
X_1191_ _0136_ _0850_ _0851_ net25 _0709_ VPWR VGND sg13g2_a22oi_1
XFILLER_33_821 VPWR VGND sg13g2_fill_2
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_32_375 VPWR VGND sg13g2_decap_8
X_0975_ VPWR _0092_ state\[68\] VGND sg13g2_inv_1
XFILLER_10_18 VPWR VGND sg13g2_decap_8
X_1527_ _0220_ _0588_ _0589_ net57 _0793_ VPWR VGND sg13g2_a22oi_1
XFILLER_19_27 VPWR VGND sg13g2_decap_8
XFILLER_27_158 VPWR VGND sg13g2_decap_8
XFILLER_43_607 VPWR VGND sg13g2_decap_4
X_1458_ VGND VPWR net86 daisychain\[74\] _0538_ net63 sg13g2_a21oi_1
X_1389_ _0759_ net118 _0485_ _0486_ VPWR VGND sg13g2_a21o_1
XFILLER_23_364 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_3_769 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_15_810 VPWR VGND sg13g2_decap_8
XFILLER_15_821 VPWR VGND sg13g2_fill_2
XFILLER_18_158 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_14_342 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_42_662 VPWR VGND sg13g2_decap_8
XFILLER_42_673 VPWR VGND sg13g2_fill_2
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
X_1312_ net159 VPWR _0428_ VGND net113 state\[39\] sg13g2_o21ai_1
X_1243_ _0149_ _0889_ _0890_ net31 _0722_ VPWR VGND sg13g2_a22oi_1
X_1174_ VGND VPWR net71 daisychain\[3\] _0839_ net31 sg13g2_a21oi_1
XFILLER_20_323 VPWR VGND sg13g2_decap_4
XFILLER_32_172 VPWR VGND sg13g2_decap_8
X_0958_ VPWR _0074_ state\[51\] VGND sg13g2_inv_1
XFILLER_15_139 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_11_312 VPWR VGND sg13g2_decap_8
XFILLER_11_389 VPWR VGND sg13g2_decap_8
XFILLER_30_109 VPWR VGND sg13g2_decap_8
XFILLER_3_511 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_decap_4
XFILLER_36_91 VPWR VGND sg13g2_decap_8
X_1930_ net189 VGND VPWR _0262_ state\[6\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_30_643 VPWR VGND sg13g2_fill_2
XFILLER_30_654 VPWR VGND sg13g2_decap_4
X_1861_ net219 VGND VPWR _0193_ daisychain\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1792_ _0684_ VPWR _0380_ VGND net141 _0027_ sg13g2_o21ai_1
XFILLER_29_209 VPWR VGND sg13g2_decap_8
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_25_437 VPWR VGND sg13g2_fill_2
XFILLER_37_231 VPWR VGND sg13g2_decap_8
XFILLER_38_754 VPWR VGND sg13g2_fill_1
X_1226_ VGND VPWR net71 daisychain\[16\] _0878_ net32 sg13g2_a21oi_1
X_1157_ net137 net3 _0826_ VPWR VGND sg13g2_nor2_1
XFILLER_20_175 VPWR VGND sg13g2_decap_8
X_1088_ VPWR _0757_ daisychain\[56\] VGND sg13g2_inv_1
XFILLER_4_319 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_44_713 VPWR VGND sg13g2_decap_4
XFILLER_11_186 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_39_507 VPWR VGND sg13g2_decap_8
XFILLER_3_385 VPWR VGND sg13g2_decap_8
X_2060_ state\[120\] net7 VPWR VGND sg13g2_buf_1
X_1011_ VPWR _0005_ state\[104\] VGND sg13g2_inv_1
XFILLER_34_245 VPWR VGND sg13g2_decap_8
X_1913_ net186 VGND VPWR _0245_ daisychain\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_7_691 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
X_1844_ net207 VGND VPWR _0176_ daisychain\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1775_ _0633_ VPWR _0363_ VGND net151 _0008_ sg13g2_o21ai_1
XFILLER_25_201 VPWR VGND sg13g2_decap_8
X_1209_ _0714_ net96 _0864_ _0865_ VPWR VGND sg13g2_a21o_1
XFILLER_21_484 VPWR VGND sg13g2_fill_2
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_16_223 VPWR VGND sg13g2_decap_8
XFILLER_44_532 VPWR VGND sg13g2_fill_2
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_12_440 VPWR VGND sg13g2_fill_2
XFILLER_31_237 VPWR VGND sg13g2_decap_8
XFILLER_32_705 VPWR VGND sg13g2_fill_2
XFILLER_32_727 VPWR VGND sg13g2_decap_4
XFILLER_40_771 VPWR VGND sg13g2_decap_8
XFILLER_44_587 VPWR VGND sg13g2_fill_2
XFILLER_33_81 VPWR VGND sg13g2_decap_8
XFILLER_8_466 VPWR VGND sg13g2_decap_8
X_1560_ net170 VPWR _0614_ VGND net123 state\[101\] sg13g2_o21ai_1
XFILLER_39_315 VPWR VGND sg13g2_decap_8
XFILLER_3_182 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
X_1491_ _0211_ _0561_ _0562_ net58 _0784_ VPWR VGND sg13g2_a22oi_1
XFILLER_22_215 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
X_2043_ net187 VGND VPWR _0375_ state\[119\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_30_270 VPWR VGND sg13g2_decap_8
XFILLER_31_771 VPWR VGND sg13g2_fill_2
X_1827_ net204 VGND VPWR _0159_ daisychain\[31\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
X_1758_ _0582_ VPWR _0346_ VGND net173 _0117_ sg13g2_o21ai_1
X_1689_ _0889_ VPWR _0277_ VGND net143 _0041_ sg13g2_o21ai_1
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_46_808 VPWR VGND sg13g2_decap_8
XFILLER_26_543 VPWR VGND sg13g2_fill_1
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_21_292 VPWR VGND sg13g2_decap_4
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_37_808 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_49_657 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
X_0991_ VPWR _0110_ state\[84\] VGND sg13g2_inv_1
XFILLER_9_731 VPWR VGND sg13g2_decap_8
XFILLER_4_480 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
Xfanout209 net214 net209 VPWR VGND sg13g2_buf_1
X_1612_ net151 VPWR _0653_ VGND net104 state\[114\] sg13g2_o21ai_1
X_1543_ _0224_ _0600_ _0601_ net42 _0797_ VPWR VGND sg13g2_a22oi_1
X_1474_ VGND VPWR net87 daisychain\[78\] _0550_ net61 sg13g2_a21oi_1
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
X_2026_ net215 VGND VPWR _0358_ state\[102\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_14_535 VPWR VGND sg13g2_decap_8
XFILLER_14_83 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_30_60 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
X_1190_ VGND VPWR net68 daisychain\[7\] _0851_ net25 sg13g2_a21oi_1
XFILLER_20_505 VPWR VGND sg13g2_decap_4
XFILLER_32_354 VPWR VGND sg13g2_decap_8
XFILLER_32_398 VPWR VGND sg13g2_decap_4
X_0974_ VPWR _0091_ state\[67\] VGND sg13g2_inv_1
XFILLER_9_594 VPWR VGND sg13g2_decap_8
X_1526_ VGND VPWR net84 daisychain\[91\] _0589_ net59 sg13g2_a21oi_1
X_1457_ _0776_ net130 _0536_ _0537_ VPWR VGND sg13g2_a21o_1
XFILLER_27_137 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
X_1388_ net164 VPWR _0485_ VGND net117 state\[58\] sg13g2_o21ai_1
X_2009_ net223 VGND VPWR _0341_ state\[85\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_14_321 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_14_398 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_531 VPWR VGND sg13g2_fill_1
XFILLER_6_575 VPWR VGND sg13g2_fill_1
X_1311_ _0166_ _0426_ _0427_ net48 _0739_ VPWR VGND sg13g2_a22oi_1
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_37_468 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
X_1242_ VGND VPWR net74 daisychain\[20\] _0890_ net31 sg13g2_a21oi_1
X_1173_ _0705_ net97 _0837_ _0838_ VPWR VGND sg13g2_a21o_1
XFILLER_17_181 VPWR VGND sg13g2_decap_8
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_33_641 VPWR VGND sg13g2_decap_8
XFILLER_45_490 VPWR VGND sg13g2_decap_8
XFILLER_20_368 VPWR VGND sg13g2_fill_1
XFILLER_20_379 VPWR VGND sg13g2_decap_4
X_0957_ VPWR _0073_ state\[50\] VGND sg13g2_inv_1
X_1509_ _0789_ net124 _0575_ _0576_ VPWR VGND sg13g2_a21o_1
XFILLER_15_118 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_23_184 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_8
XFILLER_3_567 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_14_195 VPWR VGND sg13g2_decap_8
XFILLER_15_663 VPWR VGND sg13g2_fill_1
XFILLER_30_633 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
X_1860_ net219 VGND VPWR _0192_ daisychain\[64\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_6_361 VPWR VGND sg13g2_decap_8
X_1791_ _0681_ VPWR _0379_ VGND net138 _0026_ sg13g2_o21ai_1
XFILLER_38_722 VPWR VGND sg13g2_decap_8
XFILLER_37_210 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_2_1__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_1225_ _0718_ net98 _0876_ _0877_ VPWR VGND sg13g2_a21o_1
X_1156_ _0701_ net104 _0824_ _0825_ VPWR VGND sg13g2_a21o_1
X_1087_ VPWR _0756_ daisychain\[55\] VGND sg13g2_inv_1
XFILLER_20_154 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
X_1989_ net224 VGND VPWR _0321_ state\[65\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_12_622 VPWR VGND sg13g2_fill_2
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_8_659 VPWR VGND sg13g2_fill_1
XFILLER_21_8 VPWR VGND sg13g2_decap_8
XFILLER_3_364 VPWR VGND sg13g2_decap_8
XFILLER_19_265 VPWR VGND sg13g2_decap_8
XFILLER_19_276 VPWR VGND sg13g2_fill_2
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_35_703 VPWR VGND sg13g2_fill_2
XFILLER_47_574 VPWR VGND sg13g2_decap_4
XFILLER_47_91 VPWR VGND sg13g2_decap_8
X_1010_ VPWR _0004_ state\[103\] VGND sg13g2_inv_1
XFILLER_30_452 VPWR VGND sg13g2_fill_1
XFILLER_8_74 VPWR VGND sg13g2_decap_8
X_1912_ net186 VGND VPWR _0244_ daisychain\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1843_ net207 VGND VPWR _0175_ daisychain\[47\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_6_clk clknet_2_3__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_1774_ _0630_ VPWR _0362_ VGND net152 _0007_ sg13g2_o21ai_1
XFILLER_27_39 VPWR VGND sg13g2_fill_1
X_1208_ net142 VPWR _0864_ VGND net96 state\[13\] sg13g2_o21ai_1
XFILLER_25_257 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
X_1139_ VPWR _0808_ daisychain\[107\] VGND sg13g2_inv_1
XFILLER_21_452 VPWR VGND sg13g2_fill_1
XFILLER_5_618 VPWR VGND sg13g2_decap_4
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_16_202 VPWR VGND sg13g2_decap_8
XFILLER_17_769 VPWR VGND sg13g2_decap_8
XFILLER_17_83 VPWR VGND sg13g2_decap_8
XFILLER_44_511 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_fill_1
XFILLER_16_279 VPWR VGND sg13g2_decap_8
XFILLER_31_216 VPWR VGND sg13g2_decap_8
XFILLER_33_60 VPWR VGND sg13g2_decap_8
XFILLER_44_599 VPWR VGND sg13g2_fill_2
XFILLER_8_445 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_1490_ VGND VPWR net84 daisychain\[82\] _0562_ net58 sg13g2_a21oi_1
XFILLER_12_4 VPWR VGND sg13g2_decap_4
X_2042_ net187 VGND VPWR _0374_ state\[118\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_35_588 VPWR VGND sg13g2_decap_4
XFILLER_47_371 VPWR VGND sg13g2_decap_8
X_1826_ net204 VGND VPWR _0158_ daisychain\[30\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1757_ _0579_ VPWR _0345_ VGND net155 _0115_ sg13g2_o21ai_1
X_1688_ _0886_ VPWR _0276_ VGND net147 _0040_ sg13g2_o21ai_1
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_13_249 VPWR VGND sg13g2_decap_8
XFILLER_21_271 VPWR VGND sg13g2_decap_8
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_49_603 VPWR VGND sg13g2_decap_8
XFILLER_49_636 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_fill_1
XFILLER_32_547 VPWR VGND sg13g2_decap_4
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_12_293 VPWR VGND sg13g2_decap_8
XFILLER_13_761 VPWR VGND sg13g2_fill_2
XFILLER_8_242 VPWR VGND sg13g2_decap_8
X_1611_ _0241_ _0651_ _0652_ net37 _0814_ VPWR VGND sg13g2_a22oi_1
X_0990_ VPWR _0109_ state\[83\] VGND sg13g2_inv_1
XFILLER_5_53 VPWR VGND sg13g2_decap_8
X_1542_ VGND VPWR net76 daisychain\[95\] _0601_ net42 sg13g2_a21oi_1
X_1473_ _0780_ net128 _0548_ _0549_ VPWR VGND sg13g2_a21o_1
XFILLER_36_820 VPWR VGND sg13g2_fill_2
XFILLER_39_168 VPWR VGND sg13g2_decap_8
X_2025_ net215 VGND VPWR _0357_ state\[101\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_23_503 VPWR VGND sg13g2_fill_2
XFILLER_23_536 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_4
XFILLER_35_385 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
X_1809_ net189 VGND VPWR _0141_ daisychain\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_46_639 VPWR VGND sg13g2_decap_8
XFILLER_10_786 VPWR VGND sg13g2_fill_2
XFILLER_14_62 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_6_702 VPWR VGND sg13g2_fill_1
XFILLER_6_735 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_6_779 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_17_363 VPWR VGND sg13g2_decap_8
XFILLER_17_374 VPWR VGND sg13g2_fill_1
XFILLER_20_528 VPWR VGND sg13g2_decap_8
XFILLER_32_333 VPWR VGND sg13g2_decap_8
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_45_683 VPWR VGND sg13g2_decap_8
X_0973_ VPWR _0090_ state\[66\] VGND sg13g2_inv_1
X_1525_ _0793_ net124 _0587_ _0588_ VPWR VGND sg13g2_a21o_1
X_1456_ net178 VPWR _0536_ VGND net131 state\[75\] sg13g2_o21ai_1
X_1387_ _0185_ _0483_ _0484_ net52 _0758_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
X_2008_ net220 VGND VPWR _0340_ state\[84\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_3_716 VPWR VGND sg13g2_fill_2
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_14_300 VPWR VGND sg13g2_decap_8
XFILLER_14_377 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
Xheichips25_pudding VPWR VGND uio_oe[0] sg13g2_tiehi
X_1310_ VGND VPWR net80 daisychain\[37\] _0427_ net48 sg13g2_a21oi_1
X_1241_ _0722_ net101 _0888_ _0889_ VPWR VGND sg13g2_a21o_1
XFILLER_17_160 VPWR VGND sg13g2_decap_8
XFILLER_24_119 VPWR VGND sg13g2_decap_4
XFILLER_37_447 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
X_1172_ net143 VPWR _0837_ VGND net97 state\[4\] sg13g2_o21ai_1
XFILLER_20_358 VPWR VGND sg13g2_decap_4
XFILLER_32_130 VPWR VGND sg13g2_decap_8
X_0956_ VPWR _0071_ state\[49\] VGND sg13g2_inv_1
XFILLER_28_403 VPWR VGND sg13g2_fill_1
XFILLER_28_414 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
X_1508_ net171 VPWR _0575_ VGND net124 state\[88\] sg13g2_o21ai_1
X_1439_ _0198_ _0522_ _0523_ net64 _0771_ VPWR VGND sg13g2_a22oi_1
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_7_329 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_546 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_14_174 VPWR VGND sg13g2_decap_8
XFILLER_30_667 VPWR VGND sg13g2_fill_1
XFILLER_30_678 VPWR VGND sg13g2_fill_2
XFILLER_42_483 VPWR VGND sg13g2_decap_8
X_1790_ _0678_ VPWR _0378_ VGND net138 _0025_ sg13g2_o21ai_1
XFILLER_6_340 VPWR VGND sg13g2_decap_8
X_1224_ net145 VPWR _0876_ VGND net98 state\[17\] sg13g2_o21ai_1
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_38_767 VPWR VGND sg13g2_decap_8
XFILLER_38_778 VPWR VGND sg13g2_fill_1
X_1155_ net150 VPWR _0824_ VGND net104 state\[0\] sg13g2_o21ai_1
X_1086_ VPWR _0755_ daisychain\[54\] VGND sg13g2_inv_1
XFILLER_20_100 VPWR VGND sg13g2_fill_1
XFILLER_20_133 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
X_1988_ net224 VGND VPWR _0320_ state\[64\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_0939_ VPWR _0053_ state\[32\] VGND sg13g2_inv_1
XFILLER_28_200 VPWR VGND sg13g2_decap_8
XFILLER_28_277 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_24_461 VPWR VGND sg13g2_fill_2
XFILLER_22_62 VPWR VGND sg13g2_fill_1
XFILLER_22_95 VPWR VGND sg13g2_fill_1
XFILLER_3_343 VPWR VGND sg13g2_decap_8
XFILLER_4_822 VPWR VGND sg13g2_fill_1
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_14_8 VPWR VGND sg13g2_fill_1
Xfanout190 net226 net190 VPWR VGND sg13g2_buf_1
XFILLER_19_244 VPWR VGND sg13g2_decap_8
XFILLER_19_288 VPWR VGND sg13g2_decap_8
XFILLER_34_203 VPWR VGND sg13g2_decap_8
XFILLER_35_737 VPWR VGND sg13g2_fill_1
XFILLER_35_759 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_fill_2
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_42_280 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
X_1911_ net196 VGND VPWR _0243_ daisychain\[115\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1842_ net207 VGND VPWR _0174_ daisychain\[46\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1773_ _0627_ VPWR _0361_ VGND net153 _0006_ sg13g2_o21ai_1
XFILLER_38_553 VPWR VGND sg13g2_fill_2
XFILLER_38_575 VPWR VGND sg13g2_fill_2
X_1207_ _0140_ _0862_ _0863_ net26 _0713_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_236 VPWR VGND sg13g2_decap_8
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
X_1138_ VPWR _0807_ daisychain\[106\] VGND sg13g2_inv_1
X_1069_ VPWR _0738_ daisychain\[37\] VGND sg13g2_inv_1
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_16_258 VPWR VGND sg13g2_decap_8
XFILLER_17_62 VPWR VGND sg13g2_decap_8
XFILLER_17_726 VPWR VGND sg13g2_fill_2
XFILLER_32_707 VPWR VGND sg13g2_fill_1
XFILLER_8_424 VPWR VGND sg13g2_decap_8
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
X_2041_ net186 VGND VPWR _0373_ state\[117\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_7_490 VPWR VGND sg13g2_decap_8
X_1825_ net191 VGND VPWR _0157_ daisychain\[29\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1756_ _0576_ VPWR _0344_ VGND net171 _0114_ sg13g2_o21ai_1
XFILLER_38_28 VPWR VGND sg13g2_decap_8
X_1687_ _0883_ VPWR _0275_ VGND net146 _0038_ sg13g2_o21ai_1
XFILLER_26_501 VPWR VGND sg13g2_fill_1
XFILLER_38_350 VPWR VGND sg13g2_decap_8
XFILLER_41_504 VPWR VGND sg13g2_decap_8
XFILLER_13_228 VPWR VGND sg13g2_decap_8
XFILLER_21_250 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_9_700 VPWR VGND sg13g2_fill_1
XFILLER_12_272 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
XFILLER_8_298 VPWR VGND sg13g2_decap_8
X_1610_ VGND VPWR net75 daisychain\[112\] _0652_ net37 sg13g2_a21oi_1
XFILLER_9_788 VPWR VGND sg13g2_fill_2
XFILLER_9_777 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
X_1541_ _0797_ net109 _0599_ _0600_ VPWR VGND sg13g2_a21o_1
X_1472_ net175 VPWR _0548_ VGND net128 state\[79\] sg13g2_o21ai_1
XFILLER_35_364 VPWR VGND sg13g2_decap_8
XFILLER_39_147 VPWR VGND sg13g2_decap_8
X_2024_ net216 VGND VPWR _0356_ state\[100\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1808_ net189 VGND VPWR _0140_ daisychain\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1739_ _0525_ VPWR _0327_ VGND net179 _0096_ sg13g2_o21ai_1
XFILLER_26_342 VPWR VGND sg13g2_decap_8
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_14_41 VPWR VGND sg13g2_decap_8
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_30_95 VPWR VGND sg13g2_decap_8
XFILLER_17_342 VPWR VGND sg13g2_decap_8
XFILLER_45_662 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_32_312 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_decap_4
XFILLER_44_161 VPWR VGND sg13g2_decap_8
X_0972_ VPWR _0089_ state\[65\] VGND sg13g2_inv_1
XFILLER_9_552 VPWR VGND sg13g2_fill_2
X_1524_ net172 VPWR _0587_ VGND net125 state\[92\] sg13g2_o21ai_1
X_1455_ _0202_ _0534_ _0535_ net63 _0775_ VPWR VGND sg13g2_a22oi_1
X_1386_ VGND VPWR net81 daisychain\[56\] _0484_ net52 sg13g2_a21oi_1
XFILLER_35_161 VPWR VGND sg13g2_decap_8
X_2007_ net217 VGND VPWR _0339_ state\[83\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_33_109 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_14_356 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
XFILLER_10_551 VPWR VGND sg13g2_decap_8
XFILLER_6_522 VPWR VGND sg13g2_decap_8
XFILLER_6_566 VPWR VGND sg13g2_fill_2
XFILLER_6_588 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
X_1240_ net147 VPWR _0888_ VGND net101 state\[21\] sg13g2_o21ai_1
X_1171_ _0131_ _0835_ _0836_ net35 _0704_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_37_426 VPWR VGND sg13g2_decap_8
XFILLER_32_186 VPWR VGND sg13g2_decap_8
X_0955_ VPWR _0070_ state\[48\] VGND sg13g2_inv_1
XFILLER_9_382 VPWR VGND sg13g2_decap_8
X_1507_ _0215_ _0573_ _0574_ net59 _0788_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_448 VPWR VGND sg13g2_fill_2
XFILLER_46_28 VPWR VGND sg13g2_decap_8
X_1438_ VGND VPWR net88 daisychain\[69\] _0523_ net64 sg13g2_a21oi_1
X_1369_ _0754_ net119 _0470_ _0471_ VPWR VGND sg13g2_a21o_1
XFILLER_11_326 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_3_525 VPWR VGND sg13g2_decap_8
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xdac dac/VbiasP[1] dac/Iout dac/VbiasP[0] dac/VcascP[1] dac/VcascP[0] state\[64\]
+ _0088_ state\[65\] _0089_ state\[66\] _0090_ state\[67\] _0091_ state\[68\] _0092_
+ state\[69\] _0093_ state\[70\] _0095_ state\[71\] _0096_ state\[72\] _0097_ digitalen.g\[2\].u.OUTP
+ digitalen.g\[2\].u.OUTN state\[73\] _0098_ state\[74\] _0099_ state\[75\] _0100_
+ state\[76\] _0101_ state\[77\] _0102_ state\[78\] _0103_ state\[79\] _0104_ state\[80\]
+ _0106_ state\[81\] _0107_ state\[82\] _0108_ state\[83\] _0109_ state\[84\] _0110_
+ state\[85\] _0111_ state\[86\] _0112_ state\[87\] _0113_ state\[88\] _0114_ state\[89\]
+ _0115_ state\[90\] _0117_ state\[91\] _0118_ state\[92\] _0119_ state\[93\] _0120_
+ state\[94\] _0121_ state\[95\] _0122_ state\[96\] _0123_ state\[97\] _0124_ state\[98\]
+ _0125_ state\[99\] _0126_ state\[100\] _0001_ state\[101\] _0002_ state\[102\] _0003_
+ state\[103\] _0004_ state\[104\] _0005_ state\[105\] _0006_ state\[106\] _0007_
+ state\[107\] _0008_ state\[108\] _0009_ state\[109\] _0010_ state\[110\] _0012_
+ state\[111\] _0013_ state\[112\] _0014_ state\[113\] _0015_ state\[114\] _0016_
+ state\[115\] _0017_ state\[116\] _0018_ state\[117\] _0019_ state\[118\] _0020_
+ state\[119\] _0021_ state\[120\] _0023_ state\[121\] _0024_ state\[122\] _0025_
+ digitalen.g\[3\].u.OUTP digitalen.g\[3\].u.OUTN state\[123\] _0026_ state\[124\]
+ _0027_ state\[125\] _0028_ state\[126\] _0029_ state\[127\] _0030_ state\[0\] _0000_
+ state\[1\] _0039_ state\[2\] _0050_ state\[3\] _0061_ state\[4\] _0072_ state\[5\]
+ _0083_ state\[6\] digitalen.g\[0\].u.OUTP digitalen.g\[0\].u.OUTN _0094_ state\[7\]
+ _0105_ state\[8\] _0116_ state\[9\] _0127_ state\[10\] _0011_ state\[11\] _0022_
+ state\[12\] _0031_ state\[13\] _0032_ state\[14\] _0033_ state\[15\] _0034_ state\[16\]
+ _0035_ state\[17\] _0036_ state\[18\] _0037_ state\[19\] _0038_ state\[20\] _0040_
+ state\[21\] _0041_ state\[22\] _0042_ state\[23\] _0043_ state\[24\] _0044_ state\[25\]
+ _0045_ state\[26\] _0046_ state\[27\] _0047_ state\[28\] _0048_ state\[29\] _0049_
+ state\[30\] _0051_ state\[31\] _0052_ state\[33\] _0054_ state\[32\] _0053_ state\[34\]
+ _0055_ state\[35\] _0056_ state\[36\] _0057_ state\[37\] _0058_ state\[38\] _0059_
+ state\[39\] _0060_ state\[40\] _0062_ state\[41\] _0063_ state\[42\] _0064_ state\[43\]
+ _0065_ state\[44\] _0066_ state\[45\] _0067_ state\[46\] _0068_ state\[47\] _0069_
+ state\[48\] _0070_ state\[49\] _0071_ state\[50\] _0073_ state\[51\] _0074_ state\[52\]
+ _0075_ state\[53\] _0076_ state\[54\] _0077_ state\[55\] _0078_ state\[56\] _0079_
+ state\[57\] _0080_ state\[58\] _0081_ state\[59\] _0082_ state\[60\] _0084_ state\[61\]
+ _0085_ state\[62\] _0086_ state\[63\] _0087_ digitalen.g\[1\].u.OUTP digitalen.g\[1\].u.OUTN
+ VGND VPWR dac128module
XFILLER_34_429 VPWR VGND sg13g2_fill_2
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_14_153 VPWR VGND sg13g2_decap_8
XFILLER_15_698 VPWR VGND sg13g2_fill_2
XFILLER_30_624 VPWR VGND sg13g2_decap_4
XFILLER_42_462 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_decap_8
XFILLER_37_245 VPWR VGND sg13g2_decap_8
X_1223_ _0144_ _0874_ _0875_ net32 _0717_ VPWR VGND sg13g2_a22oi_1
X_1154_ VPWR _0823_ daisychain\[122\] VGND sg13g2_inv_1
XFILLER_20_112 VPWR VGND sg13g2_decap_8
X_1085_ VPWR _0754_ daisychain\[53\] VGND sg13g2_inv_1
XFILLER_20_189 VPWR VGND sg13g2_decap_8
X_1987_ net213 VGND VPWR _0319_ state\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0938_ VPWR _0052_ state\[31\] VGND sg13g2_inv_1
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_28_256 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_44_705 VPWR VGND sg13g2_fill_2
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_12_624 VPWR VGND sg13g2_fill_1
XFILLER_12_679 VPWR VGND sg13g2_decap_8
XFILLER_24_473 VPWR VGND sg13g2_fill_1
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_8_628 VPWR VGND sg13g2_decap_4
XFILLER_8_639 VPWR VGND sg13g2_fill_1
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_3_322 VPWR VGND sg13g2_decap_8
XFILLER_19_223 VPWR VGND sg13g2_decap_8
XFILLER_35_705 VPWR VGND sg13g2_fill_1
XFILLER_3_399 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_decap_8
Xfanout180 net181 net180 VPWR VGND sg13g2_buf_1
Xfanout191 net195 net191 VPWR VGND sg13g2_buf_1
XFILLER_15_462 VPWR VGND sg13g2_decap_4
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_43_782 VPWR VGND sg13g2_decap_4
X_1910_ net196 VGND VPWR _0242_ daisychain\[114\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_30_443 VPWR VGND sg13g2_fill_2
XFILLER_30_465 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
X_1841_ net205 VGND VPWR _0173_ daisychain\[45\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1772_ _0624_ VPWR _0360_ VGND net153 _0005_ sg13g2_o21ai_1
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_25_215 VPWR VGND sg13g2_decap_8
X_1206_ VGND VPWR net68 daisychain\[11\] _0863_ net26 sg13g2_a21oi_1
X_1137_ VPWR _0806_ daisychain\[105\] VGND sg13g2_inv_1
XFILLER_21_410 VPWR VGND sg13g2_decap_4
XFILLER_21_432 VPWR VGND sg13g2_decap_8
XFILLER_21_443 VPWR VGND sg13g2_fill_1
XFILLER_21_465 VPWR VGND sg13g2_fill_2
XFILLER_33_270 VPWR VGND sg13g2_decap_8
X_1068_ VPWR _0737_ daisychain\[36\] VGND sg13g2_inv_1
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_29_532 VPWR VGND sg13g2_fill_2
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_16_237 VPWR VGND sg13g2_decap_8
XFILLER_17_41 VPWR VGND sg13g2_decap_8
XFILLER_17_738 VPWR VGND sg13g2_decap_4
XFILLER_40_730 VPWR VGND sg13g2_decap_8
XFILLER_33_95 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_3_196 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_35_546 VPWR VGND sg13g2_fill_1
XFILLER_39_329 VPWR VGND sg13g2_decap_8
X_2040_ net198 VGND VPWR _0372_ state\[116\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_229 VPWR VGND sg13g2_decap_8
XFILLER_30_284 VPWR VGND sg13g2_decap_8
X_1824_ net191 VGND VPWR _0156_ daisychain\[28\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1755_ _0573_ VPWR _0343_ VGND net173 _0113_ sg13g2_o21ai_1
X_1686_ _0880_ VPWR _0274_ VGND net145 _0037_ sg13g2_o21ai_1
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_26_524 VPWR VGND sg13g2_decap_8
XFILLER_26_535 VPWR VGND sg13g2_fill_2
XFILLER_34_590 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_4
XFILLER_12_251 VPWR VGND sg13g2_decap_8
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
X_1540_ net154 VPWR _0599_ VGND net109 state\[96\] sg13g2_o21ai_1
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
X_1471_ _0206_ _0546_ _0547_ net61 _0779_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_343 VPWR VGND sg13g2_decap_8
XFILLER_36_822 VPWR VGND sg13g2_fill_1
XFILLER_48_660 VPWR VGND sg13g2_fill_1
X_2023_ net200 VGND VPWR _0355_ state\[99\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1807_ net185 VGND VPWR _0139_ daisychain\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_49_39 VPWR VGND sg13g2_decap_8
X_1738_ _0522_ VPWR _0326_ VGND net179 _0095_ sg13g2_o21ai_1
X_1669_ _0829_ VPWR _0257_ VGND net143 _0039_ sg13g2_o21ai_1
XFILLER_14_20 VPWR VGND sg13g2_decap_8
XFILLER_26_387 VPWR VGND sg13g2_decap_8
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_10_755 VPWR VGND sg13g2_decap_8
XFILLER_14_97 VPWR VGND sg13g2_decap_8
XFILLER_30_74 VPWR VGND sg13g2_decap_8
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_6_715 VPWR VGND sg13g2_fill_1
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_17_321 VPWR VGND sg13g2_decap_8
XFILLER_18_811 VPWR VGND sg13g2_decap_8
XFILLER_18_822 VPWR VGND sg13g2_fill_1
XFILLER_29_181 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_13_560 VPWR VGND sg13g2_decap_8
XFILLER_32_368 VPWR VGND sg13g2_decap_8
X_0971_ VPWR _0088_ state\[64\] VGND sg13g2_inv_1
XFILLER_4_291 VPWR VGND sg13g2_decap_8
X_1523_ _0219_ _0585_ _0586_ net59 _0792_ VPWR VGND sg13g2_a22oi_1
X_1454_ VGND VPWR net86 daisychain\[73\] _0535_ net65 sg13g2_a21oi_1
XFILLER_48_490 VPWR VGND sg13g2_decap_8
X_1385_ _0758_ net117 _0482_ _0483_ VPWR VGND sg13g2_a21o_1
XFILLER_23_357 VPWR VGND sg13g2_decap_8
XFILLER_35_140 VPWR VGND sg13g2_decap_8
X_2006_ net225 VGND VPWR _0338_ state\[82\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_3_718 VPWR VGND sg13g2_fill_1
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_39_490 VPWR VGND sg13g2_decap_4
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_14_335 VPWR VGND sg13g2_decap_8
XFILLER_22_390 VPWR VGND sg13g2_fill_1
XFILLER_25_85 VPWR VGND sg13g2_decap_4
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_6_501 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_fill_2
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
X_1170_ VGND VPWR net71 daisychain\[2\] _0836_ net35 sg13g2_a21oi_1
XFILLER_17_195 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_20_316 VPWR VGND sg13g2_decap_8
X_0954_ VPWR _0069_ state\[47\] VGND sg13g2_inv_1
XFILLER_9_361 VPWR VGND sg13g2_decap_8
X_1506_ VGND VPWR net85 daisychain\[86\] _0574_ net59 sg13g2_a21oi_1
X_1437_ _0771_ net132 _0521_ _0522_ VPWR VGND sg13g2_a21o_1
XFILLER_28_438 VPWR VGND sg13g2_fill_2
X_1368_ net165 VPWR _0470_ VGND net118 state\[53\] sg13g2_o21ai_1
X_1299_ _0163_ _0417_ _0418_ net36 _0736_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_305 VPWR VGND sg13g2_decap_8
XFILLER_23_198 VPWR VGND sg13g2_decap_8
XFILLER_36_493 VPWR VGND sg13g2_fill_2
XFILLER_11_32 VPWR VGND sg13g2_decap_8
XFILLER_3_504 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_14_132 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_fill_1
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_42_441 VPWR VGND sg13g2_decap_8
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_fill_1
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_18_460 VPWR VGND sg13g2_decap_4
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
X_1222_ VGND VPWR net71 daisychain\[15\] _0875_ net30 sg13g2_a21oi_1
X_1153_ VPWR _0822_ daisychain\[121\] VGND sg13g2_inv_1
X_1084_ VPWR _0753_ daisychain\[52\] VGND sg13g2_inv_1
XFILLER_33_452 VPWR VGND sg13g2_fill_1
X_1986_ net213 VGND VPWR _0318_ state\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_20_168 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_9_clk clknet_2_0__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_0937_ VPWR _0051_ state\[30\] VGND sg13g2_inv_1
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_44_717 VPWR VGND sg13g2_fill_1
XFILLER_44_728 VPWR VGND sg13g2_decap_4
XFILLER_11_102 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_20_680 VPWR VGND sg13g2_fill_1
XFILLER_22_20 VPWR VGND sg13g2_decap_8
XFILLER_22_31 VPWR VGND sg13g2_fill_1
XFILLER_3_301 VPWR VGND sg13g2_decap_8
XFILLER_3_378 VPWR VGND sg13g2_decap_8
XFILLER_19_202 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
Xfanout170 net174 net170 VPWR VGND sg13g2_buf_1
Xfanout181 net182 net181 VPWR VGND sg13g2_buf_1
Xfanout192 net195 net192 VPWR VGND sg13g2_buf_1
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
X_1840_ net205 VGND VPWR _0172_ daisychain\[44\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_6_172 VPWR VGND sg13g2_decap_8
XFILLER_7_684 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_1771_ _0621_ VPWR _0359_ VGND net156 _0004_ sg13g2_o21ai_1
X_1205_ _0713_ net93 _0861_ _0862_ VPWR VGND sg13g2_a21o_1
X_1136_ VPWR _0805_ daisychain\[104\] VGND sg13g2_inv_1
X_1067_ VPWR _0736_ daisychain\[35\] VGND sg13g2_inv_1
X_1969_ net211 VGND VPWR _0301_ state\[45\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_8
XFILLER_17_20 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_12_433 VPWR VGND sg13g2_decap_8
XFILLER_16_216 VPWR VGND sg13g2_decap_8
XFILLER_17_97 VPWR VGND sg13g2_decap_8
XFILLER_24_282 VPWR VGND sg13g2_decap_8
XFILLER_44_525 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_decap_8
XFILLER_8_459 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_48_820 VPWR VGND sg13g2_fill_2
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_15_293 VPWR VGND sg13g2_decap_8
XFILLER_22_208 VPWR VGND sg13g2_decap_8
XFILLER_30_263 VPWR VGND sg13g2_decap_8
XFILLER_31_786 VPWR VGND sg13g2_fill_1
X_1823_ net191 VGND VPWR _0155_ daisychain\[27\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1754_ _0570_ VPWR _0342_ VGND net172 _0112_ sg13g2_o21ai_1
X_1685_ _0877_ VPWR _0273_ VGND net145 _0036_ sg13g2_o21ai_1
XFILLER_38_385 VPWR VGND sg13g2_decap_8
X_1119_ VPWR _0788_ daisychain\[87\] VGND sg13g2_inv_1
XFILLER_21_285 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_12_230 VPWR VGND sg13g2_decap_8
XFILLER_13_720 VPWR VGND sg13g2_fill_2
XFILLER_40_572 VPWR VGND sg13g2_decap_8
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_9_724 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_8
X_1470_ VGND VPWR net87 daisychain\[77\] _0547_ net61 sg13g2_a21oi_1
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_35_399 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
X_2022_ net201 VGND VPWR _0354_ state\[98\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1806_ net185 VGND VPWR _0138_ daisychain\[10\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
X_1737_ _0519_ VPWR _0325_ VGND net179 _0093_ sg13g2_o21ai_1
X_1668_ _0825_ VPWR _0256_ VGND net150 _0000_ sg13g2_o21ai_1
X_1599_ _0238_ _0642_ _0643_ net40 _0811_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_14_76 VPWR VGND sg13g2_decap_8
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_17_300 VPWR VGND sg13g2_decap_8
XFILLER_29_160 VPWR VGND sg13g2_decap_8
XFILLER_32_347 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
XFILLER_45_697 VPWR VGND sg13g2_decap_4
XFILLER_20_509 VPWR VGND sg13g2_fill_1
X_0970_ VPWR _0087_ state\[63\] VGND sg13g2_inv_1
XFILLER_9_587 VPWR VGND sg13g2_decap_8
XFILLER_4_270 VPWR VGND sg13g2_decap_8
X_1522_ VGND VPWR net84 daisychain\[90\] _0586_ net57 sg13g2_a21oi_1
X_1453_ _0775_ net130 _0533_ _0534_ VPWR VGND sg13g2_a21o_1
XFILLER_27_108 VPWR VGND sg13g2_fill_2
X_2005_ net215 VGND VPWR _0337_ state\[81\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1384_ net164 VPWR _0482_ VGND net117 state\[57\] sg13g2_o21ai_1
XFILLER_23_303 VPWR VGND sg13g2_decap_4
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_14_314 VPWR VGND sg13g2_decap_8
XFILLER_42_601 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_4
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_2_730 VPWR VGND sg13g2_decap_4
XFILLER_18_642 VPWR VGND sg13g2_fill_1
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_37_406 VPWR VGND sg13g2_fill_1
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_17_174 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_decap_8
X_0953_ VPWR _0068_ state\[46\] VGND sg13g2_inv_1
XFILLER_9_340 VPWR VGND sg13g2_decap_8
X_1505_ _0788_ net126 _0572_ _0573_ VPWR VGND sg13g2_a21o_1
X_1436_ net178 VPWR _0521_ VGND net132 state\[70\] sg13g2_o21ai_1
X_1367_ _0180_ _0468_ _0469_ net51 _0753_ VPWR VGND sg13g2_a22oi_1
X_1298_ VGND VPWR net73 daisychain\[34\] _0418_ net34 sg13g2_a21oi_1
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_14_111 VPWR VGND sg13g2_decap_8
XFILLER_14_188 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_42_420 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_30_648 VPWR VGND sg13g2_fill_2
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_2_593 VPWR VGND sg13g2_fill_2
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_1221_ _0717_ net98 _0873_ _0874_ VPWR VGND sg13g2_a21o_1
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_38_715 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
X_1152_ VPWR _0821_ daisychain\[120\] VGND sg13g2_inv_1
X_1083_ VPWR _0752_ daisychain\[51\] VGND sg13g2_inv_1
XFILLER_20_147 VPWR VGND sg13g2_decap_8
X_1985_ net213 VGND VPWR _0317_ state\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_0936_ VPWR _0049_ state\[29\] VGND sg13g2_inv_1
XFILLER_28_214 VPWR VGND sg13g2_decap_8
X_1419_ _0193_ _0507_ _0508_ net62 _0766_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_44_707 VPWR VGND sg13g2_fill_1
XFILLER_11_158 VPWR VGND sg13g2_decap_8
XFILLER_3_357 VPWR VGND sg13g2_decap_8
XFILLER_19_258 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_578 VPWR VGND sg13g2_fill_1
XFILLER_47_84 VPWR VGND sg13g2_decap_8
Xfanout160 net169 net160 VPWR VGND sg13g2_buf_1
Xfanout171 net173 net171 VPWR VGND sg13g2_buf_1
Xfanout182 net4 net182 VPWR VGND sg13g2_buf_1
Xfanout193 net195 net193 VPWR VGND sg13g2_buf_1
XFILLER_15_442 VPWR VGND sg13g2_fill_1
XFILLER_27_291 VPWR VGND sg13g2_decap_8
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
X_1770_ _0618_ VPWR _0358_ VGND net170 _0003_ sg13g2_o21ai_1
XFILLER_6_151 VPWR VGND sg13g2_decap_8
XFILLER_38_534 VPWR VGND sg13g2_fill_2
X_1204_ net142 VPWR _0861_ VGND net96 state\[12\] sg13g2_o21ai_1
XFILLER_18_291 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[0\].u.inv1 VPWR digitalen.g\[0\].u.OUTN net6 VGND sg13g2_inv_1
X_1135_ VPWR _0804_ daisychain\[103\] VGND sg13g2_inv_1
X_1066_ VPWR _0735_ daisychain\[34\] VGND sg13g2_inv_1
XFILLER_21_489 VPWR VGND sg13g2_fill_1
X_1968_ net211 VGND VPWR _0300_ state\[44\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1899_ net200 VGND VPWR _0231_ daisychain\[103\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_0919_ VPWR _0031_ state\[12\] VGND sg13g2_inv_1
XFILLER_29_534 VPWR VGND sg13g2_fill_1
XFILLER_44_504 VPWR VGND sg13g2_decap_8
XFILLER_12_412 VPWR VGND sg13g2_decap_8
XFILLER_12_456 VPWR VGND sg13g2_fill_1
XFILLER_17_76 VPWR VGND sg13g2_decap_8
XFILLER_24_261 VPWR VGND sg13g2_decap_8
XFILLER_31_209 VPWR VGND sg13g2_decap_8
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_40_765 VPWR VGND sg13g2_fill_2
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_8_438 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_1
XFILLER_16_762 VPWR VGND sg13g2_fill_1
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_15_272 VPWR VGND sg13g2_decap_8
XFILLER_30_242 VPWR VGND sg13g2_decap_8
X_1822_ net191 VGND VPWR _0154_ daisychain\[26\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1753_ _0567_ VPWR _0341_ VGND net172 _0111_ sg13g2_o21ai_1
X_1684_ _0874_ VPWR _0272_ VGND net142 _0035_ sg13g2_o21ai_1
XFILLER_38_364 VPWR VGND sg13g2_decap_8
XFILLER_21_264 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_fill_2
X_1118_ VPWR _0787_ daisychain\[86\] VGND sg13g2_inv_1
X_1049_ VPWR _0718_ daisychain\[17\] VGND sg13g2_inv_1
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_29_342 VPWR VGND sg13g2_fill_2
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
XFILLER_12_286 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_36_813 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
X_2021_ net202 VGND VPWR _0353_ state\[97\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_35_378 VPWR VGND sg13g2_decap_8
X_1805_ net185 VGND VPWR _0137_ daisychain\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1736_ _0516_ VPWR _0324_ VGND net178 _0092_ sg13g2_o21ai_1
X_1667_ _0255_ _0693_ _0694_ net24 _0700_ VPWR VGND sg13g2_a22oi_1
X_1598_ VGND VPWR net77 daisychain\[109\] _0643_ net40 sg13g2_a21oi_1
XFILLER_26_356 VPWR VGND sg13g2_decap_4
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_39_695 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
XFILLER_42_816 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_fill_1
XFILLER_10_768 VPWR VGND sg13g2_fill_1
XFILLER_10_779 VPWR VGND sg13g2_decap_8
XFILLER_14_55 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_6_728 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_17_356 VPWR VGND sg13g2_decap_8
XFILLER_32_326 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_45_676 VPWR VGND sg13g2_decap_8
XFILLER_13_573 VPWR VGND sg13g2_fill_1
XFILLER_40_392 VPWR VGND sg13g2_decap_8
X_1521_ _0792_ net126 _0584_ _0585_ VPWR VGND sg13g2_a21o_1
X_1452_ net178 VPWR _0533_ VGND net131 state\[74\] sg13g2_o21ai_1
X_1383_ _0184_ _0480_ _0481_ net50 _0757_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_610 VPWR VGND sg13g2_decap_4
X_2004_ net215 VGND VPWR _0336_ state\[80\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_35_175 VPWR VGND sg13g2_decap_8
X_1719_ _0465_ VPWR _0307_ VGND net167 _0074_ sg13g2_o21ai_1
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_4
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_42_657 VPWR VGND sg13g2_fill_1
XFILLER_22_381 VPWR VGND sg13g2_fill_2
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_17_153 VPWR VGND sg13g2_decap_8
XFILLER_18_687 VPWR VGND sg13g2_decap_4
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_32_123 VPWR VGND sg13g2_decap_8
XFILLER_33_635 VPWR VGND sg13g2_fill_1
XFILLER_33_679 VPWR VGND sg13g2_fill_2
X_0952_ VPWR _0067_ state\[45\] VGND sg13g2_inv_1
X_1504_ net172 VPWR _0572_ VGND net125 state\[87\] sg13g2_o21ai_1
XFILLER_9_396 VPWR VGND sg13g2_decap_8
XFILLER_28_407 VPWR VGND sg13g2_decap_8
X_1435_ _0197_ _0519_ _0520_ net64 _0770_ VPWR VGND sg13g2_a22oi_1
X_1366_ VGND VPWR net81 daisychain\[51\] _0469_ net51 sg13g2_a21oi_1
XFILLER_23_101 VPWR VGND sg13g2_fill_2
X_1297_ _0736_ net103 _0416_ _0417_ VPWR VGND sg13g2_a21o_1
XFILLER_11_67 VPWR VGND sg13g2_decap_8
XFILLER_3_539 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_14_167 VPWR VGND sg13g2_decap_8
XFILLER_30_605 VPWR VGND sg13g2_decap_4
XFILLER_42_476 VPWR VGND sg13g2_decap_8
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
X_1220_ net142 VPWR _0873_ VGND net96 state\[16\] sg13g2_o21ai_1
X_1151_ VPWR _0820_ daisychain\[119\] VGND sg13g2_inv_1
XFILLER_18_440 VPWR VGND sg13g2_fill_1
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_46_782 VPWR VGND sg13g2_decap_4
X_1082_ VPWR _0751_ daisychain\[50\] VGND sg13g2_inv_1
XFILLER_20_126 VPWR VGND sg13g2_decap_8
XFILLER_33_487 VPWR VGND sg13g2_decap_4
X_1984_ net210 VGND VPWR _0316_ state\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_0935_ VPWR _0048_ state\[28\] VGND sg13g2_inv_1
XFILLER_9_193 VPWR VGND sg13g2_decap_8
X_1418_ VGND VPWR net87 daisychain\[64\] _0508_ net62 sg13g2_a21oi_1
X_1349_ _0749_ net116 _0455_ _0456_ VPWR VGND sg13g2_a21o_1
XFILLER_11_137 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_3_336 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
Xfanout150 net151 net150 VPWR VGND sg13g2_buf_1
Xfanout161 net169 net161 VPWR VGND sg13g2_buf_1
Xfanout172 net173 net172 VPWR VGND sg13g2_buf_1
Xfanout183 net227 net183 VPWR VGND sg13g2_buf_1
XFILLER_15_454 VPWR VGND sg13g2_fill_2
XFILLER_19_237 VPWR VGND sg13g2_decap_8
XFILLER_27_270 VPWR VGND sg13g2_decap_8
XFILLER_43_752 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
Xfanout194 net195 net194 VPWR VGND sg13g2_buf_1
XFILLER_30_413 VPWR VGND sg13g2_fill_2
XFILLER_30_479 VPWR VGND sg13g2_decap_8
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_6_130 VPWR VGND sg13g2_decap_8
XFILLER_33_4 VPWR VGND sg13g2_decap_8
XFILLER_38_546 VPWR VGND sg13g2_decap_8
X_1203_ _0139_ _0859_ _0860_ net26 _0712_ VPWR VGND sg13g2_a22oi_1
X_1134_ VPWR _0803_ daisychain\[102\] VGND sg13g2_inv_1
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_25_229 VPWR VGND sg13g2_decap_8
XFILLER_33_284 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[0\].u.inv2 VPWR digitalen.g\[0\].u.OUTP digitalen.g\[0\].u.OUTN VGND
+ sg13g2_inv_1
X_1065_ VPWR _0734_ daisychain\[33\] VGND sg13g2_inv_1
X_1967_ net211 VGND VPWR _0299_ state\[43\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1898_ net199 VGND VPWR _0230_ daisychain\[102\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_0918_ VPWR _0022_ state\[11\] VGND sg13g2_inv_1
XFILLER_17_55 VPWR VGND sg13g2_decap_8
XFILLER_24_240 VPWR VGND sg13g2_decap_8
XFILLER_33_32 VPWR VGND sg13g2_decap_8
XFILLER_40_744 VPWR VGND sg13g2_fill_2
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_fill_1
XFILLER_15_251 VPWR VGND sg13g2_decap_8
XFILLER_30_221 VPWR VGND sg13g2_decap_8
XFILLER_30_298 VPWR VGND sg13g2_decap_8
XFILLER_7_483 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_2_0__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_1821_ net191 VGND VPWR _0153_ daisychain\[25\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1752_ _0564_ VPWR _0340_ VGND net172 _0110_ sg13g2_o21ai_1
X_1683_ _0871_ VPWR _0271_ VGND net143 _0034_ sg13g2_o21ai_1
XFILLER_38_343 VPWR VGND sg13g2_decap_8
X_1117_ VPWR _0786_ daisychain\[85\] VGND sg13g2_inv_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_21_243 VPWR VGND sg13g2_decap_8
X_1048_ VPWR _0717_ daisychain\[16\] VGND sg13g2_inv_1
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_321 VPWR VGND sg13g2_decap_8
XFILLER_17_527 VPWR VGND sg13g2_fill_2
XFILLER_32_508 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_12_265 VPWR VGND sg13g2_decap_8
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
X_2020_ net202 VGND VPWR _0352_ state\[96\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_35_357 VPWR VGND sg13g2_decap_8
XFILLER_7_280 VPWR VGND sg13g2_decap_8
X_1804_ net185 VGND VPWR _0136_ daisychain\[8\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1735_ _0513_ VPWR _0323_ VGND net178 _0091_ sg13g2_o21ai_1
X_1666_ VGND VPWR net70 daisychain\[126\] _0694_ net24 sg13g2_a21oi_1
X_1597_ _0811_ net107 _0641_ _0642_ VPWR VGND sg13g2_a21o_1
XFILLER_38_140 VPWR VGND sg13g2_decap_8
XFILLER_14_34 VPWR VGND sg13g2_decap_8
XFILLER_22_530 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_30_88 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_17_335 VPWR VGND sg13g2_decap_8
XFILLER_29_195 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_32_305 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_44_154 VPWR VGND sg13g2_decap_8
X_1520_ net172 VPWR _0584_ VGND net126 state\[91\] sg13g2_o21ai_1
X_1451_ _0201_ _0531_ _0532_ net65 _0774_ VPWR VGND sg13g2_a22oi_1
X_1382_ VGND VPWR net81 daisychain\[55\] _0481_ net50 sg13g2_a21oi_1
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_36_622 VPWR VGND sg13g2_fill_2
XFILLER_36_644 VPWR VGND sg13g2_fill_2
X_2003_ net219 VGND VPWR _0335_ state\[79\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_1718_ _0462_ VPWR _0306_ VGND net167 _0073_ sg13g2_o21ai_1
X_1649_ net90 _0695_ _0680_ _0681_ VPWR VGND sg13g2_a21o_1
XFILLER_14_349 VPWR VGND sg13g2_decap_8
XFILLER_15_817 VPWR VGND sg13g2_decap_4
XFILLER_22_360 VPWR VGND sg13g2_decap_8
XFILLER_25_44 VPWR VGND sg13g2_decap_4
XFILLER_26_132 VPWR VGND sg13g2_fill_1
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_42_669 VPWR VGND sg13g2_decap_4
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_6_515 VPWR VGND sg13g2_decap_8
XFILLER_6_559 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_fill_1
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_17_132 VPWR VGND sg13g2_decap_8
XFILLER_18_611 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_37_419 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_41_680 VPWR VGND sg13g2_decap_4
XFILLER_41_691 VPWR VGND sg13g2_fill_2
X_0951_ VPWR _0066_ state\[44\] VGND sg13g2_inv_1
XFILLER_9_375 VPWR VGND sg13g2_decap_8
X_1503_ _0214_ _0570_ _0571_ net58 _0787_ VPWR VGND sg13g2_a22oi_1
X_1434_ VGND VPWR net86 daisychain\[68\] _0520_ net64 sg13g2_a21oi_1
X_1365_ _0753_ net118 _0467_ _0468_ VPWR VGND sg13g2_a21o_1
X_1296_ net161 VPWR _0416_ VGND net102 state\[35\] sg13g2_o21ai_1
XFILLER_11_319 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_11_46 VPWR VGND sg13g2_decap_8
XFILLER_32_691 VPWR VGND sg13g2_fill_2
XFILLER_3_518 VPWR VGND sg13g2_decap_8
XFILLER_27_485 VPWR VGND sg13g2_fill_2
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_14_146 VPWR VGND sg13g2_decap_8
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_42_455 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_2_595 VPWR VGND sg13g2_fill_1
XFILLER_37_238 VPWR VGND sg13g2_decap_8
X_1150_ VPWR _0819_ daisychain\[118\] VGND sg13g2_inv_1
XFILLER_20_105 VPWR VGND sg13g2_decap_8
X_1081_ VPWR _0750_ daisychain\[49\] VGND sg13g2_inv_1
X_1983_ net210 VGND VPWR _0315_ state\[59\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_0934_ VPWR _0047_ state\[27\] VGND sg13g2_inv_1
XFILLER_9_172 VPWR VGND sg13g2_decap_8
X_1417_ _0766_ net129 _0506_ _0507_ VPWR VGND sg13g2_a21o_1
XFILLER_28_249 VPWR VGND sg13g2_decap_8
XFILLER_37_772 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_decap_8
X_1348_ net162 VPWR _0455_ VGND net116 state\[48\] sg13g2_o21ai_1
X_1279_ _0158_ _0402_ _0403_ net45 _0731_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_116 VPWR VGND sg13g2_decap_8
XFILLER_20_661 VPWR VGND sg13g2_decap_8
XFILLER_3_315 VPWR VGND sg13g2_decap_8
XFILLER_19_216 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
Xfanout140 net141 net140 VPWR VGND sg13g2_buf_1
Xfanout151 net152 net151 VPWR VGND sg13g2_buf_1
Xfanout162 net169 net162 VPWR VGND sg13g2_buf_1
Xfanout173 net174 net173 VPWR VGND sg13g2_buf_1
Xfanout184 net227 net184 VPWR VGND sg13g2_buf_1
Xfanout195 net226 net195 VPWR VGND sg13g2_buf_1
XFILLER_15_466 VPWR VGND sg13g2_fill_2
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_43_786 VPWR VGND sg13g2_fill_2
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_11_694 VPWR VGND sg13g2_fill_2
XFILLER_30_458 VPWR VGND sg13g2_decap_8
XFILLER_7_621 VPWR VGND sg13g2_decap_4
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_6_186 VPWR VGND sg13g2_decap_8
XFILLER_7_698 VPWR VGND sg13g2_fill_2
XFILLER_25_208 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_fill_2
X_1202_ VGND VPWR net68 daisychain\[10\] _0860_ net26 sg13g2_a21oi_1
X_1133_ VPWR _0802_ daisychain\[101\] VGND sg13g2_inv_1
X_1064_ VPWR _0733_ daisychain\[32\] VGND sg13g2_inv_1
XFILLER_21_403 VPWR VGND sg13g2_decap_8
XFILLER_21_414 VPWR VGND sg13g2_fill_1
XFILLER_21_425 VPWR VGND sg13g2_decap_8
XFILLER_21_458 VPWR VGND sg13g2_decap_8
XFILLER_33_263 VPWR VGND sg13g2_decap_8
XFILLER_34_742 VPWR VGND sg13g2_fill_1
X_1966_ net205 VGND VPWR _0298_ state\[42\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1897_ net215 VGND VPWR _0229_ daisychain\[101\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_0917_ VPWR _0011_ state\[10\] VGND sg13g2_inv_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_4
XFILLER_29_525 VPWR VGND sg13g2_fill_2
XFILLER_17_34 VPWR VGND sg13g2_decap_8
XFILLER_24_296 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_decap_8
XFILLER_40_767 VPWR VGND sg13g2_fill_1
XFILLER_40_778 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_35_528 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_15_230 VPWR VGND sg13g2_decap_8
XFILLER_30_200 VPWR VGND sg13g2_decap_8
XFILLER_31_767 VPWR VGND sg13g2_decap_4
XFILLER_47_399 VPWR VGND sg13g2_decap_8
X_1820_ net194 VGND VPWR _0152_ daisychain\[24\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_30_277 VPWR VGND sg13g2_decap_8
XFILLER_7_462 VPWR VGND sg13g2_decap_8
X_1751_ _0561_ VPWR _0339_ VGND net172 _0109_ sg13g2_o21ai_1
X_1682_ _0868_ VPWR _0270_ VGND net143 _0033_ sg13g2_o21ai_1
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_38_399 VPWR VGND sg13g2_decap_8
X_1116_ VPWR _0785_ daisychain\[84\] VGND sg13g2_inv_1
X_1047_ VPWR _0716_ daisychain\[15\] VGND sg13g2_inv_1
XFILLER_21_222 VPWR VGND sg13g2_decap_8
XFILLER_34_583 VPWR VGND sg13g2_decap_8
X_1949_ net194 VGND VPWR _0281_ state\[25\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_29_300 VPWR VGND sg13g2_decap_8
XFILLER_29_344 VPWR VGND sg13g2_fill_1
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_12_244 VPWR VGND sg13g2_decap_8
XFILLER_13_756 VPWR VGND sg13g2_fill_1
XFILLER_13_767 VPWR VGND sg13g2_decap_4
XFILLER_40_531 VPWR VGND sg13g2_fill_2
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_40_586 VPWR VGND sg13g2_fill_2
XFILLER_4_410 VPWR VGND sg13g2_decap_8
XFILLER_0_671 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
X_1803_ net185 VGND VPWR _0135_ daisychain\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1734_ _0510_ VPWR _0322_ VGND net176 _0090_ sg13g2_o21ai_1
X_1665_ _0700_ net91 _0692_ _0693_ VPWR VGND sg13g2_a21o_1
X_1596_ net153 VPWR _0641_ VGND net107 state\[110\] sg13g2_o21ai_1
XFILLER_14_13 VPWR VGND sg13g2_decap_8
XFILLER_26_369 VPWR VGND sg13g2_decap_8
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_30_67 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_17_314 VPWR VGND sg13g2_decap_8
XFILLER_18_804 VPWR VGND sg13g2_decap_8
XFILLER_29_174 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_45_623 VPWR VGND sg13g2_decap_8
XFILLER_13_553 VPWR VGND sg13g2_decap_8
XFILLER_25_380 VPWR VGND sg13g2_fill_2
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_decap_8
X_1450_ VGND VPWR net86 daisychain\[72\] _0532_ net63 sg13g2_a21oi_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
X_1381_ _0757_ net117 _0479_ _0480_ VPWR VGND sg13g2_a21o_1
XFILLER_16_391 VPWR VGND sg13g2_decap_4
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
X_2002_ net219 VGND VPWR _0334_ state\[78\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1717_ _0459_ VPWR _0305_ VGND net167 _0071_ sg13g2_o21ai_1
X_1648_ net138 VPWR _0680_ VGND net90 state\[123\] sg13g2_o21ai_1
X_1579_ _0233_ _0627_ _0628_ net40 _0806_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_111 VPWR VGND sg13g2_decap_8
XFILLER_39_483 VPWR VGND sg13g2_decap_8
XFILLER_14_328 VPWR VGND sg13g2_decap_8
XFILLER_22_394 VPWR VGND sg13g2_decap_8
XFILLER_25_89 VPWR VGND sg13g2_fill_1
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_42_615 VPWR VGND sg13g2_decap_4
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_17_111 VPWR VGND sg13g2_decap_8
XFILLER_17_188 VPWR VGND sg13g2_decap_8
XFILLER_33_648 VPWR VGND sg13g2_decap_4
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_45_497 VPWR VGND sg13g2_decap_8
XFILLER_13_361 VPWR VGND sg13g2_decap_8
XFILLER_20_309 VPWR VGND sg13g2_decap_8
XFILLER_32_158 VPWR VGND sg13g2_decap_8
X_0950_ VPWR _0065_ state\[43\] VGND sg13g2_inv_1
XFILLER_9_354 VPWR VGND sg13g2_decap_8
X_1502_ VGND VPWR net84 daisychain\[85\] _0571_ net58 sg13g2_a21oi_1
X_1433_ _0770_ net131 _0518_ _0519_ VPWR VGND sg13g2_a21o_1
XFILLER_48_280 VPWR VGND sg13g2_decap_8
X_1364_ net164 VPWR _0467_ VGND net118 state\[52\] sg13g2_o21ai_1
X_1295_ _0162_ _0414_ _0415_ net36 _0735_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_810 VPWR VGND sg13g2_fill_1
XFILLER_23_103 VPWR VGND sg13g2_fill_1
XFILLER_11_25 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_decap_8
XFILLER_15_659 VPWR VGND sg13g2_decap_4
XFILLER_27_431 VPWR VGND sg13g2_fill_1
XFILLER_27_464 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_42_434 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_11_821 VPWR VGND sg13g2_fill_2
XFILLER_22_180 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_18_453 VPWR VGND sg13g2_decap_8
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_38_729 VPWR VGND sg13g2_fill_1
X_1080_ VPWR _0749_ daisychain\[48\] VGND sg13g2_inv_1
XFILLER_18_464 VPWR VGND sg13g2_fill_2
XFILLER_45_294 VPWR VGND sg13g2_decap_8
X_1982_ net209 VGND VPWR _0314_ state\[58\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_0933_ VPWR _0046_ state\[26\] VGND sg13g2_inv_1
XFILLER_9_151 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_1416_ net175 VPWR _0506_ VGND net129 state\[65\] sg13g2_o21ai_1
X_1347_ _0175_ _0453_ _0454_ net49 _0748_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
X_1278_ VGND VPWR net72 daisychain\[29\] _0403_ net33 sg13g2_a21oi_1
XFILLER_22_13 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
Xfanout130 net133 net130 VPWR VGND sg13g2_buf_1
Xfanout141 net182 net141 VPWR VGND sg13g2_buf_1
Xfanout152 net157 net152 VPWR VGND sg13g2_buf_1
Xfanout163 net166 net163 VPWR VGND sg13g2_buf_1
Xfanout174 net181 net174 VPWR VGND sg13g2_buf_1
Xfanout185 net187 net185 VPWR VGND sg13g2_buf_1
Xfanout196 net198 net196 VPWR VGND sg13g2_buf_1
XFILLER_15_412 VPWR VGND sg13g2_decap_8
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_12_90 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_2_382 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
X_1201_ _0712_ net93 _0858_ _0859_ VPWR VGND sg13g2_a21o_1
XFILLER_19_4 VPWR VGND sg13g2_decap_4
X_1132_ VPWR _0801_ daisychain\[100\] VGND sg13g2_inv_1
X_1063_ VPWR _0732_ daisychain\[31\] VGND sg13g2_inv_1
XFILLER_33_242 VPWR VGND sg13g2_decap_8
X_1965_ net205 VGND VPWR _0297_ state\[41\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_0916_ VPWR _0127_ state\[9\] VGND sg13g2_inv_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_1896_ net216 VGND VPWR _0228_ daisychain\[100\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_17_13 VPWR VGND sg13g2_decap_8
XFILLER_29_504 VPWR VGND sg13g2_fill_2
XFILLER_12_426 VPWR VGND sg13g2_decap_8
XFILLER_16_209 VPWR VGND sg13g2_decap_8
XFILLER_24_275 VPWR VGND sg13g2_decap_8
XFILLER_40_724 VPWR VGND sg13g2_fill_2
XFILLER_44_518 VPWR VGND sg13g2_decap_8
XFILLER_12_448 VPWR VGND sg13g2_decap_4
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_15_286 VPWR VGND sg13g2_decap_8
XFILLER_30_256 VPWR VGND sg13g2_decap_8
X_1750_ _0558_ VPWR _0338_ VGND net174 _0108_ sg13g2_o21ai_1
XFILLER_7_441 VPWR VGND sg13g2_decap_8
X_1681_ _0865_ VPWR _0269_ VGND net142 _0032_ sg13g2_o21ai_1
XFILLER_38_301 VPWR VGND sg13g2_decap_8
XFILLER_21_201 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_decap_8
X_1115_ VPWR _0784_ daisychain\[83\] VGND sg13g2_inv_1
X_1046_ VPWR _0715_ daisychain\[14\] VGND sg13g2_inv_1
XFILLER_21_278 VPWR VGND sg13g2_decap_8
X_1948_ net194 VGND VPWR _0280_ state\[24\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1879_ net217 VGND VPWR _0211_ daisychain\[83\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_1_628 VPWR VGND sg13g2_fill_2
XFILLER_17_529 VPWR VGND sg13g2_fill_1
XFILLER_28_67 VPWR VGND sg13g2_decap_4
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_12_223 VPWR VGND sg13g2_decap_8
XFILLER_13_702 VPWR VGND sg13g2_decap_8
XFILLER_13_713 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_9_717 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_0_650 VPWR VGND sg13g2_decap_8
XFILLER_16_551 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_392 VPWR VGND sg13g2_decap_8
X_1802_ net186 VGND VPWR _0134_ daisychain\[6\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1733_ _0507_ VPWR _0321_ VGND net176 _0089_ sg13g2_o21ai_1
X_1664_ net137 VPWR _0692_ VGND net91 state\[127\] sg13g2_o21ai_1
X_1595_ _0237_ _0639_ _0640_ net40 _0810_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_14_69 VPWR VGND sg13g2_decap_8
XFILLER_34_392 VPWR VGND sg13g2_decap_8
XFILLER_41_329 VPWR VGND sg13g2_decap_8
X_1029_ VPWR _0025_ state\[122\] VGND sg13g2_inv_1
XFILLER_30_46 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_13_510 VPWR VGND sg13g2_decap_8
XFILLER_29_153 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_4_263 VPWR VGND sg13g2_decap_8
X_1380_ net164 VPWR _0479_ VGND net117 state\[56\] sg13g2_o21ai_1
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_36_646 VPWR VGND sg13g2_fill_1
XFILLER_48_462 VPWR VGND sg13g2_decap_8
X_2001_ net219 VGND VPWR _0333_ state\[77\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_16_370 VPWR VGND sg13g2_decap_8
XFILLER_23_307 VPWR VGND sg13g2_fill_1
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_44_690 VPWR VGND sg13g2_fill_2
X_1716_ _0456_ VPWR _0304_ VGND net162 _0070_ sg13g2_o21ai_1
XFILLER_6_81 VPWR VGND sg13g2_decap_8
X_1647_ _0250_ _0678_ _0679_ net23 _0823_ VPWR VGND sg13g2_a22oi_1
X_1578_ VGND VPWR net77 daisychain\[104\] _0628_ net40 sg13g2_a21oi_1
XFILLER_14_307 VPWR VGND sg13g2_decap_8
XFILLER_39_462 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_723 VPWR VGND sg13g2_decap_8
XFILLER_2_734 VPWR VGND sg13g2_fill_2
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_18_624 VPWR VGND sg13g2_decap_4
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_17_167 VPWR VGND sg13g2_decap_8
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_33_627 VPWR VGND sg13g2_fill_1
XFILLER_45_476 VPWR VGND sg13g2_decap_8
XFILLER_15_90 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
XFILLER_49_4 VPWR VGND sg13g2_decap_8
X_1501_ _0787_ net125 _0569_ _0570_ VPWR VGND sg13g2_a21o_1
X_1432_ net178 VPWR _0518_ VGND net131 state\[69\] sg13g2_o21ai_1
X_1363_ _0179_ _0465_ _0466_ net54 _0752_ VPWR VGND sg13g2_a22oi_1
X_1294_ VGND VPWR net73 daisychain\[33\] _0415_ net33 sg13g2_a21oi_1
XFILLER_31_181 VPWR VGND sg13g2_decap_8
XFILLER_32_671 VPWR VGND sg13g2_decap_4
Xdigitalen.g\[3\].u.inv1 VPWR digitalen.g\[3\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_14_104 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_2_586 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_46_741 VPWR VGND sg13g2_fill_2
XFILLER_18_498 VPWR VGND sg13g2_fill_2
XFILLER_41_490 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_9_130 VPWR VGND sg13g2_decap_8
X_1981_ net209 VGND VPWR _0313_ state\[57\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_0932_ VPWR _0045_ state\[25\] VGND sg13g2_inv_1
XFILLER_28_207 VPWR VGND sg13g2_decap_8
X_1415_ _0192_ _0504_ _0505_ net61 _0765_ VPWR VGND sg13g2_a22oi_1
X_1346_ VGND VPWR net80 daisychain\[46\] _0454_ net48 sg13g2_a21oi_1
XFILLER_24_457 VPWR VGND sg13g2_decap_4
XFILLER_36_273 VPWR VGND sg13g2_decap_8
X_1277_ _0731_ net112 _0401_ _0402_ VPWR VGND sg13g2_a21o_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xfanout120 net122 net120 VPWR VGND sg13g2_buf_1
Xfanout131 net133 net131 VPWR VGND sg13g2_buf_1
XFILLER_47_77 VPWR VGND sg13g2_decap_8
Xfanout142 net144 net142 VPWR VGND sg13g2_buf_1
Xfanout153 net156 net153 VPWR VGND sg13g2_buf_1
Xfanout164 net166 net164 VPWR VGND sg13g2_buf_1
Xfanout175 net181 net175 VPWR VGND sg13g2_buf_1
Xfanout186 net187 net186 VPWR VGND sg13g2_buf_1
Xfanout197 net198 net197 VPWR VGND sg13g2_buf_1
XFILLER_11_641 VPWR VGND sg13g2_decap_4
XFILLER_15_435 VPWR VGND sg13g2_decap_8
XFILLER_27_284 VPWR VGND sg13g2_decap_8
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_43_733 VPWR VGND sg13g2_fill_2
XFILLER_43_766 VPWR VGND sg13g2_decap_4
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
XFILLER_26_6 VPWR VGND sg13g2_fill_1
XFILLER_2_361 VPWR VGND sg13g2_decap_8
X_1200_ net139 VPWR _0858_ VGND net93 state\[11\] sg13g2_o21ai_1
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_33_221 VPWR VGND sg13g2_decap_8
XFILLER_34_700 VPWR VGND sg13g2_fill_2
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_46_593 VPWR VGND sg13g2_fill_1
X_1131_ VPWR _0800_ daisychain\[99\] VGND sg13g2_inv_1
X_1062_ VPWR _0731_ daisychain\[30\] VGND sg13g2_inv_1
XFILLER_33_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_1964_ net206 VGND VPWR _0296_ state\[40\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1895_ net201 VGND VPWR _0227_ daisychain\[99\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0915_ VPWR _0116_ state\[8\] VGND sg13g2_inv_1
XFILLER_29_527 VPWR VGND sg13g2_fill_1
X_1329_ _0744_ net119 _0440_ _0441_ VPWR VGND sg13g2_a21o_1
XFILLER_12_405 VPWR VGND sg13g2_decap_8
XFILLER_17_69 VPWR VGND sg13g2_decap_8
XFILLER_24_254 VPWR VGND sg13g2_decap_8
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_16_755 VPWR VGND sg13g2_decap_8
XFILLER_31_703 VPWR VGND sg13g2_decap_4
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_15_265 VPWR VGND sg13g2_decap_8
XFILLER_30_235 VPWR VGND sg13g2_decap_8
XFILLER_7_420 VPWR VGND sg13g2_decap_8
XFILLER_7_497 VPWR VGND sg13g2_decap_8
X_1680_ _0862_ VPWR _0268_ VGND net144 _0031_ sg13g2_o21ai_1
XFILLER_26_508 VPWR VGND sg13g2_fill_1
XFILLER_31_4 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_clk clknet_2_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_1114_ VPWR _0783_ daisychain\[82\] VGND sg13g2_inv_1
X_1045_ VPWR _0714_ daisychain\[13\] VGND sg13g2_inv_1
XFILLER_21_257 VPWR VGND sg13g2_decap_8
X_1947_ net194 VGND VPWR _0279_ state\[23\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1878_ net217 VGND VPWR _0210_ daisychain\[82\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_335 VPWR VGND sg13g2_decap_8
XFILLER_12_202 VPWR VGND sg13g2_decap_8
XFILLER_12_279 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_fill_2
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_9_707 VPWR VGND sg13g2_fill_2
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_36_806 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_8_773 VPWR VGND sg13g2_fill_1
X_1801_ net189 VGND VPWR _0133_ daisychain\[5\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1732_ _0504_ VPWR _0320_ VGND net176 _0088_ sg13g2_o21ai_1
X_1663_ _0254_ _0690_ _0691_ net24 _0699_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_294 VPWR VGND sg13g2_decap_8
X_1594_ VGND VPWR net77 daisychain\[108\] _0640_ net40 sg13g2_a21oi_1
XFILLER_26_349 VPWR VGND sg13g2_decap_8
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_14_48 VPWR VGND sg13g2_decap_8
XFILLER_34_371 VPWR VGND sg13g2_decap_8
XFILLER_41_308 VPWR VGND sg13g2_decap_8
X_1028_ VPWR _0024_ state\[121\] VGND sg13g2_inv_1
XFILLER_30_25 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_29_132 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_17_349 VPWR VGND sg13g2_decap_8
XFILLER_25_382 VPWR VGND sg13g2_fill_1
XFILLER_32_319 VPWR VGND sg13g2_decap_8
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_45_614 VPWR VGND sg13g2_decap_4
XFILLER_45_669 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_9_548 VPWR VGND sg13g2_fill_1
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_5_765 VPWR VGND sg13g2_fill_2
XFILLER_36_614 VPWR VGND sg13g2_fill_2
XFILLER_48_441 VPWR VGND sg13g2_decap_8
X_2000_ net220 VGND VPWR _0332_ state\[76\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_8_581 VPWR VGND sg13g2_fill_2
X_1715_ _0453_ VPWR _0303_ VGND net162 _0069_ sg13g2_o21ai_1
X_1646_ VGND VPWR net70 daisychain\[121\] _0679_ net23 sg13g2_a21oi_1
XFILLER_39_441 VPWR VGND sg13g2_decap_8
X_1577_ _0806_ net107 _0626_ _0627_ VPWR VGND sg13g2_a21o_1
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_10_525 VPWR VGND sg13g2_fill_2
XFILLER_10_558 VPWR VGND sg13g2_decap_8
XFILLER_22_374 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_fill_2
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_17_146 VPWR VGND sg13g2_decap_8
XFILLER_18_636 VPWR VGND sg13g2_fill_2
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_32_116 VPWR VGND sg13g2_decap_8
XFILLER_33_617 VPWR VGND sg13g2_fill_1
XFILLER_9_312 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_31_90 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_5_573 VPWR VGND sg13g2_fill_1
X_1500_ net177 VPWR _0569_ VGND net133 state\[86\] sg13g2_o21ai_1
XFILLER_9_389 VPWR VGND sg13g2_decap_8
XFILLER_5_584 VPWR VGND sg13g2_fill_2
X_1431_ _0196_ _0516_ _0517_ net64 _0769_ VPWR VGND sg13g2_a22oi_1
X_1362_ VGND VPWR net83 daisychain\[50\] _0466_ net54 sg13g2_a21oi_1
X_1293_ _0735_ net113 _0413_ _0414_ VPWR VGND sg13g2_a21o_1
XFILLER_23_116 VPWR VGND sg13g2_fill_2
XFILLER_31_160 VPWR VGND sg13g2_decap_8
Xdigitalen.g\[3\].u.inv2 VPWR digitalen.g\[3\].u.OUTP digitalen.g\[3\].u.OUTN VGND
+ sg13g2_inv_1
X_1629_ _0819_ net94 _0665_ _0666_ VPWR VGND sg13g2_a21o_1
XFILLER_27_422 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_fill_2
XFILLER_42_469 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_18_433 VPWR VGND sg13g2_fill_2
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_46_775 VPWR VGND sg13g2_decap_8
XFILLER_46_786 VPWR VGND sg13g2_fill_2
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_20_119 VPWR VGND sg13g2_decap_8
X_1980_ net209 VGND VPWR _0312_ state\[56\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_0931_ VPWR _0044_ state\[24\] VGND sg13g2_inv_1
XFILLER_9_186 VPWR VGND sg13g2_decap_8
X_1414_ VGND VPWR net87 daisychain\[63\] _0505_ net61 sg13g2_a21oi_1
X_1345_ _0748_ net116 _0452_ _0453_ VPWR VGND sg13g2_a21o_1
X_1276_ net158 VPWR _0401_ VGND net112 state\[30\] sg13g2_o21ai_1
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_37_786 VPWR VGND sg13g2_decap_4
XFILLER_20_675 VPWR VGND sg13g2_fill_2
XFILLER_3_329 VPWR VGND sg13g2_decap_8
Xfanout110 net111 net110 VPWR VGND sg13g2_buf_1
Xfanout121 net122 net121 VPWR VGND sg13g2_buf_1
Xfanout132 net133 net132 VPWR VGND sg13g2_buf_1
Xfanout143 net144 net143 VPWR VGND sg13g2_buf_1
Xfanout154 net156 net154 VPWR VGND sg13g2_buf_1
Xfanout165 net166 net165 VPWR VGND sg13g2_buf_1
XFILLER_27_263 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
Xfanout176 net181 net176 VPWR VGND sg13g2_buf_1
Xfanout187 net227 net187 VPWR VGND sg13g2_buf_1
Xfanout198 net203 net198 VPWR VGND sg13g2_buf_1
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_30_406 VPWR VGND sg13g2_decap_8
XFILLER_42_266 VPWR VGND sg13g2_decap_8
XFILLER_7_613 VPWR VGND sg13g2_fill_2
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_38_528 VPWR VGND sg13g2_fill_1
XFILLER_38_539 VPWR VGND sg13g2_decap_8
X_1130_ VPWR _0799_ daisychain\[98\] VGND sg13g2_inv_1
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_33_200 VPWR VGND sg13g2_decap_8
XFILLER_33_277 VPWR VGND sg13g2_decap_8
X_1061_ VPWR _0730_ daisychain\[29\] VGND sg13g2_inv_1
XFILLER_14_491 VPWR VGND sg13g2_decap_4
XFILLER_21_439 VPWR VGND sg13g2_decap_4
X_1963_ net205 VGND VPWR _0295_ state\[39\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1894_ net201 VGND VPWR _0226_ daisychain\[98\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0914_ VPWR _0105_ state\[7\] VGND sg13g2_inv_1
XFILLER_17_48 VPWR VGND sg13g2_decap_8
XFILLER_37_594 VPWR VGND sg13g2_decap_4
X_1328_ net163 VPWR _0440_ VGND net119 state\[43\] sg13g2_o21ai_1
X_1259_ _0153_ _0387_ _0388_ net33 _0726_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_233 VPWR VGND sg13g2_decap_8
XFILLER_33_25 VPWR VGND sg13g2_decap_8
XFILLER_40_726 VPWR VGND sg13g2_fill_1
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_0_822 VPWR VGND sg13g2_fill_1
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_15_244 VPWR VGND sg13g2_decap_8
XFILLER_11_483 VPWR VGND sg13g2_fill_1
XFILLER_30_214 VPWR VGND sg13g2_decap_8
XFILLER_7_476 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_fill_2
XFILLER_38_336 VPWR VGND sg13g2_decap_8
X_1113_ VPWR _0782_ daisychain\[81\] VGND sg13g2_inv_1
X_1044_ VPWR _0713_ daisychain\[12\] VGND sg13g2_inv_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_21_236 VPWR VGND sg13g2_decap_8
XFILLER_34_597 VPWR VGND sg13g2_decap_4
XFILLER_9_60 VPWR VGND sg13g2_decap_8
X_1946_ net193 VGND VPWR _0278_ state\[22\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1877_ net215 VGND VPWR _0209_ daisychain\[81\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_29_314 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_12_258 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_4
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_4_424 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_0_685 VPWR VGND sg13g2_decap_4
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_fill_1
XFILLER_48_667 VPWR VGND sg13g2_fill_1
XFILLER_16_520 VPWR VGND sg13g2_decap_4
XFILLER_43_350 VPWR VGND sg13g2_decap_8
X_1800_ net189 VGND VPWR _0132_ daisychain\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_11_291 VPWR VGND sg13g2_decap_8
XFILLER_7_273 VPWR VGND sg13g2_decap_8
X_1731_ _0501_ VPWR _0319_ VGND net168 _0087_ sg13g2_o21ai_1
X_1662_ VGND VPWR net70 daisychain\[125\] _0691_ net24 sg13g2_a21oi_1
XFILLER_39_623 VPWR VGND sg13g2_decap_4
XFILLER_3_490 VPWR VGND sg13g2_decap_8
X_1593_ _0810_ net107 _0638_ _0639_ VPWR VGND sg13g2_a21o_1
XFILLER_19_380 VPWR VGND sg13g2_decap_4
XFILLER_34_350 VPWR VGND sg13g2_decap_8
XFILLER_38_133 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_230 VPWR VGND uio_oe[3] sg13g2_tiehi
X_1027_ VPWR _0023_ state\[120\] VGND sg13g2_inv_1
XFILLER_10_718 VPWR VGND sg13g2_fill_1
XFILLER_14_27 VPWR VGND sg13g2_decap_8
X_1929_ net190 VGND VPWR _0261_ state\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_17_328 VPWR VGND sg13g2_decap_8
XFILLER_18_818 VPWR VGND sg13g2_decap_4
XFILLER_29_111 VPWR VGND sg13g2_decap_8
XFILLER_29_188 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_13_567 VPWR VGND sg13g2_fill_1
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_4_221 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_29_90 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_31_342 VPWR VGND sg13g2_decap_8
XFILLER_32_810 VPWR VGND sg13g2_decap_8
XFILLER_32_821 VPWR VGND sg13g2_fill_2
XFILLER_8_571 VPWR VGND sg13g2_decap_4
X_1714_ _0450_ VPWR _0302_ VGND net162 _0068_ sg13g2_o21ai_1
X_1645_ _0823_ net90 _0677_ _0678_ VPWR VGND sg13g2_a21o_1
X_1576_ net153 VPWR _0626_ VGND net107 state\[105\] sg13g2_o21ai_1
XFILLER_39_420 VPWR VGND sg13g2_decap_8
XFILLER_22_320 VPWR VGND sg13g2_decap_4
XFILLER_26_125 VPWR VGND sg13g2_decap_8
XFILLER_35_670 VPWR VGND sg13g2_fill_1
XFILLER_22_353 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_6_508 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_17_125 VPWR VGND sg13g2_decap_8
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_13_375 VPWR VGND sg13g2_decap_8
XFILLER_25_180 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_41_684 VPWR VGND sg13g2_fill_1
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_5_552 VPWR VGND sg13g2_fill_2
X_1430_ VGND VPWR net86 daisychain\[67\] _0517_ net64 sg13g2_a21oi_1
X_1361_ _0752_ net120 _0464_ _0465_ VPWR VGND sg13g2_a21o_1
X_1292_ net158 VPWR _0413_ VGND net113 state\[34\] sg13g2_o21ai_1
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
X_1628_ net140 VPWR _0665_ VGND net94 state\[118\] sg13g2_o21ai_1
X_1559_ _0228_ _0612_ _0613_ net57 _0801_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_14_139 VPWR VGND sg13g2_decap_8
XFILLER_22_194 VPWR VGND sg13g2_decap_8
XFILLER_42_448 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_fill_2
XFILLER_26_91 VPWR VGND sg13g2_decap_4
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_46_743 VPWR VGND sg13g2_fill_1
XFILLER_13_172 VPWR VGND sg13g2_decap_8
X_0930_ VPWR _0043_ state\[23\] VGND sg13g2_inv_1
XFILLER_9_165 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_8
X_1413_ _0765_ net128 _0503_ _0504_ VPWR VGND sg13g2_a21o_1
XFILLER_36_231 VPWR VGND sg13g2_decap_8
XFILLER_37_743 VPWR VGND sg13g2_fill_2
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_49_592 VPWR VGND sg13g2_fill_1
X_1344_ net162 VPWR _0452_ VGND net115 state\[47\] sg13g2_o21ai_1
X_1275_ _0157_ _0399_ _0400_ net33 _0730_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_109 VPWR VGND sg13g2_decap_8
XFILLER_22_27 VPWR VGND sg13g2_decap_4
XFILLER_3_308 VPWR VGND sg13g2_decap_8
XFILLER_19_209 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
Xfanout100 net103 net100 VPWR VGND sg13g2_buf_1
Xfanout111 net135 net111 VPWR VGND sg13g2_buf_1
Xfanout122 net135 net122 VPWR VGND sg13g2_buf_1
Xfanout133 net134 net133 VPWR VGND sg13g2_buf_1
Xfanout144 net145 net144 VPWR VGND sg13g2_buf_1
Xfanout155 net156 net155 VPWR VGND sg13g2_buf_1
Xfanout166 net169 net166 VPWR VGND sg13g2_buf_1
Xfanout177 net180 net177 VPWR VGND sg13g2_buf_1
Xfanout188 net190 net188 VPWR VGND sg13g2_buf_1
Xfanout199 net203 net199 VPWR VGND sg13g2_buf_1
XFILLER_27_242 VPWR VGND sg13g2_decap_8
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_43_735 VPWR VGND sg13g2_fill_1
XFILLER_43_746 VPWR VGND sg13g2_fill_2
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_11_687 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
X_1060_ VPWR _0729_ daisychain\[28\] VGND sg13g2_inv_1
XFILLER_19_787 VPWR VGND sg13g2_fill_2
XFILLER_33_256 VPWR VGND sg13g2_decap_8
X_1962_ net208 VGND VPWR _0294_ state\[38\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1893_ net202 VGND VPWR _0225_ daisychain\[97\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0913_ VPWR _0094_ state\[6\] VGND sg13g2_inv_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_17_27 VPWR VGND sg13g2_decap_8
XFILLER_24_212 VPWR VGND sg13g2_decap_8
XFILLER_37_540 VPWR VGND sg13g2_decap_8
X_1327_ _0170_ _0438_ _0439_ net46 _0743_ VPWR VGND sg13g2_a22oi_1
X_1258_ VGND VPWR net72 daisychain\[24\] _0388_ net36 sg13g2_a21oi_1
X_1189_ _0709_ net92 _0849_ _0850_ VPWR VGND sg13g2_a21o_1
XFILLER_24_289 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_15_223 VPWR VGND sg13g2_decap_8
XFILLER_43_565 VPWR VGND sg13g2_fill_1
XFILLER_7_455 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_3_672 VPWR VGND sg13g2_fill_2
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_34_521 VPWR VGND sg13g2_fill_2
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
X_1112_ VPWR _0781_ daisychain\[80\] VGND sg13g2_inv_1
X_1043_ VPWR _0712_ daisychain\[11\] VGND sg13g2_inv_1
XFILLER_21_215 VPWR VGND sg13g2_decap_8
X_1945_ net193 VGND VPWR _0277_ state\[21\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1876_ net215 VGND VPWR _0208_ daisychain\[80\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_13_749 VPWR VGND sg13g2_fill_2
XFILLER_25_543 VPWR VGND sg13g2_fill_1
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_40_513 VPWR VGND sg13g2_fill_1
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_12_237 VPWR VGND sg13g2_decap_8
XFILLER_40_579 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_decap_8
XFILLER_0_664 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_16_565 VPWR VGND sg13g2_fill_2
XFILLER_16_576 VPWR VGND sg13g2_fill_2
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_8_720 VPWR VGND sg13g2_fill_2
XFILLER_11_270 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_decap_4
X_1730_ _0498_ VPWR _0318_ VGND net168 _0086_ sg13g2_o21ai_1
X_1661_ _0699_ net91 _0689_ _0690_ VPWR VGND sg13g2_a21o_1
X_1592_ net153 VPWR _0638_ VGND net107 state\[109\] sg13g2_o21ai_1
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
XFILLER_47_690 VPWR VGND sg13g2_fill_2
X_2075_ daisychain\[127\] net22 VPWR VGND sg13g2_buf_1
Xheichips25_pudding_231 VPWR VGND uio_oe[4] sg13g2_tiehi
X_1026_ VPWR _0021_ state\[119\] VGND sg13g2_inv_1
X_1928_ net188 VGND VPWR _0260_ state\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1859_ net213 VGND VPWR _0191_ daisychain\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_17_307 VPWR VGND sg13g2_decap_8
XFILLER_29_167 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_13_546 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_41_822 VPWR VGND sg13g2_fill_1
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_20_82 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_16_384 VPWR VGND sg13g2_decap_8
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_16_395 VPWR VGND sg13g2_fill_2
XFILLER_31_321 VPWR VGND sg13g2_decap_8
X_1713_ _0447_ VPWR _0301_ VGND net160 _0067_ sg13g2_o21ai_1
XFILLER_6_95 VPWR VGND sg13g2_decap_8
X_1644_ net138 VPWR _0677_ VGND net90 state\[122\] sg13g2_o21ai_1
X_1575_ _0232_ _0624_ _0625_ net40 _0805_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_104 VPWR VGND sg13g2_fill_2
XFILLER_39_476 VPWR VGND sg13g2_decap_8
XFILLER_42_608 VPWR VGND sg13g2_decap_8
XFILLER_42_619 VPWR VGND sg13g2_fill_1
X_1009_ VPWR _0003_ state\[102\] VGND sg13g2_inv_1
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_14_822 VPWR VGND sg13g2_fill_1
XFILLER_17_104 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_decap_8
X_1360_ net167 VPWR _0464_ VGND net120 state\[51\] sg13g2_o21ai_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_fill_1
XFILLER_49_774 VPWR VGND sg13g2_decap_4
XFILLER_49_796 VPWR VGND sg13g2_fill_2
X_1291_ _0161_ _0411_ _0412_ net45 _0734_ VPWR VGND sg13g2_a22oi_1
XFILLER_16_181 VPWR VGND sg13g2_decap_8
XFILLER_20_814 VPWR VGND sg13g2_decap_4
XFILLER_23_118 VPWR VGND sg13g2_fill_1
XFILLER_44_490 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
XFILLER_31_195 VPWR VGND sg13g2_decap_8
X_1627_ _0245_ _0663_ _0664_ net28 _0818_ VPWR VGND sg13g2_a22oi_1
X_1558_ VGND VPWR net77 daisychain\[99\] _0613_ net57 sg13g2_a21oi_1
X_1489_ _0784_ net125 _0560_ _0561_ VPWR VGND sg13g2_a21o_1
XFILLER_14_118 VPWR VGND sg13g2_decap_8
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_42_427 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_11_814 VPWR VGND sg13g2_decap_8
XFILLER_22_173 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_fill_2
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_46_733 VPWR VGND sg13g2_fill_2
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_18_446 VPWR VGND sg13g2_decap_8
XFILLER_26_70 VPWR VGND sg13g2_fill_1
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_46_755 VPWR VGND sg13g2_decap_8
XFILLER_14_685 VPWR VGND sg13g2_decap_4
XFILLER_42_91 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_decap_8
X_1412_ net175 VPWR _0503_ VGND net128 state\[64\] sg13g2_o21ai_1
X_1343_ _0174_ _0450_ _0451_ net48 _0747_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
X_1274_ VGND VPWR net72 daisychain\[28\] _0400_ net33 sg13g2_a21oi_1
XFILLER_20_622 VPWR VGND sg13g2_fill_1
XFILLER_32_471 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_2_0__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_0989_ VPWR _0108_ state\[82\] VGND sg13g2_inv_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
Xfanout101 net102 net101 VPWR VGND sg13g2_buf_1
Xfanout112 net113 net112 VPWR VGND sg13g2_buf_1
Xfanout123 net127 net123 VPWR VGND sg13g2_buf_1
Xfanout134 net135 net134 VPWR VGND sg13g2_buf_1
Xfanout145 net157 net145 VPWR VGND sg13g2_buf_1
Xfanout156 net157 net156 VPWR VGND sg13g2_buf_1
Xfanout167 net169 net167 VPWR VGND sg13g2_buf_1
Xfanout178 net180 net178 VPWR VGND sg13g2_buf_1
Xfanout189 net190 net189 VPWR VGND sg13g2_buf_1
XFILLER_15_405 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_decap_8
XFILLER_27_298 VPWR VGND sg13g2_decap_4
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_decap_8
XFILLER_7_615 VPWR VGND sg13g2_fill_1
XFILLER_12_83 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_19_8 VPWR VGND sg13g2_fill_1
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_46_574 VPWR VGND sg13g2_fill_2
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_33_235 VPWR VGND sg13g2_decap_8
X_1961_ net207 VGND VPWR _0293_ state\[37\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1892_ net202 VGND VPWR _0224_ daisychain\[96\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0912_ VPWR _0083_ state\[5\] VGND sg13g2_inv_1
XFILLER_6_681 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_5_clk clknet_2_3__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_1326_ VGND VPWR net79 daisychain\[41\] _0439_ net46 sg13g2_a21oi_1
XFILLER_12_419 VPWR VGND sg13g2_decap_8
XFILLER_24_268 VPWR VGND sg13g2_decap_8
X_1257_ _0726_ net99 _0386_ _0387_ VPWR VGND sg13g2_a21o_1
X_1188_ net139 VPWR _0849_ VGND net92 state\[8\] sg13g2_o21ai_1
XFILLER_15_202 VPWR VGND sg13g2_decap_8
XFILLER_15_279 VPWR VGND sg13g2_decap_8
XFILLER_16_747 VPWR VGND sg13g2_fill_2
XFILLER_30_249 VPWR VGND sg13g2_decap_8
XFILLER_7_434 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_530 VPWR VGND sg13g2_decap_8
XFILLER_34_500 VPWR VGND sg13g2_decap_4
XFILLER_34_555 VPWR VGND sg13g2_fill_1
XFILLER_46_371 VPWR VGND sg13g2_decap_8
X_1111_ VPWR _0780_ daisychain\[79\] VGND sg13g2_inv_1
X_1042_ VPWR _0711_ daisychain\[10\] VGND sg13g2_inv_1
XFILLER_30_750 VPWR VGND sg13g2_fill_1
XFILLER_30_761 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_fill_1
XFILLER_30_783 VPWR VGND sg13g2_fill_2
X_1944_ net193 VGND VPWR _0276_ state\[20\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1875_ net215 VGND VPWR _0207_ daisychain\[79\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_44_308 VPWR VGND sg13g2_decap_8
X_1309_ _0739_ net113 _0425_ _0426_ VPWR VGND sg13g2_a21o_1
XFILLER_12_216 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_16_500 VPWR VGND sg13g2_decap_8
XFILLER_16_544 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_fill_2
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_fill_2
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_7_231 VPWR VGND sg13g2_decap_8
X_1660_ net137 VPWR _0689_ VGND net91 state\[126\] sg13g2_o21ai_1
X_1591_ _0236_ _0636_ _0637_ net39 _0809_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_168 VPWR VGND sg13g2_decap_8
XFILLER_34_385 VPWR VGND sg13g2_decap_8
X_2074_ daisychain\[126\] net21 VPWR VGND sg13g2_buf_1
Xheichips25_pudding_232 VPWR VGND uio_oe[5] sg13g2_tiehi
X_1025_ VPWR _0020_ state\[118\] VGND sg13g2_inv_1
XFILLER_30_39 VPWR VGND sg13g2_decap_8
X_1927_ net193 VGND VPWR _0259_ state\[3\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1858_ net212 VGND VPWR _0190_ daisychain\[62\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1789_ _0675_ VPWR _0377_ VGND net137 _0024_ sg13g2_o21ai_1
XFILLER_25_330 VPWR VGND sg13g2_decap_8
XFILLER_29_146 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_16_363 VPWR VGND sg13g2_decap_8
XFILLER_31_300 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND _0007_ sg13g2_antennanp
X_1712_ _0444_ VPWR _0300_ VGND net163 _0066_ sg13g2_o21ai_1
X_1643_ _0249_ _0675_ _0676_ net23 _0822_ VPWR VGND sg13g2_a22oi_1
XFILLER_6_74 VPWR VGND sg13g2_decap_8
X_1574_ VGND VPWR net77 daisychain\[103\] _0625_ net43 sg13g2_a21oi_1
XFILLER_39_455 VPWR VGND sg13g2_decap_8
XFILLER_22_388 VPWR VGND sg13g2_fill_2
XFILLER_34_182 VPWR VGND sg13g2_decap_8
XFILLER_35_683 VPWR VGND sg13g2_fill_2
XFILLER_41_119 VPWR VGND sg13g2_decap_8
X_1008_ VPWR _0002_ state\[101\] VGND sg13g2_inv_1
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_13_333 VPWR VGND sg13g2_decap_8
XFILLER_18_628 VPWR VGND sg13g2_fill_1
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_15_83 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_5_543 VPWR VGND sg13g2_decap_4
XFILLER_5_554 VPWR VGND sg13g2_fill_1
XFILLER_17_650 VPWR VGND sg13g2_fill_1
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_49_742 VPWR VGND sg13g2_decap_8
X_1290_ VGND VPWR net79 daisychain\[32\] _0412_ net45 sg13g2_a21oi_1
XFILLER_16_160 VPWR VGND sg13g2_decap_8
XFILLER_31_174 VPWR VGND sg13g2_decap_8
XFILLER_32_664 VPWR VGND sg13g2_fill_2
X_1626_ VGND VPWR net69 daisychain\[116\] _0664_ net27 sg13g2_a21oi_1
XFILLER_39_252 VPWR VGND sg13g2_decap_8
X_1557_ _0801_ net124 _0611_ _0612_ VPWR VGND sg13g2_a21o_1
X_1488_ net172 VPWR _0560_ VGND net125 state\[83\] sg13g2_o21ai_1
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
XFILLER_22_152 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_46_712 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_41_483 VPWR VGND sg13g2_decap_8
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
XFILLER_49_550 VPWR VGND sg13g2_decap_8
X_1411_ _0191_ _0501_ _0502_ net55 _0764_ VPWR VGND sg13g2_a22oi_1
X_1342_ VGND VPWR net80 daisychain\[45\] _0451_ net47 sg13g2_a21oi_1
X_1273_ _0730_ net100 _0398_ _0399_ VPWR VGND sg13g2_a21o_1
XFILLER_36_266 VPWR VGND sg13g2_decap_8
X_0988_ VPWR _0107_ state\[81\] VGND sg13g2_inv_1
Xfanout102 net103 net102 VPWR VGND sg13g2_buf_1
Xfanout113 net116 net113 VPWR VGND sg13g2_buf_1
X_1609_ _0814_ net104 _0650_ _0651_ VPWR VGND sg13g2_a21o_1
XFILLER_27_200 VPWR VGND sg13g2_decap_8
Xfanout124 net126 net124 VPWR VGND sg13g2_buf_1
Xfanout135 net136 net135 VPWR VGND sg13g2_buf_1
Xfanout146 net149 net146 VPWR VGND sg13g2_buf_1
Xfanout157 net182 net157 VPWR VGND sg13g2_buf_1
Xfanout168 net169 net168 VPWR VGND sg13g2_buf_1
Xfanout179 net180 net179 VPWR VGND sg13g2_buf_1
XFILLER_11_623 VPWR VGND sg13g2_decap_8
XFILLER_15_428 VPWR VGND sg13g2_decap_8
XFILLER_27_277 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_43_726 VPWR VGND sg13g2_decap_8
XFILLER_43_748 VPWR VGND sg13g2_fill_1
XFILLER_43_759 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_11_645 VPWR VGND sg13g2_fill_1
XFILLER_12_62 VPWR VGND sg13g2_decap_8
XFILLER_6_137 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_33_214 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
X_1960_ net207 VGND VPWR _0292_ state\[36\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1891_ net202 VGND VPWR _0223_ daisychain\[95\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0911_ VPWR _0072_ state\[4\] VGND sg13g2_inv_1
XFILLER_29_509 VPWR VGND sg13g2_fill_2
X_1325_ _0743_ net114 _0437_ _0438_ VPWR VGND sg13g2_a21o_1
X_1256_ net146 VPWR _0386_ VGND net99 state\[25\] sg13g2_o21ai_1
XFILLER_24_247 VPWR VGND sg13g2_decap_8
XFILLER_33_39 VPWR VGND sg13g2_decap_8
X_1187_ _0135_ _0847_ _0848_ net26 _0708_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_431 VPWR VGND sg13g2_decap_8
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_11_431 VPWR VGND sg13g2_decap_4
XFILLER_11_464 VPWR VGND sg13g2_fill_1
XFILLER_15_258 VPWR VGND sg13g2_decap_8
XFILLER_30_228 VPWR VGND sg13g2_decap_8
XFILLER_31_707 VPWR VGND sg13g2_fill_2
XFILLER_7_413 VPWR VGND sg13g2_decap_8
XFILLER_3_641 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_3_674 VPWR VGND sg13g2_fill_1
XFILLER_48_91 VPWR VGND sg13g2_decap_8
X_1110_ VPWR _0779_ daisychain\[78\] VGND sg13g2_inv_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
X_1041_ VPWR _0710_ daisychain\[9\] VGND sg13g2_inv_1
XFILLER_30_740 VPWR VGND sg13g2_fill_2
X_1943_ net191 VGND VPWR _0275_ state\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1874_ net219 VGND VPWR _0206_ daisychain\[78\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_29_328 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
X_1308_ net161 VPWR _0425_ VGND net115 state\[38\] sg13g2_o21ai_1
X_1239_ _0148_ _0886_ _0887_ net35 _0721_ VPWR VGND sg13g2_a22oi_1
XFILLER_40_504 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_4_438 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_fill_1
XFILLER_16_567 VPWR VGND sg13g2_fill_1
XFILLER_16_578 VPWR VGND sg13g2_fill_1
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_12_751 VPWR VGND sg13g2_fill_1
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_8_722 VPWR VGND sg13g2_fill_1
XFILLER_8_766 VPWR VGND sg13g2_decap_8
XFILLER_8_777 VPWR VGND sg13g2_decap_4
XFILLER_7_287 VPWR VGND sg13g2_decap_8
X_1590_ VGND VPWR net75 daisychain\[107\] _0637_ net38 sg13g2_a21oi_1
XFILLER_19_361 VPWR VGND sg13g2_fill_2
XFILLER_22_4 VPWR VGND sg13g2_fill_1
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_39_659 VPWR VGND sg13g2_fill_1
X_2073_ daisychain\[125\] net20 VPWR VGND sg13g2_buf_1
X_1024_ VPWR _0019_ state\[117\] VGND sg13g2_inv_1
XFILLER_22_537 VPWR VGND sg13g2_fill_1
XFILLER_34_364 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_233 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_30_18 VPWR VGND sg13g2_decap_8
X_1926_ net193 VGND VPWR _0258_ state\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1857_ net212 VGND VPWR _0189_ daisychain\[61\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1788_ _0672_ VPWR _0376_ VGND net141 _0023_ sg13g2_o21ai_1
XFILLER_29_125 VPWR VGND sg13g2_decap_8
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_45_618 VPWR VGND sg13g2_fill_2
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_9_519 VPWR VGND sg13g2_fill_2
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_5_758 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_16_342 VPWR VGND sg13g2_decap_8
XFILLER_31_356 VPWR VGND sg13g2_decap_4
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_44_662 VPWR VGND sg13g2_fill_1
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XANTENNA_2 VPWR VGND _0012_ sg13g2_antennanp
XFILLER_12_581 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
X_1711_ _0441_ VPWR _0299_ VGND net163 _0065_ sg13g2_o21ai_1
X_1642_ VGND VPWR net70 daisychain\[120\] _0676_ net23 sg13g2_a21oi_1
XFILLER_39_434 VPWR VGND sg13g2_decap_8
X_1573_ _0805_ net107 _0623_ _0624_ VPWR VGND sg13g2_a21o_1
XFILLER_34_161 VPWR VGND sg13g2_decap_8
X_1007_ VPWR _0001_ state\[100\] VGND sg13g2_inv_1
XFILLER_22_367 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
X_1909_ net196 VGND VPWR _0241_ daisychain\[113\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_18_618 VPWR VGND sg13g2_fill_2
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_15_62 VPWR VGND sg13g2_decap_8
XFILLER_17_139 VPWR VGND sg13g2_decap_8
XFILLER_25_194 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_41_632 VPWR VGND sg13g2_fill_2
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_31_83 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_566 VPWR VGND sg13g2_decap_8
XFILLER_5_577 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_31_153 VPWR VGND sg13g2_decap_8
XFILLER_32_698 VPWR VGND sg13g2_decap_8
XFILLER_8_382 VPWR VGND sg13g2_decap_8
X_1625_ _0818_ net94 _0662_ _0663_ VPWR VGND sg13g2_a21o_1
X_1556_ net171 VPWR _0611_ VGND net124 state\[100\] sg13g2_o21ai_1
XFILLER_27_415 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_39_231 VPWR VGND sg13g2_decap_8
X_1487_ _0210_ _0558_ _0559_ net60 _0783_ VPWR VGND sg13g2_a22oi_1
X_2039_ net196 VGND VPWR _0371_ state\[115\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_18_426 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_fill_1
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_41_462 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_5_396 VPWR VGND sg13g2_decap_8
X_1410_ VGND VPWR net83 daisychain\[62\] _0502_ net55 sg13g2_a21oi_1
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
X_1341_ _0747_ net115 _0449_ _0450_ VPWR VGND sg13g2_a21o_1
X_1272_ net146 VPWR _0398_ VGND net100 state\[29\] sg13g2_o21ai_1
XFILLER_17_492 VPWR VGND sg13g2_fill_2
XFILLER_32_440 VPWR VGND sg13g2_fill_2
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_37_779 VPWR VGND sg13g2_decap_8
XFILLER_20_657 VPWR VGND sg13g2_fill_1
XFILLER_20_668 VPWR VGND sg13g2_decap_8
X_0987_ VPWR _0106_ state\[80\] VGND sg13g2_inv_1
XFILLER_9_691 VPWR VGND sg13g2_decap_8
Xfanout103 net111 net103 VPWR VGND sg13g2_buf_1
Xfanout114 net116 net114 VPWR VGND sg13g2_buf_1
Xfanout125 net126 net125 VPWR VGND sg13g2_buf_1
Xfanout136 net5 net136 VPWR VGND sg13g2_buf_1
Xfanout147 net148 net147 VPWR VGND sg13g2_buf_1
X_1608_ net150 VPWR _0650_ VGND net104 state\[113\] sg13g2_o21ai_1
X_1539_ _0223_ _0597_ _0598_ net43 _0796_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_256 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
Xfanout158 net160 net158 VPWR VGND sg13g2_buf_1
Xfanout169 net182 net169 VPWR VGND sg13g2_buf_1
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_7_606 VPWR VGND sg13g2_decap_8
XFILLER_12_41 VPWR VGND sg13g2_decap_8
XFILLER_3_801 VPWR VGND sg13g2_fill_1
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_14_484 VPWR VGND sg13g2_decap_8
XFILLER_14_495 VPWR VGND sg13g2_fill_1
XFILLER_42_782 VPWR VGND sg13g2_decap_8
X_1890_ net201 VGND VPWR _0222_ daisychain\[94\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_0910_ VPWR _0061_ state\[3\] VGND sg13g2_inv_1
XFILLER_5_193 VPWR VGND sg13g2_decap_8
X_1324_ net159 VPWR _0437_ VGND net114 state\[42\] sg13g2_o21ai_1
X_1255_ _0152_ _0384_ _0385_ net36 _0725_ VPWR VGND sg13g2_a22oi_1
X_1186_ VGND VPWR net68 daisychain\[6\] _0848_ net25 sg13g2_a21oi_1
XFILLER_24_226 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_33_760 VPWR VGND sg13g2_decap_8
XFILLER_37_598 VPWR VGND sg13g2_fill_1
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_15_237 VPWR VGND sg13g2_decap_8
XFILLER_16_749 VPWR VGND sg13g2_fill_1
XFILLER_11_410 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_decap_8
XFILLER_23_51 VPWR VGND sg13g2_decap_8
XFILLER_30_207 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_3_631 VPWR VGND sg13g2_fill_1
XFILLER_7_469 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_fill_2
XFILLER_19_543 VPWR VGND sg13g2_fill_1
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_4
XFILLER_48_70 VPWR VGND sg13g2_decap_8
X_1040_ VPWR _0709_ daisychain\[8\] VGND sg13g2_inv_1
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_21_229 VPWR VGND sg13g2_decap_8
X_1942_ net190 VGND VPWR _0274_ state\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_30_785 VPWR VGND sg13g2_fill_1
XFILLER_30_796 VPWR VGND sg13g2_fill_1
XFILLER_6_480 VPWR VGND sg13g2_decap_8
X_1873_ net219 VGND VPWR _0205_ daisychain\[77\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_29_307 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_8
X_1307_ _0165_ _0423_ _0424_ net48 _0738_ VPWR VGND sg13g2_a22oi_1
X_1238_ VGND VPWR net72 daisychain\[19\] _0887_ net34 sg13g2_a21oi_1
X_1169_ _0704_ net102 _0834_ _0835_ VPWR VGND sg13g2_a21o_1
XFILLER_20_273 VPWR VGND sg13g2_decap_4
XFILLER_20_295 VPWR VGND sg13g2_fill_1
XFILLER_4_417 VPWR VGND sg13g2_decap_8
XFILLER_0_678 VPWR VGND sg13g2_decap_4
XFILLER_28_351 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_fill_2
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_28_362 VPWR VGND sg13g2_fill_1
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_44_822 VPWR VGND sg13g2_fill_1
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_4
XFILLER_19_373 VPWR VGND sg13g2_fill_2
XFILLER_19_384 VPWR VGND sg13g2_fill_2
XFILLER_34_343 VPWR VGND sg13g2_decap_8
XFILLER_38_126 VPWR VGND sg13g2_decap_8
X_2072_ daisychain\[124\] net19 VPWR VGND sg13g2_buf_1
X_1023_ VPWR _0018_ state\[116\] VGND sg13g2_inv_1
XFILLER_30_571 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_234 VPWR VGND uio_oe[7] sg13g2_tiehi
X_1925_ net188 VGND VPWR _0257_ state\[1\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_30_593 VPWR VGND sg13g2_fill_2
X_1856_ net209 VGND VPWR _0188_ daisychain\[60\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1787_ _0669_ VPWR _0375_ VGND net141 _0021_ sg13g2_o21ai_1
XFILLER_29_104 VPWR VGND sg13g2_decap_8
XFILLER_39_28 VPWR VGND sg13g2_decap_8
XFILLER_13_527 VPWR VGND sg13g2_fill_2
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_20_41 VPWR VGND sg13g2_decap_8
XFILLER_20_96 VPWR VGND sg13g2_decap_4
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_16_321 VPWR VGND sg13g2_decap_8
XFILLER_17_822 VPWR VGND sg13g2_fill_1
XFILLER_29_83 VPWR VGND sg13g2_decap_8
XFILLER_44_641 VPWR VGND sg13g2_fill_1
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_31_335 VPWR VGND sg13g2_decap_8
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_8_520 VPWR VGND sg13g2_decap_8
XFILLER_8_531 VPWR VGND sg13g2_fill_1
XANTENNA_3 VPWR VGND _0047_ sg13g2_antennanp
XFILLER_6_32 VPWR VGND sg13g2_decap_8
XFILLER_8_564 VPWR VGND sg13g2_decap_8
XFILLER_8_575 VPWR VGND sg13g2_fill_2
XFILLER_8_586 VPWR VGND sg13g2_fill_2
X_1710_ _0438_ VPWR _0298_ VGND net159 _0064_ sg13g2_o21ai_1
X_1641_ _0822_ net90 _0674_ _0675_ VPWR VGND sg13g2_a21o_1
X_1572_ net156 VPWR _0623_ VGND net107 state\[104\] sg13g2_o21ai_1
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_3_280 VPWR VGND sg13g2_decap_8
XFILLER_19_181 VPWR VGND sg13g2_decap_8
XFILLER_22_313 VPWR VGND sg13g2_decap_8
XFILLER_26_118 VPWR VGND sg13g2_decap_8
XFILLER_34_140 VPWR VGND sg13g2_decap_8
XFILLER_35_685 VPWR VGND sg13g2_fill_1
XFILLER_35_696 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
X_1006_ VPWR _0126_ state\[99\] VGND sg13g2_inv_1
XFILLER_22_346 VPWR VGND sg13g2_decap_8
X_1908_ net196 VGND VPWR _0240_ daisychain\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1839_ net205 VGND VPWR _0171_ daisychain\[43\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_17_118 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_13_368 VPWR VGND sg13g2_decap_8
XFILLER_15_41 VPWR VGND sg13g2_decap_8
XFILLER_25_173 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_31_62 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_fill_2
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_16_195 VPWR VGND sg13g2_decap_8
XFILLER_20_806 VPWR VGND sg13g2_decap_4
XFILLER_31_132 VPWR VGND sg13g2_decap_8
XFILLER_32_655 VPWR VGND sg13g2_fill_2
XFILLER_8_361 VPWR VGND sg13g2_decap_8
X_1624_ net140 VPWR _0662_ VGND net94 state\[117\] sg13g2_o21ai_1
X_1555_ _0227_ _0609_ _0610_ net41 _0800_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
X_1486_ VGND VPWR net85 daisychain\[81\] _0559_ net60 sg13g2_a21oi_1
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_35_482 VPWR VGND sg13g2_decap_4
X_2038_ net198 VGND VPWR _0370_ state\[114\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_22_187 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_14_622 VPWR VGND sg13g2_decap_8
XFILLER_26_84 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_46_747 VPWR VGND sg13g2_fill_1
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_9_158 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_decap_8
X_1340_ net162 VPWR _0449_ VGND net115 state\[46\] sg13g2_o21ai_1
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
XFILLER_49_596 VPWR VGND sg13g2_decap_8
X_1271_ _0156_ _0396_ _0397_ net33 _0729_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_603 VPWR VGND sg13g2_fill_1
XFILLER_45_791 VPWR VGND sg13g2_fill_2
XFILLER_32_485 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_0986_ VPWR _0104_ state\[79\] VGND sg13g2_inv_1
XFILLER_47_28 VPWR VGND sg13g2_decap_8
Xfanout104 net105 net104 VPWR VGND sg13g2_buf_1
Xfanout115 net116 net115 VPWR VGND sg13g2_buf_1
Xfanout126 net127 net126 VPWR VGND sg13g2_buf_1
Xfanout137 net138 net137 VPWR VGND sg13g2_buf_1
Xfanout148 net149 net148 VPWR VGND sg13g2_buf_1
Xfanout159 net160 net159 VPWR VGND sg13g2_buf_1
X_1607_ _0240_ _0648_ _0649_ net37 _0813_ VPWR VGND sg13g2_a22oi_1
X_1538_ VGND VPWR net76 daisychain\[94\] _0598_ net41 sg13g2_a21oi_1
X_1469_ _0779_ net128 _0545_ _0546_ VPWR VGND sg13g2_a21o_1
XFILLER_15_419 VPWR VGND sg13g2_decap_4
XFILLER_27_235 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_12_20 VPWR VGND sg13g2_decap_8
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_97 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_18_235 VPWR VGND sg13g2_decap_8
XFILLER_33_249 VPWR VGND sg13g2_decap_8
XFILLER_42_761 VPWR VGND sg13g2_decap_8
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_6_695 VPWR VGND sg13g2_decap_8
X_1323_ _0169_ _0435_ _0436_ net46 _0742_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_205 VPWR VGND sg13g2_decap_8
XFILLER_49_382 VPWR VGND sg13g2_decap_8
X_1254_ VGND VPWR net73 daisychain\[23\] _0385_ net35 sg13g2_a21oi_1
X_1185_ _0708_ net92 _0846_ _0847_ VPWR VGND sg13g2_a21o_1
XFILLER_18_791 VPWR VGND sg13g2_fill_1
X_0969_ VPWR _0086_ state\[62\] VGND sg13g2_inv_1
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_15_216 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_fill_2
XFILLER_11_499 VPWR VGND sg13g2_decap_8
XFILLER_23_282 VPWR VGND sg13g2_decap_8
XFILLER_7_448 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_514 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_14_293 VPWR VGND sg13g2_decap_8
XFILLER_21_208 VPWR VGND sg13g2_decap_8
XFILLER_30_742 VPWR VGND sg13g2_fill_1
XFILLER_42_580 VPWR VGND sg13g2_decap_8
X_1941_ net190 VGND VPWR _0273_ state\[17\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1872_ net220 VGND VPWR _0204_ daisychain\[76\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_1306_ VGND VPWR net80 daisychain\[36\] _0424_ net48 sg13g2_a21oi_1
XFILLER_25_536 VPWR VGND sg13g2_decap_8
XFILLER_37_385 VPWR VGND sg13g2_decap_8
X_1237_ _0721_ net101 _0885_ _0886_ VPWR VGND sg13g2_a21o_1
X_1168_ net147 VPWR _0834_ VGND net101 state\[3\] sg13g2_o21ai_1
X_1099_ VPWR _0768_ daisychain\[67\] VGND sg13g2_inv_1
XFILLER_20_252 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_613 VPWR VGND sg13g2_fill_1
XFILLER_0_657 VPWR VGND sg13g2_decap_8
XFILLER_16_514 VPWR VGND sg13g2_fill_2
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_28_374 VPWR VGND sg13g2_decap_4
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_16_558 VPWR VGND sg13g2_fill_1
XFILLER_28_396 VPWR VGND sg13g2_decap_8
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_8_713 VPWR VGND sg13g2_decap_8
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_12_786 VPWR VGND sg13g2_decap_4
XFILLER_7_245 VPWR VGND sg13g2_decap_8
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_3_462 VPWR VGND sg13g2_decap_8
XFILLER_22_517 VPWR VGND sg13g2_fill_2
XFILLER_34_322 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
X_2071_ daisychain\[123\] net18 VPWR VGND sg13g2_buf_1
X_1022_ VPWR _0017_ state\[115\] VGND sg13g2_inv_1
XFILLER_34_399 VPWR VGND sg13g2_decap_4
X_1924_ net196 VGND VPWR _0256_ state\[0\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1855_ net209 VGND VPWR _0187_ daisychain\[59\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1786_ _0666_ VPWR _0374_ VGND net141 _0020_ sg13g2_o21ai_1
XFILLER_25_300 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_13_506 VPWR VGND sg13g2_fill_1
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_20_20 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_20_64 VPWR VGND sg13g2_fill_1
XFILLER_20_75 VPWR VGND sg13g2_decap_8
XFILLER_29_62 VPWR VGND sg13g2_decap_8
XFILLER_16_300 VPWR VGND sg13g2_decap_8
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_32_804 VPWR VGND sg13g2_fill_2
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_16_377 VPWR VGND sg13g2_decap_8
XFILLER_31_314 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND _0112_ sg13g2_antennanp
XFILLER_4_782 VPWR VGND sg13g2_fill_1
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
X_1640_ net138 VPWR _0674_ VGND net90 state\[121\] sg13g2_o21ai_1
X_1571_ _0231_ _0621_ _0622_ net43 _0804_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_469 VPWR VGND sg13g2_decap_8
XFILLER_19_160 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_decap_8
X_1005_ VPWR _0125_ state\[98\] VGND sg13g2_inv_1
XFILLER_10_509 VPWR VGND sg13g2_fill_2
XFILLER_30_380 VPWR VGND sg13g2_decap_8
X_1907_ net197 VGND VPWR _0239_ daisychain\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1838_ net205 VGND VPWR _0170_ daisychain\[42\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1769_ _0615_ VPWR _0357_ VGND net170 _0002_ sg13g2_o21ai_1
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_20 VPWR VGND sg13g2_decap_8
XFILLER_15_97 VPWR VGND sg13g2_decap_8
XFILLER_21_391 VPWR VGND sg13g2_decap_8
XFILLER_25_152 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_31_41 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_1_774 VPWR VGND sg13g2_decap_4
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_49_756 VPWR VGND sg13g2_decap_8
XFILLER_49_778 VPWR VGND sg13g2_fill_2
XFILLER_16_174 VPWR VGND sg13g2_decap_8
XFILLER_31_111 VPWR VGND sg13g2_decap_8
XFILLER_32_601 VPWR VGND sg13g2_fill_1
XFILLER_44_483 VPWR VGND sg13g2_decap_8
XFILLER_12_391 VPWR VGND sg13g2_decap_8
XFILLER_20_818 VPWR VGND sg13g2_fill_2
XFILLER_31_188 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
X_1623_ _0244_ _0660_ _0661_ net27 _0817_ VPWR VGND sg13g2_a22oi_1
X_1554_ VGND VPWR net77 daisychain\[98\] _0610_ net41 sg13g2_a21oi_1
X_1485_ _0783_ net127 _0557_ _0558_ VPWR VGND sg13g2_a21o_1
.ends

