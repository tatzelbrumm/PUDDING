** sch_path: /home/user/PUDDING/schematic/Pmirrors_top.sch
**.subckt Pmirrors_top VDD Iout Vbiasp
*+ VcascodeP[255],VcascodeP[254],VcascodeP[253],VcascodeP[252],VcascodeP[251],VcascodeP[250],VcascodeP[249],VcascodeP[248],VcascodeP[247],VcascodeP[246],VcascodeP[245],VcascodeP[244],VcascodeP[243],VcascodeP[242],VcascodeP[241],VcascodeP[240],VcascodeP[239],VcascodeP[238],VcascodeP[237],VcascodeP[236],VcascodeP[235],VcascodeP[234],VcascodeP[233],VcascodeP[232],VcascodeP[231],VcascodeP[230],VcascodeP[229],VcascodeP[228],VcascodeP[227],VcascodeP[226],VcascodeP[225],VcascodeP[224],VcascodeP[223],VcascodeP[222],VcascodeP[221],VcascodeP[220],VcascodeP[219],VcascodeP[218],VcascodeP[217],VcascodeP[216],VcascodeP[215],VcascodeP[214],VcascodeP[213],VcascodeP[212],VcascodeP[211],VcascodeP[210],VcascodeP[209],VcascodeP[208],VcascodeP[207],VcascodeP[206],VcascodeP[205],VcascodeP[204],VcascodeP[203],VcascodeP[202],VcascodeP[201],VcascodeP[200],VcascodeP[199],VcascodeP[198],VcascodeP[197],VcascodeP[196],VcascodeP[195],VcascodeP[194],VcascodeP[193],VcascodeP[192],VcascodeP[191],VcascodeP[190],VcascodeP[189],VcascodeP[188],VcascodeP[187],VcascodeP[186],VcascodeP[185],VcascodeP[184],VcascodeP[183],VcascodeP[182],VcascodeP[181],VcascodeP[180],VcascodeP[179],VcascodeP[178],VcascodeP[177],VcascodeP[176],VcascodeP[175],VcascodeP[174],VcascodeP[173],VcascodeP[172],VcascodeP[171],VcascodeP[170],VcascodeP[169],VcascodeP[168],VcascodeP[167],VcascodeP[166],VcascodeP[165],VcascodeP[164],VcascodeP[163],VcascodeP[162],VcascodeP[161],VcascodeP[160],VcascodeP[159],VcascodeP[158],VcascodeP[157],VcascodeP[156],VcascodeP[155],VcascodeP[154],VcascodeP[153],VcascodeP[152],VcascodeP[151],VcascodeP[150],VcascodeP[149],VcascodeP[148],VcascodeP[147],VcascodeP[146],VcascodeP[145],VcascodeP[144],VcascodeP[143],VcascodeP[142],VcascodeP[141],VcascodeP[140],VcascodeP[139],VcascodeP[138],VcascodeP[137],VcascodeP[136],VcascodeP[135],VcascodeP[134],VcascodeP[133],VcascodeP[132],VcascodeP[131],VcascodeP[130],VcascodeP[129],VcascodeP[128],VcascodeP[127],VcascodeP[126],VcascodeP[125],VcascodeP[124],VcascodeP[123],VcascodeP[122],VcascodeP[121],VcascodeP[120],VcascodeP[119],VcascodeP[118],VcascodeP[117],VcascodeP[116],VcascodeP[115],VcascodeP[114],VcascodeP[113],VcascodeP[112],VcascodeP[111],VcascodeP[110],VcascodeP[109],VcascodeP[108],VcascodeP[107],VcascodeP[106],VcascodeP[105],VcascodeP[104],VcascodeP[103],VcascodeP[102],VcascodeP[101],VcascodeP[100],VcascodeP[99],VcascodeP[98],VcascodeP[97],VcascodeP[96],VcascodeP[95],VcascodeP[94],VcascodeP[93],VcascodeP[92],VcascodeP[91],VcascodeP[90],VcascodeP[89],VcascodeP[88],VcascodeP[87],VcascodeP[86],VcascodeP[85],VcascodeP[84],VcascodeP[83],VcascodeP[82],VcascodeP[81],VcascodeP[80],VcascodeP[79],VcascodeP[78],VcascodeP[77],VcascodeP[76],VcascodeP[75],VcascodeP[74],VcascodeP[73],VcascodeP[72],VcascodeP[71],VcascodeP[70],VcascodeP[69],VcascodeP[68],VcascodeP[67],VcascodeP[66],VcascodeP[65],VcascodeP[64],VcascodeP[63],VcascodeP[62],VcascodeP[61],VcascodeP[60],VcascodeP[59],VcascodeP[58],VcascodeP[57],VcascodeP[56],VcascodeP[55],VcascodeP[54],VcascodeP[53],VcascodeP[52],VcascodeP[51],VcascodeP[50],VcascodeP[49],VcascodeP[48],VcascodeP[47],VcascodeP[46],VcascodeP[45],VcascodeP[44],VcascodeP[43],VcascodeP[42],VcascodeP[41],VcascodeP[40],VcascodeP[39],VcascodeP[38],VcascodeP[37],VcascodeP[36],VcascodeP[35],VcascodeP[34],VcascodeP[33],VcascodeP[32],VcascodeP[31],VcascodeP[30],VcascodeP[29],VcascodeP[28],VcascodeP[27],VcascodeP[26],VcascodeP[25],VcascodeP[24],VcascodeP[23],VcascodeP[22],VcascodeP[21],VcascodeP[20],VcascodeP[19],VcascodeP[18],VcascodeP[17],VcascodeP[16],VcascodeP[15],VcascodeP[14],VcascodeP[13],VcascodeP[12],VcascodeP[11],VcascodeP[10],VcascodeP[9],VcascodeP[8],VcascodeP[7],VcascodeP[6],VcascodeP[5],VcascodeP[4],VcascodeP[3],VcascodeP[2],VcascodeP[1],VcascodeP[0]
*.ipin Vbiasp
*.ipin VDD
*.ipin
*+ VcascodeP[255],VcascodeP[254],VcascodeP[253],VcascodeP[252],VcascodeP[251],VcascodeP[250],VcascodeP[249],VcascodeP[248],VcascodeP[247],VcascodeP[246],VcascodeP[245],VcascodeP[244],VcascodeP[243],VcascodeP[242],VcascodeP[241],VcascodeP[240],VcascodeP[239],VcascodeP[238],VcascodeP[237],VcascodeP[236],VcascodeP[235],VcascodeP[234],VcascodeP[233],VcascodeP[232],VcascodeP[231],VcascodeP[230],VcascodeP[229],VcascodeP[228],VcascodeP[227],VcascodeP[226],VcascodeP[225],VcascodeP[224],VcascodeP[223],VcascodeP[222],VcascodeP[221],VcascodeP[220],VcascodeP[219],VcascodeP[218],VcascodeP[217],VcascodeP[216],VcascodeP[215],VcascodeP[214],VcascodeP[213],VcascodeP[212],VcascodeP[211],VcascodeP[210],VcascodeP[209],VcascodeP[208],VcascodeP[207],VcascodeP[206],VcascodeP[205],VcascodeP[204],VcascodeP[203],VcascodeP[202],VcascodeP[201],VcascodeP[200],VcascodeP[199],VcascodeP[198],VcascodeP[197],VcascodeP[196],VcascodeP[195],VcascodeP[194],VcascodeP[193],VcascodeP[192],VcascodeP[191],VcascodeP[190],VcascodeP[189],VcascodeP[188],VcascodeP[187],VcascodeP[186],VcascodeP[185],VcascodeP[184],VcascodeP[183],VcascodeP[182],VcascodeP[181],VcascodeP[180],VcascodeP[179],VcascodeP[178],VcascodeP[177],VcascodeP[176],VcascodeP[175],VcascodeP[174],VcascodeP[173],VcascodeP[172],VcascodeP[171],VcascodeP[170],VcascodeP[169],VcascodeP[168],VcascodeP[167],VcascodeP[166],VcascodeP[165],VcascodeP[164],VcascodeP[163],VcascodeP[162],VcascodeP[161],VcascodeP[160],VcascodeP[159],VcascodeP[158],VcascodeP[157],VcascodeP[156],VcascodeP[155],VcascodeP[154],VcascodeP[153],VcascodeP[152],VcascodeP[151],VcascodeP[150],VcascodeP[149],VcascodeP[148],VcascodeP[147],VcascodeP[146],VcascodeP[145],VcascodeP[144],VcascodeP[143],VcascodeP[142],VcascodeP[141],VcascodeP[140],VcascodeP[139],VcascodeP[138],VcascodeP[137],VcascodeP[136],VcascodeP[135],VcascodeP[134],VcascodeP[133],VcascodeP[132],VcascodeP[131],VcascodeP[130],VcascodeP[129],VcascodeP[128],VcascodeP[127],VcascodeP[126],VcascodeP[125],VcascodeP[124],VcascodeP[123],VcascodeP[122],VcascodeP[121],VcascodeP[120],VcascodeP[119],VcascodeP[118],VcascodeP[117],VcascodeP[116],VcascodeP[115],VcascodeP[114],VcascodeP[113],VcascodeP[112],VcascodeP[111],VcascodeP[110],VcascodeP[109],VcascodeP[108],VcascodeP[107],VcascodeP[106],VcascodeP[105],VcascodeP[104],VcascodeP[103],VcascodeP[102],VcascodeP[101],VcascodeP[100],VcascodeP[99],VcascodeP[98],VcascodeP[97],VcascodeP[96],VcascodeP[95],VcascodeP[94],VcascodeP[93],VcascodeP[92],VcascodeP[91],VcascodeP[90],VcascodeP[89],VcascodeP[88],VcascodeP[87],VcascodeP[86],VcascodeP[85],VcascodeP[84],VcascodeP[83],VcascodeP[82],VcascodeP[81],VcascodeP[80],VcascodeP[79],VcascodeP[78],VcascodeP[77],VcascodeP[76],VcascodeP[75],VcascodeP[74],VcascodeP[73],VcascodeP[72],VcascodeP[71],VcascodeP[70],VcascodeP[69],VcascodeP[68],VcascodeP[67],VcascodeP[66],VcascodeP[65],VcascodeP[64],VcascodeP[63],VcascodeP[62],VcascodeP[61],VcascodeP[60],VcascodeP[59],VcascodeP[58],VcascodeP[57],VcascodeP[56],VcascodeP[55],VcascodeP[54],VcascodeP[53],VcascodeP[52],VcascodeP[51],VcascodeP[50],VcascodeP[49],VcascodeP[48],VcascodeP[47],VcascodeP[46],VcascodeP[45],VcascodeP[44],VcascodeP[43],VcascodeP[42],VcascodeP[41],VcascodeP[40],VcascodeP[39],VcascodeP[38],VcascodeP[37],VcascodeP[36],VcascodeP[35],VcascodeP[34],VcascodeP[33],VcascodeP[32],VcascodeP[31],VcascodeP[30],VcascodeP[29],VcascodeP[28],VcascodeP[27],VcascodeP[26],VcascodeP[25],VcascodeP[24],VcascodeP[23],VcascodeP[22],VcascodeP[21],VcascodeP[20],VcascodeP[19],VcascodeP[18],VcascodeP[17],VcascodeP[16],VcascodeP[15],VcascodeP[14],VcascodeP[13],VcascodeP[12],VcascodeP[11],VcascodeP[10],VcascodeP[9],VcascodeP[8],VcascodeP[7],VcascodeP[6],VcascodeP[5],VcascodeP[4],VcascodeP[3],VcascodeP[2],VcascodeP[1],VcascodeP[0]
*.opin Iout
XI_MIRROR[255] VDD Vbiasp VcascodeP[255] Iout Pmirror_StdCell
XI_MIRROR[254] VDD Vbiasp VcascodeP[254] Iout Pmirror_StdCell
XI_MIRROR[253] VDD Vbiasp VcascodeP[253] Iout Pmirror_StdCell
XI_MIRROR[252] VDD Vbiasp VcascodeP[252] Iout Pmirror_StdCell
XI_MIRROR[251] VDD Vbiasp VcascodeP[251] Iout Pmirror_StdCell
XI_MIRROR[250] VDD Vbiasp VcascodeP[250] Iout Pmirror_StdCell
XI_MIRROR[249] VDD Vbiasp VcascodeP[249] Iout Pmirror_StdCell
XI_MIRROR[248] VDD Vbiasp VcascodeP[248] Iout Pmirror_StdCell
XI_MIRROR[247] VDD Vbiasp VcascodeP[247] Iout Pmirror_StdCell
XI_MIRROR[246] VDD Vbiasp VcascodeP[246] Iout Pmirror_StdCell
XI_MIRROR[245] VDD Vbiasp VcascodeP[245] Iout Pmirror_StdCell
XI_MIRROR[244] VDD Vbiasp VcascodeP[244] Iout Pmirror_StdCell
XI_MIRROR[243] VDD Vbiasp VcascodeP[243] Iout Pmirror_StdCell
XI_MIRROR[242] VDD Vbiasp VcascodeP[242] Iout Pmirror_StdCell
XI_MIRROR[241] VDD Vbiasp VcascodeP[241] Iout Pmirror_StdCell
XI_MIRROR[240] VDD Vbiasp VcascodeP[240] Iout Pmirror_StdCell
XI_MIRROR[239] VDD Vbiasp VcascodeP[239] Iout Pmirror_StdCell
XI_MIRROR[238] VDD Vbiasp VcascodeP[238] Iout Pmirror_StdCell
XI_MIRROR[237] VDD Vbiasp VcascodeP[237] Iout Pmirror_StdCell
XI_MIRROR[236] VDD Vbiasp VcascodeP[236] Iout Pmirror_StdCell
XI_MIRROR[235] VDD Vbiasp VcascodeP[235] Iout Pmirror_StdCell
XI_MIRROR[234] VDD Vbiasp VcascodeP[234] Iout Pmirror_StdCell
XI_MIRROR[233] VDD Vbiasp VcascodeP[233] Iout Pmirror_StdCell
XI_MIRROR[232] VDD Vbiasp VcascodeP[232] Iout Pmirror_StdCell
XI_MIRROR[231] VDD Vbiasp VcascodeP[231] Iout Pmirror_StdCell
XI_MIRROR[230] VDD Vbiasp VcascodeP[230] Iout Pmirror_StdCell
XI_MIRROR[229] VDD Vbiasp VcascodeP[229] Iout Pmirror_StdCell
XI_MIRROR[228] VDD Vbiasp VcascodeP[228] Iout Pmirror_StdCell
XI_MIRROR[227] VDD Vbiasp VcascodeP[227] Iout Pmirror_StdCell
XI_MIRROR[226] VDD Vbiasp VcascodeP[226] Iout Pmirror_StdCell
XI_MIRROR[225] VDD Vbiasp VcascodeP[225] Iout Pmirror_StdCell
XI_MIRROR[224] VDD Vbiasp VcascodeP[224] Iout Pmirror_StdCell
XI_MIRROR[223] VDD Vbiasp VcascodeP[223] Iout Pmirror_StdCell
XI_MIRROR[222] VDD Vbiasp VcascodeP[222] Iout Pmirror_StdCell
XI_MIRROR[221] VDD Vbiasp VcascodeP[221] Iout Pmirror_StdCell
XI_MIRROR[220] VDD Vbiasp VcascodeP[220] Iout Pmirror_StdCell
XI_MIRROR[219] VDD Vbiasp VcascodeP[219] Iout Pmirror_StdCell
XI_MIRROR[218] VDD Vbiasp VcascodeP[218] Iout Pmirror_StdCell
XI_MIRROR[217] VDD Vbiasp VcascodeP[217] Iout Pmirror_StdCell
XI_MIRROR[216] VDD Vbiasp VcascodeP[216] Iout Pmirror_StdCell
XI_MIRROR[215] VDD Vbiasp VcascodeP[215] Iout Pmirror_StdCell
XI_MIRROR[214] VDD Vbiasp VcascodeP[214] Iout Pmirror_StdCell
XI_MIRROR[213] VDD Vbiasp VcascodeP[213] Iout Pmirror_StdCell
XI_MIRROR[212] VDD Vbiasp VcascodeP[212] Iout Pmirror_StdCell
XI_MIRROR[211] VDD Vbiasp VcascodeP[211] Iout Pmirror_StdCell
XI_MIRROR[210] VDD Vbiasp VcascodeP[210] Iout Pmirror_StdCell
XI_MIRROR[209] VDD Vbiasp VcascodeP[209] Iout Pmirror_StdCell
XI_MIRROR[208] VDD Vbiasp VcascodeP[208] Iout Pmirror_StdCell
XI_MIRROR[207] VDD Vbiasp VcascodeP[207] Iout Pmirror_StdCell
XI_MIRROR[206] VDD Vbiasp VcascodeP[206] Iout Pmirror_StdCell
XI_MIRROR[205] VDD Vbiasp VcascodeP[205] Iout Pmirror_StdCell
XI_MIRROR[204] VDD Vbiasp VcascodeP[204] Iout Pmirror_StdCell
XI_MIRROR[203] VDD Vbiasp VcascodeP[203] Iout Pmirror_StdCell
XI_MIRROR[202] VDD Vbiasp VcascodeP[202] Iout Pmirror_StdCell
XI_MIRROR[201] VDD Vbiasp VcascodeP[201] Iout Pmirror_StdCell
XI_MIRROR[200] VDD Vbiasp VcascodeP[200] Iout Pmirror_StdCell
XI_MIRROR[199] VDD Vbiasp VcascodeP[199] Iout Pmirror_StdCell
XI_MIRROR[198] VDD Vbiasp VcascodeP[198] Iout Pmirror_StdCell
XI_MIRROR[197] VDD Vbiasp VcascodeP[197] Iout Pmirror_StdCell
XI_MIRROR[196] VDD Vbiasp VcascodeP[196] Iout Pmirror_StdCell
XI_MIRROR[195] VDD Vbiasp VcascodeP[195] Iout Pmirror_StdCell
XI_MIRROR[194] VDD Vbiasp VcascodeP[194] Iout Pmirror_StdCell
XI_MIRROR[193] VDD Vbiasp VcascodeP[193] Iout Pmirror_StdCell
XI_MIRROR[192] VDD Vbiasp VcascodeP[192] Iout Pmirror_StdCell
XI_MIRROR[191] VDD Vbiasp VcascodeP[191] Iout Pmirror_StdCell
XI_MIRROR[190] VDD Vbiasp VcascodeP[190] Iout Pmirror_StdCell
XI_MIRROR[189] VDD Vbiasp VcascodeP[189] Iout Pmirror_StdCell
XI_MIRROR[188] VDD Vbiasp VcascodeP[188] Iout Pmirror_StdCell
XI_MIRROR[187] VDD Vbiasp VcascodeP[187] Iout Pmirror_StdCell
XI_MIRROR[186] VDD Vbiasp VcascodeP[186] Iout Pmirror_StdCell
XI_MIRROR[185] VDD Vbiasp VcascodeP[185] Iout Pmirror_StdCell
XI_MIRROR[184] VDD Vbiasp VcascodeP[184] Iout Pmirror_StdCell
XI_MIRROR[183] VDD Vbiasp VcascodeP[183] Iout Pmirror_StdCell
XI_MIRROR[182] VDD Vbiasp VcascodeP[182] Iout Pmirror_StdCell
XI_MIRROR[181] VDD Vbiasp VcascodeP[181] Iout Pmirror_StdCell
XI_MIRROR[180] VDD Vbiasp VcascodeP[180] Iout Pmirror_StdCell
XI_MIRROR[179] VDD Vbiasp VcascodeP[179] Iout Pmirror_StdCell
XI_MIRROR[178] VDD Vbiasp VcascodeP[178] Iout Pmirror_StdCell
XI_MIRROR[177] VDD Vbiasp VcascodeP[177] Iout Pmirror_StdCell
XI_MIRROR[176] VDD Vbiasp VcascodeP[176] Iout Pmirror_StdCell
XI_MIRROR[175] VDD Vbiasp VcascodeP[175] Iout Pmirror_StdCell
XI_MIRROR[174] VDD Vbiasp VcascodeP[174] Iout Pmirror_StdCell
XI_MIRROR[173] VDD Vbiasp VcascodeP[173] Iout Pmirror_StdCell
XI_MIRROR[172] VDD Vbiasp VcascodeP[172] Iout Pmirror_StdCell
XI_MIRROR[171] VDD Vbiasp VcascodeP[171] Iout Pmirror_StdCell
XI_MIRROR[170] VDD Vbiasp VcascodeP[170] Iout Pmirror_StdCell
XI_MIRROR[169] VDD Vbiasp VcascodeP[169] Iout Pmirror_StdCell
XI_MIRROR[168] VDD Vbiasp VcascodeP[168] Iout Pmirror_StdCell
XI_MIRROR[167] VDD Vbiasp VcascodeP[167] Iout Pmirror_StdCell
XI_MIRROR[166] VDD Vbiasp VcascodeP[166] Iout Pmirror_StdCell
XI_MIRROR[165] VDD Vbiasp VcascodeP[165] Iout Pmirror_StdCell
XI_MIRROR[164] VDD Vbiasp VcascodeP[164] Iout Pmirror_StdCell
XI_MIRROR[163] VDD Vbiasp VcascodeP[163] Iout Pmirror_StdCell
XI_MIRROR[162] VDD Vbiasp VcascodeP[162] Iout Pmirror_StdCell
XI_MIRROR[161] VDD Vbiasp VcascodeP[161] Iout Pmirror_StdCell
XI_MIRROR[160] VDD Vbiasp VcascodeP[160] Iout Pmirror_StdCell
XI_MIRROR[159] VDD Vbiasp VcascodeP[159] Iout Pmirror_StdCell
XI_MIRROR[158] VDD Vbiasp VcascodeP[158] Iout Pmirror_StdCell
XI_MIRROR[157] VDD Vbiasp VcascodeP[157] Iout Pmirror_StdCell
XI_MIRROR[156] VDD Vbiasp VcascodeP[156] Iout Pmirror_StdCell
XI_MIRROR[155] VDD Vbiasp VcascodeP[155] Iout Pmirror_StdCell
XI_MIRROR[154] VDD Vbiasp VcascodeP[154] Iout Pmirror_StdCell
XI_MIRROR[153] VDD Vbiasp VcascodeP[153] Iout Pmirror_StdCell
XI_MIRROR[152] VDD Vbiasp VcascodeP[152] Iout Pmirror_StdCell
XI_MIRROR[151] VDD Vbiasp VcascodeP[151] Iout Pmirror_StdCell
XI_MIRROR[150] VDD Vbiasp VcascodeP[150] Iout Pmirror_StdCell
XI_MIRROR[149] VDD Vbiasp VcascodeP[149] Iout Pmirror_StdCell
XI_MIRROR[148] VDD Vbiasp VcascodeP[148] Iout Pmirror_StdCell
XI_MIRROR[147] VDD Vbiasp VcascodeP[147] Iout Pmirror_StdCell
XI_MIRROR[146] VDD Vbiasp VcascodeP[146] Iout Pmirror_StdCell
XI_MIRROR[145] VDD Vbiasp VcascodeP[145] Iout Pmirror_StdCell
XI_MIRROR[144] VDD Vbiasp VcascodeP[144] Iout Pmirror_StdCell
XI_MIRROR[143] VDD Vbiasp VcascodeP[143] Iout Pmirror_StdCell
XI_MIRROR[142] VDD Vbiasp VcascodeP[142] Iout Pmirror_StdCell
XI_MIRROR[141] VDD Vbiasp VcascodeP[141] Iout Pmirror_StdCell
XI_MIRROR[140] VDD Vbiasp VcascodeP[140] Iout Pmirror_StdCell
XI_MIRROR[139] VDD Vbiasp VcascodeP[139] Iout Pmirror_StdCell
XI_MIRROR[138] VDD Vbiasp VcascodeP[138] Iout Pmirror_StdCell
XI_MIRROR[137] VDD Vbiasp VcascodeP[137] Iout Pmirror_StdCell
XI_MIRROR[136] VDD Vbiasp VcascodeP[136] Iout Pmirror_StdCell
XI_MIRROR[135] VDD Vbiasp VcascodeP[135] Iout Pmirror_StdCell
XI_MIRROR[134] VDD Vbiasp VcascodeP[134] Iout Pmirror_StdCell
XI_MIRROR[133] VDD Vbiasp VcascodeP[133] Iout Pmirror_StdCell
XI_MIRROR[132] VDD Vbiasp VcascodeP[132] Iout Pmirror_StdCell
XI_MIRROR[131] VDD Vbiasp VcascodeP[131] Iout Pmirror_StdCell
XI_MIRROR[130] VDD Vbiasp VcascodeP[130] Iout Pmirror_StdCell
XI_MIRROR[129] VDD Vbiasp VcascodeP[129] Iout Pmirror_StdCell
XI_MIRROR[128] VDD Vbiasp VcascodeP[128] Iout Pmirror_StdCell
XI_MIRROR[127] VDD Vbiasp VcascodeP[127] Iout Pmirror_StdCell
XI_MIRROR[126] VDD Vbiasp VcascodeP[126] Iout Pmirror_StdCell
XI_MIRROR[125] VDD Vbiasp VcascodeP[125] Iout Pmirror_StdCell
XI_MIRROR[124] VDD Vbiasp VcascodeP[124] Iout Pmirror_StdCell
XI_MIRROR[123] VDD Vbiasp VcascodeP[123] Iout Pmirror_StdCell
XI_MIRROR[122] VDD Vbiasp VcascodeP[122] Iout Pmirror_StdCell
XI_MIRROR[121] VDD Vbiasp VcascodeP[121] Iout Pmirror_StdCell
XI_MIRROR[120] VDD Vbiasp VcascodeP[120] Iout Pmirror_StdCell
XI_MIRROR[119] VDD Vbiasp VcascodeP[119] Iout Pmirror_StdCell
XI_MIRROR[118] VDD Vbiasp VcascodeP[118] Iout Pmirror_StdCell
XI_MIRROR[117] VDD Vbiasp VcascodeP[117] Iout Pmirror_StdCell
XI_MIRROR[116] VDD Vbiasp VcascodeP[116] Iout Pmirror_StdCell
XI_MIRROR[115] VDD Vbiasp VcascodeP[115] Iout Pmirror_StdCell
XI_MIRROR[114] VDD Vbiasp VcascodeP[114] Iout Pmirror_StdCell
XI_MIRROR[113] VDD Vbiasp VcascodeP[113] Iout Pmirror_StdCell
XI_MIRROR[112] VDD Vbiasp VcascodeP[112] Iout Pmirror_StdCell
XI_MIRROR[111] VDD Vbiasp VcascodeP[111] Iout Pmirror_StdCell
XI_MIRROR[110] VDD Vbiasp VcascodeP[110] Iout Pmirror_StdCell
XI_MIRROR[109] VDD Vbiasp VcascodeP[109] Iout Pmirror_StdCell
XI_MIRROR[108] VDD Vbiasp VcascodeP[108] Iout Pmirror_StdCell
XI_MIRROR[107] VDD Vbiasp VcascodeP[107] Iout Pmirror_StdCell
XI_MIRROR[106] VDD Vbiasp VcascodeP[106] Iout Pmirror_StdCell
XI_MIRROR[105] VDD Vbiasp VcascodeP[105] Iout Pmirror_StdCell
XI_MIRROR[104] VDD Vbiasp VcascodeP[104] Iout Pmirror_StdCell
XI_MIRROR[103] VDD Vbiasp VcascodeP[103] Iout Pmirror_StdCell
XI_MIRROR[102] VDD Vbiasp VcascodeP[102] Iout Pmirror_StdCell
XI_MIRROR[101] VDD Vbiasp VcascodeP[101] Iout Pmirror_StdCell
XI_MIRROR[100] VDD Vbiasp VcascodeP[100] Iout Pmirror_StdCell
XI_MIRROR[99] VDD Vbiasp VcascodeP[99] Iout Pmirror_StdCell
XI_MIRROR[98] VDD Vbiasp VcascodeP[98] Iout Pmirror_StdCell
XI_MIRROR[97] VDD Vbiasp VcascodeP[97] Iout Pmirror_StdCell
XI_MIRROR[96] VDD Vbiasp VcascodeP[96] Iout Pmirror_StdCell
XI_MIRROR[95] VDD Vbiasp VcascodeP[95] Iout Pmirror_StdCell
XI_MIRROR[94] VDD Vbiasp VcascodeP[94] Iout Pmirror_StdCell
XI_MIRROR[93] VDD Vbiasp VcascodeP[93] Iout Pmirror_StdCell
XI_MIRROR[92] VDD Vbiasp VcascodeP[92] Iout Pmirror_StdCell
XI_MIRROR[91] VDD Vbiasp VcascodeP[91] Iout Pmirror_StdCell
XI_MIRROR[90] VDD Vbiasp VcascodeP[90] Iout Pmirror_StdCell
XI_MIRROR[89] VDD Vbiasp VcascodeP[89] Iout Pmirror_StdCell
XI_MIRROR[88] VDD Vbiasp VcascodeP[88] Iout Pmirror_StdCell
XI_MIRROR[87] VDD Vbiasp VcascodeP[87] Iout Pmirror_StdCell
XI_MIRROR[86] VDD Vbiasp VcascodeP[86] Iout Pmirror_StdCell
XI_MIRROR[85] VDD Vbiasp VcascodeP[85] Iout Pmirror_StdCell
XI_MIRROR[84] VDD Vbiasp VcascodeP[84] Iout Pmirror_StdCell
XI_MIRROR[83] VDD Vbiasp VcascodeP[83] Iout Pmirror_StdCell
XI_MIRROR[82] VDD Vbiasp VcascodeP[82] Iout Pmirror_StdCell
XI_MIRROR[81] VDD Vbiasp VcascodeP[81] Iout Pmirror_StdCell
XI_MIRROR[80] VDD Vbiasp VcascodeP[80] Iout Pmirror_StdCell
XI_MIRROR[79] VDD Vbiasp VcascodeP[79] Iout Pmirror_StdCell
XI_MIRROR[78] VDD Vbiasp VcascodeP[78] Iout Pmirror_StdCell
XI_MIRROR[77] VDD Vbiasp VcascodeP[77] Iout Pmirror_StdCell
XI_MIRROR[76] VDD Vbiasp VcascodeP[76] Iout Pmirror_StdCell
XI_MIRROR[75] VDD Vbiasp VcascodeP[75] Iout Pmirror_StdCell
XI_MIRROR[74] VDD Vbiasp VcascodeP[74] Iout Pmirror_StdCell
XI_MIRROR[73] VDD Vbiasp VcascodeP[73] Iout Pmirror_StdCell
XI_MIRROR[72] VDD Vbiasp VcascodeP[72] Iout Pmirror_StdCell
XI_MIRROR[71] VDD Vbiasp VcascodeP[71] Iout Pmirror_StdCell
XI_MIRROR[70] VDD Vbiasp VcascodeP[70] Iout Pmirror_StdCell
XI_MIRROR[69] VDD Vbiasp VcascodeP[69] Iout Pmirror_StdCell
XI_MIRROR[68] VDD Vbiasp VcascodeP[68] Iout Pmirror_StdCell
XI_MIRROR[67] VDD Vbiasp VcascodeP[67] Iout Pmirror_StdCell
XI_MIRROR[66] VDD Vbiasp VcascodeP[66] Iout Pmirror_StdCell
XI_MIRROR[65] VDD Vbiasp VcascodeP[65] Iout Pmirror_StdCell
XI_MIRROR[64] VDD Vbiasp VcascodeP[64] Iout Pmirror_StdCell
XI_MIRROR[63] VDD Vbiasp VcascodeP[63] Iout Pmirror_StdCell
XI_MIRROR[62] VDD Vbiasp VcascodeP[62] Iout Pmirror_StdCell
XI_MIRROR[61] VDD Vbiasp VcascodeP[61] Iout Pmirror_StdCell
XI_MIRROR[60] VDD Vbiasp VcascodeP[60] Iout Pmirror_StdCell
XI_MIRROR[59] VDD Vbiasp VcascodeP[59] Iout Pmirror_StdCell
XI_MIRROR[58] VDD Vbiasp VcascodeP[58] Iout Pmirror_StdCell
XI_MIRROR[57] VDD Vbiasp VcascodeP[57] Iout Pmirror_StdCell
XI_MIRROR[56] VDD Vbiasp VcascodeP[56] Iout Pmirror_StdCell
XI_MIRROR[55] VDD Vbiasp VcascodeP[55] Iout Pmirror_StdCell
XI_MIRROR[54] VDD Vbiasp VcascodeP[54] Iout Pmirror_StdCell
XI_MIRROR[53] VDD Vbiasp VcascodeP[53] Iout Pmirror_StdCell
XI_MIRROR[52] VDD Vbiasp VcascodeP[52] Iout Pmirror_StdCell
XI_MIRROR[51] VDD Vbiasp VcascodeP[51] Iout Pmirror_StdCell
XI_MIRROR[50] VDD Vbiasp VcascodeP[50] Iout Pmirror_StdCell
XI_MIRROR[49] VDD Vbiasp VcascodeP[49] Iout Pmirror_StdCell
XI_MIRROR[48] VDD Vbiasp VcascodeP[48] Iout Pmirror_StdCell
XI_MIRROR[47] VDD Vbiasp VcascodeP[47] Iout Pmirror_StdCell
XI_MIRROR[46] VDD Vbiasp VcascodeP[46] Iout Pmirror_StdCell
XI_MIRROR[45] VDD Vbiasp VcascodeP[45] Iout Pmirror_StdCell
XI_MIRROR[44] VDD Vbiasp VcascodeP[44] Iout Pmirror_StdCell
XI_MIRROR[43] VDD Vbiasp VcascodeP[43] Iout Pmirror_StdCell
XI_MIRROR[42] VDD Vbiasp VcascodeP[42] Iout Pmirror_StdCell
XI_MIRROR[41] VDD Vbiasp VcascodeP[41] Iout Pmirror_StdCell
XI_MIRROR[40] VDD Vbiasp VcascodeP[40] Iout Pmirror_StdCell
XI_MIRROR[39] VDD Vbiasp VcascodeP[39] Iout Pmirror_StdCell
XI_MIRROR[38] VDD Vbiasp VcascodeP[38] Iout Pmirror_StdCell
XI_MIRROR[37] VDD Vbiasp VcascodeP[37] Iout Pmirror_StdCell
XI_MIRROR[36] VDD Vbiasp VcascodeP[36] Iout Pmirror_StdCell
XI_MIRROR[35] VDD Vbiasp VcascodeP[35] Iout Pmirror_StdCell
XI_MIRROR[34] VDD Vbiasp VcascodeP[34] Iout Pmirror_StdCell
XI_MIRROR[33] VDD Vbiasp VcascodeP[33] Iout Pmirror_StdCell
XI_MIRROR[32] VDD Vbiasp VcascodeP[32] Iout Pmirror_StdCell
XI_MIRROR[31] VDD Vbiasp VcascodeP[31] Iout Pmirror_StdCell
XI_MIRROR[30] VDD Vbiasp VcascodeP[30] Iout Pmirror_StdCell
XI_MIRROR[29] VDD Vbiasp VcascodeP[29] Iout Pmirror_StdCell
XI_MIRROR[28] VDD Vbiasp VcascodeP[28] Iout Pmirror_StdCell
XI_MIRROR[27] VDD Vbiasp VcascodeP[27] Iout Pmirror_StdCell
XI_MIRROR[26] VDD Vbiasp VcascodeP[26] Iout Pmirror_StdCell
XI_MIRROR[25] VDD Vbiasp VcascodeP[25] Iout Pmirror_StdCell
XI_MIRROR[24] VDD Vbiasp VcascodeP[24] Iout Pmirror_StdCell
XI_MIRROR[23] VDD Vbiasp VcascodeP[23] Iout Pmirror_StdCell
XI_MIRROR[22] VDD Vbiasp VcascodeP[22] Iout Pmirror_StdCell
XI_MIRROR[21] VDD Vbiasp VcascodeP[21] Iout Pmirror_StdCell
XI_MIRROR[20] VDD Vbiasp VcascodeP[20] Iout Pmirror_StdCell
XI_MIRROR[19] VDD Vbiasp VcascodeP[19] Iout Pmirror_StdCell
XI_MIRROR[18] VDD Vbiasp VcascodeP[18] Iout Pmirror_StdCell
XI_MIRROR[17] VDD Vbiasp VcascodeP[17] Iout Pmirror_StdCell
XI_MIRROR[16] VDD Vbiasp VcascodeP[16] Iout Pmirror_StdCell
XI_MIRROR[15] VDD Vbiasp VcascodeP[15] Iout Pmirror_StdCell
XI_MIRROR[14] VDD Vbiasp VcascodeP[14] Iout Pmirror_StdCell
XI_MIRROR[13] VDD Vbiasp VcascodeP[13] Iout Pmirror_StdCell
XI_MIRROR[12] VDD Vbiasp VcascodeP[12] Iout Pmirror_StdCell
XI_MIRROR[11] VDD Vbiasp VcascodeP[11] Iout Pmirror_StdCell
XI_MIRROR[10] VDD Vbiasp VcascodeP[10] Iout Pmirror_StdCell
XI_MIRROR[9] VDD Vbiasp VcascodeP[9] Iout Pmirror_StdCell
XI_MIRROR[8] VDD Vbiasp VcascodeP[8] Iout Pmirror_StdCell
XI_MIRROR[7] VDD Vbiasp VcascodeP[7] Iout Pmirror_StdCell
XI_MIRROR[6] VDD Vbiasp VcascodeP[6] Iout Pmirror_StdCell
XI_MIRROR[5] VDD Vbiasp VcascodeP[5] Iout Pmirror_StdCell
XI_MIRROR[4] VDD Vbiasp VcascodeP[4] Iout Pmirror_StdCell
XI_MIRROR[3] VDD Vbiasp VcascodeP[3] Iout Pmirror_StdCell
XI_MIRROR[2] VDD Vbiasp VcascodeP[2] Iout Pmirror_StdCell
XI_MIRROR[1] VDD Vbiasp VcascodeP[1] Iout Pmirror_StdCell
XI_MIRROR[0] VDD Vbiasp VcascodeP[0] Iout Pmirror_StdCell
**.ends

* expanding   symbol:  /home/user/PUDDING/schematic/Pmirror_StdCell.sym # of pins=4
** sym_path: /home/user/PUDDING/schematic/Pmirror_StdCell.sym
** sch_path: /home/user/PUDDING/schematic/Pmirror_StdCell.sch
.subckt Pmirror_StdCell VDD VbiasP VcascodeP Iout
*.ipin VcascodeP
*.ipin VbiasP
*.opin Iout
*.ipin VDD
XM2 net1 VbiasP VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 Iout VcascodeP net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends

.end
