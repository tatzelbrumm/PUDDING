magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771122832
<< metal1 >>
rect -70 61 70 70
rect -70 -61 -61 61
rect 61 -61 70 61
rect -70 -70 70 -61
<< via1 >>
rect -61 -61 61 61
<< metal2 >>
rect -70 61 70 70
rect -70 -61 -61 61
rect 61 -61 70 61
rect -70 -70 70 -61
<< via2 >>
rect -61 -61 61 61
<< metal3 >>
rect -70 61 70 70
rect -70 -61 -61 61
rect 61 -61 70 61
rect -70 -70 70 -61
<< end >>
